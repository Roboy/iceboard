// Verilog netlist produced by program LSE :  version Diamond Version 0.0.0
// Netlist written on Fri Oct  4 18:55:36 2019
//
// Verilog Description of module TinyFPGA_B
//

module TinyFPGA_B (CLK, LED, USBPU, PIN_1, PIN_2, PIN_3, PIN_4, 
            PIN_5, PIN_6, PIN_7, PIN_8, PIN_9, PIN_10, PIN_11, 
            PIN_12, PIN_13, PIN_14, PIN_15, PIN_16, PIN_17, PIN_18, 
            PIN_19, PIN_20, PIN_21, PIN_22, PIN_23, PIN_24) /* synthesis syn_preserve=0, syn_noprune=0, syn_module_defined=1 */ ;   // verilog/TinyFPGA_B.v(2[8:18])
    input CLK;   // verilog/TinyFPGA_B.v(3[9:12])
    output LED;   // verilog/TinyFPGA_B.v(4[10:13])
    output USBPU;   // verilog/TinyFPGA_B.v(5[10:15])
    input PIN_1 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(6[9:14])
    input PIN_2 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(7[9:14])
    input PIN_3 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(8[9:14])
    input PIN_4 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(9[9:14])
    input PIN_5 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(10[9:14])
    output PIN_6 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(11[9:14])
    output PIN_7 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(12[9:14])
    output PIN_8 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(13[9:14])
    output PIN_9 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(14[9:14])
    output PIN_10 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(15[9:15])
    output PIN_11 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(16[9:15])
    inout PIN_12 /* synthesis black_box_pad_pin=1 */ ;   // verilog/TinyFPGA_B.v(17[9:15])
    input PIN_13 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(18[9:15])
    input PIN_14 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(19[9:15])
    input PIN_15 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(20[9:15])
    input PIN_16 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(21[9:15])
    input PIN_17 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(22[9:15])
    input PIN_18 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(23[9:15])
    input PIN_19 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(24[9:15])
    inout PIN_20 /* synthesis black_box_pad_pin=1 */ ;   // verilog/TinyFPGA_B.v(25[9:15])
    inout PIN_21 /* synthesis black_box_pad_pin=1 */ ;   // verilog/TinyFPGA_B.v(26[9:15])
    inout PIN_22 /* synthesis black_box_pad_pin=1 */ ;   // verilog/TinyFPGA_B.v(27[9:15])
    input PIN_23 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(28[9:15])
    input PIN_24 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(29[9:15])
    
    wire clk32MHz /* synthesis SET_AS_NETWORK=clk32MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(34[8:16])
    
    wire GND_net, VCC_net, CLK_c, LED_c, PIN_6_c_0, PIN_7_c_1, PIN_8_c_2, 
        PIN_9_c_3, PIN_10_c_4, PIN_11_c_5, PIN_13_c, PIN_18_c_1, PIN_19_c_0, 
        PIN_23_c_1, PIN_24_c_0, tx_o, tx_enable;
    wire [23:0]encoder0_position;   // verilog/TinyFPGA_B.v(55[22:39])
    wire [23:0]encoder1_position;   // verilog/TinyFPGA_B.v(56[22:39])
    wire [23:0]displacement;   // verilog/TinyFPGA_B.v(57[21:33])
    wire [23:0]setpoint;   // verilog/TinyFPGA_B.v(58[22:30])
    
    wire n45634;
    wire [23:0]Kp;   // verilog/TinyFPGA_B.v(59[22:24])
    wire [23:0]Ki;   // verilog/TinyFPGA_B.v(60[22:24])
    wire [23:0]Kd;   // verilog/TinyFPGA_B.v(61[22:24])
    wire [7:0]control_mode;   // verilog/TinyFPGA_B.v(62[14:26])
    wire [23:0]PWMLimit;   // verilog/TinyFPGA_B.v(63[22:30])
    wire [23:0]IntegralLimit;   // verilog/TinyFPGA_B.v(64[22:35])
    wire [23:0]deadband;   // verilog/TinyFPGA_B.v(65[22:30])
    wire [23:0]gearBoxRatio;   // verilog/TinyFPGA_B.v(66[22:34])
    
    wire hall1, hall2, hall3;
    wire [23:0]pwm;   // verilog/TinyFPGA_B.v(74[10:13])
    wire [31:0]motor_state;   // verilog/TinyFPGA_B.v(134[22:33])
    
    wire PIN_13_N_26, n45172, n44550, n34801, n2281;
    wire [31:0]motor_state_23__N_27;
    wire [24:0]displacement_23__N_93;
    wire [23:0]displacement_23__N_1;
    
    wire n45181, n34800, n34479, n34799, n34478, n34798, n34477, 
        n34476, n34475, rx_data_ready;
    wire [7:0]rx_data;   // verilog/coms.v(89[13:20])
    wire [7:0]\data_in[3] ;   // verilog/coms.v(93[12:19])
    wire [7:0]\data_in[2] ;   // verilog/coms.v(93[12:19])
    wire [7:0]\data_in[1] ;   // verilog/coms.v(93[12:19])
    wire [7:0]\data_in[0] ;   // verilog/coms.v(93[12:19])
    
    wire n34797, n46887, n34474, n34796;
    wire [7:0]\data_in_frame[21] ;   // verilog/coms.v(94[12:25])
    wire [7:0]\data_in_frame[19] ;   // verilog/coms.v(94[12:25])
    wire [7:0]\data_in_frame[18] ;   // verilog/coms.v(94[12:25])
    wire [7:0]\data_in_frame[17] ;   // verilog/coms.v(94[12:25])
    wire [7:0]\data_in_frame[13] ;   // verilog/coms.v(94[12:25])
    wire [7:0]\data_in_frame[12] ;   // verilog/coms.v(94[12:25])
    wire [7:0]\data_in_frame[11] ;   // verilog/coms.v(94[12:25])
    wire [7:0]\data_in_frame[10] ;   // verilog/coms.v(94[12:25])
    wire [7:0]\data_in_frame[9] ;   // verilog/coms.v(94[12:25])
    wire [7:0]\data_in_frame[8] ;   // verilog/coms.v(94[12:25])
    wire [7:0]\data_in_frame[7] ;   // verilog/coms.v(94[12:25])
    wire [7:0]\data_in_frame[6] ;   // verilog/coms.v(94[12:25])
    wire [7:0]\data_in_frame[5] ;   // verilog/coms.v(94[12:25])
    wire [7:0]\data_in_frame[4] ;   // verilog/coms.v(94[12:25])
    wire [7:0]\data_in_frame[3] ;   // verilog/coms.v(94[12:25])
    wire [7:0]\data_in_frame[2] ;   // verilog/coms.v(94[12:25])
    wire [7:0]\data_in_frame[1] ;   // verilog/coms.v(94[12:25])
    wire [7:0]\data_out_frame[22] ;   // verilog/coms.v(95[12:26])
    wire [7:0]\data_out_frame[21] ;   // verilog/coms.v(95[12:26])
    wire [7:0]\data_out_frame[20] ;   // verilog/coms.v(95[12:26])
    wire [7:0]\data_out_frame[19] ;   // verilog/coms.v(95[12:26])
    wire [7:0]\data_out_frame[18] ;   // verilog/coms.v(95[12:26])
    wire [7:0]\data_out_frame[5] ;   // verilog/coms.v(95[12:26])
    
    wire n34795, n45739, n45215;
    wire [7:0]\data_out_frame[0] ;   // verilog/coms.v(95[12:26])
    wire [7:0]byte_transmit_counter;   // verilog/coms.v(100[12:33])
    
    wire n27220, n34794, n249, n248, n34793, n34792, n34791, n34790, 
        n34789, n45162, n34788, n45160, n45156, n34787, n45154, 
        n34786, n45655, n34785, n34784, n34783, n45150, n45148, 
        n34782, n34781, n34780, n34779, n34778, n6, n4, n2, 
        n34777, n34776, n34775, n34774, n24158, n2280, n44526, 
        n2279, n35122, n35121, n35120, n35119, n35118, n34773, 
        n34772, n34771, n34770, n34769, n34768, n34767, n34766, 
        n46083, n46203, n34765, n34764, n34763, n34762, n34761, 
        n34760, n34759, n34758, n35117, n34757, n34756, n34755, 
        n34754, n34753, n35116, n34752, n34751, n45140, n34750, 
        n35115, n44517, n45138, n44493, n34749, n34748, n4_adj_3956, 
        n45134, n35114, n35113, n35112, n35111, n35110, n35109, 
        n27212, n35108, n35107, n35106, n34747, n24172, n24171, 
        n35105, n6929, n34746, n24120, n24119, n24118, n22463, 
        n24117, n2_adj_3957, n22460, n34745, n24116, n24115, n24114, 
        n34744, n22457, n22454, n34743, n2_adj_3958, n22451, n45106, 
        n34742, n34741, n34740, n34739, n35104, n35103, n34738, 
        n22448, n40216, n45658, n45091, n35102, n35101, n35100, 
        n35099, n34737, n22445, n34736, n34735, n34734, n35098, 
        n34733, n46109, n34732, n34731, n35097, n35096, n35095, 
        n35094, n22442, n35093, n35092, n24113, n35091, n35090, 
        n35089, n22439, n35088, n35087, n35086, n35085, n35084, 
        n35083, n35082, n35081, n35080, n35079, n35078, n22436, 
        n35077, n24112, n24111, n22433, n24110, n22430, n24109, 
        n22427, n24108, n24107, n22424, n45059, n2278, n2277, 
        n2250, n2249, n2248, n2247, n2246, n2245, n2244, n2243, 
        n2242, n2241, n2240, n2239, n2238, n44486, n24106, n24105, 
        n24104, n24103, n24102, n24101, n22421, n24100, n24099, 
        n24098, n24097, n24096, n24095, n22418, n40207, n24094, 
        n24093, n24149, n24150, n24151, n46201, n45041, n27725, 
        n34700, n34699, n34698, n34697, n34696, n34695, n34694, 
        Kp_23__N_516, n45021, n45690, n22415, n24092, n25455, n44470, 
        n44468, n28231, n28263, n24091, n22412, n24090, n24089, 
        n35010, n35009, n35008, n35007, n24144, n35006, n35005, 
        n35004, n35003, n1, n44464, n44462, n45478, n35002, n35001, 
        n35000, n34999, n34998, n34997, n34996, n34995, n34994, 
        n34993, n34992, n23930, n23929, n23928, n23927, n23926, 
        n23925, n23924, n23923, n23914, n23913, n23912, n23911, 
        n23910, n23909, n23908, n23907, n23898, n23897, n23896, 
        n23895, n23894, n23893, n23892, n23891, n23866, n23865, 
        n23864, n23863, n23862, n23861, n23860, n23859, n23850, 
        n23849, n23848, n23847, n23846, n23845, n23844, n23843, 
        n23834, n23833, n23832, n23831, n23830, n23829, n23828, 
        n23827, n224, n45480, n40211, n6834, n34991, n99, n98, 
        n97, n96, n95, n94, n93, n92, n91, n90, n89, n88, 
        n87, n86, n85, n84, n83, n82, n81, n80, n79, n78, 
        n77, n75, n74, n73, n72, n71, n70, n69, n68, n67, 
        n66, n65, n64, n63, n62, n61, n60, n59, n58, n57, 
        n56, n55, n54, n53, n25, n24, n23, n22, n21, n20, 
        n19, n18, n17, n16, n15, n14, n13, n12, n11, n10, 
        n9, n8, n7, n6_adj_3959, n5, n4_adj_3960, n3, n23802, 
        n23801, n23800, n23799, n23798, n23797, n23796, n23795, 
        n23786, n23785, n23784, n23783, n23782, n23781, n23780, 
        n23779, n34990, n34989, n34988, n24140, n34987, n34986, 
        n45649, n34985, n34984, n15_adj_3961, n34983, n34982, n34981, 
        n34980, n34979, n34978, n34977, n34976, n15_adj_3962, n34975, 
        n34974, n7023, n6998, n6974, n6951, n4034, n34973, n34972, 
        n15_adj_3963, n3815, n3814, n3813, n3812, n3811, n3810, 
        n3809, n3808, n3807, n3806, n3805, n3804, n3803, n3802, 
        n3801, n3800, n3799, n3798, n3797, n3796, n3795, n3794, 
        n3793, n3792, n34971, n34970, n24146, n46199, n24081, 
        n24147, n24148, n44973, n34969, n34968, n34315, n34967, 
        n34966, n34965, n34964, n24157, n34963, n34962, n34961, 
        n34960, n34959, n2227;
    wire [31:0]\PID_CONTROLLER.err ;   // verilog/motorControl.v(30[23:26])
    wire [31:0]\PID_CONTROLLER.err_prev ;   // verilog/motorControl.v(31[23:31])
    
    wire n24139, n24138;
    wire [31:0]\PID_CONTROLLER.result ;   // verilog/motorControl.v(32[23:29])
    wire [8:0]pwm_count;   // verilog/motorControl.v(62[13:22])
    
    wire n34958, n24163, n24162, n24161, n24160, n24159, n24088, 
        n25_adj_3964, n24_adj_3965, n23_adj_3966, n22_adj_3967, n21_adj_3968, 
        n20_adj_3969, n19_adj_3970, n18_adj_3971, n17_adj_3972, n16_adj_3973, 
        n15_adj_3974, n14_adj_3975, n13_adj_3976, n12_adj_3977, n11_adj_3978, 
        n10_adj_3979, n9_adj_3980, n8_adj_3981, n7_adj_3982, n6_adj_3983, 
        n34957, n44964, n44430, n24137;
    wire [31:0]pwm_23__N_2960;
    
    wire pwm_23__N_2957, n387, n24136, n414, n415, n421, n22409, 
        n44422, n455, n456, n457, n458, n459, n460, n461, n462, 
        n463, n464, n467, n468, n469, n470, n471, n34956, n34955, 
        n34954, n4_adj_3984, n34953, n34952, n4_adj_3985, n2237, 
        n2236, n34951, n2235, n2234, n2233, n34950, n22406, n2228, 
        n2229, n34949, n34948, n45716, n34314, n8_adj_3986, n34947, 
        n44407, n853, n855, n856, n857, n859, n860, n861, n862, 
        n863, n864, n865, n866, n867, n868, n869, n870, n871, 
        n872, n873, n874, n875, n34946, n4_adj_3987, n34313, n34312, 
        n40892, n22_adj_3988, n34311, n6_adj_3989, quadA_debounced, 
        quadB_debounced, count_enable, n34945, n34944, n34943, n34942, 
        n34941, n34940, n34939, n34938, n34937, n34936, n34935, 
        n34934, n34933, n34932, n34931, quadA_debounced_adj_3990, 
        quadB_debounced_adj_3991, count_enable_adj_3992, n34930, n2300, 
        n2299, n2298, n2297, n2296, n34929, n34928, n34927, n34926, 
        n2311, n46044, r_Rx_Data;
    wire [2:0]r_Bit_Index;   // verilog/uart_rx.v(33[17:28])
    wire [2:0]r_SM_Main;   // verilog/uart_rx.v(36[17:26])
    
    wire n34925, n34924, n4_adj_3993, n46090, n24087, n24086, n24085, 
        n34923, n34922, n23770, n23769, n2232;
    wire [2:0]r_SM_Main_adj_4397;   // verilog/uart_tx.v(31[16:25])
    wire [8:0]r_Clock_Count_adj_4398;   // verilog/uart_tx.v(32[16:29])
    wire [2:0]r_Bit_Index_adj_4399;   // verilog/uart_tx.v(33[16:27])
    
    wire n34921, n34920, n34919, n34918, n2231, n2295, n2230, 
        n313, n314, n315, n24084, n24083, n24082, n45642, n23768, 
        n23767, n23766, n23765, n23764, n23763, n23762, n23761, 
        n23760, n44391, n2294, n316, n317, n318, n319, n320, 
        n2293, n2292, n2291, n2290, n2289, n2288, n2287, n34917, 
        n4012, n34916, n34915, n2286, n2285, n2284, n34914, n2283;
    wire [1:0]reg_B;   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(142[19:24])
    
    wire n40890;
    wire [1:0]reg_B_adj_4406;   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(142[19:24])
    
    wire n2282, n44385, n6908, n34913, n34912, n34911, n34910, 
        n34909, n34908, n34907, n34906, n34905, n34904, n34903, 
        n34902, n34901, n34900, n34899, n34898, n34897, n34896, 
        n34895, n34894, n34893, n3_adj_4000, n34892, n34891, n44381, 
        n369, n370, n371, n372, n373, n374, n375, n376, n377, 
        n378, n379, n380, n381, n382, n383, n384, n385, n386, 
        n387_adj_4001, n388, n389, n390, n391, n392, n393, n34890, 
        n34889, n34888, n34887, n46197, n40894, n510, n533, n534, 
        n558, n648, n649, n671, n672, n6851, n40227, n783, n784, 
        n785, n806, n807, n45812, n914, n915, n916, n917, n918, 
        n938, n939, n1043, n1044, n1045, n1046, n1047, n1048, 
        n1067, n1068, n23562, n1169, n1170, n1171, n1172, n1173, 
        n1174, n1175, n1193, n1194, n1292, n1293, n1294, n1295, 
        n1296, n1297, n1298, n1299, n23560, n1316, n1317, n6869, 
        n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419, 
        n1420, n1436, n1437, n34855, n40225, n45548, n1529, n1530, 
        n1531, n1532, n1533, n1534, n1535, n1536, n1537, n1538, 
        n1553, n1554, n34854, n34853, n6739, n6740, n6741, n6742, 
        n6743, n6744, n6745, n6746, n6747, n6748, n6749, n1643, 
        n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, 
        n1652, n1653, n1667, n1668, n1754, n1755, n1756, n1757, 
        n1758, n1759, n1760, n1761, n1762, n1763, n1764, n1765, 
        n1778, n1779, n34852, n34851, n34850, n45855, n34849, 
        n34848, n34847, n1862, n1863, n1864, n1865, n1866, n1867, 
        n1868, n1869, n1870, n1871, n1872, n1873, n1874, n34846, 
        n1886, n1887, n34845, n6837, n6838, n6839, n6840, n6841, 
        n6842, n6843, n6844, n6845, n6846, n6847, n6848, n6849, 
        n6850, n34844, n1967, n1968, n1969, n1970, n1971, n1972, 
        n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, 
        n1991, n1992, n6854, n6855, n6856, n6857, n6858, n6859, 
        n6860, n6861, n6862, n6863, n6864, n6865, n6866, n6867, 
        n6868, n2069, n2070, n2071, n2072, n2073, n2074, n2075, 
        n2076, n2077, n2078, n2079, n2080, n2081, n2082, n2083, 
        n2093, n2094, n44785, n6872, n6873, n6874, n6875, n6876, 
        n6877, n6878, n6879, n6880, n6881, n6882, n6883, n6884, 
        n6885, n6886, n6887, n34843, n2168, n2169, n2170, n2171, 
        n2172, n2173, n2174, n2175, n2176, n2177, n2178, n2179, 
        n2180, n2181, n2182, n2183, n5822, n2192, n2193, n6891, 
        n6892, n6893, n6894, n6895, n6896, n6897, n6898, n6899, 
        n6900, n6901, n6902, n6903, n6904, n6905, n6906, n6907, 
        n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, 
        n2272, n2273, n2274, n2275, n2276, n2277_adj_4002, n2278_adj_4003, 
        n2279_adj_4004, n2280_adj_4005, n2288_adj_4006, n2289_adj_4007, 
        n30, n6911, n6912, n6913, n6914, n6915, n6916, n6917, 
        n6918, n6919, n6920, n6921, n6922, n6923, n6924, n6925, 
        n6926, n6927, n6928, n6214, n2357, n2358, n2359, n2360, 
        n2361, n2362, n2363, n2364, n2365, n2366, n2367, n2368, 
        n2369, n2370, n2371, n2372, n2373, n2374, n28, n2381, 
        n2382, n6932, n6933, n6934, n6935, n6936, n6937, n6938, 
        n6939, n6940, n6941, n6942, n6943, n6944, n6945, n6946, 
        n6947, n6948, n6949, n6950, n26, n25_adj_4008, n2447, 
        n2448, n2449, n2450, n2451, n2452, n2453, n2454, n2455, 
        n2456, n2457, n2458, n2459, n2460, n2461, n2462, n2463, 
        n2464, n2465, n2471, n2472, n45822, n6954, n6955, n6956, 
        n6957, n6958, n6959, n6960, n6961, n6962, n6963, n6964, 
        n6965, n6966, n6967, n6968, n6969, n6970, n6971, n6972, 
        n6973, n6575, n44771, n2534, n2535, n2536, n2537, n2538, 
        n2539, n2540, n2541, n2542, n2543, n2544, n2545, n2546, 
        n2547, n2548, n2549, n2550, n2551, n2552, n2553, n2558, 
        n2559, n34842, n44769, n6977, n6978, n6979, n6980, n6981, 
        n6982, n6983, n6984, n6985, n6986, n6987, n6988, n6989, 
        n6990, n6991, n6992, n6993, n6994, n6995, n6996, n6997, 
        n5823, n2618, n2619, n2620, n2621, n2622, n2623, n2624, 
        n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632, 
        n2633, n2634, n2635, n2636, n2637, n2638, n2642, n2643, 
        n7001, n7002, n7003, n7004, n7005, n7006, n7007, n7008, 
        n7009, n7010, n7011, n7012, n7013, n7014, n7015, n7016, 
        n7017, n7018, n7019, n7020, n7021, n7022, n2699, n2700, 
        n2701, n2702, n2703, n2704, n2705, n2706, n2707, n2708, 
        n2709, n2710, n2711, n2712, n2713, n2714, n2715, n2716, 
        n2717, n2718, n2719, n2720, n2723, n2724, n34841, n44765, 
        n2777, n2798, n2799, n2801, n2802, n21_adj_4009, n23759, 
        n23758, n23757, n23756, n23755, n23754, n23753, n23752, 
        n23751, n23749, n23748, n23747, n23746, n23745, n23744, 
        n23743, n23742, n23741, n23740, n23739, n23738, n23737, 
        n23736, n23735, n23734, n23733, n23732, n23731, n44761, 
        n6215, n23730, n46088, n34840, n34839, n34838, n34837, 
        n6576, n6646, n5824, n45568, n6216, n40218, n2_adj_4010, 
        n6577, n22403, n6686, n6647, n5825, n34262, n34261, n34260, 
        n34259, n6217, n34258, n34257, n34256, n34255, n34254, 
        n34253, n34252, n34251, n6578, n45572, n6726, n6687, n6648, 
        n5826, n34250, n34249, n34248, n34247, n34246, n34245, 
        n34244, n34243, n34242, n34241, n45674, n11_adj_4011, n13_adj_4012, 
        n11_adj_4013, n13_adj_4014, n11_adj_4015, n13_adj_4016, n44367, 
        n11_adj_4017, n13_adj_4018, n6833, n34240, n4_adj_4019, n6_adj_4020, 
        n8_adj_4021, n9_adj_4022, n11_adj_4023, n13_adj_4024, n15_adj_4025, 
        n23729, n23728, n23727, n23726, n23725, n23724, n23723, 
        n23721, n23720, n23719, n23718, n23717, n23716, n23715, 
        n23714, n23713, n23712, n23711, n23710, n23709, n23708, 
        n23707, n23706, n23705, n23704, n23703, n23702, n23701, 
        n23700, n23699, n23698, n23695, n23665, n23664, n23663, 
        n23662, n23661, n45861, n23660, n23659, n23658, n23655, 
        n23652, n23649, n23645, n23644, n23642, n23639, n23636, 
        n23633, n23630, n23627, n23624, n44365, n6888, n40222, 
        n44721, n6218, n45830, n6579, n6780, n6727, n6688, n6649, 
        n5827, n44710, n6219, n44705, n6580, n6821, n6781, n6728, 
        n6689, n6650, n6220, n4_adj_4026, n6_adj_4027, n8_adj_4028, 
        n9_adj_4029, n16_adj_4030, n5019, n6792, n6832, n44696, 
        n44694, n45586, n6581, n6822, n6782, n6729, n6690, n6651, 
        n2_adj_4031, n3_adj_4032, n4_adj_4033, n5_adj_4034, n6_adj_4035, 
        n7_adj_4036, n8_adj_4037, n9_adj_4038, n10_adj_4039, n11_adj_4040, 
        n12_adj_4041, n13_adj_4042, n14_adj_4043, n15_adj_4044, n16_adj_4045, 
        n17_adj_4046, n18_adj_4047, n19_adj_4048, n20_adj_4049, n21_adj_4050, 
        n22_adj_4051, n23_adj_4052, n24_adj_4053, n25_adj_4054, n2_adj_4055, 
        n3_adj_4056, n4_adj_4057, n5_adj_4058, n6_adj_4059, n7_adj_4060, 
        n8_adj_4061, n9_adj_4062, n10_adj_4063, n11_adj_4064, n12_adj_4065, 
        n13_adj_4066, n14_adj_4067, n15_adj_4068, n16_adj_4069, n17_adj_4070, 
        n18_adj_4071, n19_adj_4072, n20_adj_4073, n21_adj_4074, n22_adj_4075, 
        n23_adj_4076, n24_adj_4077, n25_adj_4078, n6582, n6823, n6783, 
        n6730, n6691, n6652, n44348, n45588, n6824, n45857, n6784, 
        n6731, n6692, n6653, n44346, n46, n40213, n6825, n6785, 
        n44340, n6732, n44, n45506, n6693, n6654, n44332, n44678, 
        n42, n24269, n24268, n24267, n24266, n24265, n24264, n24263, 
        n24262, n40209, n24260, n24259, n24258, n24257, n24256, 
        n24255, n24254, n24253, n24252, n24251, n6826, n6786, 
        n6733, n6694, n40, n42_adj_4079, n44_adj_4080, n45, n24250, 
        n24249, n24248, n24247, n24246, n24245, n24244, n24243, 
        n24242, n24241, n24240, n24239, n24238, n24237, n44326, 
        n38, n40_adj_4081, n42_adj_4082, n43, n45510, n45890, n24231, 
        n24229, n24227, n24226, n24225, n24224, n24223, n39110, 
        n24220, n24219, n24218, n6827, n6787, n6734, n6695, n24217, 
        n24216, n36, n38_adj_4083, n40_adj_4084, n41, n45944, n24215, 
        n24214, n24213, n24212, n24211, n46084, n24208, n24207, 
        n24206, n24205, n24204, n24203, n24202, n24201, n24200, 
        n24199, n34, n36_adj_4085, n38_adj_4086, n39, n41_adj_4087, 
        n43_adj_4088, n44_adj_4089, n45_adj_4090, n45512, n24198, 
        n24197, n24196, n24195, n24194, n24193, n24192, n24191, 
        n24190, n24189, n24188, n24187, n24186, n24185, n24184, 
        n24183, n6828, n6788, n6735, n32, n34_adj_4091, n37, n39_adj_4092, 
        n41_adj_4093, n45884, n43_adj_4094, n45514, n45882, n24078, 
        n23600, n24079, n23599, n30_adj_4095, n31, n32_adj_4096, 
        n33, n34_adj_4097, n35, n37_adj_4098, n39_adj_4099, n45880, 
        n41_adj_4100, n42_adj_4101, n43_adj_4102, n45_adj_4103, n46085, 
        n24077, n24076, n24075, n23595, n24074, n23594, n24072, 
        n23593, n24073, n23592, n6829, n6789, n28_adj_4104, n29, 
        n30_adj_4105, n31_adj_4106, n32_adj_4107, n33_adj_4108, n35_adj_4109, 
        n37_adj_4110, n45878, n39_adj_4111, n40_adj_4112, n41_adj_4113, 
        n43_adj_4114, n45648, n45876, n46066, n23591, n24071, n6736, 
        n24070, n23589, n24069, n23588, n24068, n23587, n24067, 
        n44318, n26_adj_4115, n27, n28_adj_4116, n29_adj_4117, n30_adj_4118, 
        n31_adj_4119, n33_adj_4120, n35_adj_4121, n45874, n37_adj_4122, 
        n38_adj_4123, n39_adj_4124, n41_adj_4125, n46087, n23477, 
        n24066, n23471, n24063, n24135, n24134, n24133, n24_adj_4126, 
        n25_adj_4127, n26_adj_4128, n27_adj_4129, n28_adj_4130, n29_adj_4131, 
        n30_adj_4132, n31_adj_4133, n32_adj_4134, n33_adj_4135, n35_adj_4136, 
        n36_adj_4137, n37_adj_4138, n39_adj_4139, n41_adj_4140, n45744, 
        n43_adj_4141, n44_adj_4142, n45_adj_4143, n45746, n24132, 
        n24131, n24130, n24129, n23458, n44666, n44314, n22_adj_4144, 
        n23_adj_4145, n24_adj_4146, n25_adj_4147, n26_adj_4148, n27_adj_4149, 
        n28_adj_4150, n29_adj_4151, n30_adj_4152, n31_adj_4153, n33_adj_4154, 
        n34_adj_4155, n35_adj_4156, n37_adj_4157, n39_adj_4158, n41_adj_4159, 
        n42_adj_4160, n43_adj_4161, n46048, n6830, n6790, n44312, 
        n20_adj_4162, n21_adj_4163, n22_adj_4164, n23_adj_4165, n24_adj_4166, 
        n25_adj_4167, n26_adj_4168, n27_adj_4169, n28_adj_4170, n29_adj_4171, 
        n31_adj_4172, n32_adj_4173, n33_adj_4174, n35_adj_4175, n37_adj_4176, 
        n45866, n39_adj_4177, n41_adj_4178, n46168, n46095, n44308, 
        n18_adj_4179, n19_adj_4180, n20_adj_4181, n21_adj_4182, n22_adj_4183, 
        n23_adj_4184, n24_adj_4185, n25_adj_4186, n26_adj_4187, n27_adj_4188, 
        n29_adj_4189, n30_adj_4190, n31_adj_4191, n33_adj_4192, n35_adj_4193, 
        n45762, n37_adj_4194, n46097, n39_adj_4195, n41_adj_4196, 
        n43_adj_4197, n45_adj_4198, n45764, n46068, n44662, n23430, 
        n16_adj_4199, n17_adj_4200, n18_adj_4201, n19_adj_4202, n20_adj_4203, 
        n21_adj_4204, n22_adj_4205, n23_adj_4206, n25_adj_4207, n27_adj_4208, 
        n28_adj_4209, n29_adj_4210, n31_adj_4211, n33_adj_4212, n35_adj_4213, 
        n37_adj_4214, n39_adj_4215, n41_adj_4216, n43_adj_4217, n46164, 
        n23585, n14_adj_4218, n16_adj_4219, n17_adj_4220, n18_adj_4221, 
        n19_adj_4222, n20_adj_4223, n21_adj_4224, n22_adj_4225, n23_adj_4226, 
        n25_adj_4227, n26_adj_4228, n27_adj_4229, n29_adj_4230, n31_adj_4231, 
        n45904, n33_adj_4232, n45644, n35_adj_4233, n37_adj_4234, 
        n39_adj_4235, n40_adj_4236, n41_adj_4237, n43_adj_4238, n45_adj_4239, 
        n46070, n12_adj_4240, n14_adj_4241, n15_adj_4242, n16_adj_4243, 
        n17_adj_4244, n18_adj_4245, n19_adj_4246, n20_adj_4247, n21_adj_4248, 
        n23_adj_4249, n24_adj_4250, n25_adj_4251, n27_adj_4252, n29_adj_4253, 
        n46040, n31_adj_4254, n33_adj_4255, n35_adj_4256, n37_adj_4257, 
        n38_adj_4258, n39_adj_4259, n41_adj_4260, n43_adj_4261, n46016, 
        n46205, n6831, n6791, n10_adj_4262, n12_adj_4263, n13_adj_4264, 
        n14_adj_4265, n15_adj_4266, n16_adj_4267, n17_adj_4268, n18_adj_4269, 
        n19_adj_4270, n21_adj_4271, n22_adj_4272, n23_adj_4273, n25_adj_4274, 
        n27_adj_4275, n29_adj_4276, n45638, n31_adj_4277, n33_adj_4278, 
        n35_adj_4279, n36_adj_4280, n37_adj_4281, n39_adj_4282, n41_adj_4283, 
        n46200, n6750, n23584, n8_adj_4284, n10_adj_4285, n11_adj_4286, 
        n12_adj_4287, n13_adj_4288, n14_adj_4289, n15_adj_4290, n16_adj_4291, 
        n17_adj_4292, n19_adj_4293, n20_adj_4294, n21_adj_4295, n23_adj_4296, 
        n25_adj_4297, n45173, n27_adj_4298, n29_adj_4299, n31_adj_4300, 
        n45860, n33_adj_4301, n34_adj_4302, n35_adj_4303, n37_adj_4304, 
        n39_adj_4305, n45774, n46099, n45776, n44296, n6_adj_4306, 
        n8_adj_4307, n9_adj_4308, n10_adj_4309, n11_adj_4310, n12_adj_4311, 
        n13_adj_4312, n14_adj_4313, n15_adj_4314, n17_adj_4315, n19_adj_4316, 
        n21_adj_4317, n23_adj_4318, n45780, n25_adj_4319, n45856, 
        n27_adj_4320, n29_adj_4321, n45854, n31_adj_4322, n32_adj_4323, 
        n33_adj_4324, n35_adj_4325, n37_adj_4326, n46101, n46046, 
        n45850, n4_adj_4327, n6_adj_4328, n7_adj_4329, n8_adj_4330, 
        n9_adj_4331, n10_adj_4332, n11_adj_4333, n12_adj_4334, n13_adj_4335, 
        n15_adj_4336, n16_adj_4337, n17_adj_4338, n19_adj_4339, n21_adj_4340, 
        n45848, n23_adj_4341, n24_adj_4342, n25_adj_4343, n27_adj_4344, 
        n45846, n29_adj_4345, n30_adj_4346, n31_adj_4347, n33_adj_4348, 
        n35_adj_4349, n45796, n37_adj_4350, n45970, n39_adj_4351, 
        n40_adj_4352, n41_adj_4353, n43_adj_4354, n45_adj_4355, n45972, 
        n45836, n46082, n44656, n44654, n10_adj_4356, n24128, n44291, 
        n23583, n24141, n23582, n45849, n23399, n24142, n23581, 
        n24143, n23580, n45847, n44634, n44626, n44622, n44618, 
        n44616, n22338, n45654, n44287, n44285, n45444, n44153, 
        n41998, n41767, n46050, n22466, n45684, n44281, n44134, 
        n44133, n24080, n1_adj_4357, n24127, n24126, n24125, n24145, 
        n24124, n24170, n24164, n22371, n24123, n24165, n44268, 
        n44257, n17_adj_4358, n44255, n44253, n44249, n44247, n44245, 
        n44243, n34836, n34835, n34834, n34833, n22471, n21_adj_4359, 
        n34832, n34831, n34830, n34829, n44229, n34828, n34827, 
        n34826, n34825, n34824, n34823, n34822, n34821, n34820, 
        n34819, n24156, n24166, n34818, n34817, n24155, n24167, 
        n24122, n24168, n24121, n24169, n34816, n34815, n34814, 
        n34813, n34812, n34811, n34810, n34809, n34808, n34807, 
        n34806, n34805, n34804, n34803, n34802, n44117, n45653, 
        n44115, n44113, n44111, n44109, n45652, n5_adj_4360, n44225, 
        n44223, n44221, n44217, n44075, n44211, n46081, n44074, 
        n45714, n46193, n46191, n46185, n46184, n46204, n46169, 
        n46165, n46155, n46186, n46147, n46192, n46190, n46188, 
        n46152, n41887, n44203, n46110, n46108, n45504, n46166, 
        n46104, n46096, n46092, n46049, n46047, n46045, n46041, 
        n46039, n46091, n46037, n46031, n46027, n46025, n46023, 
        n46093, n46019, n44201, n44199, n45643, n46202, n45961, 
        n45955, n44197, n46089, n45941, n45940, n45526, n45920, 
        n46036, n45907, n46038, n45903, n45901, n46042, n45897, 
        n45891, n45639, n45887, n45885, n45883, n45881, n45879, 
        n45875, n44195, n45629, n45793, n45791, n45783, n45779, 
        n45771, n45530, n45766, n45628, n45377, n45351, n45347, 
        n45335, n45550, n46195, n45297, n45259, n45635, n45735, 
        n45733, n45729, n45886;
    
    VCC i2 (.Y(VCC_net));
    SB_IO hall1_input (.PACKAGE_PIN(PIN_20), .LATCH_INPUT_VALUE(GND_net), 
          .INPUT_CLK(GND_net), .OUTPUT_CLK(GND_net), .OUTPUT_ENABLE(GND_net), 
          .D_OUT_1(GND_net), .D_OUT_0(GND_net), .D_IN_0(hall1)) /* synthesis lattice_noprune=1, syn_instantiated=1 */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam hall1_input.PIN_TYPE = 6'b000001;
    defparam hall1_input.PULLUP = 1'b1;
    defparam hall1_input.NEG_TRIGGER = 1'b0;
    defparam hall1_input.IO_STANDARD = "SB_LVCMOS";
    SB_IO hall2_input (.PACKAGE_PIN(PIN_21), .LATCH_INPUT_VALUE(GND_net), 
          .INPUT_CLK(GND_net), .OUTPUT_CLK(GND_net), .OUTPUT_ENABLE(GND_net), 
          .D_OUT_1(GND_net), .D_OUT_0(GND_net), .D_IN_0(hall2)) /* synthesis lattice_noprune=1, syn_instantiated=1 */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam hall2_input.PIN_TYPE = 6'b000001;
    defparam hall2_input.PULLUP = 1'b1;
    defparam hall2_input.NEG_TRIGGER = 1'b0;
    defparam hall2_input.IO_STANDARD = "SB_LVCMOS";
    SB_IO hall3_input (.PACKAGE_PIN(PIN_22), .LATCH_INPUT_VALUE(GND_net), 
          .INPUT_CLK(GND_net), .OUTPUT_CLK(GND_net), .OUTPUT_ENABLE(GND_net), 
          .D_OUT_1(GND_net), .D_OUT_0(GND_net), .D_IN_0(hall3)) /* synthesis lattice_noprune=1, syn_instantiated=1 */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam hall3_input.PIN_TYPE = 6'b000001;
    defparam hall3_input.PULLUP = 1'b1;
    defparam hall3_input.NEG_TRIGGER = 1'b0;
    defparam hall3_input.IO_STANDARD = "SB_LVCMOS";
    SB_IO tx_output (.PACKAGE_PIN(PIN_12), .LATCH_INPUT_VALUE(GND_net), 
          .INPUT_CLK(GND_net), .OUTPUT_CLK(GND_net), .OUTPUT_ENABLE(tx_enable), 
          .D_OUT_1(GND_net), .D_OUT_0(tx_o)) /* synthesis lattice_noprune=1, syn_instantiated=1 */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam tx_output.PIN_TYPE = 6'b101001;
    defparam tx_output.PULLUP = 1'b1;
    defparam tx_output.NEG_TRIGGER = 1'b0;
    defparam tx_output.IO_STANDARD = "SB_LVCMOS";
    motorControl control (.\Kd[3] (Kd[3]), .GND_net(GND_net), .\motor_state[15] (motor_state[15]), 
            .\Kp[6] (Kp[6]), .\PID_CONTROLLER.err[18] (\PID_CONTROLLER.err [18]), 
            .\Kd[4] (Kd[4]), .\motor_state[14] (motor_state[14]), .\motor_state[13] (motor_state[13]), 
            .\motor_state[12] (motor_state[12]), .\motor_state[11] (motor_state[11]), 
            .\motor_state[10] (motor_state[10]), .\motor_state[9] (motor_state[9]), 
            .\motor_state[8] (motor_state[8]), .\Kd[5] (Kd[5]), .\motor_state[7] (motor_state[7]), 
            .\Kd[6] (Kd[6]), .\motor_state[6] (motor_state[6]), .\Kd[1] (Kd[1]), 
            .\motor_state[5] (motor_state[5]), .\Kd[0] (Kd[0]), .\motor_state[4] (motor_state[4]), 
            .\motor_state[3] (motor_state[3]), .\Kd[7] (Kd[7]), .\motor_state[2] (motor_state[2]), 
            .\Kd[2] (Kd[2]), .\motor_state[1] (motor_state[1]), .\Kp[7] (Kp[7]), 
            .\motor_state[0] (motor_state[0]), .VCC_net(VCC_net), .\PID_CONTROLLER.err_prev[31] (\PID_CONTROLLER.err_prev [31]), 
            .\PID_CONTROLLER.err_prev[23] (\PID_CONTROLLER.err_prev [23]), 
            .\PID_CONTROLLER.err_prev[22] (\PID_CONTROLLER.err_prev [22]), 
            .\PID_CONTROLLER.err_prev[21] (\PID_CONTROLLER.err_prev [21]), 
            .\Kp[1] (Kp[1]), .\PID_CONTROLLER.err[6] (\PID_CONTROLLER.err [6]), 
            .\PID_CONTROLLER.err_prev[20] (\PID_CONTROLLER.err_prev [20]), 
            .\PID_CONTROLLER.err_prev[19] (\PID_CONTROLLER.err_prev [19]), 
            .\Kp[0] (Kp[0]), .\PID_CONTROLLER.err[7] (\PID_CONTROLLER.err [7]), 
            .\Kp[2] (Kp[2]), .\Kp[3] (Kp[3]), .\Kp[4] (Kp[4]), .\PID_CONTROLLER.err_prev[18] (\PID_CONTROLLER.err_prev [18]), 
            .\PID_CONTROLLER.err_prev[17] (\PID_CONTROLLER.err_prev [17]), 
            .\Kp[5] (Kp[5]), .\PID_CONTROLLER.err_prev[16] (\PID_CONTROLLER.err_prev [16]), 
            .\PID_CONTROLLER.err[9] (\PID_CONTROLLER.err [9]), .\PID_CONTROLLER.err[8] (\PID_CONTROLLER.err [8]), 
            .\PID_CONTROLLER.err[5] (\PID_CONTROLLER.err [5]), .\PID_CONTROLLER.err[4] (\PID_CONTROLLER.err [4]), 
            .\PID_CONTROLLER.err[3] (\PID_CONTROLLER.err [3]), .\PID_CONTROLLER.err[2] (\PID_CONTROLLER.err [2]), 
            .\PID_CONTROLLER.err[1] (\PID_CONTROLLER.err [1]), .\PID_CONTROLLER.err[0] (\PID_CONTROLLER.err [0]), 
            .pwm_count({pwm_count}), .\PID_CONTROLLER.err[31] (\PID_CONTROLLER.err [31]), 
            .n24227(n24227), .pwm({pwm}), .clk32MHz(clk32MHz), .n24226(n24226), 
            .n24225(n24225), .n24224(n24224), .n24223(n24223), .n39110(n39110), 
            .n24220(n24220), .n24219(n24219), .n24218(n24218), .n24217(n24217), 
            .n24216(n24216), .n24215(n24215), .n24214(n24214), .n24213(n24213), 
            .n24212(n24212), .n24211(n24211), .n24208(n24208), .n24207(n24207), 
            .n24206(n24206), .n24205(n24205), .n24172(n24172), .\PID_CONTROLLER.err[16] (\PID_CONTROLLER.err [16]), 
            .\PID_CONTROLLER.err_prev[15] (\PID_CONTROLLER.err_prev [15]), 
            .\PID_CONTROLLER.err[17] (\PID_CONTROLLER.err [17]), .\PID_CONTROLLER.err[21] (\PID_CONTROLLER.err [21]), 
            .\Ki[5] (Ki[5]), .\Ki[6] (Ki[6]), .\Ki[7] (Ki[7]), .\PID_CONTROLLER.err_prev[14] (\PID_CONTROLLER.err_prev [14]), 
            .\PID_CONTROLLER.err_prev[13] (\PID_CONTROLLER.err_prev [13]), 
            .\PID_CONTROLLER.err_prev[12] (\PID_CONTROLLER.err_prev [12]), 
            .\PID_CONTROLLER.err[19] (\PID_CONTROLLER.err [19]), .\PID_CONTROLLER.err_prev[11] (\PID_CONTROLLER.err_prev [11]), 
            .\PID_CONTROLLER.err[20] (\PID_CONTROLLER.err [20]), .\PID_CONTROLLER.err[22] (\PID_CONTROLLER.err [22]), 
            .\PID_CONTROLLER.err[23] (\PID_CONTROLLER.err [23]), .PIN_7_c_1(PIN_7_c_1), 
            .setpoint({setpoint}), .\PID_CONTROLLER.err[10] (\PID_CONTROLLER.err [10]), 
            .PIN_6_c_0(PIN_6_c_0), .\PID_CONTROLLER.err_prev[10] (\PID_CONTROLLER.err_prev [10]), 
            .\PID_CONTROLLER.err[11] (\PID_CONTROLLER.err [11]), .\PID_CONTROLLER.err_prev[9] (\PID_CONTROLLER.err_prev [9]), 
            .\PID_CONTROLLER.err_prev[8] (\PID_CONTROLLER.err_prev [8]), .\PID_CONTROLLER.err_prev[7] (\PID_CONTROLLER.err_prev [7]), 
            .\PID_CONTROLLER.err_prev[6] (\PID_CONTROLLER.err_prev [6]), .\PID_CONTROLLER.err_prev[5] (\PID_CONTROLLER.err_prev [5]), 
            .\PWMLimit[3] (PWMLimit[3]), .\PWMLimit[2] (PWMLimit[2]), .\Ki[0] (Ki[0]), 
            .\PID_CONTROLLER.err_prev[4] (\PID_CONTROLLER.err_prev [4]), .\Ki[1] (Ki[1]), 
            .\Ki[2] (Ki[2]), .\PID_CONTROLLER.err_prev[3] (\PID_CONTROLLER.err_prev [3]), 
            .\Ki[3] (Ki[3]), .hall1(hall1), .hall2(hall2), .\Ki[4] (Ki[4]), 
            .\PID_CONTROLLER.err_prev[2] (\PID_CONTROLLER.err_prev [2]), .\PID_CONTROLLER.err_prev[1] (\PID_CONTROLLER.err_prev [1]), 
            .n421(n421), .n44153(n44153), .\PID_CONTROLLER.err_prev[0] (\PID_CONTROLLER.err_prev [0]), 
            .hall3(hall3), .n44109(n44109), .n44111(n44111), .n44117(n44117), 
            .n44113(n44113), .n44115(n44115), .n25(n25_adj_4008), .n30(n30), 
            .n26(n26), .n853(n853), .n21(n21_adj_4009), .n855(n855), 
            .n856(n856), .n857(n857), .n859(n859), .n860(n860), .n861(n861), 
            .n862(n862), .n863(n863), .n864(n864), .n865(n865), .n866(n866), 
            .n867(n867), .n868(n868), .n869(n869), .n870(n870), .n871(n871), 
            .n872(n872), .n873(n873), .n874(n874), .n875(n875), .n44074(n44074), 
            .n414(n414), .n415(n415), .n45714(n45714), .\pwm_23__N_2960[6] (pwm_23__N_2960[6]), 
            .\pwm_23__N_2960[5] (pwm_23__N_2960[5]), .\PID_CONTROLLER.err[12] (\PID_CONTROLLER.err [12]), 
            .\PID_CONTROLLER.err[13] (\PID_CONTROLLER.err [13]), .\PID_CONTROLLER.err[14] (\PID_CONTROLLER.err [14]), 
            .n23746(n23746), .n23745(n23745), .n23744(n23744), .n23743(n23743), 
            .n23742(n23742), .n23741(n23741), .n23740(n23740), .n23739(n23739), 
            .n23738(n23738), .n23737(n23737), .n23736(n23736), .n23735(n23735), 
            .n23734(n23734), .n23733(n23733), .n23732(n23732), .n23731(n23731), 
            .n23730(n23730), .n23729(n23729), .n23728(n23728), .n23727(n23727), 
            .n23726(n23726), .n23725(n23725), .n23724(n23724), .n23723(n23723), 
            .\motor_state[23] (motor_state[23]), .\PID_CONTROLLER.result[5] (\PID_CONTROLLER.result [5]), 
            .\PID_CONTROLLER.result[6] (\PID_CONTROLLER.result [6]), .PIN_8_c_2(PIN_8_c_2), 
            .PIN_9_c_3(PIN_9_c_3), .PIN_10_c_4(PIN_10_c_4), .PIN_11_c_5(PIN_11_c_5), 
            .\motor_state[22] (motor_state[22]), .\PID_CONTROLLER.err[15] (\PID_CONTROLLER.err [15]), 
            .\motor_state[21] (motor_state[21]), .\motor_state[20] (motor_state[20]), 
            .\motor_state[19] (motor_state[19]), .\motor_state[18] (motor_state[18]), 
            .\motor_state[17] (motor_state[17]), .\motor_state[16] (motor_state[16]), 
            .n23589(n23589), .n471(n471), .n470(n470), .n469(n469), 
            .n468(n468), .n467(n467), .pwm_23__N_2957(pwm_23__N_2957), 
            .n1(n1), .\PWMLimit[5] (PWMLimit[5]), .n387(n387), .n27212(n27212), 
            .\PWMLimit[6] (PWMLimit[6]), .n464(n464), .n463(n463), .n462(n462), 
            .n461(n461), .n460(n460), .n459(n459), .n458(n458), .n457(n457), 
            .n456(n456), .n455(n455), .\PWMLimit[9] (PWMLimit[9]), .n11(n11_adj_4017), 
            .n13(n13_adj_4018), .\deadband[3] (deadband[3]), .\deadband[7] (deadband[7]), 
            .\deadband[4] (deadband[4]), .\deadband[8] (deadband[8]), .\deadband[9] (deadband[9]), 
            .n13_adj_10(n13_adj_4012), .n11_adj_11(n11_adj_4011), .\deadband[2] (deadband[2]), 
            .\deadband[0] (deadband[0]), .\deadband[1] (deadband[1]), .n16(n16_adj_4030), 
            .\PWMLimit[7] (PWMLimit[7]), .\PWMLimit[4] (PWMLimit[4]), .n41887(n41887), 
            .\PWMLimit[0] (PWMLimit[0]), .\PWMLimit[1] (PWMLimit[1]), .n11_adj_12(n11_adj_4015), 
            .n13_adj_13(n13_adj_4016), .\PWMLimit[8] (PWMLimit[8]), .n11_adj_14(n11_adj_4013), 
            .n13_adj_15(n13_adj_4014), .\deadband[5] (deadband[5]), .\deadband[6] (deadband[6]), 
            .IntegralLimit({IntegralLimit})) /* synthesis lattice_noprune=1, syn_preserve=0, syn_module_defined=1, syn_noprune=0 */ ;   // verilog/TinyFPGA_B.v(143[16] 159[4])
    SB_IO PIN_10_pad (.PACKAGE_PIN(PIN_10), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(PIN_10_c_4)) /* synthesis IO_FF_OUT=TRUE */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam PIN_10_pad.PIN_TYPE = 6'b011001;
    defparam PIN_10_pad.PULLUP = 1'b0;
    defparam PIN_10_pad.NEG_TRIGGER = 1'b0;
    defparam PIN_10_pad.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 i10479_3_lut (.I0(\data_in_frame[5] [1]), .I1(rx_data[1]), .I2(n40218), 
            .I3(GND_net), .O(n23897));   // verilog/coms.v(126[12] 289[6])
    defparam i10479_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 add_2999_19_lut (.I0(GND_net), .I1(n2264), .I2(n83), .I3(n34855), 
            .O(n6891)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2999_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2999_18_lut (.I0(GND_net), .I1(n2265), .I2(n84), .I3(n34854), 
            .O(n6892)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2999_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2999_18 (.CI(n34854), .I0(n2265), .I1(n84), .CO(n34855));
    SB_LUT4 add_2999_17_lut (.I0(GND_net), .I1(n2266), .I2(n85), .I3(n34853), 
            .O(n6893)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2999_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2999_17 (.CI(n34853), .I0(n2266), .I1(n85), .CO(n34854));
    SB_LUT4 add_2999_16_lut (.I0(GND_net), .I1(n2267), .I2(n86), .I3(n34852), 
            .O(n6894)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2999_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2999_16 (.CI(n34852), .I0(n2267), .I1(n86), .CO(n34853));
    SB_LUT4 add_2999_15_lut (.I0(GND_net), .I1(n2268), .I2(n87), .I3(n34851), 
            .O(n6895)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2999_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2999_15 (.CI(n34851), .I0(n2268), .I1(n87), .CO(n34852));
    SB_LUT4 add_2999_14_lut (.I0(GND_net), .I1(n2269), .I2(n88), .I3(n34850), 
            .O(n6896)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2999_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2999_14 (.CI(n34850), .I0(n2269), .I1(n88), .CO(n34851));
    SB_LUT4 div_11_unary_minus_2_add_3_25_lut (.I0(encoder0_position[23]), 
            .I1(GND_net), .I2(n2_adj_4055), .I3(n35122), .O(n224)) /* synthesis syn_instantiated=1 */ ;
    defparam div_11_unary_minus_2_add_3_25_lut.LUT_INIT = 16'h8228;
    SB_LUT4 add_2999_13_lut (.I0(GND_net), .I1(n2270), .I2(n89), .I3(n34849), 
            .O(n6897)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2999_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2999_13 (.CI(n34849), .I0(n2270), .I1(n89), .CO(n34850));
    SB_LUT4 div_11_unary_minus_2_add_3_24_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n3_adj_4056), .I3(n35121), .O(n3)) /* synthesis syn_instantiated=1 */ ;
    defparam div_11_unary_minus_2_add_3_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2999_12_lut (.I0(GND_net), .I1(n2271), .I2(n90), .I3(n34848), 
            .O(n6898)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2999_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2999_12 (.CI(n34848), .I0(n2271), .I1(n90), .CO(n34849));
    SB_CARRY div_11_unary_minus_2_add_3_24 (.CI(n35121), .I0(GND_net), .I1(n3_adj_4056), 
            .CO(n35122));
    SB_LUT4 add_2999_11_lut (.I0(GND_net), .I1(n2272), .I2(n91), .I3(n34847), 
            .O(n6899)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2999_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2999_11 (.CI(n34847), .I0(n2272), .I1(n91), .CO(n34848));
    SB_LUT4 div_11_unary_minus_2_add_3_23_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n4_adj_4057), .I3(n35120), .O(n4_adj_3960)) /* synthesis syn_instantiated=1 */ ;
    defparam div_11_unary_minus_2_add_3_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2999_10_lut (.I0(GND_net), .I1(n2273), .I2(n92), .I3(n34846), 
            .O(n6900)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2999_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2999_10 (.CI(n34846), .I0(n2273), .I1(n92), .CO(n34847));
    SB_CARRY div_11_unary_minus_2_add_3_23 (.CI(n35120), .I0(GND_net), .I1(n4_adj_4057), 
            .CO(n35121));
    SB_LUT4 add_2999_9_lut (.I0(GND_net), .I1(n2274), .I2(n93), .I3(n34845), 
            .O(n6901)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2999_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2999_9 (.CI(n34845), .I0(n2274), .I1(n93), .CO(n34846));
    SB_LUT4 div_11_unary_minus_2_add_3_22_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n5_adj_4058), .I3(n35119), .O(n5)) /* synthesis syn_instantiated=1 */ ;
    defparam div_11_unary_minus_2_add_3_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2999_8_lut (.I0(GND_net), .I1(n2275), .I2(n94), .I3(n34844), 
            .O(n6902)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2999_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2999_8 (.CI(n34844), .I0(n2275), .I1(n94), .CO(n34845));
    SB_LUT4 add_2999_7_lut (.I0(GND_net), .I1(n2276), .I2(n95), .I3(n34843), 
            .O(n6903)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2999_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2999_7 (.CI(n34843), .I0(n2276), .I1(n95), .CO(n34844));
    SB_CARRY div_11_unary_minus_2_add_3_22 (.CI(n35119), .I0(GND_net), .I1(n5_adj_4058), 
            .CO(n35120));
    SB_LUT4 add_2999_6_lut (.I0(GND_net), .I1(n2277_adj_4002), .I2(n96), 
            .I3(n34842), .O(n6904)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2999_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_11_unary_minus_2_add_3_21_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n6_adj_4059), .I3(n35118), .O(n6_adj_3959)) /* synthesis syn_instantiated=1 */ ;
    defparam div_11_unary_minus_2_add_3_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY div_11_unary_minus_2_add_3_21 (.CI(n35118), .I0(GND_net), .I1(n6_adj_4059), 
            .CO(n35119));
    SB_CARRY add_2999_6 (.CI(n34842), .I0(n2277_adj_4002), .I1(n96), .CO(n34843));
    SB_LUT4 add_2999_5_lut (.I0(GND_net), .I1(n2278_adj_4003), .I2(n97), 
            .I3(n34841), .O(n6905)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2999_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_11_unary_minus_2_add_3_20_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n7_adj_4060), .I3(n35117), .O(n7)) /* synthesis syn_instantiated=1 */ ;
    defparam div_11_unary_minus_2_add_3_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2999_5 (.CI(n34841), .I0(n2278_adj_4003), .I1(n97), .CO(n34842));
    SB_LUT4 add_2999_4_lut (.I0(GND_net), .I1(n2279_adj_4004), .I2(n98), 
            .I3(n34840), .O(n6906)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2999_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY div_11_unary_minus_2_add_3_20 (.CI(n35117), .I0(GND_net), .I1(n7_adj_4060), 
            .CO(n35118));
    SB_LUT4 i10480_3_lut (.I0(\data_in_frame[5] [0]), .I1(rx_data[0]), .I2(n40218), 
            .I3(GND_net), .O(n23898));   // verilog/coms.v(126[12] 289[6])
    defparam i10480_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY add_2999_4 (.CI(n34840), .I0(n2279_adj_4004), .I1(n98), .CO(n34841));
    SB_LUT4 div_11_unary_minus_2_add_3_19_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n8_adj_4061), .I3(n35116), .O(n8)) /* synthesis syn_instantiated=1 */ ;
    defparam div_11_unary_minus_2_add_3_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY div_11_unary_minus_2_add_3_19 (.CI(n35116), .I0(GND_net), .I1(n8_adj_4061), 
            .CO(n35117));
    SB_LUT4 add_2999_3_lut (.I0(GND_net), .I1(n2280_adj_4005), .I2(n99), 
            .I3(n34839), .O(n6907)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2999_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_11_unary_minus_2_add_3_18_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n9_adj_4062), .I3(n35115), .O(n9)) /* synthesis syn_instantiated=1 */ ;
    defparam div_11_unary_minus_2_add_3_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2999_3 (.CI(n34839), .I0(n2280_adj_4005), .I1(n99), .CO(n34840));
    SB_CARRY div_11_unary_minus_2_add_3_18 (.CI(n35115), .I0(GND_net), .I1(n9_adj_4062), 
            .CO(n35116));
    SB_LUT4 add_2999_2_lut (.I0(GND_net), .I1(n385), .I2(n558), .I3(VCC_net), 
            .O(n6908)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2999_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_11_unary_minus_2_add_3_17_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n10_adj_4063), .I3(n35114), .O(n10)) /* synthesis syn_instantiated=1 */ ;
    defparam div_11_unary_minus_2_add_3_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2999_2 (.CI(VCC_net), .I0(n385), .I1(n558), .CO(n34839));
    SB_LUT4 add_2998_18_lut (.I0(GND_net), .I1(n2168), .I2(n84), .I3(n34838), 
            .O(n6872)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2998_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY div_11_unary_minus_2_add_3_17 (.CI(n35114), .I0(GND_net), .I1(n10_adj_4063), 
            .CO(n35115));
    SB_LUT4 add_2998_17_lut (.I0(GND_net), .I1(n2169), .I2(n85), .I3(n34837), 
            .O(n6873)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2998_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_11_unary_minus_2_add_3_16_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n11_adj_4064), .I3(n35113), .O(n11)) /* synthesis syn_instantiated=1 */ ;
    defparam div_11_unary_minus_2_add_3_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2998_17 (.CI(n34837), .I0(n2169), .I1(n85), .CO(n34838));
    SB_CARRY div_11_unary_minus_2_add_3_16 (.CI(n35113), .I0(GND_net), .I1(n11_adj_4064), 
            .CO(n35114));
    SB_LUT4 add_2998_16_lut (.I0(GND_net), .I1(n2170), .I2(n86), .I3(n34836), 
            .O(n6874)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2998_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_11_unary_minus_2_add_3_15_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n12_adj_4065), .I3(n35112), .O(n12)) /* synthesis syn_instantiated=1 */ ;
    defparam div_11_unary_minus_2_add_3_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2998_16 (.CI(n34836), .I0(n2170), .I1(n86), .CO(n34837));
    SB_CARRY div_11_unary_minus_2_add_3_15 (.CI(n35112), .I0(GND_net), .I1(n12_adj_4065), 
            .CO(n35113));
    SB_LUT4 add_2998_15_lut (.I0(GND_net), .I1(n2171), .I2(n87), .I3(n34835), 
            .O(n6875)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2998_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_11_unary_minus_2_add_3_14_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n13_adj_4066), .I3(n35111), .O(n13)) /* synthesis syn_instantiated=1 */ ;
    defparam div_11_unary_minus_2_add_3_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2998_15 (.CI(n34835), .I0(n2171), .I1(n87), .CO(n34836));
    SB_CARRY div_11_unary_minus_2_add_3_14 (.CI(n35111), .I0(GND_net), .I1(n13_adj_4066), 
            .CO(n35112));
    SB_LUT4 add_2998_14_lut (.I0(GND_net), .I1(n2172), .I2(n88), .I3(n34834), 
            .O(n6876)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2998_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_11_unary_minus_2_add_3_13_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n14_adj_4067), .I3(n35110), .O(n14)) /* synthesis syn_instantiated=1 */ ;
    defparam div_11_unary_minus_2_add_3_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2998_14 (.CI(n34834), .I0(n2172), .I1(n88), .CO(n34835));
    SB_CARRY div_11_unary_minus_2_add_3_13 (.CI(n35110), .I0(GND_net), .I1(n14_adj_4067), 
            .CO(n35111));
    SB_LUT4 add_2998_13_lut (.I0(GND_net), .I1(n2173), .I2(n89), .I3(n34833), 
            .O(n6877)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2998_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_11_unary_minus_2_add_3_12_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n15_adj_4068), .I3(n35109), .O(n15)) /* synthesis syn_instantiated=1 */ ;
    defparam div_11_unary_minus_2_add_3_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2998_13 (.CI(n34833), .I0(n2173), .I1(n89), .CO(n34834));
    SB_CARRY div_11_unary_minus_2_add_3_12 (.CI(n35109), .I0(GND_net), .I1(n15_adj_4068), 
            .CO(n35110));
    SB_LUT4 add_2998_12_lut (.I0(GND_net), .I1(n2174), .I2(n90), .I3(n34832), 
            .O(n6878)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2998_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_11_unary_minus_2_add_3_11_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n16_adj_4069), .I3(n35108), .O(n16)) /* synthesis syn_instantiated=1 */ ;
    defparam div_11_unary_minus_2_add_3_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2998_12 (.CI(n34832), .I0(n2174), .I1(n90), .CO(n34833));
    SB_CARRY div_11_unary_minus_2_add_3_11 (.CI(n35108), .I0(GND_net), .I1(n16_adj_4069), 
            .CO(n35109));
    SB_LUT4 div_11_unary_minus_2_add_3_10_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n17_adj_4070), .I3(n35107), .O(n17)) /* synthesis syn_instantiated=1 */ ;
    defparam div_11_unary_minus_2_add_3_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2998_11_lut (.I0(GND_net), .I1(n2175), .I2(n91), .I3(n34831), 
            .O(n6879)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2998_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY div_11_unary_minus_2_add_3_10 (.CI(n35107), .I0(GND_net), .I1(n17_adj_4070), 
            .CO(n35108));
    SB_CARRY add_2998_11 (.CI(n34831), .I0(n2175), .I1(n91), .CO(n34832));
    SB_LUT4 add_2998_10_lut (.I0(GND_net), .I1(n2176), .I2(n92), .I3(n34830), 
            .O(n6880)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2998_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2998_10 (.CI(n34830), .I0(n2176), .I1(n92), .CO(n34831));
    SB_LUT4 div_11_unary_minus_2_add_3_9_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n18_adj_4071), .I3(n35106), .O(n18)) /* synthesis syn_instantiated=1 */ ;
    defparam div_11_unary_minus_2_add_3_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2998_9_lut (.I0(GND_net), .I1(n2177), .I2(n93), .I3(n34829), 
            .O(n6881)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2998_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2998_9 (.CI(n34829), .I0(n2177), .I1(n93), .CO(n34830));
    SB_CARRY div_11_unary_minus_2_add_3_9 (.CI(n35106), .I0(GND_net), .I1(n18_adj_4071), 
            .CO(n35107));
    SB_LUT4 add_2998_8_lut (.I0(GND_net), .I1(n2178), .I2(n94), .I3(n34828), 
            .O(n6882)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2998_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2998_8 (.CI(n34828), .I0(n2178), .I1(n94), .CO(n34829));
    SB_LUT4 div_11_unary_minus_2_add_3_8_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n19_adj_4072), .I3(n35105), .O(n19)) /* synthesis syn_instantiated=1 */ ;
    defparam div_11_unary_minus_2_add_3_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2998_7_lut (.I0(GND_net), .I1(n2179), .I2(n95), .I3(n34827), 
            .O(n6883)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2998_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2998_7 (.CI(n34827), .I0(n2179), .I1(n95), .CO(n34828));
    SB_CARRY div_11_unary_minus_2_add_3_8 (.CI(n35105), .I0(GND_net), .I1(n19_adj_4072), 
            .CO(n35106));
    SB_LUT4 add_2998_6_lut (.I0(GND_net), .I1(n2180), .I2(n96), .I3(n34826), 
            .O(n6884)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2998_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2998_6 (.CI(n34826), .I0(n2180), .I1(n96), .CO(n34827));
    SB_LUT4 div_11_unary_minus_2_add_3_7_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n20_adj_4073), .I3(n35104), .O(n20)) /* synthesis syn_instantiated=1 */ ;
    defparam div_11_unary_minus_2_add_3_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2998_5_lut (.I0(GND_net), .I1(n2181), .I2(n97), .I3(n34825), 
            .O(n6885)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2998_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2998_5 (.CI(n34825), .I0(n2181), .I1(n97), .CO(n34826));
    SB_CARRY div_11_unary_minus_2_add_3_7 (.CI(n35104), .I0(GND_net), .I1(n20_adj_4073), 
            .CO(n35105));
    SB_LUT4 add_2998_4_lut (.I0(GND_net), .I1(n2182), .I2(n98), .I3(n34824), 
            .O(n6886)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2998_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2998_4 (.CI(n34824), .I0(n2182), .I1(n98), .CO(n34825));
    SB_LUT4 div_11_unary_minus_2_add_3_6_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n21_adj_4074), .I3(n35103), .O(n21)) /* synthesis syn_instantiated=1 */ ;
    defparam div_11_unary_minus_2_add_3_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2998_3_lut (.I0(GND_net), .I1(n2183), .I2(n99), .I3(n34823), 
            .O(n6887)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2998_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2998_3 (.CI(n34823), .I0(n2183), .I1(n99), .CO(n34824));
    SB_CARRY div_11_unary_minus_2_add_3_6 (.CI(n35103), .I0(GND_net), .I1(n21_adj_4074), 
            .CO(n35104));
    SB_LUT4 add_2998_2_lut (.I0(GND_net), .I1(n384), .I2(n558), .I3(VCC_net), 
            .O(n6888)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2998_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2998_2 (.CI(VCC_net), .I0(n384), .I1(n558), .CO(n34823));
    SB_LUT4 div_11_unary_minus_2_add_3_5_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n22_adj_4075), .I3(n35102), .O(n22)) /* synthesis syn_instantiated=1 */ ;
    defparam div_11_unary_minus_2_add_3_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2997_17_lut (.I0(GND_net), .I1(n2069), .I2(n85), .I3(n34822), 
            .O(n6854)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2997_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2997_16_lut (.I0(GND_net), .I1(n2070), .I2(n86), .I3(n34821), 
            .O(n6855)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2997_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY div_11_unary_minus_2_add_3_5 (.CI(n35102), .I0(GND_net), .I1(n22_adj_4075), 
            .CO(n35103));
    SB_CARRY add_2997_16 (.CI(n34821), .I0(n2070), .I1(n86), .CO(n34822));
    SB_LUT4 add_2997_15_lut (.I0(GND_net), .I1(n2071), .I2(n87), .I3(n34820), 
            .O(n6856)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2997_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_11_unary_minus_2_add_3_4_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n23_adj_4076), .I3(n35101), .O(n23)) /* synthesis syn_instantiated=1 */ ;
    defparam div_11_unary_minus_2_add_3_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2997_15 (.CI(n34820), .I0(n2071), .I1(n87), .CO(n34821));
    SB_LUT4 add_2997_14_lut (.I0(GND_net), .I1(n2072), .I2(n88), .I3(n34819), 
            .O(n6857)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2997_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY div_11_unary_minus_2_add_3_4 (.CI(n35101), .I0(GND_net), .I1(n23_adj_4076), 
            .CO(n35102));
    SB_CARRY add_2997_14 (.CI(n34819), .I0(n2072), .I1(n88), .CO(n34820));
    SB_LUT4 add_2997_13_lut (.I0(GND_net), .I1(n2073), .I2(n89), .I3(n34818), 
            .O(n6858)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2997_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_11_unary_minus_2_add_3_3_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n24_adj_4077), .I3(n35100), .O(n24)) /* synthesis syn_instantiated=1 */ ;
    defparam div_11_unary_minus_2_add_3_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2997_13 (.CI(n34818), .I0(n2073), .I1(n89), .CO(n34819));
    SB_LUT4 add_2997_12_lut (.I0(GND_net), .I1(n2074), .I2(n90), .I3(n34817), 
            .O(n6859)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2997_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY div_11_unary_minus_2_add_3_3 (.CI(n35100), .I0(GND_net), .I1(n24_adj_4077), 
            .CO(n35101));
    SB_CARRY add_2997_12 (.CI(n34817), .I0(n2074), .I1(n90), .CO(n34818));
    SB_LUT4 add_2997_11_lut (.I0(GND_net), .I1(n2075), .I2(n91), .I3(n34816), 
            .O(n6860)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2997_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_11_unary_minus_2_add_3_2_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n25_adj_4078), .I3(VCC_net), .O(n25)) /* synthesis syn_instantiated=1 */ ;
    defparam div_11_unary_minus_2_add_3_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2997_11 (.CI(n34816), .I0(n2075), .I1(n91), .CO(n34817));
    SB_LUT4 add_2997_10_lut (.I0(GND_net), .I1(n2076), .I2(n92), .I3(n34815), 
            .O(n6861)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2997_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY div_11_unary_minus_2_add_3_2 (.CI(VCC_net), .I0(GND_net), .I1(n25_adj_4078), 
            .CO(n35100));
    SB_CARRY add_2997_10 (.CI(n34815), .I0(n2076), .I1(n92), .CO(n34816));
    SB_LUT4 add_2997_9_lut (.I0(GND_net), .I1(n2077), .I2(n93), .I3(n34814), 
            .O(n6862)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2997_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_11_unary_minus_4_add_3_25_lut (.I0(gearBoxRatio[23]), .I1(GND_net), 
            .I2(n2_adj_4031), .I3(n35099), .O(n77)) /* synthesis syn_instantiated=1 */ ;
    defparam div_11_unary_minus_4_add_3_25_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_2997_9 (.CI(n34814), .I0(n2077), .I1(n93), .CO(n34815));
    SB_LUT4 div_11_unary_minus_4_add_3_24_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n3_adj_4032), .I3(n35098), .O(n53)) /* synthesis syn_instantiated=1 */ ;
    defparam div_11_unary_minus_4_add_3_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2997_8_lut (.I0(GND_net), .I1(n2078), .I2(n94), .I3(n34813), 
            .O(n6863)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2997_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY div_11_unary_minus_4_add_3_24 (.CI(n35098), .I0(GND_net), .I1(n3_adj_4032), 
            .CO(n35099));
    SB_CARRY add_2997_8 (.CI(n34813), .I0(n2078), .I1(n94), .CO(n34814));
    SB_LUT4 add_2997_7_lut (.I0(GND_net), .I1(n2079), .I2(n95), .I3(n34812), 
            .O(n6864)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2997_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_11_unary_minus_4_add_3_23_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n4_adj_4033), .I3(n35097), .O(n54)) /* synthesis syn_instantiated=1 */ ;
    defparam div_11_unary_minus_4_add_3_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2997_7 (.CI(n34812), .I0(n2079), .I1(n95), .CO(n34813));
    SB_LUT4 add_2997_6_lut (.I0(GND_net), .I1(n2080), .I2(n96), .I3(n34811), 
            .O(n6865)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2997_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY div_11_unary_minus_4_add_3_23 (.CI(n35097), .I0(GND_net), .I1(n4_adj_4033), 
            .CO(n35098));
    SB_CARRY add_2997_6 (.CI(n34811), .I0(n2080), .I1(n96), .CO(n34812));
    SB_LUT4 add_2997_5_lut (.I0(GND_net), .I1(n2081), .I2(n97), .I3(n34810), 
            .O(n6866)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2997_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_11_unary_minus_4_add_3_22_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n5_adj_4034), .I3(n35096), .O(n55)) /* synthesis syn_instantiated=1 */ ;
    defparam div_11_unary_minus_4_add_3_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2997_5 (.CI(n34810), .I0(n2081), .I1(n97), .CO(n34811));
    SB_LUT4 add_2997_4_lut (.I0(GND_net), .I1(n2082), .I2(n98), .I3(n34809), 
            .O(n6867)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2997_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY div_11_unary_minus_4_add_3_22 (.CI(n35096), .I0(GND_net), .I1(n5_adj_4034), 
            .CO(n35097));
    SB_CARRY add_2997_4 (.CI(n34809), .I0(n2082), .I1(n98), .CO(n34810));
    SB_LUT4 add_2997_3_lut (.I0(GND_net), .I1(n2083), .I2(n99), .I3(n34808), 
            .O(n6868)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2997_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_11_unary_minus_4_add_3_21_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n6_adj_4035), .I3(n35095), .O(n56)) /* synthesis syn_instantiated=1 */ ;
    defparam div_11_unary_minus_4_add_3_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2997_3 (.CI(n34808), .I0(n2083), .I1(n99), .CO(n34809));
    SB_LUT4 add_2997_2_lut (.I0(GND_net), .I1(n383), .I2(n558), .I3(VCC_net), 
            .O(n6869)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2997_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY div_11_unary_minus_4_add_3_21 (.CI(n35095), .I0(GND_net), .I1(n6_adj_4035), 
            .CO(n35096));
    SB_CARRY add_2997_2 (.CI(VCC_net), .I0(n383), .I1(n558), .CO(n34808));
    SB_LUT4 add_2996_16_lut (.I0(GND_net), .I1(n1967), .I2(n86), .I3(n34807), 
            .O(n6837)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2996_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_11_unary_minus_4_add_3_20_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n7_adj_4036), .I3(n35094), .O(n57)) /* synthesis syn_instantiated=1 */ ;
    defparam div_11_unary_minus_4_add_3_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2996_15_lut (.I0(GND_net), .I1(n1968), .I2(n87), .I3(n34806), 
            .O(n6838)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2996_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2996_15 (.CI(n34806), .I0(n1968), .I1(n87), .CO(n34807));
    SB_CARRY div_11_unary_minus_4_add_3_20 (.CI(n35094), .I0(GND_net), .I1(n7_adj_4036), 
            .CO(n35095));
    SB_LUT4 add_2996_14_lut (.I0(GND_net), .I1(n1969), .I2(n88), .I3(n34805), 
            .O(n6839)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2996_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2996_14 (.CI(n34805), .I0(n1969), .I1(n88), .CO(n34806));
    SB_LUT4 div_11_unary_minus_4_add_3_19_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n8_adj_4037), .I3(n35093), .O(n58)) /* synthesis syn_instantiated=1 */ ;
    defparam div_11_unary_minus_4_add_3_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2996_13_lut (.I0(GND_net), .I1(n1970), .I2(n89), .I3(n34804), 
            .O(n6840)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2996_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2996_13 (.CI(n34804), .I0(n1970), .I1(n89), .CO(n34805));
    SB_CARRY div_11_unary_minus_4_add_3_19 (.CI(n35093), .I0(GND_net), .I1(n8_adj_4037), 
            .CO(n35094));
    SB_LUT4 add_2996_12_lut (.I0(GND_net), .I1(n1971), .I2(n90), .I3(n34803), 
            .O(n6841)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2996_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2996_12 (.CI(n34803), .I0(n1971), .I1(n90), .CO(n34804));
    SB_LUT4 div_11_unary_minus_4_add_3_18_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n9_adj_4038), .I3(n35092), .O(n59)) /* synthesis syn_instantiated=1 */ ;
    defparam div_11_unary_minus_4_add_3_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2996_11_lut (.I0(GND_net), .I1(n1972), .I2(n91), .I3(n34802), 
            .O(n6842)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2996_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2996_11 (.CI(n34802), .I0(n1972), .I1(n91), .CO(n34803));
    SB_CARRY div_11_unary_minus_4_add_3_18 (.CI(n35092), .I0(GND_net), .I1(n9_adj_4038), 
            .CO(n35093));
    SB_LUT4 add_2996_10_lut (.I0(GND_net), .I1(n1973), .I2(n92), .I3(n34801), 
            .O(n6843)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2996_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2996_10 (.CI(n34801), .I0(n1973), .I1(n92), .CO(n34802));
    SB_LUT4 div_11_unary_minus_4_add_3_17_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n10_adj_4039), .I3(n35091), .O(n60)) /* synthesis syn_instantiated=1 */ ;
    defparam div_11_unary_minus_4_add_3_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2996_9_lut (.I0(GND_net), .I1(n1974), .I2(n93), .I3(n34800), 
            .O(n6844)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2996_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2996_9 (.CI(n34800), .I0(n1974), .I1(n93), .CO(n34801));
    SB_CARRY div_11_unary_minus_4_add_3_17 (.CI(n35091), .I0(GND_net), .I1(n10_adj_4039), 
            .CO(n35092));
    SB_LUT4 add_2996_8_lut (.I0(GND_net), .I1(n1975), .I2(n94), .I3(n34799), 
            .O(n6845)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2996_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2996_8 (.CI(n34799), .I0(n1975), .I1(n94), .CO(n34800));
    SB_LUT4 i10489_3_lut (.I0(\data_in_frame[3] [7]), .I1(rx_data[7]), .I2(n40216), 
            .I3(GND_net), .O(n23907));   // verilog/coms.v(126[12] 289[6])
    defparam i10489_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_11_unary_minus_4_add_3_16_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n11_adj_4040), .I3(n35090), .O(n61)) /* synthesis syn_instantiated=1 */ ;
    defparam div_11_unary_minus_4_add_3_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2996_7_lut (.I0(GND_net), .I1(n1976), .I2(n95), .I3(n34798), 
            .O(n6846)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2996_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i10490_3_lut (.I0(\data_in_frame[3] [6]), .I1(rx_data[6]), .I2(n40216), 
            .I3(GND_net), .O(n23908));   // verilog/coms.v(126[12] 289[6])
    defparam i10490_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY add_2996_7 (.CI(n34798), .I0(n1976), .I1(n95), .CO(n34799));
    SB_CARRY div_11_unary_minus_4_add_3_16 (.CI(n35090), .I0(GND_net), .I1(n11_adj_4040), 
            .CO(n35091));
    SB_LUT4 add_2996_6_lut (.I0(GND_net), .I1(n1977), .I2(n96), .I3(n34797), 
            .O(n6847)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2996_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2996_6 (.CI(n34797), .I0(n1977), .I1(n96), .CO(n34798));
    SB_LUT4 div_11_unary_minus_4_add_3_15_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n12_adj_4041), .I3(n35089), .O(n62)) /* synthesis syn_instantiated=1 */ ;
    defparam div_11_unary_minus_4_add_3_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2996_5_lut (.I0(GND_net), .I1(n1978), .I2(n97), .I3(n34796), 
            .O(n6848)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2996_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2996_5 (.CI(n34796), .I0(n1978), .I1(n97), .CO(n34797));
    SB_CARRY div_11_unary_minus_4_add_3_15 (.CI(n35089), .I0(GND_net), .I1(n12_adj_4041), 
            .CO(n35090));
    SB_LUT4 add_2996_4_lut (.I0(GND_net), .I1(n1979), .I2(n98), .I3(n34795), 
            .O(n6849)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2996_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2996_4 (.CI(n34795), .I0(n1979), .I1(n98), .CO(n34796));
    SB_LUT4 div_11_unary_minus_4_add_3_14_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n13_adj_4042), .I3(n35088), .O(n63)) /* synthesis syn_instantiated=1 */ ;
    defparam div_11_unary_minus_4_add_3_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2996_3_lut (.I0(GND_net), .I1(n1980), .I2(n99), .I3(n34794), 
            .O(n6850)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2996_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2996_3 (.CI(n34794), .I0(n1980), .I1(n99), .CO(n34795));
    SB_CARRY div_11_unary_minus_4_add_3_14 (.CI(n35088), .I0(GND_net), .I1(n13_adj_4042), 
            .CO(n35089));
    SB_LUT4 add_2996_2_lut (.I0(GND_net), .I1(n382), .I2(n558), .I3(VCC_net), 
            .O(n6851)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2996_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2996_2 (.CI(VCC_net), .I0(n382), .I1(n558), .CO(n34794));
    SB_LUT4 div_11_unary_minus_4_add_3_13_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n14_adj_4043), .I3(n35087), .O(n64)) /* synthesis syn_instantiated=1 */ ;
    defparam div_11_unary_minus_4_add_3_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2995_15_lut (.I0(GND_net), .I1(n1862), .I2(n87), .I3(n34793), 
            .O(n6821)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2995_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i10491_3_lut (.I0(\data_in_frame[3] [5]), .I1(rx_data[5]), .I2(n40216), 
            .I3(GND_net), .O(n23909));   // verilog/coms.v(126[12] 289[6])
    defparam i10491_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 add_2995_14_lut (.I0(GND_net), .I1(n1863), .I2(n88), .I3(n34792), 
            .O(n6822)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2995_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY div_11_unary_minus_4_add_3_13 (.CI(n35087), .I0(GND_net), .I1(n14_adj_4043), 
            .CO(n35088));
    SB_LUT4 i10673_3_lut (.I0(\data_in[1] [1]), .I1(\data_in[2] [1]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n24091));   // verilog/coms.v(126[12] 289[6])
    defparam i10673_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_2995_14 (.CI(n34792), .I0(n1863), .I1(n88), .CO(n34793));
    SB_LUT4 add_2995_13_lut (.I0(GND_net), .I1(n1864), .I2(n89), .I3(n34791), 
            .O(n6823)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2995_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_11_unary_minus_4_add_3_12_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n15_adj_4044), .I3(n35086), .O(n65)) /* synthesis syn_instantiated=1 */ ;
    defparam div_11_unary_minus_4_add_3_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2995_13 (.CI(n34791), .I0(n1864), .I1(n89), .CO(n34792));
    SB_LUT4 add_2995_12_lut (.I0(GND_net), .I1(n1865), .I2(n90), .I3(n34790), 
            .O(n6824)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2995_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY div_11_unary_minus_4_add_3_12 (.CI(n35086), .I0(GND_net), .I1(n15_adj_4044), 
            .CO(n35087));
    SB_CARRY add_2995_12 (.CI(n34790), .I0(n1865), .I1(n90), .CO(n34791));
    SB_LUT4 add_2995_11_lut (.I0(GND_net), .I1(n1866), .I2(n91), .I3(n34789), 
            .O(n6825)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2995_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_11_unary_minus_4_add_3_11_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n16_adj_4045), .I3(n35085), .O(n66)) /* synthesis syn_instantiated=1 */ ;
    defparam div_11_unary_minus_4_add_3_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2995_11 (.CI(n34789), .I0(n1866), .I1(n91), .CO(n34790));
    SB_LUT4 add_2995_10_lut (.I0(GND_net), .I1(n1867), .I2(n92), .I3(n34788), 
            .O(n6826)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2995_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY div_11_unary_minus_4_add_3_11 (.CI(n35085), .I0(GND_net), .I1(n16_adj_4045), 
            .CO(n35086));
    SB_CARRY add_2995_10 (.CI(n34788), .I0(n1867), .I1(n92), .CO(n34789));
    SB_LUT4 add_2995_9_lut (.I0(GND_net), .I1(n1868), .I2(n93), .I3(n34787), 
            .O(n6827)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2995_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_11_unary_minus_4_add_3_10_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n17_adj_4046), .I3(n35084), .O(n67)) /* synthesis syn_instantiated=1 */ ;
    defparam div_11_unary_minus_4_add_3_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2995_9 (.CI(n34787), .I0(n1868), .I1(n93), .CO(n34788));
    SB_LUT4 div_11_unary_minus_4_inv_0_i1_1_lut (.I0(gearBoxRatio[0]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n25_adj_4054));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_unary_minus_4_inv_0_i1_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_2995_8_lut (.I0(GND_net), .I1(n1869), .I2(n94), .I3(n34786), 
            .O(n6828)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2995_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY div_11_unary_minus_4_add_3_10 (.CI(n35084), .I0(GND_net), .I1(n17_adj_4046), 
            .CO(n35085));
    SB_CARRY add_2995_8 (.CI(n34786), .I0(n1869), .I1(n94), .CO(n34787));
    SB_LUT4 add_2995_7_lut (.I0(GND_net), .I1(n1870), .I2(n95), .I3(n34785), 
            .O(n6829)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2995_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_11_unary_minus_4_add_3_9_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n18_adj_4047), .I3(n35083), .O(n68)) /* synthesis syn_instantiated=1 */ ;
    defparam div_11_unary_minus_4_add_3_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2995_7 (.CI(n34785), .I0(n1870), .I1(n95), .CO(n34786));
    SB_LUT4 add_2995_6_lut (.I0(GND_net), .I1(n1871), .I2(n96), .I3(n34784), 
            .O(n6830)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2995_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY div_11_unary_minus_4_add_3_9 (.CI(n35083), .I0(GND_net), .I1(n18_adj_4047), 
            .CO(n35084));
    SB_CARRY add_2995_6 (.CI(n34784), .I0(n1871), .I1(n96), .CO(n34785));
    SB_LUT4 add_2995_5_lut (.I0(GND_net), .I1(n1872), .I2(n97), .I3(n34783), 
            .O(n6831)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2995_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_11_unary_minus_4_add_3_8_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n19_adj_4048), .I3(n35082), .O(n69)) /* synthesis syn_instantiated=1 */ ;
    defparam div_11_unary_minus_4_add_3_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2995_5 (.CI(n34783), .I0(n1872), .I1(n97), .CO(n34784));
    SB_LUT4 add_2995_4_lut (.I0(GND_net), .I1(n1873), .I2(n98), .I3(n34782), 
            .O(n6832)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2995_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY div_11_unary_minus_4_add_3_8 (.CI(n35082), .I0(GND_net), .I1(n19_adj_4048), 
            .CO(n35083));
    SB_CARRY add_2995_4 (.CI(n34782), .I0(n1873), .I1(n98), .CO(n34783));
    SB_LUT4 i10492_3_lut (.I0(\data_in_frame[3] [4]), .I1(rx_data[4]), .I2(n40216), 
            .I3(GND_net), .O(n23910));   // verilog/coms.v(126[12] 289[6])
    defparam i10492_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_11_unary_minus_4_inv_0_i2_1_lut (.I0(gearBoxRatio[1]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n24_adj_4053));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_unary_minus_4_inv_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_11_unary_minus_4_inv_0_i3_1_lut (.I0(gearBoxRatio[2]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n23_adj_4052));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_unary_minus_4_inv_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_2995_3_lut (.I0(GND_net), .I1(n1874), .I2(n99), .I3(n34781), 
            .O(n6833)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2995_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_11_unary_minus_4_add_3_7_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n20_adj_4049), .I3(n35081), .O(n70)) /* synthesis syn_instantiated=1 */ ;
    defparam div_11_unary_minus_4_add_3_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2995_3 (.CI(n34781), .I0(n1874), .I1(n99), .CO(n34782));
    SB_LUT4 div_11_unary_minus_4_inv_0_i4_1_lut (.I0(gearBoxRatio[3]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n22_adj_4051));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_unary_minus_4_inv_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i10674_3_lut (.I0(\data_in[1] [0]), .I1(\data_in[2] [0]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n24092));   // verilog/coms.v(126[12] 289[6])
    defparam i10674_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_2995_2_lut (.I0(GND_net), .I1(n381), .I2(n558), .I3(VCC_net), 
            .O(n6834)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2995_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY div_11_unary_minus_4_add_3_7 (.CI(n35081), .I0(GND_net), .I1(n20_adj_4049), 
            .CO(n35082));
    SB_CARRY add_2995_2 (.CI(VCC_net), .I0(n381), .I1(n558), .CO(n34781));
    SB_LUT4 i10675_3_lut (.I0(\data_in[0] [7]), .I1(\data_in[1] [7]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n24093));   // verilog/coms.v(126[12] 289[6])
    defparam i10675_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_2993_14_lut (.I0(GND_net), .I1(n1754), .I2(n88), .I3(n34780), 
            .O(n6780)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2993_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i10676_3_lut (.I0(\data_in[0] [6]), .I1(\data_in[1] [6]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n24094));   // verilog/coms.v(126[12] 289[6])
    defparam i10676_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10677_3_lut (.I0(\data_in[0] [5]), .I1(\data_in[1] [5]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n24095));   // verilog/coms.v(126[12] 289[6])
    defparam i10677_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_11_unary_minus_4_add_3_6_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n21_adj_4050), .I3(n35080), .O(n71)) /* synthesis syn_instantiated=1 */ ;
    defparam div_11_unary_minus_4_add_3_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2993_13_lut (.I0(GND_net), .I1(n1755), .I2(n89), .I3(n34779), 
            .O(n6781)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2993_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_11_unary_minus_4_inv_0_i5_1_lut (.I0(gearBoxRatio[4]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n21_adj_4050));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_unary_minus_4_inv_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_2993_13 (.CI(n34779), .I0(n1755), .I1(n89), .CO(n34780));
    SB_CARRY div_11_unary_minus_4_add_3_6 (.CI(n35080), .I0(GND_net), .I1(n21_adj_4050), 
            .CO(n35081));
    SB_LUT4 add_2993_12_lut (.I0(GND_net), .I1(n1756), .I2(n90), .I3(n34778), 
            .O(n6782)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2993_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2993_12 (.CI(n34778), .I0(n1756), .I1(n90), .CO(n34779));
    SB_LUT4 i10493_3_lut (.I0(\data_in_frame[3] [3]), .I1(rx_data[3]), .I2(n40216), 
            .I3(GND_net), .O(n23911));   // verilog/coms.v(126[12] 289[6])
    defparam i10493_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_11_unary_minus_4_add_3_5_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n22_adj_4051), .I3(n35079), .O(n72)) /* synthesis syn_instantiated=1 */ ;
    defparam div_11_unary_minus_4_add_3_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2993_11_lut (.I0(GND_net), .I1(n1757), .I2(n91), .I3(n34777), 
            .O(n6783)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2993_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2993_11 (.CI(n34777), .I0(n1757), .I1(n91), .CO(n34778));
    SB_CARRY div_11_unary_minus_4_add_3_5 (.CI(n35079), .I0(GND_net), .I1(n22_adj_4051), 
            .CO(n35080));
    SB_LUT4 add_2993_10_lut (.I0(GND_net), .I1(n1758), .I2(n92), .I3(n34776), 
            .O(n6784)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2993_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2993_10 (.CI(n34776), .I0(n1758), .I1(n92), .CO(n34777));
    SB_LUT4 div_11_unary_minus_4_add_3_4_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n23_adj_4052), .I3(n35078), .O(n73)) /* synthesis syn_instantiated=1 */ ;
    defparam div_11_unary_minus_4_add_3_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2993_9_lut (.I0(GND_net), .I1(n1759), .I2(n93), .I3(n34775), 
            .O(n6785)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2993_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2993_9 (.CI(n34775), .I0(n1759), .I1(n93), .CO(n34776));
    SB_LUT4 i10678_3_lut (.I0(\data_in[0] [4]), .I1(\data_in[1] [4]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n24096));   // verilog/coms.v(126[12] 289[6])
    defparam i10678_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY div_11_unary_minus_4_add_3_4 (.CI(n35078), .I0(GND_net), .I1(n23_adj_4052), 
            .CO(n35079));
    SB_LUT4 add_2993_8_lut (.I0(GND_net), .I1(n1760), .I2(n94), .I3(n34774), 
            .O(n6786)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2993_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2993_8 (.CI(n34774), .I0(n1760), .I1(n94), .CO(n34775));
    SB_LUT4 div_11_unary_minus_4_add_3_3_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n24_adj_4053), .I3(n35077), .O(n74)) /* synthesis syn_instantiated=1 */ ;
    defparam div_11_unary_minus_4_add_3_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2993_7_lut (.I0(GND_net), .I1(n1761), .I2(n95), .I3(n34773), 
            .O(n6787)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2993_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2993_7 (.CI(n34773), .I0(n1761), .I1(n95), .CO(n34774));
    SB_CARRY div_11_unary_minus_4_add_3_3 (.CI(n35077), .I0(GND_net), .I1(n24_adj_4053), 
            .CO(n35078));
    SB_LUT4 add_2993_6_lut (.I0(GND_net), .I1(n1762), .I2(n96), .I3(n34772), 
            .O(n6788)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2993_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2993_6 (.CI(n34772), .I0(n1762), .I1(n96), .CO(n34773));
    SB_LUT4 div_11_unary_minus_4_add_3_2_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n25_adj_4054), .I3(VCC_net), .O(n75)) /* synthesis syn_instantiated=1 */ ;
    defparam div_11_unary_minus_4_add_3_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2993_5_lut (.I0(GND_net), .I1(n1763), .I2(n97), .I3(n34771), 
            .O(n6789)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2993_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2993_5 (.CI(n34771), .I0(n1763), .I1(n97), .CO(n34772));
    SB_CARRY div_11_unary_minus_4_add_3_2 (.CI(VCC_net), .I0(GND_net), .I1(n25_adj_4054), 
            .CO(n35077));
    SB_LUT4 add_2993_4_lut (.I0(GND_net), .I1(n1764), .I2(n98), .I3(n34770), 
            .O(n6790)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2993_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2993_4 (.CI(n34770), .I0(n1764), .I1(n98), .CO(n34771));
    SB_LUT4 add_2993_3_lut (.I0(GND_net), .I1(n1765), .I2(n99), .I3(n34769), 
            .O(n6791)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2993_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2993_3 (.CI(n34769), .I0(n1765), .I1(n99), .CO(n34770));
    SB_LUT4 add_2993_2_lut (.I0(GND_net), .I1(n380), .I2(n558), .I3(VCC_net), 
            .O(n6792)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2993_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2993_2 (.CI(VCC_net), .I0(n380), .I1(n558), .CO(n34769));
    SB_LUT4 add_2991_13_lut (.I0(GND_net), .I1(n1643), .I2(n89), .I3(n34768), 
            .O(n6739)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2991_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2991_12_lut (.I0(GND_net), .I1(n1644), .I2(n90), .I3(n34767), 
            .O(n6740)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2991_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2991_12 (.CI(n34767), .I0(n1644), .I1(n90), .CO(n34768));
    SB_LUT4 add_2991_11_lut (.I0(GND_net), .I1(n1645), .I2(n91), .I3(n34766), 
            .O(n6741)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2991_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2991_11 (.CI(n34766), .I0(n1645), .I1(n91), .CO(n34767));
    SB_LUT4 add_2991_10_lut (.I0(GND_net), .I1(n1646), .I2(n92), .I3(n34765), 
            .O(n6742)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2991_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2991_10 (.CI(n34765), .I0(n1646), .I1(n92), .CO(n34766));
    SB_LUT4 add_2991_9_lut (.I0(GND_net), .I1(n1647), .I2(n93), .I3(n34764), 
            .O(n6743)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2991_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2991_9 (.CI(n34764), .I0(n1647), .I1(n93), .CO(n34765));
    SB_LUT4 add_2991_8_lut (.I0(GND_net), .I1(n1648), .I2(n94), .I3(n34763), 
            .O(n6744)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2991_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2991_8 (.CI(n34763), .I0(n1648), .I1(n94), .CO(n34764));
    SB_LUT4 i10679_3_lut (.I0(\data_in[0] [3]), .I1(\data_in[1] [3]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n24097));   // verilog/coms.v(126[12] 289[6])
    defparam i10679_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_2991_7_lut (.I0(GND_net), .I1(n1649), .I2(n95), .I3(n34762), 
            .O(n6745)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2991_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2991_7 (.CI(n34762), .I0(n1649), .I1(n95), .CO(n34763));
    SB_LUT4 add_2991_6_lut (.I0(GND_net), .I1(n1650), .I2(n96), .I3(n34761), 
            .O(n6746)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2991_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2991_6 (.CI(n34761), .I0(n1650), .I1(n96), .CO(n34762));
    SB_LUT4 add_2991_5_lut (.I0(GND_net), .I1(n1651), .I2(n97), .I3(n34760), 
            .O(n6747)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2991_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i10680_3_lut (.I0(\data_in[0] [2]), .I1(\data_in[1] [2]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n24098));   // verilog/coms.v(126[12] 289[6])
    defparam i10680_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_2991_5 (.CI(n34760), .I0(n1651), .I1(n97), .CO(n34761));
    SB_LUT4 i10681_3_lut (.I0(\data_in[0] [1]), .I1(\data_in[1] [1]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n24099));   // verilog/coms.v(126[12] 289[6])
    defparam i10681_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10682_3_lut (.I0(gearBoxRatio[23]), .I1(\data_in_frame[17] [7]), 
            .I2(n23399), .I3(GND_net), .O(n24100));   // verilog/coms.v(126[12] 289[6])
    defparam i10682_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_2991_4_lut (.I0(GND_net), .I1(n1652), .I2(n98), .I3(n34759), 
            .O(n6748)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2991_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2991_4 (.CI(n34759), .I0(n1652), .I1(n98), .CO(n34760));
    SB_LUT4 add_2991_3_lut (.I0(GND_net), .I1(n1653), .I2(n99), .I3(n34758), 
            .O(n6749)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2991_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2991_3 (.CI(n34758), .I0(n1653), .I1(n99), .CO(n34759));
    SB_LUT4 add_2991_2_lut (.I0(GND_net), .I1(n379), .I2(n558), .I3(VCC_net), 
            .O(n6750)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2991_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2991_2 (.CI(VCC_net), .I0(n379), .I1(n558), .CO(n34758));
    SB_LUT4 add_2990_12_lut (.I0(GND_net), .I1(n1529), .I2(n90), .I3(n34757), 
            .O(n6726)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2990_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2990_11_lut (.I0(GND_net), .I1(n1530), .I2(n91), .I3(n34756), 
            .O(n6727)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2990_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2990_11 (.CI(n34756), .I0(n1530), .I1(n91), .CO(n34757));
    SB_LUT4 add_2990_10_lut (.I0(GND_net), .I1(n1531), .I2(n92), .I3(n34755), 
            .O(n6728)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2990_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2990_10 (.CI(n34755), .I0(n1531), .I1(n92), .CO(n34756));
    SB_LUT4 add_2990_9_lut (.I0(GND_net), .I1(n1532), .I2(n93), .I3(n34754), 
            .O(n6729)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2990_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2990_9 (.CI(n34754), .I0(n1532), .I1(n93), .CO(n34755));
    SB_LUT4 add_2990_8_lut (.I0(GND_net), .I1(n1533), .I2(n94), .I3(n34753), 
            .O(n6730)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2990_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2990_8 (.CI(n34753), .I0(n1533), .I1(n94), .CO(n34754));
    SB_LUT4 add_2990_7_lut (.I0(GND_net), .I1(n1534), .I2(n95), .I3(n34752), 
            .O(n6731)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2990_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2990_7 (.CI(n34752), .I0(n1534), .I1(n95), .CO(n34753));
    SB_LUT4 add_2990_6_lut (.I0(GND_net), .I1(n1535), .I2(n96), .I3(n34751), 
            .O(n6732)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2990_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i10683_3_lut (.I0(gearBoxRatio[22]), .I1(\data_in_frame[17] [6]), 
            .I2(n23399), .I3(GND_net), .O(n24101));   // verilog/coms.v(126[12] 289[6])
    defparam i10683_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_2990_6 (.CI(n34751), .I0(n1535), .I1(n96), .CO(n34752));
    SB_LUT4 add_2990_5_lut (.I0(GND_net), .I1(n1536), .I2(n97), .I3(n34750), 
            .O(n6733)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2990_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i10684_3_lut (.I0(gearBoxRatio[21]), .I1(\data_in_frame[17] [5]), 
            .I2(n23399), .I3(GND_net), .O(n24102));   // verilog/coms.v(126[12] 289[6])
    defparam i10684_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_2990_5 (.CI(n34750), .I0(n1536), .I1(n97), .CO(n34751));
    SB_LUT4 add_2990_4_lut (.I0(GND_net), .I1(n1537), .I2(n98), .I3(n34749), 
            .O(n6734)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2990_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2990_4 (.CI(n34749), .I0(n1537), .I1(n98), .CO(n34750));
    SB_LUT4 add_2971_8_lut (.I0(GND_net), .I1(n1043), .I2(n94), .I3(n34479), 
            .O(n6214)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2971_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2990_3_lut (.I0(GND_net), .I1(n1538), .I2(n99), .I3(n34748), 
            .O(n6735)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2990_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2990_3 (.CI(n34748), .I0(n1538), .I1(n99), .CO(n34749));
    SB_LUT4 add_2971_7_lut (.I0(GND_net), .I1(n1044), .I2(n95), .I3(n34478), 
            .O(n6215)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2971_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2971_7 (.CI(n34478), .I0(n1044), .I1(n95), .CO(n34479));
    SB_LUT4 add_2990_2_lut (.I0(GND_net), .I1(n378), .I2(n558), .I3(VCC_net), 
            .O(n6736)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2990_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2990_2 (.CI(VCC_net), .I0(n378), .I1(n558), .CO(n34748));
    SB_LUT4 add_2971_6_lut (.I0(GND_net), .I1(n1045), .I2(n96), .I3(n34477), 
            .O(n6216)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2971_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2971_6 (.CI(n34477), .I0(n1045), .I1(n96), .CO(n34478));
    SB_LUT4 add_2988_11_lut (.I0(GND_net), .I1(n1412), .I2(n91), .I3(n34747), 
            .O(n6686)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2988_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2988_10_lut (.I0(GND_net), .I1(n1413), .I2(n92), .I3(n34746), 
            .O(n6687)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2988_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2971_5_lut (.I0(GND_net), .I1(n1046), .I2(n97), .I3(n34476), 
            .O(n6217)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2971_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2971_5 (.CI(n34476), .I0(n1046), .I1(n97), .CO(n34477));
    SB_CARRY add_2988_10 (.CI(n34746), .I0(n1413), .I1(n92), .CO(n34747));
    SB_LUT4 add_2988_9_lut (.I0(GND_net), .I1(n1414), .I2(n93), .I3(n34745), 
            .O(n6688)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2988_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2971_4_lut (.I0(GND_net), .I1(n1047), .I2(n98), .I3(n34475), 
            .O(n6218)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2971_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2971_4 (.CI(n34475), .I0(n1047), .I1(n98), .CO(n34476));
    SB_CARRY add_2988_9 (.CI(n34745), .I0(n1414), .I1(n93), .CO(n34746));
    SB_LUT4 add_2988_8_lut (.I0(GND_net), .I1(n1415), .I2(n94), .I3(n34744), 
            .O(n6689)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2988_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2971_3_lut (.I0(GND_net), .I1(n1048), .I2(n99), .I3(n34474), 
            .O(n6219)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2971_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2971_3 (.CI(n34474), .I0(n1048), .I1(n99), .CO(n34475));
    SB_CARRY add_2988_8 (.CI(n34744), .I0(n1415), .I1(n94), .CO(n34745));
    SB_LUT4 add_2988_7_lut (.I0(GND_net), .I1(n1416), .I2(n95), .I3(n34743), 
            .O(n6690)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2988_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2971_2_lut (.I0(GND_net), .I1(n374), .I2(n558), .I3(VCC_net), 
            .O(n6220)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2971_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2971_2 (.CI(VCC_net), .I0(n374), .I1(n558), .CO(n34474));
    SB_CARRY add_2988_7 (.CI(n34743), .I0(n1416), .I1(n95), .CO(n34744));
    SB_LUT4 add_2988_6_lut (.I0(GND_net), .I1(n1417), .I2(n96), .I3(n34742), 
            .O(n6691)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2988_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2988_6 (.CI(n34742), .I0(n1417), .I1(n96), .CO(n34743));
    SB_LUT4 div_11_unary_minus_4_inv_0_i6_1_lut (.I0(gearBoxRatio[5]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n20_adj_4049));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_unary_minus_4_inv_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_2988_5_lut (.I0(GND_net), .I1(n1418), .I2(n97), .I3(n34741), 
            .O(n6692)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2988_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_11_unary_minus_4_inv_0_i7_1_lut (.I0(gearBoxRatio[6]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n19_adj_4048));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_unary_minus_4_inv_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_2988_5 (.CI(n34741), .I0(n1418), .I1(n97), .CO(n34742));
    SB_LUT4 add_2988_4_lut (.I0(GND_net), .I1(n1419), .I2(n98), .I3(n34740), 
            .O(n6693)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2988_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2988_4 (.CI(n34740), .I0(n1419), .I1(n98), .CO(n34741));
    SB_LUT4 add_2988_3_lut (.I0(GND_net), .I1(n1420), .I2(n99), .I3(n34739), 
            .O(n6694)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2988_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2988_3 (.CI(n34739), .I0(n1420), .I1(n99), .CO(n34740));
    SB_LUT4 add_2988_2_lut (.I0(GND_net), .I1(n377), .I2(n558), .I3(VCC_net), 
            .O(n6695)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2988_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2988_2 (.CI(VCC_net), .I0(n377), .I1(n558), .CO(n34739));
    SB_LUT4 add_2986_10_lut (.I0(GND_net), .I1(n1292), .I2(n92), .I3(n34738), 
            .O(n6646)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2986_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2986_9_lut (.I0(GND_net), .I1(n1293), .I2(n93), .I3(n34737), 
            .O(n6647)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2986_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2986_9 (.CI(n34737), .I0(n1293), .I1(n93), .CO(n34738));
    SB_LUT4 add_2986_8_lut (.I0(GND_net), .I1(n1294), .I2(n94), .I3(n34736), 
            .O(n6648)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2986_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2986_8 (.CI(n34736), .I0(n1294), .I1(n94), .CO(n34737));
    SB_LUT4 add_2986_7_lut (.I0(GND_net), .I1(n1295), .I2(n95), .I3(n34735), 
            .O(n6649)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2986_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2986_7 (.CI(n34735), .I0(n1295), .I1(n95), .CO(n34736));
    SB_LUT4 add_2986_6_lut (.I0(GND_net), .I1(n1296), .I2(n96), .I3(n34734), 
            .O(n6650)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2986_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2986_6 (.CI(n34734), .I0(n1296), .I1(n96), .CO(n34735));
    SB_LUT4 add_2986_5_lut (.I0(GND_net), .I1(n1297), .I2(n97), .I3(n34733), 
            .O(n6651)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2986_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2986_5 (.CI(n34733), .I0(n1297), .I1(n97), .CO(n34734));
    SB_LUT4 add_2986_4_lut (.I0(GND_net), .I1(n1298), .I2(n98), .I3(n34732), 
            .O(n6652)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2986_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2986_4 (.CI(n34732), .I0(n1298), .I1(n98), .CO(n34733));
    SB_LUT4 div_11_unary_minus_4_inv_0_i8_1_lut (.I0(gearBoxRatio[7]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n18_adj_4047));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_unary_minus_4_inv_0_i8_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_2986_3_lut (.I0(GND_net), .I1(n1299), .I2(n99), .I3(n34731), 
            .O(n6653)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2986_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2986_3 (.CI(n34731), .I0(n1299), .I1(n99), .CO(n34732));
    SB_LUT4 add_2986_2_lut (.I0(GND_net), .I1(n376), .I2(n558), .I3(VCC_net), 
            .O(n6654)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2986_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2986_2 (.CI(VCC_net), .I0(n376), .I1(n558), .CO(n34731));
    SB_LUT4 i10685_3_lut (.I0(gearBoxRatio[20]), .I1(\data_in_frame[17] [4]), 
            .I2(n23399), .I3(GND_net), .O(n24103));   // verilog/coms.v(126[12] 289[6])
    defparam i10685_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10686_3_lut (.I0(gearBoxRatio[19]), .I1(\data_in_frame[17] [3]), 
            .I2(n23399), .I3(GND_net), .O(n24104));   // verilog/coms.v(126[12] 289[6])
    defparam i10686_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10494_3_lut (.I0(\data_in_frame[3] [2]), .I1(rx_data[2]), .I2(n40216), 
            .I3(GND_net), .O(n23912));   // verilog/coms.v(126[12] 289[6])
    defparam i10494_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_11_unary_minus_4_inv_0_i9_1_lut (.I0(gearBoxRatio[8]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n17_adj_4046));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_unary_minus_4_inv_0_i9_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i10687_3_lut (.I0(gearBoxRatio[18]), .I1(\data_in_frame[17] [2]), 
            .I2(n23399), .I3(GND_net), .O(n24105));   // verilog/coms.v(126[12] 289[6])
    defparam i10687_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_11_unary_minus_4_inv_0_i10_1_lut (.I0(gearBoxRatio[9]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n16_adj_4045));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_unary_minus_4_inv_0_i10_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i10688_3_lut (.I0(gearBoxRatio[17]), .I1(\data_in_frame[17] [1]), 
            .I2(n23399), .I3(GND_net), .O(n24106));   // verilog/coms.v(126[12] 289[6])
    defparam i10688_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_11_unary_minus_4_inv_0_i11_1_lut (.I0(gearBoxRatio[10]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n15_adj_4044));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_unary_minus_4_inv_0_i11_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i10495_3_lut (.I0(\data_in_frame[3] [1]), .I1(rx_data[1]), .I2(n40216), 
            .I3(GND_net), .O(n23913));   // verilog/coms.v(126[12] 289[6])
    defparam i10495_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_11_unary_minus_4_inv_0_i12_1_lut (.I0(gearBoxRatio[11]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n14_adj_4043));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_unary_minus_4_inv_0_i12_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_11_unary_minus_4_inv_0_i13_1_lut (.I0(gearBoxRatio[12]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n13_adj_4042));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_unary_minus_4_inv_0_i13_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i10737_3_lut (.I0(IntegralLimit[15]), .I1(\data_in_frame[9] [7]), 
            .I2(n23399), .I3(GND_net), .O(n24155));   // verilog/coms.v(126[12] 289[6])
    defparam i10737_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_11_unary_minus_4_inv_0_i14_1_lut (.I0(gearBoxRatio[13]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n12_adj_4041));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_unary_minus_4_inv_0_i14_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i10496_3_lut (.I0(\data_in_frame[3] [0]), .I1(rx_data[0]), .I2(n40216), 
            .I3(GND_net), .O(n23914));   // verilog/coms.v(126[12] 289[6])
    defparam i10496_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_11_unary_minus_4_inv_0_i15_1_lut (.I0(gearBoxRatio[14]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n11_adj_4040));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_unary_minus_4_inv_0_i15_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i10689_3_lut (.I0(gearBoxRatio[16]), .I1(\data_in_frame[17] [0]), 
            .I2(n23399), .I3(GND_net), .O(n24107));   // verilog/coms.v(126[12] 289[6])
    defparam i10689_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_11_unary_minus_4_inv_0_i16_1_lut (.I0(gearBoxRatio[15]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n10_adj_4039));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_unary_minus_4_inv_0_i16_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i10690_3_lut (.I0(gearBoxRatio[15]), .I1(\data_in_frame[18] [7]), 
            .I2(n23399), .I3(GND_net), .O(n24108));   // verilog/coms.v(126[12] 289[6])
    defparam i10690_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_11_unary_minus_4_inv_0_i17_1_lut (.I0(gearBoxRatio[16]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n9_adj_4038));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_unary_minus_4_inv_0_i17_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_11_unary_minus_4_inv_0_i18_1_lut (.I0(gearBoxRatio[17]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n8_adj_4037));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_unary_minus_4_inv_0_i18_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i10691_3_lut (.I0(gearBoxRatio[14]), .I1(\data_in_frame[18] [6]), 
            .I2(n23399), .I3(GND_net), .O(n24109));   // verilog/coms.v(126[12] 289[6])
    defparam i10691_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_11_unary_minus_4_inv_0_i19_1_lut (.I0(gearBoxRatio[18]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n7_adj_4036));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_unary_minus_4_inv_0_i19_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_11_unary_minus_4_inv_0_i20_1_lut (.I0(gearBoxRatio[19]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_4035));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_unary_minus_4_inv_0_i20_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_11_unary_minus_4_inv_0_i21_1_lut (.I0(gearBoxRatio[20]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n5_adj_4034));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_unary_minus_4_inv_0_i21_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_11_unary_minus_4_inv_0_i22_1_lut (.I0(gearBoxRatio[21]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n4_adj_4033));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_unary_minus_4_inv_0_i22_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_11_unary_minus_4_inv_0_i23_1_lut (.I0(gearBoxRatio[22]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_4032));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_unary_minus_4_inv_0_i23_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_11_unary_minus_4_inv_0_i24_1_lut (.I0(gearBoxRatio[23]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n2_adj_4031));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_unary_minus_4_inv_0_i24_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_11_unary_minus_2_inv_0_i1_1_lut (.I0(encoder0_position[0]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n25_adj_4078));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_unary_minus_2_inv_0_i1_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_11_unary_minus_2_inv_0_i2_1_lut (.I0(encoder0_position[1]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n24_adj_4077));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_unary_minus_2_inv_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_11_unary_minus_2_inv_0_i3_1_lut (.I0(encoder0_position[2]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n23_adj_4076));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_unary_minus_2_inv_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_11_unary_minus_2_inv_0_i4_1_lut (.I0(encoder0_position[3]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n22_adj_4075));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_unary_minus_2_inv_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_11_unary_minus_2_inv_0_i5_1_lut (.I0(encoder0_position[4]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n21_adj_4074));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_unary_minus_2_inv_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_11_unary_minus_2_inv_0_i6_1_lut (.I0(encoder0_position[5]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n20_adj_4073));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_unary_minus_2_inv_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_11_unary_minus_2_inv_0_i7_1_lut (.I0(encoder0_position[6]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n19_adj_4072));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_unary_minus_2_inv_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_11_unary_minus_2_inv_0_i8_1_lut (.I0(encoder0_position[7]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n18_adj_4071));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_unary_minus_2_inv_0_i8_1_lut.LUT_INIT = 16'h5555;
    SB_IO PIN_18_pad (.PACKAGE_PIN(PIN_18), .OUTPUT_ENABLE(VCC_net), .D_IN_0(PIN_18_c_1)) /* synthesis IO_FF_IN=TRUE */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam PIN_18_pad.PIN_TYPE = 6'b000001;
    defparam PIN_18_pad.PULLUP = 1'b0;
    defparam PIN_18_pad.NEG_TRIGGER = 1'b0;
    defparam PIN_18_pad.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 div_11_unary_minus_2_inv_0_i9_1_lut (.I0(encoder0_position[8]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n17_adj_4070));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_unary_minus_2_inv_0_i9_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_11_unary_minus_2_inv_0_i10_1_lut (.I0(encoder0_position[9]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n16_adj_4069));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_unary_minus_2_inv_0_i10_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i10505_3_lut (.I0(\data_in_frame[1] [7]), .I1(rx_data[7]), .I2(n40213), 
            .I3(GND_net), .O(n23923));   // verilog/coms.v(126[12] 289[6])
    defparam i10505_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i10506_3_lut (.I0(\data_in_frame[1] [6]), .I1(rx_data[6]), .I2(n40213), 
            .I3(GND_net), .O(n23924));   // verilog/coms.v(126[12] 289[6])
    defparam i10506_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i10507_3_lut (.I0(\data_in_frame[1] [5]), .I1(rx_data[5]), .I2(n40213), 
            .I3(GND_net), .O(n23925));   // verilog/coms.v(126[12] 289[6])
    defparam i10507_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_11_unary_minus_2_inv_0_i11_1_lut (.I0(encoder0_position[10]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n15_adj_4068));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_unary_minus_2_inv_0_i11_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mux_22_i1_4_lut (.I0(encoder1_position[0]), .I1(displacement[0]), 
            .I2(n15_adj_3962), .I3(n15_adj_3963), .O(motor_state_23__N_27[0]));   // verilog/TinyFPGA_B.v(138[5] 141[10])
    defparam mux_22_i1_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_21_i1_3_lut (.I0(encoder0_position[0]), .I1(motor_state_23__N_27[0]), 
            .I2(n15_adj_3961), .I3(GND_net), .O(motor_state[0]));   // verilog/TinyFPGA_B.v(137[5] 141[10])
    defparam mux_21_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10508_3_lut (.I0(\data_in_frame[1] [4]), .I1(rx_data[4]), .I2(n40213), 
            .I3(GND_net), .O(n23926));   // verilog/coms.v(126[12] 289[6])
    defparam i10508_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i10509_3_lut (.I0(\data_in_frame[1] [3]), .I1(rx_data[3]), .I2(n40213), 
            .I3(GND_net), .O(n23927));   // verilog/coms.v(126[12] 289[6])
    defparam i10509_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mux_22_i2_4_lut (.I0(encoder1_position[1]), .I1(displacement[1]), 
            .I2(n15_adj_3962), .I3(n15_adj_3963), .O(motor_state_23__N_27[1]));   // verilog/TinyFPGA_B.v(138[5] 141[10])
    defparam mux_22_i2_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i10510_3_lut (.I0(\data_in_frame[1] [2]), .I1(rx_data[2]), .I2(n40213), 
            .I3(GND_net), .O(n23928));   // verilog/coms.v(126[12] 289[6])
    defparam i10510_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mux_21_i2_3_lut (.I0(encoder0_position[1]), .I1(motor_state_23__N_27[1]), 
            .I2(n15_adj_3961), .I3(GND_net), .O(motor_state[1]));   // verilog/TinyFPGA_B.v(137[5] 141[10])
    defparam mux_21_i2_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_11_unary_minus_2_inv_0_i12_1_lut (.I0(encoder0_position[11]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n14_adj_4067));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_unary_minus_2_inv_0_i12_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i10511_3_lut (.I0(\data_in_frame[1] [1]), .I1(rx_data[1]), .I2(n40213), 
            .I3(GND_net), .O(n23929));   // verilog/coms.v(126[12] 289[6])
    defparam i10511_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mux_22_i3_4_lut (.I0(encoder1_position[2]), .I1(displacement[2]), 
            .I2(n15_adj_3962), .I3(n15_adj_3963), .O(motor_state_23__N_27[2]));   // verilog/TinyFPGA_B.v(138[5] 141[10])
    defparam mux_22_i3_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_21_i3_3_lut (.I0(encoder0_position[2]), .I1(motor_state_23__N_27[2]), 
            .I2(n15_adj_3961), .I3(GND_net), .O(motor_state[2]));   // verilog/TinyFPGA_B.v(137[5] 141[10])
    defparam mux_21_i3_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10512_3_lut (.I0(\data_in_frame[1] [0]), .I1(rx_data[0]), .I2(n40213), 
            .I3(GND_net), .O(n23930));   // verilog/coms.v(126[12] 289[6])
    defparam i10512_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mux_22_i4_4_lut (.I0(encoder1_position[3]), .I1(displacement[3]), 
            .I2(n15_adj_3962), .I3(n15_adj_3963), .O(motor_state_23__N_27[3]));   // verilog/TinyFPGA_B.v(138[5] 141[10])
    defparam mux_22_i4_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_21_i4_3_lut (.I0(encoder0_position[3]), .I1(motor_state_23__N_27[3]), 
            .I2(n15_adj_3961), .I3(GND_net), .O(motor_state[3]));   // verilog/TinyFPGA_B.v(137[5] 141[10])
    defparam mux_21_i4_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_11_unary_minus_2_inv_0_i13_1_lut (.I0(encoder0_position[12]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n13_adj_4066));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_unary_minus_2_inv_0_i13_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i10738_3_lut (.I0(IntegralLimit[14]), .I1(\data_in_frame[9] [6]), 
            .I2(n23399), .I3(GND_net), .O(n24156));   // verilog/coms.v(126[12] 289[6])
    defparam i10738_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_22_i5_4_lut (.I0(encoder1_position[4]), .I1(displacement[4]), 
            .I2(n15_adj_3962), .I3(n15_adj_3963), .O(motor_state_23__N_27[4]));   // verilog/TinyFPGA_B.v(138[5] 141[10])
    defparam mux_22_i5_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_21_i5_3_lut (.I0(encoder0_position[4]), .I1(motor_state_23__N_27[4]), 
            .I2(n15_adj_3961), .I3(GND_net), .O(motor_state[4]));   // verilog/TinyFPGA_B.v(137[5] 141[10])
    defparam mux_21_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_11_unary_minus_2_inv_0_i14_1_lut (.I0(encoder0_position[13]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n12_adj_4065));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_unary_minus_2_inv_0_i14_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mux_22_i6_4_lut (.I0(encoder1_position[5]), .I1(displacement[5]), 
            .I2(n15_adj_3962), .I3(n15_adj_3963), .O(motor_state_23__N_27[5]));   // verilog/TinyFPGA_B.v(138[5] 141[10])
    defparam mux_22_i6_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_21_i6_3_lut (.I0(encoder0_position[5]), .I1(motor_state_23__N_27[5]), 
            .I2(n15_adj_3961), .I3(GND_net), .O(motor_state[5]));   // verilog/TinyFPGA_B.v(137[5] 141[10])
    defparam mux_21_i6_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_11_unary_minus_2_inv_0_i15_1_lut (.I0(encoder0_position[14]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n11_adj_4064));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_unary_minus_2_inv_0_i15_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mux_22_i7_4_lut (.I0(encoder1_position[6]), .I1(displacement[6]), 
            .I2(n15_adj_3962), .I3(n15_adj_3963), .O(motor_state_23__N_27[6]));   // verilog/TinyFPGA_B.v(138[5] 141[10])
    defparam mux_22_i7_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_21_i7_3_lut (.I0(encoder0_position[6]), .I1(motor_state_23__N_27[6]), 
            .I2(n15_adj_3961), .I3(GND_net), .O(motor_state[6]));   // verilog/TinyFPGA_B.v(137[5] 141[10])
    defparam mux_21_i7_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10692_3_lut (.I0(gearBoxRatio[13]), .I1(\data_in_frame[18] [5]), 
            .I2(n23399), .I3(GND_net), .O(n24110));   // verilog/coms.v(126[12] 289[6])
    defparam i10692_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10693_3_lut (.I0(gearBoxRatio[12]), .I1(\data_in_frame[18] [4]), 
            .I2(n23399), .I3(GND_net), .O(n24111));   // verilog/coms.v(126[12] 289[6])
    defparam i10693_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF displacement_i0 (.Q(displacement[0]), .C(clk32MHz), .D(displacement_23__N_1[0]));   // verilog/TinyFPGA_B.v(161[10] 163[6])
    SB_LUT4 i10694_3_lut (.I0(gearBoxRatio[11]), .I1(\data_in_frame[18] [3]), 
            .I2(n23399), .I3(GND_net), .O(n24112));   // verilog/coms.v(126[12] 289[6])
    defparam i10694_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_11_unary_minus_2_inv_0_i16_1_lut (.I0(encoder0_position[15]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n10_adj_4063));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_unary_minus_2_inv_0_i16_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_11_mux_3_i7_3_lut (.I0(encoder0_position[6]), .I1(n19), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n385));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_mux_3_i7_3_lut.LUT_INIT = 16'hcaca;
    SB_IO PIN_13_pad (.PACKAGE_PIN(PIN_13), .OUTPUT_ENABLE(VCC_net), .D_IN_0(PIN_13_c));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam PIN_13_pad.PIN_TYPE = 6'b000001;
    defparam PIN_13_pad.PULLUP = 1'b0;
    defparam PIN_13_pad.NEG_TRIGGER = 1'b0;
    defparam PIN_13_pad.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 div_11_unary_minus_2_inv_0_i17_1_lut (.I0(encoder0_position[16]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n9_adj_4062));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_unary_minus_2_inv_0_i17_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mux_22_i8_4_lut (.I0(encoder1_position[7]), .I1(displacement[7]), 
            .I2(n15_adj_3962), .I3(n15_adj_3963), .O(motor_state_23__N_27[7]));   // verilog/TinyFPGA_B.v(138[5] 141[10])
    defparam mux_22_i8_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_21_i8_3_lut (.I0(encoder0_position[7]), .I1(motor_state_23__N_27[7]), 
            .I2(n15_adj_3961), .I3(GND_net), .O(motor_state[7]));   // verilog/TinyFPGA_B.v(137[5] 141[10])
    defparam mux_21_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_11_i1475_3_lut (.I0(n384), .I1(n6888), .I2(n2192), .I3(GND_net), 
            .O(n2280_adj_4005));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1475_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i10695_3_lut (.I0(gearBoxRatio[10]), .I1(\data_in_frame[18] [2]), 
            .I2(n23399), .I3(GND_net), .O(n24113));   // verilog/coms.v(126[12] 289[6])
    defparam i10695_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_11_unary_minus_2_inv_0_i18_1_lut (.I0(encoder0_position[17]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n8_adj_4061));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_unary_minus_2_inv_0_i18_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i10696_3_lut (.I0(gearBoxRatio[9]), .I1(\data_in_frame[18] [1]), 
            .I2(n23399), .I3(GND_net), .O(n24114));   // verilog/coms.v(126[12] 289[6])
    defparam i10696_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10697_3_lut (.I0(gearBoxRatio[8]), .I1(\data_in_frame[18] [0]), 
            .I2(n23399), .I3(GND_net), .O(n24115));   // verilog/coms.v(126[12] 289[6])
    defparam i10697_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10698_3_lut (.I0(gearBoxRatio[7]), .I1(\data_in_frame[19] [7]), 
            .I2(n23399), .I3(GND_net), .O(n24116));   // verilog/coms.v(126[12] 289[6])
    defparam i10698_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_22_i9_4_lut (.I0(encoder1_position[8]), .I1(displacement[8]), 
            .I2(n15_adj_3962), .I3(n15_adj_3963), .O(motor_state_23__N_27[8]));   // verilog/TinyFPGA_B.v(138[5] 141[10])
    defparam mux_22_i9_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_21_i9_3_lut (.I0(encoder0_position[8]), .I1(motor_state_23__N_27[8]), 
            .I2(n15_adj_3961), .I3(GND_net), .O(motor_state[8]));   // verilog/TinyFPGA_B.v(137[5] 141[10])
    defparam mux_21_i9_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10739_3_lut (.I0(IntegralLimit[13]), .I1(\data_in_frame[9] [5]), 
            .I2(n23399), .I3(GND_net), .O(n24157));   // verilog/coms.v(126[12] 289[6])
    defparam i10739_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10699_3_lut (.I0(gearBoxRatio[6]), .I1(\data_in_frame[19] [6]), 
            .I2(n23399), .I3(GND_net), .O(n24117));   // verilog/coms.v(126[12] 289[6])
    defparam i10699_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10745_3_lut (.I0(IntegralLimit[7]), .I1(\data_in_frame[10] [7]), 
            .I2(n23399), .I3(GND_net), .O(n24163));   // verilog/coms.v(126[12] 289[6])
    defparam i10745_3_lut.LUT_INIT = 16'hcaca;
    SB_IO CLK_pad (.PACKAGE_PIN(CLK), .OUTPUT_ENABLE(VCC_net), .D_IN_0(CLK_c));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam CLK_pad.PIN_TYPE = 6'b000001;
    defparam CLK_pad.PULLUP = 1'b0;
    defparam CLK_pad.NEG_TRIGGER = 1'b0;
    defparam CLK_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO PIN_11_pad (.PACKAGE_PIN(PIN_11), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(PIN_11_c_5)) /* synthesis IO_FF_OUT=TRUE */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam PIN_11_pad.PIN_TYPE = 6'b011001;
    defparam PIN_11_pad.PULLUP = 1'b0;
    defparam PIN_11_pad.NEG_TRIGGER = 1'b0;
    defparam PIN_11_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO PIN_23_pad (.PACKAGE_PIN(PIN_23), .OUTPUT_ENABLE(VCC_net), .D_IN_0(PIN_23_c_1)) /* synthesis IO_FF_IN=TRUE */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam PIN_23_pad.PIN_TYPE = 6'b000001;
    defparam PIN_23_pad.PULLUP = 1'b0;
    defparam PIN_23_pad.NEG_TRIGGER = 1'b0;
    defparam PIN_23_pad.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 i10746_3_lut (.I0(IntegralLimit[6]), .I1(\data_in_frame[10] [6]), 
            .I2(n23399), .I3(GND_net), .O(n24164));   // verilog/coms.v(126[12] 289[6])
    defparam i10746_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_11_i1474_3_lut (.I0(n2183), .I1(n6887), .I2(n2192), .I3(GND_net), 
            .O(n2279_adj_4004));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1474_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_11_unary_minus_2_inv_0_i19_1_lut (.I0(encoder0_position[18]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n7_adj_4060));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_unary_minus_2_inv_0_i19_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mux_22_i10_4_lut (.I0(encoder1_position[9]), .I1(displacement[9]), 
            .I2(n15_adj_3962), .I3(n15_adj_3963), .O(motor_state_23__N_27[9]));   // verilog/TinyFPGA_B.v(138[5] 141[10])
    defparam mux_22_i10_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 add_2983_9_lut (.I0(GND_net), .I1(n1169), .I2(n93), .I3(n34700), 
            .O(n6575)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2983_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mux_21_i10_3_lut (.I0(encoder0_position[9]), .I1(motor_state_23__N_27[9]), 
            .I2(n15_adj_3961), .I3(GND_net), .O(motor_state[9]));   // verilog/TinyFPGA_B.v(137[5] 141[10])
    defparam mux_21_i10_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_11_i1473_3_lut (.I0(n2182), .I1(n6886), .I2(n2192), .I3(GND_net), 
            .O(n2278_adj_4003));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1473_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 add_2983_8_lut (.I0(GND_net), .I1(n1170), .I2(n94), .I3(n34699), 
            .O(n6576)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2983_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2983_8 (.CI(n34699), .I0(n1170), .I1(n94), .CO(n34700));
    SB_LUT4 mux_22_i11_4_lut (.I0(encoder1_position[10]), .I1(displacement[10]), 
            .I2(n15_adj_3962), .I3(n15_adj_3963), .O(motor_state_23__N_27[10]));   // verilog/TinyFPGA_B.v(138[5] 141[10])
    defparam mux_22_i11_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_21_i11_3_lut (.I0(encoder0_position[10]), .I1(motor_state_23__N_27[10]), 
            .I2(n15_adj_3961), .I3(GND_net), .O(motor_state[10]));   // verilog/TinyFPGA_B.v(137[5] 141[10])
    defparam mux_21_i11_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_2983_7_lut (.I0(GND_net), .I1(n1171), .I2(n95), .I3(n34698), 
            .O(n6577)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2983_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_11_unary_minus_2_inv_0_i20_1_lut (.I0(encoder0_position[19]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n6_adj_4059));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_unary_minus_2_inv_0_i20_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_11_i1472_3_lut (.I0(n2181), .I1(n6885), .I2(n2192), .I3(GND_net), 
            .O(n2277_adj_4002));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1472_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY add_2983_7 (.CI(n34698), .I0(n1171), .I1(n95), .CO(n34699));
    SB_LUT4 mux_22_i12_4_lut (.I0(encoder1_position[11]), .I1(displacement[11]), 
            .I2(n15_adj_3962), .I3(n15_adj_3963), .O(motor_state_23__N_27[11]));   // verilog/TinyFPGA_B.v(138[5] 141[10])
    defparam mux_22_i12_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_21_i12_3_lut (.I0(encoder0_position[11]), .I1(motor_state_23__N_27[11]), 
            .I2(n15_adj_3961), .I3(GND_net), .O(motor_state[11]));   // verilog/TinyFPGA_B.v(137[5] 141[10])
    defparam mux_21_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_11_i1471_3_lut (.I0(n2180), .I1(n6884), .I2(n2192), .I3(GND_net), 
            .O(n2276));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1471_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 add_2983_6_lut (.I0(GND_net), .I1(n1172), .I2(n96), .I3(n34697), 
            .O(n6578)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2983_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2983_6 (.CI(n34697), .I0(n1172), .I1(n96), .CO(n34698));
    SB_IO PIN_9_pad (.PACKAGE_PIN(PIN_9), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(PIN_9_c_3)) /* synthesis IO_FF_OUT=TRUE */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam PIN_9_pad.PIN_TYPE = 6'b011001;
    defparam PIN_9_pad.PULLUP = 1'b0;
    defparam PIN_9_pad.NEG_TRIGGER = 1'b0;
    defparam PIN_9_pad.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 add_2983_5_lut (.I0(GND_net), .I1(n1173), .I2(n97), .I3(n34696), 
            .O(n6579)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2983_5_lut.LUT_INIT = 16'hC33C;
    SB_IO PIN_8_pad (.PACKAGE_PIN(PIN_8), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(PIN_8_c_2)) /* synthesis IO_FF_OUT=TRUE */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam PIN_8_pad.PIN_TYPE = 6'b011001;
    defparam PIN_8_pad.PULLUP = 1'b0;
    defparam PIN_8_pad.NEG_TRIGGER = 1'b0;
    defparam PIN_8_pad.IO_STANDARD = "SB_LVCMOS";
    SB_CARRY add_2983_5 (.CI(n34696), .I0(n1173), .I1(n97), .CO(n34697));
    SB_LUT4 add_2983_4_lut (.I0(GND_net), .I1(n1174), .I2(n98), .I3(n34695), 
            .O(n6580)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2983_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2983_4 (.CI(n34695), .I0(n1174), .I1(n98), .CO(n34696));
    SB_LUT4 add_2983_3_lut (.I0(GND_net), .I1(n1175), .I2(n99), .I3(n34694), 
            .O(n6581)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2983_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_11_i1470_3_lut (.I0(n2179), .I1(n6883), .I2(n2192), .I3(GND_net), 
            .O(n2275));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1470_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY add_2983_3 (.CI(n34694), .I0(n1175), .I1(n99), .CO(n34695));
    SB_LUT4 add_2983_2_lut (.I0(GND_net), .I1(n375), .I2(n558), .I3(VCC_net), 
            .O(n6582)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2983_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2983_2 (.CI(VCC_net), .I0(n375), .I1(n558), .CO(n34694));
    SB_LUT4 div_11_unary_minus_2_inv_0_i21_1_lut (.I0(encoder0_position[20]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n5_adj_4058));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_unary_minus_2_inv_0_i21_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_11_i1469_3_lut (.I0(n2178), .I1(n6882), .I2(n2192), .I3(GND_net), 
            .O(n2274));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1469_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_11_i1468_3_lut (.I0(n2177), .I1(n6881), .I2(n2192), .I3(GND_net), 
            .O(n2273));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1468_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_11_unary_minus_2_inv_0_i22_1_lut (.I0(encoder0_position[21]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n4_adj_4057));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_unary_minus_2_inv_0_i22_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_11_i1467_3_lut (.I0(n2176), .I1(n6880), .I2(n2192), .I3(GND_net), 
            .O(n2272));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1467_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_11_i1466_3_lut (.I0(n2175), .I1(n6879), .I2(n2192), .I3(GND_net), 
            .O(n2271));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1466_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_11_i1533_3_lut_3_lut (.I0(n2288_adj_4006), .I1(n6902), .I2(n2275), 
            .I3(GND_net), .O(n2368));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1533_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_11_unary_minus_2_inv_0_i23_1_lut (.I0(encoder0_position[22]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n3_adj_4056));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_unary_minus_2_inv_0_i23_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_11_i1522_3_lut_3_lut (.I0(n2288_adj_4006), .I1(n6891), .I2(n2264), 
            .I3(GND_net), .O(n2357));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1522_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_11_i1465_3_lut (.I0(n2174), .I1(n6878), .I2(n2192), .I3(GND_net), 
            .O(n2270));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1465_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_11_i1525_3_lut_3_lut (.I0(n2288_adj_4006), .I1(n6894), .I2(n2267), 
            .I3(GND_net), .O(n2360));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1525_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_11_unary_minus_2_inv_0_i24_1_lut (.I0(encoder0_position[23]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n2_adj_4055));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_unary_minus_2_inv_0_i24_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_11_i1464_3_lut (.I0(n2173), .I1(n6877), .I2(n2192), .I3(GND_net), 
            .O(n2269));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1464_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_11_i1523_3_lut_3_lut (.I0(n2288_adj_4006), .I1(n6892), .I2(n2265), 
            .I3(GND_net), .O(n2358));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1523_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_11_i1463_3_lut (.I0(n2172), .I1(n6876), .I2(n2192), .I3(GND_net), 
            .O(n2268));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1463_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_11_i1526_3_lut_3_lut (.I0(n2288_adj_4006), .I1(n6895), .I2(n2268), 
            .I3(GND_net), .O(n2361));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1526_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_11_i1462_3_lut (.I0(n2171), .I1(n6875), .I2(n2192), .I3(GND_net), 
            .O(n2267));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1462_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_11_i1535_3_lut_3_lut (.I0(n2288_adj_4006), .I1(n6904), .I2(n2277_adj_4002), 
            .I3(GND_net), .O(n2370));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1535_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i10740_3_lut (.I0(IntegralLimit[12]), .I1(\data_in_frame[9] [4]), 
            .I2(n23399), .I3(GND_net), .O(n24158));   // verilog/coms.v(126[12] 289[6])
    defparam i10740_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_11_i1461_3_lut (.I0(n2170), .I1(n6874), .I2(n2192), .I3(GND_net), 
            .O(n2266));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1461_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i10741_3_lut (.I0(IntegralLimit[11]), .I1(\data_in_frame[9] [3]), 
            .I2(n23399), .I3(GND_net), .O(n24159));   // verilog/coms.v(126[12] 289[6])
    defparam i10741_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_11_i1537_3_lut_3_lut (.I0(n2288_adj_4006), .I1(n6906), .I2(n2279_adj_4004), 
            .I3(GND_net), .O(n2372));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1537_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i10742_3_lut (.I0(IntegralLimit[10]), .I1(\data_in_frame[9] [2]), 
            .I2(n23399), .I3(GND_net), .O(n24160));   // verilog/coms.v(126[12] 289[6])
    defparam i10742_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_11_i1460_3_lut (.I0(n2169), .I1(n6873), .I2(n2192), .I3(GND_net), 
            .O(n2265));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1460_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i10743_3_lut (.I0(IntegralLimit[9]), .I1(\data_in_frame[9] [1]), 
            .I2(n23399), .I3(GND_net), .O(n24161));   // verilog/coms.v(126[12] 289[6])
    defparam i10743_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_11_mux_5_i23_3_lut (.I0(gearBoxRatio[22]), .I1(n53), .I2(gearBoxRatio[23]), 
            .I3(GND_net), .O(n78));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_mux_5_i23_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 div_11_i1536_3_lut_3_lut (.I0(n2288_adj_4006), .I1(n6905), .I2(n2278_adj_4003), 
            .I3(GND_net), .O(n2371));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1536_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i1_2_lut (.I0(n78), .I1(n77), .I2(GND_net), .I3(GND_net), 
            .O(n22463));
    defparam i1_2_lut.LUT_INIT = 16'hdddd;
    SB_LUT4 div_11_mux_5_i22_3_lut (.I0(gearBoxRatio[21]), .I1(n54), .I2(gearBoxRatio[23]), 
            .I3(GND_net), .O(n79));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_mux_5_i22_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 div_11_mux_5_i21_3_lut (.I0(gearBoxRatio[20]), .I1(n55), .I2(gearBoxRatio[23]), 
            .I3(GND_net), .O(n80));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_mux_5_i21_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 div_11_mux_5_i20_3_lut (.I0(gearBoxRatio[19]), .I1(n56), .I2(gearBoxRatio[23]), 
            .I3(GND_net), .O(n81));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_mux_5_i20_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 div_11_i1530_3_lut_3_lut (.I0(n2288_adj_4006), .I1(n6899), .I2(n2272), 
            .I3(GND_net), .O(n2365));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1530_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i1_2_lut_adj_1449 (.I0(n81), .I1(n22457), .I2(GND_net), .I3(GND_net), 
            .O(n22454));
    defparam i1_2_lut_adj_1449.LUT_INIT = 16'hdddd;
    SB_LUT4 div_11_mux_5_i19_3_lut (.I0(gearBoxRatio[18]), .I1(n57), .I2(gearBoxRatio[23]), 
            .I3(GND_net), .O(n82));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_mux_5_i19_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 div_11_i1532_3_lut_3_lut (.I0(n2288_adj_4006), .I1(n6901), .I2(n2274), 
            .I3(GND_net), .O(n2367));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1532_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_11_mux_5_i17_3_lut (.I0(gearBoxRatio[16]), .I1(n59), .I2(gearBoxRatio[23]), 
            .I3(GND_net), .O(n84));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_mux_5_i17_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 div_11_i1531_3_lut_3_lut (.I0(n2288_adj_4006), .I1(n6900), .I2(n2273), 
            .I3(GND_net), .O(n2366));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1531_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_11_i1404_3_lut (.I0(n2079), .I1(n6864), .I2(n2093), .I3(GND_net), 
            .O(n2178));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1404_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_11_i1524_3_lut_3_lut (.I0(n2288_adj_4006), .I1(n6893), .I2(n2266), 
            .I3(GND_net), .O(n2359));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1524_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_11_i1398_3_lut (.I0(n2073), .I1(n6858), .I2(n2093), .I3(GND_net), 
            .O(n2172));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1398_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_11_LessThan_1417_i39_2_lut (.I0(n2172), .I1(n88), .I2(GND_net), 
            .I3(GND_net), .O(n39_adj_4195));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1417_i39_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_11_i1395_3_lut (.I0(n2070), .I1(n6855), .I2(n2093), .I3(GND_net), 
            .O(n2169));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1395_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_11_i1539_3_lut_3_lut (.I0(n2288_adj_4006), .I1(n6908), .I2(n385), 
            .I3(GND_net), .O(n2374));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1539_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_11_LessThan_1417_i45_2_lut (.I0(n2169), .I1(n85), .I2(GND_net), 
            .I3(GND_net), .O(n45_adj_4198));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1417_i45_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_11_i1396_3_lut (.I0(n2071), .I1(n6856), .I2(n2093), .I3(GND_net), 
            .O(n2170));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1396_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_11_i1534_3_lut_3_lut (.I0(n2288_adj_4006), .I1(n6903), .I2(n2276), 
            .I3(GND_net), .O(n2369));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1534_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_11_i1529_3_lut_3_lut (.I0(n2288_adj_4006), .I1(n6898), .I2(n2271), 
            .I3(GND_net), .O(n2364));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1529_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_11_LessThan_1417_i43_2_lut (.I0(n2170), .I1(n86), .I2(GND_net), 
            .I3(GND_net), .O(n43_adj_4197));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1417_i43_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_11_i1402_3_lut (.I0(n2077), .I1(n6862), .I2(n2093), .I3(GND_net), 
            .O(n2176));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1402_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_11_i1528_3_lut_3_lut (.I0(n2288_adj_4006), .I1(n6897), .I2(n2270), 
            .I3(GND_net), .O(n2363));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1528_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_11_i1403_3_lut (.I0(n2078), .I1(n6863), .I2(n2093), .I3(GND_net), 
            .O(n2177));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1403_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_11_LessThan_1417_i29_2_lut (.I0(n2177), .I1(n93), .I2(GND_net), 
            .I3(GND_net), .O(n29_adj_4189));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1417_i29_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_11_LessThan_1417_i31_2_lut (.I0(n2176), .I1(n92), .I2(GND_net), 
            .I3(GND_net), .O(n31_adj_4191));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1417_i31_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_11_i1397_3_lut (.I0(n2072), .I1(n6857), .I2(n2093), .I3(GND_net), 
            .O(n2171));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1397_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_11_i1527_3_lut_3_lut (.I0(n2288_adj_4006), .I1(n6896), .I2(n2269), 
            .I3(GND_net), .O(n2362));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1527_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_11_i1538_3_lut_3_lut (.I0(n2288_adj_4006), .I1(n6907), .I2(n2280_adj_4005), 
            .I3(GND_net), .O(n2373));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1538_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_11_LessThan_1417_i41_2_lut (.I0(n2171), .I1(n87), .I2(GND_net), 
            .I3(GND_net), .O(n41_adj_4196));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1417_i41_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_11_i1408_3_lut (.I0(n2083), .I1(n6868), .I2(n2093), .I3(GND_net), 
            .O(n2182));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1408_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_11_i1595_3_lut_3_lut (.I0(n2381), .I1(n6923), .I2(n2369), 
            .I3(GND_net), .O(n2459));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1595_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_11_i1409_3_lut (.I0(n383), .I1(n6869), .I2(n2093), .I3(GND_net), 
            .O(n2183));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1409_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_11_mux_3_i8_3_lut (.I0(encoder0_position[7]), .I1(n18), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n384));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_mux_3_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_11_i1583_3_lut_3_lut (.I0(n2381), .I1(n6911), .I2(n2357), 
            .I3(GND_net), .O(n2447));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1583_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_11_i1584_3_lut_3_lut (.I0(n2381), .I1(n6912), .I2(n2358), 
            .I3(GND_net), .O(n2448));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1584_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_11_i1399_3_lut (.I0(n2074), .I1(n6859), .I2(n2093), .I3(GND_net), 
            .O(n2173));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1399_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_11_i1401_3_lut (.I0(n2076), .I1(n6861), .I2(n2093), .I3(GND_net), 
            .O(n2175));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1401_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_11_i1587_3_lut_3_lut (.I0(n2381), .I1(n6915), .I2(n2361), 
            .I3(GND_net), .O(n2451));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1587_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_11_i1400_3_lut (.I0(n2075), .I1(n6860), .I2(n2093), .I3(GND_net), 
            .O(n2174));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1400_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_11_i1588_3_lut_3_lut (.I0(n2381), .I1(n6916), .I2(n2362), 
            .I3(GND_net), .O(n2452));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1588_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i10744_3_lut (.I0(IntegralLimit[8]), .I1(\data_in_frame[9] [0]), 
            .I2(n23399), .I3(GND_net), .O(n24162));   // verilog/coms.v(126[12] 289[6])
    defparam i10744_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_11_LessThan_1417_i33_2_lut (.I0(n2175), .I1(n91), .I2(GND_net), 
            .I3(GND_net), .O(n33_adj_4192));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1417_i33_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_11_LessThan_1417_i35_2_lut (.I0(n2174), .I1(n90), .I2(GND_net), 
            .I3(GND_net), .O(n35_adj_4193));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1417_i35_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_11_LessThan_1417_i37_2_lut (.I0(n2173), .I1(n89), .I2(GND_net), 
            .I3(GND_net), .O(n37_adj_4194));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1417_i37_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i10667_3_lut (.I0(\data_in[1] [7]), .I1(\data_in[2] [7]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n24085));   // verilog/coms.v(126[12] 289[6])
    defparam i10667_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_11_i1406_3_lut (.I0(n2081), .I1(n6866), .I2(n2093), .I3(GND_net), 
            .O(n2180));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1406_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_11_i1407_3_lut (.I0(n2082), .I1(n6867), .I2(n2093), .I3(GND_net), 
            .O(n2181));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1407_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 PIN_13_I_0_1_lut (.I0(PIN_13_c), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(PIN_13_N_26));   // verilog/TinyFPGA_B.v(73[10:15])
    defparam PIN_13_I_0_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_11_i1585_3_lut_3_lut (.I0(n2381), .I1(n6913), .I2(n2359), 
            .I3(GND_net), .O(n2449));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1585_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i10706_3_lut (.I0(Kd[6]), .I1(\data_in_frame[4] [6]), .I2(n23399), 
            .I3(GND_net), .O(n24124));   // verilog/coms.v(126[12] 289[6])
    defparam i10706_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_11_LessThan_1417_i21_2_lut (.I0(n2181), .I1(n97), .I2(GND_net), 
            .I3(GND_net), .O(n21_adj_4182));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1417_i21_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i10718_3_lut (.I0(Ki[1]), .I1(\data_in_frame[3] [1]), .I2(n23399), 
            .I3(GND_net), .O(n24136));   // verilog/coms.v(126[12] 289[6])
    defparam i10718_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_11_LessThan_1417_i23_2_lut (.I0(n2180), .I1(n96), .I2(GND_net), 
            .I3(GND_net), .O(n23_adj_4184));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1417_i23_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_11_i1327_3_lut (.I0(n1967), .I1(n6837), .I2(n1991), .I3(GND_net), 
            .O(n2069));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1327_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i10719_3_lut (.I0(Kp[7]), .I1(\data_in_frame[2] [7]), .I2(n23399), 
            .I3(GND_net), .O(n24137));   // verilog/coms.v(126[12] 289[6])
    defparam i10719_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_11_i1328_3_lut (.I0(n1968), .I1(n6838), .I2(n1991), .I3(GND_net), 
            .O(n2070));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1328_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i10668_3_lut (.I0(\data_in[1] [6]), .I1(\data_in[2] [6]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n24086));   // verilog/coms.v(126[12] 289[6])
    defparam i10668_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_11_i1329_3_lut (.I0(n1969), .I1(n6839), .I2(n1991), .I3(GND_net), 
            .O(n2071));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1329_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_11_i1586_3_lut_3_lut (.I0(n2381), .I1(n6914), .I2(n2360), 
            .I3(GND_net), .O(n2450));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1586_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_11_i1601_3_lut_3_lut (.I0(n2381), .I1(n6929), .I2(n386), 
            .I3(GND_net), .O(n2465));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1601_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_11_i1330_3_lut (.I0(n1970), .I1(n6840), .I2(n1991), .I3(GND_net), 
            .O(n2072));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1330_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_11_LessThan_1350_i41_2_lut (.I0(n2072), .I1(n88), .I2(GND_net), 
            .I3(GND_net), .O(n41_adj_4178));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1350_i41_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_11_i1332_3_lut (.I0(n1972), .I1(n6842), .I2(n1991), .I3(GND_net), 
            .O(n2074));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1332_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_11_i1597_3_lut_3_lut (.I0(n2381), .I1(n6925), .I2(n2371), 
            .I3(GND_net), .O(n2461));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1597_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_11_LessThan_1350_i37_2_lut (.I0(n2074), .I1(n90), .I2(GND_net), 
            .I3(GND_net), .O(n37_adj_4176));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1350_i37_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_11_i1331_3_lut (.I0(n1971), .I1(n6841), .I2(n1991), .I3(GND_net), 
            .O(n2073));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1331_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_11_i1598_3_lut_3_lut (.I0(n2381), .I1(n6926), .I2(n2372), 
            .I3(GND_net), .O(n2462));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1598_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_11_LessThan_1350_i39_2_lut (.I0(n2073), .I1(n89), .I2(GND_net), 
            .I3(GND_net), .O(n39_adj_4177));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1350_i39_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_11_i1594_3_lut_3_lut (.I0(n2381), .I1(n6922), .I2(n2368), 
            .I3(GND_net), .O(n2458));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1594_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_11_i1333_3_lut (.I0(n1973), .I1(n6843), .I2(n1991), .I3(GND_net), 
            .O(n2075));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1333_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 LessThan_542_i9_2_lut (.I0(pwm_count[4]), .I1(n872), .I2(GND_net), 
            .I3(GND_net), .O(n9_adj_4029));   // verilog/motorControl.v(86[28:44])
    defparam LessThan_542_i9_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_11_LessThan_1350_i35_2_lut (.I0(n2075), .I1(n91), .I2(GND_net), 
            .I3(GND_net), .O(n35_adj_4175));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1350_i35_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_11_i1341_3_lut (.I0(n382), .I1(n6851), .I2(n1991), .I3(GND_net), 
            .O(n2083));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1341_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 LessThan_542_i4_3_lut (.I0(n44074), .I1(n875), .I2(pwm_count[1]), 
            .I3(GND_net), .O(n4_adj_4026));   // verilog/motorControl.v(86[28:44])
    defparam LessThan_542_i4_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_11_mux_3_i9_3_lut (.I0(encoder0_position[8]), .I1(n17), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n383));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_mux_3_i9_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_11_mux_3_i12_3_lut (.I0(encoder0_position[11]), .I1(n14), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n380));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_mux_3_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_542_i8_3_lut (.I0(n6_adj_4027), .I1(n872), .I2(n9_adj_4029), 
            .I3(GND_net), .O(n8_adj_4028));   // verilog/motorControl.v(86[28:44])
    defparam LessThan_542_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_11_i1199_3_lut (.I0(n380), .I1(n6792), .I2(n1778), .I3(GND_net), 
            .O(n1874));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1199_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_11_i1270_3_lut (.I0(n1874), .I1(n6833), .I2(n1886), .I3(GND_net), 
            .O(n1979));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1270_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i30643_4_lut (.I0(n8_adj_4028), .I1(n4_adj_4026), .I2(n9_adj_4029), 
            .I3(n44486), .O(n46164));   // verilog/motorControl.v(86[28:44])
    defparam i30643_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i30644_3_lut (.I0(n46164), .I1(n871), .I2(pwm_count[5]), .I3(GND_net), 
            .O(n46165));   // verilog/motorControl.v(86[28:44])
    defparam i30644_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_11_i1593_3_lut_3_lut (.I0(n2381), .I1(n6921), .I2(n2367), 
            .I3(GND_net), .O(n2457));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1593_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_11_i1337_3_lut (.I0(n1977), .I1(n6847), .I2(n1991), .I3(GND_net), 
            .O(n2079));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1337_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i7_2_lut (.I0(\data_in_frame[7] [6]), .I1(\data_in_frame[7] [7]), 
            .I2(GND_net), .I3(GND_net), .O(Kp_23__N_516));   // verilog/coms.v(94[12:25])
    defparam i7_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i30587_3_lut (.I0(n46165), .I1(n870), .I2(pwm_count[6]), .I3(GND_net), 
            .O(n46108));   // verilog/motorControl.v(86[28:44])
    defparam i30587_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i30542_3_lut (.I0(n46108), .I1(n869), .I2(pwm_count[7]), .I3(GND_net), 
            .O(n16_adj_4030));   // verilog/motorControl.v(86[28:44])
    defparam i30542_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i12_4_lut (.I0(n857), .I1(n855), .I2(n865), .I3(n866), .O(n28));
    defparam i12_4_lut.LUT_INIT = 16'hfffe;
    SB_IO PIN_7_pad (.PACKAGE_PIN(PIN_7), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(PIN_7_c_1)) /* synthesis IO_FF_OUT=TRUE */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam PIN_7_pad.PIN_TYPE = 6'b011001;
    defparam PIN_7_pad.PULLUP = 1'b0;
    defparam PIN_7_pad.NEG_TRIGGER = 1'b0;
    defparam PIN_7_pad.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 div_11_i1592_3_lut_3_lut (.I0(n2381), .I1(n6920), .I2(n2366), 
            .I3(GND_net), .O(n2456));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1592_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 LessThan_542_i18_3_lut (.I0(n16_adj_4030), .I1(n868), .I2(pwm_count[8]), 
            .I3(GND_net), .O(n2311));   // verilog/motorControl.v(86[28:44])
    defparam LessThan_542_i18_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_11_i1339_3_lut (.I0(n1979), .I1(n6849), .I2(n1991), .I3(GND_net), 
            .O(n2081));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1339_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i10_4_lut (.I0(n861), .I1(n856), .I2(n859), .I3(n860), .O(n26));
    defparam i10_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i14_4_lut (.I0(n21_adj_4009), .I1(n28), .I2(n862), .I3(n853), 
            .O(n30));
    defparam i14_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 div_11_LessThan_1350_i23_2_lut (.I0(n2081), .I1(n97), .I2(GND_net), 
            .I3(GND_net), .O(n23_adj_4165));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1350_i23_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i9_4_lut (.I0(n2311), .I1(n864), .I2(n863), .I3(n867), .O(n25_adj_4008));
    defparam i9_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 div_11_LessThan_1350_i25_2_lut (.I0(n2080), .I1(n96), .I2(GND_net), 
            .I3(GND_net), .O(n25_adj_4167));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1350_i25_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_11_LessThan_1350_i27_2_lut (.I0(n2079), .I1(n95), .I2(GND_net), 
            .I3(GND_net), .O(n27_adj_4169));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1350_i27_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_11_i1591_3_lut_3_lut (.I0(n2381), .I1(n6919), .I2(n2365), 
            .I3(GND_net), .O(n2455));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1591_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_11_mux_3_i15_3_lut (.I0(encoder0_position[14]), .I1(n11), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n377));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_mux_3_i15_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_11_i971_3_lut (.I0(n377), .I1(n6695), .I2(n1436), .I3(GND_net), 
            .O(n1538));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i971_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_11_i1590_3_lut_3_lut (.I0(n2381), .I1(n6918), .I2(n2364), 
            .I3(GND_net), .O(n2454));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1590_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_11_i1048_3_lut (.I0(n1538), .I1(n6735), .I2(n1553), .I3(GND_net), 
            .O(n1652));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1048_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 add_3005_25_lut (.I0(n249), .I1(n46887), .I2(n248), .I3(n35010), 
            .O(displacement_23__N_93[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3005_25_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 div_11_i1589_3_lut_3_lut (.I0(n2381), .I1(n6917), .I2(n2363), 
            .I3(GND_net), .O(n2453));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1589_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_11_i1596_3_lut_3_lut (.I0(n2381), .I1(n6924), .I2(n2370), 
            .I3(GND_net), .O(n2460));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1596_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_11_i1600_3_lut_3_lut (.I0(n2381), .I1(n6928), .I2(n2374), 
            .I3(GND_net), .O(n2464));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1600_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_11_i1123_3_lut (.I0(n1652), .I1(n6748), .I2(n1667), .I3(GND_net), 
            .O(n1763));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1123_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_11_i1196_3_lut (.I0(n1763), .I1(n6789), .I2(n1778), .I3(GND_net), 
            .O(n1871));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1196_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_11_i1267_3_lut (.I0(n1871), .I1(n6830), .I2(n1886), .I3(GND_net), 
            .O(n1976));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1267_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 add_3005_24_lut (.I0(n393), .I1(n46887), .I2(n392), .I3(n35009), 
            .O(displacement_23__N_93[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3005_24_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_3005_24 (.CI(n35009), .I0(n46887), .I1(n392), .CO(n35010));
    SB_LUT4 add_3005_23_lut (.I0(n534), .I1(n46887), .I2(n533), .I3(n35008), 
            .O(displacement_23__N_93[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3005_23_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_3005_23 (.CI(n35008), .I0(n46887), .I1(n533), .CO(n35009));
    SB_LUT4 add_3005_22_lut (.I0(n672), .I1(n46887), .I2(n671), .I3(n35007), 
            .O(displacement_23__N_93[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3005_22_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 div_11_i1599_3_lut_3_lut (.I0(n2381), .I1(n6927), .I2(n2373), 
            .I3(GND_net), .O(n2463));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1599_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_11_i1335_3_lut (.I0(n1975), .I1(n6845), .I2(n1991), .I3(GND_net), 
            .O(n2077));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1335_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY add_3005_22 (.CI(n35007), .I0(n46887), .I1(n671), .CO(n35008));
    SB_LUT4 add_3005_21_lut (.I0(n807), .I1(n46887), .I2(n806), .I3(n35006), 
            .O(displacement_23__N_93[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3005_21_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_3005_21 (.CI(n35006), .I0(n46887), .I1(n806), .CO(n35007));
    SB_LUT4 LessThan_539_i15_2_lut (.I0(pwm_count[7]), .I1(pwm[7]), .I2(GND_net), 
            .I3(GND_net), .O(n15_adj_4025));   // verilog/motorControl.v(65[19:32])
    defparam LessThan_539_i15_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_3005_20_lut (.I0(n939), .I1(n46887), .I2(n938), .I3(n35005), 
            .O(displacement_23__N_93[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3005_20_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 add_2958_7_lut (.I0(GND_net), .I1(n914), .I2(n95), .I3(n34315), 
            .O(n5822)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2958_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_11_mux_3_i17_3_lut (.I0(encoder0_position[16]), .I1(n9), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n375));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_mux_3_i17_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_2958_6_lut (.I0(GND_net), .I1(n915), .I2(n96), .I3(n34314), 
            .O(n5823)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2958_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2958_6 (.CI(n34314), .I0(n915), .I1(n96), .CO(n34315));
    SB_CARRY add_3005_20 (.CI(n35005), .I0(n46887), .I1(n938), .CO(n35006));
    SB_LUT4 add_2958_5_lut (.I0(GND_net), .I1(n916), .I2(n97), .I3(n34313), 
            .O(n5824)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2958_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2958_5 (.CI(n34313), .I0(n916), .I1(n97), .CO(n34314));
    SB_LUT4 add_3005_19_lut (.I0(n1068), .I1(n46887), .I2(n1067), .I3(n35004), 
            .O(displacement_23__N_93[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3005_19_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 add_2958_4_lut (.I0(GND_net), .I1(n917), .I2(n98), .I3(n34312), 
            .O(n5825)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2958_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3005_19 (.CI(n35004), .I0(n46887), .I1(n1067), .CO(n35005));
    SB_CARRY add_2958_4 (.CI(n34312), .I0(n917), .I1(n98), .CO(n34313));
    SB_LUT4 add_2958_3_lut (.I0(GND_net), .I1(n918), .I2(n99), .I3(n34311), 
            .O(n5826)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2958_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3005_18_lut (.I0(n1194), .I1(n46887), .I2(n1193), .I3(n35003), 
            .O(displacement_23__N_93[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3005_18_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_2958_3 (.CI(n34311), .I0(n918), .I1(n99), .CO(n34312));
    SB_LUT4 add_2958_2_lut (.I0(GND_net), .I1(n373), .I2(n558), .I3(VCC_net), 
            .O(n5827)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2958_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_11_i1658_3_lut_3_lut (.I0(n2471), .I1(n6948), .I2(n2463), 
            .I3(GND_net), .O(n2550));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1658_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_CARRY add_2958_2 (.CI(VCC_net), .I0(n373), .I1(n558), .CO(n34311));
    SB_CARRY add_3005_18 (.CI(n35003), .I0(n46887), .I1(n1193), .CO(n35004));
    SB_LUT4 div_11_i809_3_lut (.I0(n375), .I1(n6582), .I2(n1193), .I3(GND_net), 
            .O(n1299));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i809_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 LessThan_539_i9_2_lut (.I0(pwm_count[4]), .I1(pwm[4]), .I2(GND_net), 
            .I3(GND_net), .O(n9_adj_4022));   // verilog/motorControl.v(65[19:32])
    defparam LessThan_539_i9_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_3005_17_lut (.I0(n1317), .I1(n46887), .I2(n1316), .I3(n35002), 
            .O(displacement_23__N_93[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3005_17_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_3005_17 (.CI(n35002), .I0(n46887), .I1(n1316), .CO(n35003));
    SB_LUT4 add_3005_16_lut (.I0(n1437), .I1(n46887), .I2(n1436), .I3(n35001), 
            .O(displacement_23__N_93[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3005_16_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_3005_16 (.CI(n35001), .I0(n46887), .I1(n1436), .CO(n35002));
    SB_LUT4 add_3005_15_lut (.I0(n1554), .I1(n46887), .I2(n1553), .I3(n35000), 
            .O(displacement_23__N_93[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3005_15_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 div_11_i1642_3_lut_3_lut (.I0(n2471), .I1(n6932), .I2(n2447), 
            .I3(GND_net), .O(n2534));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1642_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_11_i890_3_lut (.I0(n1299), .I1(n6653), .I2(n1316), .I3(GND_net), 
            .O(n1419));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i890_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY add_3005_15 (.CI(n35000), .I0(n46887), .I1(n1553), .CO(n35001));
    SB_LUT4 add_3005_14_lut (.I0(n1668), .I1(n46887), .I2(n1667), .I3(n34999), 
            .O(displacement_23__N_93[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3005_14_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 LessThan_539_i11_2_lut (.I0(pwm_count[5]), .I1(pwm[5]), .I2(GND_net), 
            .I3(GND_net), .O(n11_adj_4023));   // verilog/motorControl.v(65[19:32])
    defparam LessThan_539_i11_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_3005_14 (.CI(n34999), .I0(n46887), .I1(n1667), .CO(n35000));
    SB_LUT4 add_3005_13_lut (.I0(n1779), .I1(n46887), .I2(n1778), .I3(n34998), 
            .O(displacement_23__N_93[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3005_13_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 LessThan_539_i13_2_lut (.I0(pwm_count[6]), .I1(pwm[6]), .I2(GND_net), 
            .I3(GND_net), .O(n13_adj_4024));   // verilog/motorControl.v(65[19:32])
    defparam LessThan_539_i13_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_3005_13 (.CI(n34998), .I0(n46887), .I1(n1778), .CO(n34999));
    SB_LUT4 div_11_i969_3_lut (.I0(n1419), .I1(n6693), .I2(n1436), .I3(GND_net), 
            .O(n1536));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i969_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_11_i1046_3_lut (.I0(n1536), .I1(n6733), .I2(n1553), .I3(GND_net), 
            .O(n1650));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1046_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 LessThan_539_i4_4_lut (.I0(pwm_count[0]), .I1(pwm[1]), .I2(pwm_count[1]), 
            .I3(pwm[0]), .O(n4_adj_4019));   // verilog/motorControl.v(65[19:32])
    defparam LessThan_539_i4_4_lut.LUT_INIT = 16'h4d0c;
    SB_LUT4 i30133_3_lut (.I0(n4_adj_4019), .I1(pwm[5]), .I2(n11_adj_4023), 
            .I3(GND_net), .O(n45654));   // verilog/motorControl.v(65[19:32])
    defparam i30133_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_11_i1121_3_lut (.I0(n1650), .I1(n6746), .I2(n1667), .I3(GND_net), 
            .O(n1761));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1121_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 add_3005_12_lut (.I0(n1887), .I1(n46887), .I2(n1886), .I3(n34997), 
            .O(displacement_23__N_93[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3005_12_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_3005_12 (.CI(n34997), .I0(n46887), .I1(n1886), .CO(n34998));
    SB_LUT4 add_3005_11_lut (.I0(n1992), .I1(n46887), .I2(n1991), .I3(n34996), 
            .O(displacement_23__N_93[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3005_11_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_3005_11 (.CI(n34996), .I0(n46887), .I1(n1991), .CO(n34997));
    SB_LUT4 div_11_i1194_3_lut (.I0(n1761), .I1(n6787), .I2(n1778), .I3(GND_net), 
            .O(n1869));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1194_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_11_i1643_3_lut_3_lut (.I0(n2471), .I1(n6933), .I2(n2448), 
            .I3(GND_net), .O(n2535));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1643_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i30134_3_lut (.I0(n45654), .I1(pwm[6]), .I2(n13_adj_4024), 
            .I3(GND_net), .O(n45655));   // verilog/motorControl.v(65[19:32])
    defparam i30134_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_11_mux_3_i16_3_lut (.I0(encoder0_position[15]), .I1(n10), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n376));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_mux_3_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_11_i1644_3_lut_3_lut (.I0(n2471), .I1(n6934), .I2(n2449), 
            .I3(GND_net), .O(n2536));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1644_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 add_3005_10_lut (.I0(n2094), .I1(n46887), .I2(n2093), .I3(n34995), 
            .O(displacement_23__N_93[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3005_10_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 div_11_i891_3_lut (.I0(n376), .I1(n6654), .I2(n1316), .I3(GND_net), 
            .O(n1420));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i891_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY add_3005_10 (.CI(n34995), .I0(n46887), .I1(n2093), .CO(n34996));
    SB_LUT4 add_3005_9_lut (.I0(n2193), .I1(n46887), .I2(n2192), .I3(n34994), 
            .O(displacement_23__N_93[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3005_9_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_3005_9 (.CI(n34994), .I0(n46887), .I1(n2192), .CO(n34995));
    SB_LUT4 add_3005_8_lut (.I0(n2289_adj_4007), .I1(n46887), .I2(n2288_adj_4006), 
            .I3(n34993), .O(displacement_23__N_93[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3005_8_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 div_11_i1647_3_lut_3_lut (.I0(n2471), .I1(n6937), .I2(n2452), 
            .I3(GND_net), .O(n2539));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1647_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_CARRY add_3005_8 (.CI(n34993), .I0(n46887), .I1(n2288_adj_4006), 
            .CO(n34994));
    SB_LUT4 div_11_i970_3_lut (.I0(n1420), .I1(n6694), .I2(n1436), .I3(GND_net), 
            .O(n1537));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i970_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_11_i1047_3_lut (.I0(n1537), .I1(n6734), .I2(n1553), .I3(GND_net), 
            .O(n1651));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1047_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_11_i1122_3_lut (.I0(n1651), .I1(n6747), .I2(n1667), .I3(GND_net), 
            .O(n1762));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1122_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_11_i1195_3_lut (.I0(n1762), .I1(n6788), .I2(n1778), .I3(GND_net), 
            .O(n1870));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1195_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_11_i1266_3_lut (.I0(n1870), .I1(n6829), .I2(n1886), .I3(GND_net), 
            .O(n1975));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1266_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_11_i1258_3_lut (.I0(n1862), .I1(n6821), .I2(n1886), .I3(GND_net), 
            .O(n1967));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1258_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_11_i1645_3_lut_3_lut (.I0(n2471), .I1(n6935), .I2(n2450), 
            .I3(GND_net), .O(n2537));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1645_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_11_i1259_3_lut (.I0(n1863), .I1(n6822), .I2(n1886), .I3(GND_net), 
            .O(n1968));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1259_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_11_mux_3_i22_3_lut (.I0(encoder0_position[21]), .I1(n4_adj_3960), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n370));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_mux_3_i22_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_11_i1648_3_lut_3_lut (.I0(n2471), .I1(n6938), .I2(n2453), 
            .I3(GND_net), .O(n2540));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1648_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i20157_2_lut (.I0(n371), .I1(n558), .I2(GND_net), .I3(GND_net), 
            .O(n2));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i20157_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i29194_3_lut (.I0(n370), .I1(n558), .I2(n533), .I3(GND_net), 
            .O(n649));
    defparam i29194_3_lut.LUT_INIT = 16'ha9a9;
    SB_LUT4 div_11_i460_4_lut (.I0(n649), .I1(n2), .I2(n671), .I3(n99), 
            .O(n784));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i460_4_lut.LUT_INIT = 16'ha9a6;
    SB_LUT4 div_11_i549_4_lut (.I0(n784), .I1(n4_adj_3993), .I2(n806), 
            .I3(n98), .O(n916));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i549_4_lut.LUT_INIT = 16'ha9a6;
    SB_LUT4 div_11_i636_3_lut (.I0(n916), .I1(n5824), .I2(n938), .I3(GND_net), 
            .O(n1045));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i636_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_11_i721_3_lut (.I0(n1045), .I1(n6216), .I2(n1067), .I3(GND_net), 
            .O(n1171));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i721_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 add_3005_7_lut (.I0(n2382), .I1(n46887), .I2(n2381), .I3(n34992), 
            .O(displacement_23__N_93[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3005_7_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 div_11_i804_3_lut (.I0(n1171), .I1(n6577), .I2(n1193), .I3(GND_net), 
            .O(n1294));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i804_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i29652_4_lut (.I0(n13_adj_4024), .I1(n11_adj_4023), .I2(n9_adj_4022), 
            .I3(n44526), .O(n45173));
    defparam i29652_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 div_11_i885_3_lut (.I0(n1294), .I1(n6648), .I2(n1316), .I3(GND_net), 
            .O(n1414));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i885_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_11_i964_3_lut (.I0(n1414), .I1(n6688), .I2(n1436), .I3(GND_net), 
            .O(n1531));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i964_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_11_i1661_3_lut_3_lut (.I0(n2471), .I1(n6951), .I2(n387_adj_4001), 
            .I3(GND_net), .O(n2553));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1661_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_11_i1041_3_lut (.I0(n1531), .I1(n6728), .I2(n1553), .I3(GND_net), 
            .O(n1645));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1041_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i28888_3_lut_4_lut (.I0(n1418), .I1(n97), .I2(n98), .I3(n1419), 
            .O(n44407));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i28888_3_lut_4_lut.LUT_INIT = 16'hf99f;
    SB_LUT4 div_11_i1116_3_lut (.I0(n1645), .I1(n6741), .I2(n1667), .I3(GND_net), 
            .O(n1756));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1116_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 LessThan_539_i8_3_lut (.I0(n6_adj_4020), .I1(pwm[4]), .I2(n9_adj_4022), 
            .I3(GND_net), .O(n8_adj_4021));   // verilog/motorControl.v(65[19:32])
    defparam LessThan_539_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_11_i1189_3_lut (.I0(n1756), .I1(n6782), .I2(n1778), .I3(GND_net), 
            .O(n1864));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1189_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_11_i1646_3_lut_3_lut (.I0(n2471), .I1(n6936), .I2(n2451), 
            .I3(GND_net), .O(n2538));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1646_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_11_i1260_3_lut (.I0(n1864), .I1(n6823), .I2(n1886), .I3(GND_net), 
            .O(n1969));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1260_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_11_LessThan_1281_i43_2_lut (.I0(n1969), .I1(n88), .I2(GND_net), 
            .I3(GND_net), .O(n43_adj_4161));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1281_i43_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_11_mux_3_i21_3_lut (.I0(encoder0_position[20]), .I1(n5), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n371));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_mux_3_i21_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_11_i1650_3_lut_3_lut (.I0(n2471), .I1(n6940), .I2(n2455), 
            .I3(GND_net), .O(n2542));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1650_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i20189_2_lut (.I0(n372), .I1(n558), .I2(GND_net), .I3(GND_net), 
            .O(n2_adj_4010));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i20189_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i29186_3_lut (.I0(n371), .I1(n558), .I2(n671), .I3(GND_net), 
            .O(n785));
    defparam i29186_3_lut.LUT_INIT = 16'ha9a9;
    SB_LUT4 div_11_i550_4_lut (.I0(n785), .I1(n2_adj_4010), .I2(n806), 
            .I3(n99), .O(n917));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i550_4_lut.LUT_INIT = 16'ha9a6;
    SB_LUT4 div_11_i637_3_lut (.I0(n917), .I1(n5825), .I2(n938), .I3(GND_net), 
            .O(n1046));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i637_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_11_i722_3_lut (.I0(n1046), .I1(n6217), .I2(n1067), .I3(GND_net), 
            .O(n1172));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i722_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY add_3005_7 (.CI(n34992), .I0(n46887), .I1(n2381), .CO(n34993));
    SB_LUT4 add_3005_6_lut (.I0(n2472), .I1(n46887), .I2(n2471), .I3(n34991), 
            .O(displacement_23__N_93[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3005_6_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_3005_6 (.CI(n34991), .I0(n46887), .I1(n2471), .CO(n34992));
    SB_LUT4 add_3005_5_lut (.I0(n2559), .I1(n46887), .I2(n2558), .I3(n34990), 
            .O(displacement_23__N_93[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3005_5_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_3005_5 (.CI(n34990), .I0(n46887), .I1(n2558), .CO(n34991));
    SB_LUT4 i29585_3_lut (.I0(n45655), .I1(pwm[7]), .I2(n15_adj_4025), 
            .I3(GND_net), .O(n45106));   // verilog/motorControl.v(65[19:32])
    defparam i29585_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_3005_4_lut (.I0(n2643), .I1(n46887), .I2(n2642), .I3(n34989), 
            .O(displacement_23__N_93[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3005_4_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_3005_4 (.CI(n34989), .I0(n46887), .I1(n2642), .CO(n34990));
    SB_LUT4 add_3005_3_lut (.I0(n2724), .I1(n46887), .I2(n2723), .I3(n34988), 
            .O(displacement_23__N_93[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3005_3_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_3005_3 (.CI(n34988), .I0(n46887), .I1(n2723), .CO(n34989));
    SB_LUT4 add_3005_2_lut (.I0(n2802), .I1(n46887), .I2(n2801), .I3(VCC_net), 
            .O(displacement_23__N_93[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3005_2_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 div_11_i805_3_lut (.I0(n1172), .I1(n6578), .I2(n1193), .I3(GND_net), 
            .O(n1295));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i805_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY add_3005_2 (.CI(VCC_net), .I0(n46887), .I1(n2801), .CO(n34988));
    SB_LUT4 add_3004_25_lut (.I0(GND_net), .I1(n2699), .I2(n78), .I3(n34987), 
            .O(n7001)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3004_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3004_24_lut (.I0(GND_net), .I1(n2700), .I2(n79), .I3(n34986), 
            .O(n7002)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3004_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_11_i886_3_lut (.I0(n1295), .I1(n6649), .I2(n1316), .I3(GND_net), 
            .O(n1415));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i886_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_11_i1651_3_lut_3_lut (.I0(n2471), .I1(n6941), .I2(n2456), 
            .I3(GND_net), .O(n2543));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1651_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_DFF displacement_i23 (.Q(displacement[23]), .C(clk32MHz), .D(displacement_23__N_1[23]));   // verilog/TinyFPGA_B.v(161[10] 163[6])
    SB_DFF displacement_i22 (.Q(displacement[22]), .C(clk32MHz), .D(displacement_23__N_1[22]));   // verilog/TinyFPGA_B.v(161[10] 163[6])
    SB_CARRY add_3004_24 (.CI(n34986), .I0(n2700), .I1(n79), .CO(n34987));
    SB_LUT4 add_3004_23_lut (.I0(GND_net), .I1(n2701), .I2(n80), .I3(n34985), 
            .O(n7003)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3004_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i30193_4_lut (.I0(n45106), .I1(n8_adj_4021), .I2(n15_adj_4025), 
            .I3(n45173), .O(n45714));   // verilog/motorControl.v(65[19:32])
    defparam i30193_4_lut.LUT_INIT = 16'haaac;
    SB_CARRY add_3004_23 (.CI(n34985), .I0(n2701), .I1(n80), .CO(n34986));
    SB_LUT4 add_3004_22_lut (.I0(GND_net), .I1(n2702), .I2(n81), .I3(n34984), 
            .O(n7004)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3004_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3004_22 (.CI(n34984), .I0(n2702), .I1(n81), .CO(n34985));
    SB_LUT4 add_3004_21_lut (.I0(GND_net), .I1(n2703), .I2(n82), .I3(n34983), 
            .O(n7005)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3004_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_11_i965_3_lut (.I0(n1415), .I1(n6689), .I2(n1436), .I3(GND_net), 
            .O(n1532));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i965_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY add_3004_21 (.CI(n34983), .I0(n2703), .I1(n82), .CO(n34984));
    SB_LUT4 div_11_i1660_3_lut_3_lut (.I0(n2471), .I1(n6950), .I2(n2465), 
            .I3(GND_net), .O(n2552));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1660_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_11_i1042_3_lut (.I0(n1532), .I1(n6729), .I2(n1553), .I3(GND_net), 
            .O(n1646));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1042_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 add_3004_20_lut (.I0(GND_net), .I1(n2704), .I2(n83), .I3(n34982), 
            .O(n7006)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3004_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3004_20 (.CI(n34982), .I0(n2704), .I1(n83), .CO(n34983));
    SB_LUT4 add_3004_19_lut (.I0(GND_net), .I1(n2705), .I2(n84), .I3(n34981), 
            .O(n7007)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3004_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3004_19 (.CI(n34981), .I0(n2705), .I1(n84), .CO(n34982));
    SB_LUT4 div_11_i1117_3_lut (.I0(n1646), .I1(n6742), .I2(n1667), .I3(GND_net), 
            .O(n1757));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1117_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 add_3004_18_lut (.I0(GND_net), .I1(n2706), .I2(n85), .I3(n34980), 
            .O(n7008)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3004_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3004_18 (.CI(n34980), .I0(n2706), .I1(n85), .CO(n34981));
    SB_LUT4 add_3004_17_lut (.I0(GND_net), .I1(n2707), .I2(n86), .I3(n34979), 
            .O(n7009)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3004_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3004_17 (.CI(n34979), .I0(n2707), .I1(n86), .CO(n34980));
    SB_LUT4 div_11_i1655_3_lut_3_lut (.I0(n2471), .I1(n6945), .I2(n2460), 
            .I3(GND_net), .O(n2547));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1655_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_11_i1649_3_lut_3_lut (.I0(n2471), .I1(n6939), .I2(n2454), 
            .I3(GND_net), .O(n2541));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1649_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_11_i1190_3_lut (.I0(n1757), .I1(n6783), .I2(n1778), .I3(GND_net), 
            .O(n1865));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1190_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_11_i1261_3_lut (.I0(n1865), .I1(n6824), .I2(n1886), .I3(GND_net), 
            .O(n1970));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1261_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 add_3004_16_lut (.I0(GND_net), .I1(n2708), .I2(n87), .I3(n34978), 
            .O(n7010)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3004_16_lut.LUT_INIT = 16'hC33C;
    SB_DFF displacement_i21 (.Q(displacement[21]), .C(clk32MHz), .D(displacement_23__N_1[21]));   // verilog/TinyFPGA_B.v(161[10] 163[6])
    SB_DFF displacement_i20 (.Q(displacement[20]), .C(clk32MHz), .D(displacement_23__N_1[20]));   // verilog/TinyFPGA_B.v(161[10] 163[6])
    SB_DFF displacement_i19 (.Q(displacement[19]), .C(clk32MHz), .D(displacement_23__N_1[19]));   // verilog/TinyFPGA_B.v(161[10] 163[6])
    SB_DFF displacement_i18 (.Q(displacement[18]), .C(clk32MHz), .D(displacement_23__N_1[18]));   // verilog/TinyFPGA_B.v(161[10] 163[6])
    SB_DFF displacement_i17 (.Q(displacement[17]), .C(clk32MHz), .D(displacement_23__N_1[17]));   // verilog/TinyFPGA_B.v(161[10] 163[6])
    SB_DFF displacement_i16 (.Q(displacement[16]), .C(clk32MHz), .D(displacement_23__N_1[16]));   // verilog/TinyFPGA_B.v(161[10] 163[6])
    SB_DFF displacement_i15 (.Q(displacement[15]), .C(clk32MHz), .D(displacement_23__N_1[15]));   // verilog/TinyFPGA_B.v(161[10] 163[6])
    SB_DFF displacement_i14 (.Q(displacement[14]), .C(clk32MHz), .D(displacement_23__N_1[14]));   // verilog/TinyFPGA_B.v(161[10] 163[6])
    SB_DFF displacement_i13 (.Q(displacement[13]), .C(clk32MHz), .D(displacement_23__N_1[13]));   // verilog/TinyFPGA_B.v(161[10] 163[6])
    SB_DFF displacement_i12 (.Q(displacement[12]), .C(clk32MHz), .D(displacement_23__N_1[12]));   // verilog/TinyFPGA_B.v(161[10] 163[6])
    SB_DFF displacement_i11 (.Q(displacement[11]), .C(clk32MHz), .D(displacement_23__N_1[11]));   // verilog/TinyFPGA_B.v(161[10] 163[6])
    SB_DFF displacement_i10 (.Q(displacement[10]), .C(clk32MHz), .D(displacement_23__N_1[10]));   // verilog/TinyFPGA_B.v(161[10] 163[6])
    SB_DFF displacement_i9 (.Q(displacement[9]), .C(clk32MHz), .D(displacement_23__N_1[9]));   // verilog/TinyFPGA_B.v(161[10] 163[6])
    SB_DFF displacement_i8 (.Q(displacement[8]), .C(clk32MHz), .D(displacement_23__N_1[8]));   // verilog/TinyFPGA_B.v(161[10] 163[6])
    SB_DFF displacement_i7 (.Q(displacement[7]), .C(clk32MHz), .D(displacement_23__N_1[7]));   // verilog/TinyFPGA_B.v(161[10] 163[6])
    SB_DFF displacement_i6 (.Q(displacement[6]), .C(clk32MHz), .D(displacement_23__N_1[6]));   // verilog/TinyFPGA_B.v(161[10] 163[6])
    SB_DFF displacement_i5 (.Q(displacement[5]), .C(clk32MHz), .D(displacement_23__N_1[5]));   // verilog/TinyFPGA_B.v(161[10] 163[6])
    SB_DFF displacement_i4 (.Q(displacement[4]), .C(clk32MHz), .D(displacement_23__N_1[4]));   // verilog/TinyFPGA_B.v(161[10] 163[6])
    SB_DFF displacement_i3 (.Q(displacement[3]), .C(clk32MHz), .D(displacement_23__N_1[3]));   // verilog/TinyFPGA_B.v(161[10] 163[6])
    SB_DFF displacement_i2 (.Q(displacement[2]), .C(clk32MHz), .D(displacement_23__N_1[2]));   // verilog/TinyFPGA_B.v(161[10] 163[6])
    SB_DFF displacement_i1 (.Q(displacement[1]), .C(clk32MHz), .D(displacement_23__N_1[1]));   // verilog/TinyFPGA_B.v(161[10] 163[6])
    SB_CARRY add_3004_16 (.CI(n34978), .I0(n2708), .I1(n87), .CO(n34979));
    SB_LUT4 div_11_LessThan_1281_i41_2_lut (.I0(n1970), .I1(n89), .I2(GND_net), 
            .I3(GND_net), .O(n41_adj_4159));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1281_i41_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 add_3004_15_lut (.I0(GND_net), .I1(n2709), .I2(n88), .I3(n34977), 
            .O(n7011)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3004_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3004_15 (.CI(n34977), .I0(n2709), .I1(n88), .CO(n34978));
    SB_LUT4 add_3004_14_lut (.I0(GND_net), .I1(n2710), .I2(n89), .I3(n34976), 
            .O(n7012)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3004_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3004_14 (.CI(n34976), .I0(n2710), .I1(n89), .CO(n34977));
    SB_LUT4 div_11_mux_3_i20_3_lut (.I0(encoder0_position[19]), .I1(n6_adj_3959), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n372));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_mux_3_i20_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_3004_13_lut (.I0(GND_net), .I1(n2711), .I2(n90), .I3(n34975), 
            .O(n7013)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3004_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3004_13 (.CI(n34975), .I0(n2711), .I1(n90), .CO(n34976));
    SB_LUT4 i29183_3_lut (.I0(n372), .I1(n558), .I2(n806), .I3(GND_net), 
            .O(n918));
    defparam i29183_3_lut.LUT_INIT = 16'ha9a9;
    SB_LUT4 add_3004_12_lut (.I0(GND_net), .I1(n2712), .I2(n91), .I3(n34974), 
            .O(n7014)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3004_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_11_i1654_3_lut_3_lut (.I0(n2471), .I1(n6944), .I2(n2459), 
            .I3(GND_net), .O(n2546));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1654_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_CARRY add_3004_12 (.CI(n34974), .I0(n2712), .I1(n91), .CO(n34975));
    SB_LUT4 add_3004_11_lut (.I0(GND_net), .I1(n2713), .I2(n92), .I3(n34973), 
            .O(n7015)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3004_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3004_11 (.CI(n34973), .I0(n2713), .I1(n92), .CO(n34974));
    SB_LUT4 add_3004_10_lut (.I0(GND_net), .I1(n2714), .I2(n93), .I3(n34972), 
            .O(n7016)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3004_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_11_LessThan_906_i34_3_lut_3_lut (.I0(n1418), .I1(n97), .I2(n98), 
            .I3(GND_net), .O(n34_adj_4091));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_906_i34_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 div_11_i638_3_lut (.I0(n918), .I1(n5826), .I2(n938), .I3(GND_net), 
            .O(n1047));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i638_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY add_3004_10 (.CI(n34972), .I0(n2714), .I1(n93), .CO(n34973));
    SB_LUT4 add_3004_9_lut (.I0(GND_net), .I1(n2715), .I2(n94), .I3(n34971), 
            .O(n7017)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3004_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3004_9 (.CI(n34971), .I0(n2715), .I1(n94), .CO(n34972));
    SB_LUT4 add_3004_8_lut (.I0(GND_net), .I1(n2716), .I2(n95), .I3(n34970), 
            .O(n7018)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3004_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_11_i723_3_lut (.I0(n1047), .I1(n6218), .I2(n1067), .I3(GND_net), 
            .O(n1173));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i723_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY add_3004_8 (.CI(n34970), .I0(n2716), .I1(n95), .CO(n34971));
    SB_LUT4 div_11_i806_3_lut (.I0(n1173), .I1(n6579), .I2(n1193), .I3(GND_net), 
            .O(n1296));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i806_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 add_3004_7_lut (.I0(GND_net), .I1(n2717), .I2(n96), .I3(n34969), 
            .O(n7019)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3004_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3004_7 (.CI(n34969), .I0(n2717), .I1(n96), .CO(n34970));
    SB_LUT4 add_3004_6_lut (.I0(GND_net), .I1(n2718), .I2(n97), .I3(n34968), 
            .O(n7020)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3004_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_11_i1653_3_lut_3_lut (.I0(n2471), .I1(n6943), .I2(n2458), 
            .I3(GND_net), .O(n2545));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1653_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_CARRY add_3004_6 (.CI(n34968), .I0(n2718), .I1(n97), .CO(n34969));
    SB_LUT4 div_11_i887_3_lut (.I0(n1296), .I1(n6650), .I2(n1316), .I3(GND_net), 
            .O(n1416));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i887_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 add_3004_5_lut (.I0(GND_net), .I1(n2719), .I2(n98), .I3(n34967), 
            .O(n7021)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3004_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3004_5 (.CI(n34967), .I0(n2719), .I1(n98), .CO(n34968));
    SB_LUT4 add_3004_4_lut (.I0(GND_net), .I1(n2720), .I2(n99), .I3(n34966), 
            .O(n7022)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3004_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_11_i966_3_lut (.I0(n1416), .I1(n6690), .I2(n1436), .I3(GND_net), 
            .O(n1533));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i966_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY add_3004_4 (.CI(n34966), .I0(n2720), .I1(n99), .CO(n34967));
    SB_LUT4 add_3004_3_lut (.I0(GND_net), .I1(n390), .I2(n558), .I3(n34965), 
            .O(n7023)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3004_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3004_3 (.CI(n34965), .I0(n390), .I1(n558), .CO(n34966));
    SB_CARRY add_3004_2 (.CI(VCC_net), .I0(n391), .I1(VCC_net), .CO(n34965));
    SB_LUT4 div_11_i1043_3_lut (.I0(n1533), .I1(n6730), .I2(n1553), .I3(GND_net), 
            .O(n1647));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1043_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_11_i1118_3_lut (.I0(n1647), .I1(n6743), .I2(n1667), .I3(GND_net), 
            .O(n1758));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1118_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 add_3003_23_lut (.I0(GND_net), .I1(n2618), .I2(n79), .I3(n34964), 
            .O(n6977)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3003_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_11_i1652_3_lut_3_lut (.I0(n2471), .I1(n6942), .I2(n2457), 
            .I3(GND_net), .O(n2544));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1652_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_11_i1191_3_lut (.I0(n1758), .I1(n6784), .I2(n1778), .I3(GND_net), 
            .O(n1866));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1191_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 add_3003_22_lut (.I0(GND_net), .I1(n2619), .I2(n80), .I3(n34963), 
            .O(n6978)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3003_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_11_i1262_3_lut (.I0(n1866), .I1(n6825), .I2(n1886), .I3(GND_net), 
            .O(n1971));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1262_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY add_3003_22 (.CI(n34963), .I0(n2619), .I1(n80), .CO(n34964));
    SB_LUT4 add_3003_21_lut (.I0(GND_net), .I1(n2620), .I2(n81), .I3(n34962), 
            .O(n6979)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3003_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3003_21 (.CI(n34962), .I0(n2620), .I1(n81), .CO(n34963));
    SB_LUT4 div_11_LessThan_1281_i39_2_lut (.I0(n1971), .I1(n90), .I2(GND_net), 
            .I3(GND_net), .O(n39_adj_4158));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1281_i39_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_11_mux_5_i11_3_lut (.I0(gearBoxRatio[10]), .I1(n65), .I2(gearBoxRatio[23]), 
            .I3(GND_net), .O(n90));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_mux_5_i11_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 div_11_mux_3_i19_3_lut (.I0(encoder0_position[18]), .I1(n7), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n373));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_mux_3_i19_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_3003_20_lut (.I0(GND_net), .I1(n2621), .I2(n82), .I3(n34961), 
            .O(n6980)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3003_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3003_20 (.CI(n34961), .I0(n2621), .I1(n82), .CO(n34962));
    SB_LUT4 div_11_i639_3_lut (.I0(n373), .I1(n5827), .I2(n938), .I3(GND_net), 
            .O(n1048));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i639_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 add_3003_19_lut (.I0(GND_net), .I1(n2622), .I2(n83), .I3(n34960), 
            .O(n6981)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3003_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3003_19 (.CI(n34960), .I0(n2622), .I1(n83), .CO(n34961));
    SB_LUT4 add_3003_18_lut (.I0(GND_net), .I1(n2623), .I2(n84), .I3(n34959), 
            .O(n6982)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3003_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3003_18 (.CI(n34959), .I0(n2623), .I1(n84), .CO(n34960));
    SB_LUT4 div_11_i724_3_lut (.I0(n1048), .I1(n6219), .I2(n1067), .I3(GND_net), 
            .O(n1174));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i724_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 add_3003_17_lut (.I0(GND_net), .I1(n2624), .I2(n85), .I3(n34958), 
            .O(n6983)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3003_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3003_17 (.CI(n34958), .I0(n2624), .I1(n85), .CO(n34959));
    SB_LUT4 div_11_i1659_3_lut_3_lut (.I0(n2471), .I1(n6949), .I2(n2464), 
            .I3(GND_net), .O(n2551));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1659_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 add_3003_16_lut (.I0(GND_net), .I1(n2625), .I2(n86), .I3(n34957), 
            .O(n6984)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3003_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3003_16 (.CI(n34957), .I0(n2625), .I1(n86), .CO(n34958));
    SB_LUT4 add_3003_15_lut (.I0(GND_net), .I1(n2626), .I2(n87), .I3(n34956), 
            .O(n6985)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3003_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_11_i807_3_lut (.I0(n1174), .I1(n6580), .I2(n1193), .I3(GND_net), 
            .O(n1297));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i807_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY add_3003_15 (.CI(n34956), .I0(n2626), .I1(n87), .CO(n34957));
    SB_LUT4 add_3003_14_lut (.I0(GND_net), .I1(n2627), .I2(n88), .I3(n34955), 
            .O(n6986)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3003_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3003_14 (.CI(n34955), .I0(n2627), .I1(n88), .CO(n34956));
    SB_LUT4 div_11_i888_3_lut (.I0(n1297), .I1(n6651), .I2(n1316), .I3(GND_net), 
            .O(n1417));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i888_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_11_i967_3_lut (.I0(n1417), .I1(n6691), .I2(n1436), .I3(GND_net), 
            .O(n1534));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i967_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_11_i1044_3_lut (.I0(n1534), .I1(n6731), .I2(n1553), .I3(GND_net), 
            .O(n1648));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1044_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 add_3003_13_lut (.I0(GND_net), .I1(n2628), .I2(n89), .I3(n34954), 
            .O(n6987)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3003_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3003_13 (.CI(n34954), .I0(n2628), .I1(n89), .CO(n34955));
    SB_LUT4 add_3003_12_lut (.I0(GND_net), .I1(n2629), .I2(n90), .I3(n34953), 
            .O(n6988)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3003_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_11_i1119_3_lut (.I0(n1648), .I1(n6744), .I2(n1667), .I3(GND_net), 
            .O(n1759));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1119_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY add_3003_12 (.CI(n34953), .I0(n2629), .I1(n90), .CO(n34954));
    SB_LUT4 div_11_i1656_3_lut_3_lut (.I0(n2471), .I1(n6946), .I2(n2461), 
            .I3(GND_net), .O(n2548));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1656_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 add_3003_11_lut (.I0(GND_net), .I1(n2630), .I2(n91), .I3(n34952), 
            .O(n6989)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3003_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_11_i1192_3_lut (.I0(n1759), .I1(n6785), .I2(n1778), .I3(GND_net), 
            .O(n1867));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1192_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY add_3003_11 (.CI(n34952), .I0(n2630), .I1(n91), .CO(n34953));
    SB_LUT4 i28903_3_lut_4_lut (.I0(n1297), .I1(n97), .I2(n98), .I3(n1298), 
            .O(n44422));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i28903_3_lut_4_lut.LUT_INIT = 16'hf99f;
    SB_LUT4 add_3003_10_lut (.I0(GND_net), .I1(n2631), .I2(n92), .I3(n34951), 
            .O(n6990)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3003_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3003_10 (.CI(n34951), .I0(n2631), .I1(n92), .CO(n34952));
    SB_LUT4 add_3003_9_lut (.I0(GND_net), .I1(n2632), .I2(n93), .I3(n34950), 
            .O(n6991)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3003_9_lut.LUT_INIT = 16'hC33C;
    SB_IO PIN_6_pad (.PACKAGE_PIN(PIN_6), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(PIN_6_c_0)) /* synthesis IO_FF_OUT=TRUE */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam PIN_6_pad.PIN_TYPE = 6'b011001;
    defparam PIN_6_pad.PULLUP = 1'b0;
    defparam PIN_6_pad.NEG_TRIGGER = 1'b0;
    defparam PIN_6_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO USBPU_pad (.PACKAGE_PIN(USBPU), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(GND_net));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam USBPU_pad.PIN_TYPE = 6'b011001;
    defparam USBPU_pad.PULLUP = 1'b0;
    defparam USBPU_pad.NEG_TRIGGER = 1'b0;
    defparam USBPU_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO LED_pad (.PACKAGE_PIN(LED), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(LED_c)) /* synthesis IO_FF_OUT=TRUE */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam LED_pad.PIN_TYPE = 6'b011001;
    defparam LED_pad.PULLUP = 1'b0;
    defparam LED_pad.NEG_TRIGGER = 1'b0;
    defparam LED_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO PIN_24_pad (.PACKAGE_PIN(PIN_24), .OUTPUT_ENABLE(VCC_net), .D_IN_0(PIN_24_c_0)) /* synthesis IO_FF_IN=TRUE */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam PIN_24_pad.PIN_TYPE = 6'b000001;
    defparam PIN_24_pad.PULLUP = 1'b0;
    defparam PIN_24_pad.NEG_TRIGGER = 1'b0;
    defparam PIN_24_pad.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 div_11_i1657_3_lut_3_lut (.I0(n2471), .I1(n6947), .I2(n2462), 
            .I3(GND_net), .O(n2549));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1657_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_11_i1707_3_lut_3_lut (.I0(n2558), .I1(n6962), .I2(n2542), 
            .I3(GND_net), .O(n2626));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1707_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_11_i1263_3_lut (.I0(n1867), .I1(n6826), .I2(n1886), .I3(GND_net), 
            .O(n1972));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1263_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY add_3003_9 (.CI(n34950), .I0(n2632), .I1(n93), .CO(n34951));
    SB_LUT4 div_11_i1699_3_lut_3_lut (.I0(n2558), .I1(n6954), .I2(n2534), 
            .I3(GND_net), .O(n2618));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1699_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_11_LessThan_1281_i37_2_lut (.I0(n1972), .I1(n91), .I2(GND_net), 
            .I3(GND_net), .O(n37_adj_4157));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1281_i37_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_11_mux_3_i14_3_lut (.I0(encoder0_position[13]), .I1(n12), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n378));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_mux_3_i14_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_11_i1049_3_lut (.I0(n378), .I1(n6736), .I2(n1553), .I3(GND_net), 
            .O(n1653));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1049_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_11_i1124_3_lut (.I0(n1653), .I1(n6749), .I2(n1667), .I3(GND_net), 
            .O(n1764));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1124_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_11_i1700_3_lut_3_lut (.I0(n2558), .I1(n6955), .I2(n2535), 
            .I3(GND_net), .O(n2619));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1700_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_11_LessThan_825_i36_3_lut_3_lut (.I0(n1297), .I1(n97), .I2(n98), 
            .I3(GND_net), .O(n36_adj_4085));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_825_i36_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 div_11_i1701_3_lut_3_lut (.I0(n2558), .I1(n6956), .I2(n2536), 
            .I3(GND_net), .O(n2620));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1701_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 add_3003_8_lut (.I0(GND_net), .I1(n2633), .I2(n94), .I3(n34949), 
            .O(n6992)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3003_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3003_8 (.CI(n34949), .I0(n2633), .I1(n94), .CO(n34950));
    SB_LUT4 div_11_i1702_3_lut_3_lut (.I0(n2558), .I1(n6957), .I2(n2537), 
            .I3(GND_net), .O(n2621));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1702_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 add_3003_7_lut (.I0(GND_net), .I1(n2634), .I2(n95), .I3(n34948), 
            .O(n6993)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3003_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3003_7 (.CI(n34948), .I0(n2634), .I1(n95), .CO(n34949));
    SB_LUT4 div_11_i1705_3_lut_3_lut (.I0(n2558), .I1(n6960), .I2(n2540), 
            .I3(GND_net), .O(n2624));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1705_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_11_i1197_3_lut (.I0(n1764), .I1(n6790), .I2(n1778), .I3(GND_net), 
            .O(n1872));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1197_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 add_3003_6_lut (.I0(GND_net), .I1(n2635), .I2(n96), .I3(n34947), 
            .O(n6994)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3003_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3003_6 (.CI(n34947), .I0(n2635), .I1(n96), .CO(n34948));
    SB_LUT4 div_11_i1268_3_lut (.I0(n1872), .I1(n6831), .I2(n1886), .I3(GND_net), 
            .O(n1977));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1268_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 add_3003_5_lut (.I0(GND_net), .I1(n2636), .I2(n97), .I3(n34946), 
            .O(n6995)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3003_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_11_LessThan_1281_i27_2_lut (.I0(n1977), .I1(n96), .I2(GND_net), 
            .I3(GND_net), .O(n27_adj_4149));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1281_i27_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_11_i1703_3_lut_3_lut (.I0(n2558), .I1(n6958), .I2(n2538), 
            .I3(GND_net), .O(n2622));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1703_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_CARRY add_3003_5 (.CI(n34946), .I0(n2636), .I1(n97), .CO(n34947));
    SB_LUT4 div_11_mux_3_i13_3_lut (.I0(encoder0_position[12]), .I1(n13), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n379));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_mux_3_i13_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_11_i1125_3_lut (.I0(n379), .I1(n6750), .I2(n1667), .I3(GND_net), 
            .O(n1765));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1125_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 add_3003_4_lut (.I0(GND_net), .I1(n2637), .I2(n98), .I3(n34945), 
            .O(n6996)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3003_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3003_4 (.CI(n34945), .I0(n2637), .I1(n98), .CO(n34946));
    SB_LUT4 add_3003_3_lut (.I0(GND_net), .I1(n2638), .I2(n99), .I3(n34944), 
            .O(n6997)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3003_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3003_3 (.CI(n34944), .I0(n2638), .I1(n99), .CO(n34945));
    SB_LUT4 div_11_i1198_3_lut (.I0(n1765), .I1(n6791), .I2(n1778), .I3(GND_net), 
            .O(n1873));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1198_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 add_3003_2_lut (.I0(GND_net), .I1(n389), .I2(n558), .I3(VCC_net), 
            .O(n6998)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3003_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3003_2 (.CI(VCC_net), .I0(n389), .I1(n558), .CO(n34944));
    SB_LUT4 add_3002_22_lut (.I0(GND_net), .I1(n2534), .I2(n80), .I3(n34943), 
            .O(n6954)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3002_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_11_i1269_3_lut (.I0(n1873), .I1(n6832), .I2(n1886), .I3(GND_net), 
            .O(n1978));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1269_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 displacement_23__I_0_add_2_25_lut (.I0(GND_net), .I1(displacement_23__N_93[23]), 
            .I2(n3_adj_4000), .I3(n34262), .O(displacement_23__N_1[23])) /* synthesis syn_instantiated=1 */ ;
    defparam displacement_23__I_0_add_2_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3002_21_lut (.I0(GND_net), .I1(n2535), .I2(n81), .I3(n34942), 
            .O(n6955)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3002_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 displacement_23__I_0_add_2_24_lut (.I0(GND_net), .I1(displacement_23__N_93[22]), 
            .I2(n3_adj_4000), .I3(n34261), .O(displacement_23__N_1[22])) /* synthesis syn_instantiated=1 */ ;
    defparam displacement_23__I_0_add_2_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY displacement_23__I_0_add_2_24 (.CI(n34261), .I0(displacement_23__N_93[22]), 
            .I1(n3_adj_4000), .CO(n34262));
    SB_LUT4 displacement_23__I_0_add_2_23_lut (.I0(GND_net), .I1(displacement_23__N_93[21]), 
            .I2(n3_adj_4000), .I3(n34260), .O(displacement_23__N_1[21])) /* synthesis syn_instantiated=1 */ ;
    defparam displacement_23__I_0_add_2_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_11_LessThan_1281_i25_2_lut (.I0(n1978), .I1(n97), .I2(GND_net), 
            .I3(GND_net), .O(n25_adj_4147));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1281_i25_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_11_mux_3_i18_3_lut (.I0(encoder0_position[17]), .I1(n8), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n374));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_mux_3_i18_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_11_i725_3_lut (.I0(n374), .I1(n6220), .I2(n1067), .I3(GND_net), 
            .O(n1175));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i725_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY add_3002_21 (.CI(n34942), .I0(n2535), .I1(n81), .CO(n34943));
    SB_CARRY displacement_23__I_0_add_2_23 (.CI(n34260), .I0(displacement_23__N_93[21]), 
            .I1(n3_adj_4000), .CO(n34261));
    SB_LUT4 displacement_23__I_0_add_2_22_lut (.I0(GND_net), .I1(displacement_23__N_93[20]), 
            .I2(n3_adj_4000), .I3(n34259), .O(displacement_23__N_1[20])) /* synthesis syn_instantiated=1 */ ;
    defparam displacement_23__I_0_add_2_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3002_20_lut (.I0(GND_net), .I1(n2536), .I2(n82), .I3(n34941), 
            .O(n6956)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3002_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_11_i1706_3_lut_3_lut (.I0(n2558), .I1(n6961), .I2(n2541), 
            .I3(GND_net), .O(n2625));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1706_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_11_i808_3_lut (.I0(n1175), .I1(n6581), .I2(n1193), .I3(GND_net), 
            .O(n1298));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i808_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_11_i889_3_lut (.I0(n1298), .I1(n6652), .I2(n1316), .I3(GND_net), 
            .O(n1418));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i889_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_11_i1719_3_lut_3_lut (.I0(n2558), .I1(n6974), .I2(n388), 
            .I3(GND_net), .O(n2638));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1719_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_CARRY displacement_23__I_0_add_2_22 (.CI(n34259), .I0(displacement_23__N_93[20]), 
            .I1(n3_adj_4000), .CO(n34260));
    SB_LUT4 displacement_23__I_0_add_2_21_lut (.I0(GND_net), .I1(displacement_23__N_93[19]), 
            .I2(n6_adj_3983), .I3(n34258), .O(displacement_23__N_1[19])) /* synthesis syn_instantiated=1 */ ;
    defparam displacement_23__I_0_add_2_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3002_20 (.CI(n34941), .I0(n2536), .I1(n82), .CO(n34942));
    SB_LUT4 div_11_i968_3_lut (.I0(n1418), .I1(n6692), .I2(n1436), .I3(GND_net), 
            .O(n1535));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i968_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_11_i1045_3_lut (.I0(n1535), .I1(n6732), .I2(n1553), .I3(GND_net), 
            .O(n1649));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1045_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 add_3002_19_lut (.I0(GND_net), .I1(n2537), .I2(n83), .I3(n34940), 
            .O(n6957)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3002_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3002_19 (.CI(n34940), .I0(n2537), .I1(n83), .CO(n34941));
    SB_LUT4 div_11_i1120_3_lut (.I0(n1649), .I1(n6745), .I2(n1667), .I3(GND_net), 
            .O(n1760));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1120_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 add_3002_18_lut (.I0(GND_net), .I1(n2538), .I2(n84), .I3(n34939), 
            .O(n6958)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3002_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_11_i1193_3_lut (.I0(n1760), .I1(n6786), .I2(n1778), .I3(GND_net), 
            .O(n1868));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1193_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY add_3002_18 (.CI(n34939), .I0(n2538), .I1(n84), .CO(n34940));
    SB_LUT4 div_11_i1264_3_lut (.I0(n1868), .I1(n6827), .I2(n1886), .I3(GND_net), 
            .O(n1973));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1264_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_11_LessThan_1281_i35_2_lut (.I0(n1973), .I1(n92), .I2(GND_net), 
            .I3(GND_net), .O(n35_adj_4156));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1281_i35_2_lut.LUT_INIT = 16'h9999;
    SB_CARRY displacement_23__I_0_add_2_21 (.CI(n34258), .I0(displacement_23__N_93[19]), 
            .I1(n6_adj_3983), .CO(n34259));
    SB_LUT4 displacement_23__I_0_add_2_20_lut (.I0(GND_net), .I1(displacement_23__N_93[18]), 
            .I2(n7_adj_3982), .I3(n34257), .O(displacement_23__N_1[18])) /* synthesis syn_instantiated=1 */ ;
    defparam displacement_23__I_0_add_2_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3002_17_lut (.I0(GND_net), .I1(n2539), .I2(n85), .I3(n34938), 
            .O(n6959)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3002_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY displacement_23__I_0_add_2_20 (.CI(n34257), .I0(displacement_23__N_93[18]), 
            .I1(n7_adj_3982), .CO(n34258));
    SB_LUT4 displacement_23__I_0_add_2_19_lut (.I0(GND_net), .I1(displacement_23__N_93[17]), 
            .I2(n8_adj_3981), .I3(n34256), .O(displacement_23__N_1[17])) /* synthesis syn_instantiated=1 */ ;
    defparam displacement_23__I_0_add_2_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_11_mux_5_i10_3_lut (.I0(gearBoxRatio[9]), .I1(n66), .I2(gearBoxRatio[23]), 
            .I3(GND_net), .O(n91));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_mux_5_i10_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 i1_2_lut_adj_1450 (.I0(n92), .I1(n22424), .I2(GND_net), .I3(GND_net), 
            .O(n22421));
    defparam i1_2_lut_adj_1450.LUT_INIT = 16'hdddd;
    SB_LUT4 div_11_i1704_3_lut_3_lut (.I0(n2558), .I1(n6959), .I2(n2539), 
            .I3(GND_net), .O(n2623));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1704_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_CARRY add_3002_17 (.CI(n34938), .I0(n2539), .I1(n85), .CO(n34939));
    SB_CARRY displacement_23__I_0_add_2_19 (.CI(n34256), .I0(displacement_23__N_93[17]), 
            .I1(n8_adj_3981), .CO(n34257));
    SB_LUT4 i1_2_lut_adj_1451 (.I0(n95), .I1(n22415), .I2(GND_net), .I3(GND_net), 
            .O(n22412));
    defparam i1_2_lut_adj_1451.LUT_INIT = 16'hdddd;
    SB_LUT4 i1_2_lut_adj_1452 (.I0(n98), .I1(n22406), .I2(GND_net), .I3(GND_net), 
            .O(n22403));
    defparam i1_2_lut_adj_1452.LUT_INIT = 16'hdddd;
    SB_LUT4 i1_4_lut (.I0(n224), .I1(n99), .I2(n22403), .I3(n558), .O(n5_adj_4360));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i1_4_lut.LUT_INIT = 16'h555d;
    SB_LUT4 displacement_23__I_0_add_2_18_lut (.I0(GND_net), .I1(displacement_23__N_93[16]), 
            .I2(n9_adj_3980), .I3(n34255), .O(displacement_23__N_1[16])) /* synthesis syn_instantiated=1 */ ;
    defparam displacement_23__I_0_add_2_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY displacement_23__I_0_add_2_18 (.CI(n34255), .I0(displacement_23__N_93[16]), 
            .I1(n9_adj_3980), .CO(n34256));
    SB_LUT4 displacement_23__I_0_add_2_17_lut (.I0(GND_net), .I1(displacement_23__N_93[15]), 
            .I2(n10_adj_3979), .I3(n34254), .O(displacement_23__N_1[15])) /* synthesis syn_instantiated=1 */ ;
    defparam displacement_23__I_0_add_2_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_11_i1708_3_lut_3_lut (.I0(n2558), .I1(n6963), .I2(n2543), 
            .I3(GND_net), .O(n2627));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1708_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 add_3002_16_lut (.I0(GND_net), .I1(n2540), .I2(n86), .I3(n34937), 
            .O(n6960)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3002_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3002_16 (.CI(n34937), .I0(n2540), .I1(n86), .CO(n34938));
    SB_LUT4 add_3002_15_lut (.I0(GND_net), .I1(n2541), .I2(n87), .I3(n34936), 
            .O(n6961)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3002_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3002_15 (.CI(n34936), .I0(n2541), .I1(n87), .CO(n34937));
    SB_LUT4 add_3002_14_lut (.I0(GND_net), .I1(n2542), .I2(n88), .I3(n34935), 
            .O(n6962)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3002_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3002_14 (.CI(n34935), .I0(n2542), .I1(n88), .CO(n34936));
    SB_LUT4 add_3002_13_lut (.I0(GND_net), .I1(n2543), .I2(n89), .I3(n34934), 
            .O(n6963)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3002_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i20117_2_lut (.I0(n369), .I1(n558), .I2(GND_net), .I3(GND_net), 
            .O(n2_adj_3958));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i20117_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 div_11_i274_4_lut (.I0(n5_adj_4360), .I1(n2_adj_3958), .I2(n392), 
            .I3(n99), .O(n40890));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i274_4_lut.LUT_INIT = 16'ha9a6;
    SB_CARRY displacement_23__I_0_add_2_17 (.CI(n34254), .I0(displacement_23__N_93[15]), 
            .I1(n10_adj_3979), .CO(n34255));
    SB_CARRY add_3002_13 (.CI(n34934), .I0(n2543), .I1(n89), .CO(n34935));
    SB_LUT4 div_11_i367_4_lut (.I0(n40890), .I1(n4_adj_3956), .I2(n533), 
            .I3(n98), .O(n40892));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i367_4_lut.LUT_INIT = 16'ha9a6;
    SB_LUT4 div_11_mux_5_i5_3_lut (.I0(gearBoxRatio[4]), .I1(n71), .I2(gearBoxRatio[23]), 
            .I3(GND_net), .O(n96));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_mux_5_i5_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 i20173_3_lut (.I0(n648), .I1(n98), .I2(n4), .I3(GND_net), 
            .O(n6));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i20173_3_lut.LUT_INIT = 16'he8e8;
    SB_LUT4 div_11_i458_4_lut (.I0(n40892), .I1(n6), .I2(n671), .I3(n97), 
            .O(n40894));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i458_4_lut.LUT_INIT = 16'ha9a6;
    SB_LUT4 add_3002_12_lut (.I0(GND_net), .I1(n2544), .I2(n90), .I3(n34933), 
            .O(n6964)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3002_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_11_i1709_3_lut_3_lut (.I0(n2558), .I1(n6964), .I2(n2544), 
            .I3(GND_net), .O(n2628));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1709_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i20213_3_lut (.I0(n783), .I1(n97), .I2(n6_adj_3989), .I3(GND_net), 
            .O(n8_adj_3986));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i20213_3_lut.LUT_INIT = 16'he8e8;
    SB_LUT4 div_11_i547_4_lut (.I0(n40894), .I1(n8_adj_3986), .I2(n806), 
            .I3(n96), .O(n914));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i547_4_lut.LUT_INIT = 16'h5659;
    SB_LUT4 div_11_i634_3_lut (.I0(n914), .I1(n5822), .I2(n938), .I3(GND_net), 
            .O(n1043));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i634_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 displacement_23__I_0_add_2_16_lut (.I0(GND_net), .I1(displacement_23__N_93[14]), 
            .I2(n11_adj_3978), .I3(n34253), .O(displacement_23__N_1[14])) /* synthesis syn_instantiated=1 */ ;
    defparam displacement_23__I_0_add_2_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3002_12 (.CI(n34933), .I0(n2544), .I1(n90), .CO(n34934));
    SB_CARRY displacement_23__I_0_add_2_16 (.CI(n34253), .I0(displacement_23__N_93[14]), 
            .I1(n11_adj_3978), .CO(n34254));
    SB_LUT4 div_11_i719_3_lut (.I0(n1043), .I1(n6214), .I2(n1067), .I3(GND_net), 
            .O(n1169));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i719_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_11_i802_3_lut (.I0(n1169), .I1(n6575), .I2(n1193), .I3(GND_net), 
            .O(n1292));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i802_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_11_i1710_3_lut_3_lut (.I0(n2558), .I1(n6965), .I2(n2545), 
            .I3(GND_net), .O(n2629));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1710_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_11_i883_3_lut (.I0(n1292), .I1(n6646), .I2(n1316), .I3(GND_net), 
            .O(n1412));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i883_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 displacement_23__I_0_add_2_15_lut (.I0(GND_net), .I1(displacement_23__N_93[13]), 
            .I2(n12_adj_3977), .I3(n34252), .O(displacement_23__N_1[13])) /* synthesis syn_instantiated=1 */ ;
    defparam displacement_23__I_0_add_2_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_11_i962_3_lut (.I0(n1412), .I1(n6686), .I2(n1436), .I3(GND_net), 
            .O(n1529));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i962_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_11_i1039_3_lut (.I0(n1529), .I1(n6726), .I2(n1553), .I3(GND_net), 
            .O(n1643));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1039_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_11_i1114_3_lut (.I0(n1643), .I1(n6739), .I2(n1667), .I3(GND_net), 
            .O(n1754));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1114_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i28982_2_lut (.I0(n369), .I1(n558), .I2(GND_net), .I3(GND_net), 
            .O(n44075));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i28982_2_lut.LUT_INIT = 16'h1111;
    SB_LUT4 div_11_i1711_3_lut_3_lut (.I0(n2558), .I1(n6966), .I2(n2546), 
            .I3(GND_net), .O(n2630));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1711_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i1_4_lut_adj_1453 (.I0(n44075), .I1(n22403), .I2(n99), .I3(n5_adj_4360), 
            .O(n392));
    defparam i1_4_lut_adj_1453.LUT_INIT = 16'hefce;
    SB_LUT4 div_11_mux_3_i23_3_lut (.I0(encoder0_position[22]), .I1(n3), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n369));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_mux_3_i23_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_11_LessThan_297_i46_4_lut (.I0(n370), .I1(n99), .I2(n510), 
            .I3(n558), .O(n46));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_297_i46_4_lut.LUT_INIT = 16'h0317;
    SB_LUT4 i1_4_lut_adj_1454 (.I0(n46), .I1(n22406), .I2(n98), .I3(n40890), 
            .O(n533));
    defparam i1_4_lut_adj_1454.LUT_INIT = 16'hefce;
    SB_LUT4 i20133_2_lut (.I0(n370), .I1(n558), .I2(GND_net), .I3(GND_net), 
            .O(n2_adj_3957));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i20133_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 add_3002_11_lut (.I0(GND_net), .I1(n2545), .I2(n91), .I3(n34932), 
            .O(n6965)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3002_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_11_i1715_3_lut_3_lut (.I0(n2558), .I1(n6970), .I2(n2550), 
            .I3(GND_net), .O(n2634));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1715_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i29199_3_lut (.I0(n369), .I1(n558), .I2(n392), .I3(GND_net), 
            .O(n510));
    defparam i29199_3_lut.LUT_INIT = 16'ha9a9;
    SB_LUT4 div_11_LessThan_390_i44_4_lut (.I0(n371), .I1(n99), .I2(n649), 
            .I3(n558), .O(n44));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_390_i44_4_lut.LUT_INIT = 16'h0317;
    SB_LUT4 i29983_3_lut (.I0(n44), .I1(n98), .I2(n648), .I3(GND_net), 
            .O(n45504));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i29983_3_lut.LUT_INIT = 16'h2b2b;
    SB_LUT4 i1_4_lut_adj_1455 (.I0(n45504), .I1(n22409), .I2(n97), .I3(n40892), 
            .O(n671));
    defparam i1_4_lut_adj_1455.LUT_INIT = 16'hefce;
    SB_LUT4 div_11_i368_4_lut (.I0(n510), .I1(n2_adj_3957), .I2(n533), 
            .I3(n99), .O(n648));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i368_4_lut.LUT_INIT = 16'ha9a6;
    SB_LUT4 div_11_mux_5_i4_3_lut (.I0(gearBoxRatio[3]), .I1(n72), .I2(gearBoxRatio[23]), 
            .I3(GND_net), .O(n97));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_mux_5_i4_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 div_11_LessThan_481_i42_4_lut (.I0(n372), .I1(n99), .I2(n785), 
            .I3(n558), .O(n42));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_481_i42_4_lut.LUT_INIT = 16'h0317;
    SB_LUT4 i30419_3_lut (.I0(n42), .I1(n98), .I2(n784), .I3(GND_net), 
            .O(n45940));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i30419_3_lut.LUT_INIT = 16'h2b2b;
    SB_LUT4 i30420_3_lut (.I0(n45940), .I1(n97), .I2(n783), .I3(GND_net), 
            .O(n45941));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i30420_3_lut.LUT_INIT = 16'h2b2b;
    SB_LUT4 div_11_i1712_3_lut_3_lut (.I0(n2558), .I1(n6967), .I2(n2547), 
            .I3(GND_net), .O(n2631));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1712_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i1_4_lut_adj_1456 (.I0(n45941), .I1(n22412), .I2(n96), .I3(n40894), 
            .O(n806));
    defparam i1_4_lut_adj_1456.LUT_INIT = 16'hefce;
    SB_LUT4 i20205_3_lut (.I0(n784), .I1(n98), .I2(n4_adj_3993), .I3(GND_net), 
            .O(n6_adj_3989));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i20205_3_lut.LUT_INIT = 16'he8e8;
    SB_CARRY displacement_23__I_0_add_2_15 (.CI(n34252), .I0(displacement_23__N_93[13]), 
            .I1(n12_adj_3977), .CO(n34253));
    SB_LUT4 displacement_23__I_0_add_2_14_lut (.I0(GND_net), .I1(displacement_23__N_93[12]), 
            .I2(n13_adj_3976), .I3(n34251), .O(displacement_23__N_1[12])) /* synthesis syn_instantiated=1 */ ;
    defparam displacement_23__I_0_add_2_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3002_11 (.CI(n34932), .I0(n2545), .I1(n91), .CO(n34933));
    SB_CARRY displacement_23__I_0_add_2_14 (.CI(n34251), .I0(displacement_23__N_93[12]), 
            .I1(n13_adj_3976), .CO(n34252));
    SB_LUT4 displacement_23__I_0_add_2_13_lut (.I0(GND_net), .I1(displacement_23__N_93[11]), 
            .I2(n14_adj_3975), .I3(n34250), .O(displacement_23__N_1[11])) /* synthesis syn_instantiated=1 */ ;
    defparam displacement_23__I_0_add_2_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3002_10_lut (.I0(GND_net), .I1(n2546), .I2(n92), .I3(n34931), 
            .O(n6966)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3002_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY displacement_23__I_0_add_2_13 (.CI(n34250), .I0(displacement_23__N_93[11]), 
            .I1(n14_adj_3975), .CO(n34251));
    SB_LUT4 displacement_23__I_0_add_2_12_lut (.I0(GND_net), .I1(displacement_23__N_93[10]), 
            .I2(n15_adj_3974), .I3(n34249), .O(displacement_23__N_1[10])) /* synthesis syn_instantiated=1 */ ;
    defparam displacement_23__I_0_add_2_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3002_10 (.CI(n34931), .I0(n2546), .I1(n92), .CO(n34932));
    SB_CARRY displacement_23__I_0_add_2_12 (.CI(n34249), .I0(displacement_23__N_93[10]), 
            .I1(n15_adj_3974), .CO(n34250));
    SB_LUT4 add_3002_9_lut (.I0(GND_net), .I1(n2547), .I2(n93), .I3(n34930), 
            .O(n6967)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3002_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3002_9 (.CI(n34930), .I0(n2547), .I1(n93), .CO(n34931));
    SB_LUT4 add_3002_8_lut (.I0(GND_net), .I1(n2548), .I2(n94), .I3(n34929), 
            .O(n6968)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3002_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 displacement_23__I_0_add_2_11_lut (.I0(GND_net), .I1(displacement_23__N_93[9]), 
            .I2(n16_adj_3973), .I3(n34248), .O(displacement_23__N_1[9])) /* synthesis syn_instantiated=1 */ ;
    defparam displacement_23__I_0_add_2_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3002_8 (.CI(n34929), .I0(n2548), .I1(n94), .CO(n34930));
    SB_LUT4 add_3002_7_lut (.I0(GND_net), .I1(n2549), .I2(n95), .I3(n34928), 
            .O(n6969)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3002_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3002_7 (.CI(n34928), .I0(n2549), .I1(n95), .CO(n34929));
    SB_LUT4 add_3002_6_lut (.I0(GND_net), .I1(n2550), .I2(n96), .I3(n34927), 
            .O(n6970)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3002_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3002_6 (.CI(n34927), .I0(n2550), .I1(n96), .CO(n34928));
    SB_LUT4 add_3002_5_lut (.I0(GND_net), .I1(n2551), .I2(n97), .I3(n34926), 
            .O(n6971)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3002_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3002_5 (.CI(n34926), .I0(n2551), .I1(n97), .CO(n34927));
    SB_LUT4 add_3002_4_lut (.I0(GND_net), .I1(n2552), .I2(n98), .I3(n34925), 
            .O(n6972)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3002_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3002_4 (.CI(n34925), .I0(n2552), .I1(n98), .CO(n34926));
    SB_LUT4 add_3002_3_lut (.I0(GND_net), .I1(n2553), .I2(n99), .I3(n34924), 
            .O(n6973)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3002_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3002_3 (.CI(n34924), .I0(n2553), .I1(n99), .CO(n34925));
    SB_LUT4 add_3002_2_lut (.I0(GND_net), .I1(n388), .I2(n558), .I3(VCC_net), 
            .O(n6974)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3002_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3002_2 (.CI(VCC_net), .I0(n388), .I1(n558), .CO(n34924));
    SB_LUT4 add_3001_21_lut (.I0(GND_net), .I1(n2447), .I2(n81), .I3(n34923), 
            .O(n6932)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3001_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3001_20_lut (.I0(GND_net), .I1(n2448), .I2(n82), .I3(n34922), 
            .O(n6933)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3001_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3001_20 (.CI(n34922), .I0(n2448), .I1(n82), .CO(n34923));
    SB_LUT4 add_3001_19_lut (.I0(GND_net), .I1(n2449), .I2(n83), .I3(n34921), 
            .O(n6934)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3001_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3001_19 (.CI(n34921), .I0(n2449), .I1(n83), .CO(n34922));
    SB_IO PIN_19_pad (.PACKAGE_PIN(PIN_19), .OUTPUT_ENABLE(VCC_net), .D_IN_0(PIN_19_c_0)) /* synthesis IO_FF_IN=TRUE */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam PIN_19_pad.PIN_TYPE = 6'b000001;
    defparam PIN_19_pad.PULLUP = 1'b0;
    defparam PIN_19_pad.NEG_TRIGGER = 1'b0;
    defparam PIN_19_pad.IO_STANDARD = "SB_LVCMOS";
    SB_CARRY displacement_23__I_0_add_2_11 (.CI(n34248), .I0(displacement_23__N_93[9]), 
            .I1(n16_adj_3973), .CO(n34249));
    SB_LUT4 div_11_i459_4_lut (.I0(n648), .I1(n4), .I2(n671), .I3(n98), 
            .O(n783));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i459_4_lut.LUT_INIT = 16'ha9a6;
    SB_LUT4 add_3001_18_lut (.I0(GND_net), .I1(n2450), .I2(n84), .I3(n34920), 
            .O(n6935)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3001_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3001_18 (.CI(n34920), .I0(n2450), .I1(n84), .CO(n34921));
    SB_LUT4 add_3001_17_lut (.I0(GND_net), .I1(n2451), .I2(n85), .I3(n34919), 
            .O(n6936)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3001_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3001_17 (.CI(n34919), .I0(n2451), .I1(n85), .CO(n34920));
    SB_LUT4 add_3001_16_lut (.I0(GND_net), .I1(n2452), .I2(n86), .I3(n34918), 
            .O(n6937)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3001_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3001_16 (.CI(n34918), .I0(n2452), .I1(n86), .CO(n34919));
    SB_LUT4 add_3001_15_lut (.I0(GND_net), .I1(n2453), .I2(n87), .I3(n34917), 
            .O(n6938)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3001_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3001_15 (.CI(n34917), .I0(n2453), .I1(n87), .CO(n34918));
    SB_LUT4 add_3001_14_lut (.I0(GND_net), .I1(n2454), .I2(n88), .I3(n34916), 
            .O(n6939)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3001_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_11_i1718_3_lut_3_lut (.I0(n2558), .I1(n6973), .I2(n2553), 
            .I3(GND_net), .O(n2637));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1718_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_CARRY add_3001_14 (.CI(n34916), .I0(n2454), .I1(n88), .CO(n34917));
    SB_LUT4 add_3001_13_lut (.I0(GND_net), .I1(n2455), .I2(n89), .I3(n34915), 
            .O(n6940)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3001_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3001_13 (.CI(n34915), .I0(n2455), .I1(n89), .CO(n34916));
    SB_LUT4 add_3001_12_lut (.I0(GND_net), .I1(n2456), .I2(n90), .I3(n34914), 
            .O(n6941)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3001_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 displacement_23__I_0_add_2_10_lut (.I0(GND_net), .I1(displacement_23__N_93[8]), 
            .I2(n17_adj_3972), .I3(n34247), .O(displacement_23__N_1[8])) /* synthesis syn_instantiated=1 */ ;
    defparam displacement_23__I_0_add_2_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY displacement_23__I_0_add_2_10 (.CI(n34247), .I0(displacement_23__N_93[8]), 
            .I1(n17_adj_3972), .CO(n34248));
    SB_CARRY add_3001_12 (.CI(n34914), .I0(n2456), .I1(n90), .CO(n34915));
    SB_LUT4 add_3001_11_lut (.I0(GND_net), .I1(n2457), .I2(n91), .I3(n34913), 
            .O(n6942)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3001_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3001_11 (.CI(n34913), .I0(n2457), .I1(n91), .CO(n34914));
    SB_LUT4 displacement_23__I_0_add_2_9_lut (.I0(GND_net), .I1(displacement_23__N_93[7]), 
            .I2(n18_adj_3971), .I3(n34246), .O(displacement_23__N_1[7])) /* synthesis syn_instantiated=1 */ ;
    defparam displacement_23__I_0_add_2_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3001_10_lut (.I0(GND_net), .I1(n2458), .I2(n92), .I3(n34912), 
            .O(n6943)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3001_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3001_10 (.CI(n34912), .I0(n2458), .I1(n92), .CO(n34913));
    SB_LUT4 add_3001_9_lut (.I0(GND_net), .I1(n2459), .I2(n93), .I3(n34911), 
            .O(n6944)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3001_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3001_9 (.CI(n34911), .I0(n2459), .I1(n93), .CO(n34912));
    SB_LUT4 add_3001_8_lut (.I0(GND_net), .I1(n2460), .I2(n94), .I3(n34910), 
            .O(n6945)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3001_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3001_8 (.CI(n34910), .I0(n2460), .I1(n94), .CO(n34911));
    SB_LUT4 add_3001_7_lut (.I0(GND_net), .I1(n2461), .I2(n95), .I3(n34909), 
            .O(n6946)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3001_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3001_7 (.CI(n34909), .I0(n2461), .I1(n95), .CO(n34910));
    SB_LUT4 div_11_LessThan_570_i40_4_lut (.I0(n373), .I1(n99), .I2(n918), 
            .I3(n558), .O(n40));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_570_i40_4_lut.LUT_INIT = 16'h0317;
    SB_LUT4 add_3001_6_lut (.I0(GND_net), .I1(n2462), .I2(n96), .I3(n34908), 
            .O(n6947)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3001_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3001_6 (.CI(n34908), .I0(n2462), .I1(n96), .CO(n34909));
    SB_LUT4 add_3001_5_lut (.I0(GND_net), .I1(n2463), .I2(n97), .I3(n34907), 
            .O(n6948)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3001_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3001_5 (.CI(n34907), .I0(n2463), .I1(n97), .CO(n34908));
    SB_LUT4 add_3001_4_lut (.I0(GND_net), .I1(n2464), .I2(n98), .I3(n34906), 
            .O(n6949)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3001_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3001_4 (.CI(n34906), .I0(n2464), .I1(n98), .CO(n34907));
    SB_LUT4 add_3001_3_lut (.I0(GND_net), .I1(n2465), .I2(n99), .I3(n34905), 
            .O(n6950)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3001_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3001_3 (.CI(n34905), .I0(n2465), .I1(n99), .CO(n34906));
    SB_LUT4 add_3001_2_lut (.I0(GND_net), .I1(n387_adj_4001), .I2(n558), 
            .I3(VCC_net), .O(n6951)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3001_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3001_2 (.CI(VCC_net), .I0(n387_adj_4001), .I1(n558), 
            .CO(n34905));
    SB_LUT4 add_3000_20_lut (.I0(GND_net), .I1(n2357), .I2(n82), .I3(n34904), 
            .O(n6911)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3000_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3000_19_lut (.I0(GND_net), .I1(n2358), .I2(n83), .I3(n34903), 
            .O(n6912)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3000_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3000_19 (.CI(n34903), .I0(n2358), .I1(n83), .CO(n34904));
    SB_LUT4 add_3000_18_lut (.I0(GND_net), .I1(n2359), .I2(n84), .I3(n34902), 
            .O(n6913)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3000_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3000_18 (.CI(n34902), .I0(n2359), .I1(n84), .CO(n34903));
    SB_LUT4 add_3000_17_lut (.I0(GND_net), .I1(n2360), .I2(n85), .I3(n34901), 
            .O(n6914)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3000_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_11_LessThan_570_i44_3_lut (.I0(n42_adj_4079), .I1(n96), 
            .I2(n45), .I3(GND_net), .O(n44_adj_4080));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_570_i44_3_lut.LUT_INIT = 16'h3a3a;
    SB_CARRY add_3000_17 (.CI(n34901), .I0(n2360), .I1(n85), .CO(n34902));
    SB_LUT4 add_3000_16_lut (.I0(GND_net), .I1(n2361), .I2(n86), .I3(n34900), 
            .O(n6915)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3000_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i10669_3_lut (.I0(\data_in[1] [5]), .I1(\data_in[2] [5]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n24087));   // verilog/coms.v(126[12] 289[6])
    defparam i10669_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY displacement_23__I_0_add_2_9 (.CI(n34246), .I0(displacement_23__N_93[7]), 
            .I1(n18_adj_3971), .CO(n34247));
    SB_CARRY add_3000_16 (.CI(n34900), .I0(n2361), .I1(n86), .CO(n34901));
    SB_LUT4 add_3000_15_lut (.I0(GND_net), .I1(n2362), .I2(n87), .I3(n34899), 
            .O(n6916)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3000_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3000_15 (.CI(n34899), .I0(n2362), .I1(n87), .CO(n34900));
    SB_LUT4 add_3000_14_lut (.I0(GND_net), .I1(n2363), .I2(n88), .I3(n34898), 
            .O(n6917)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3000_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3000_14 (.CI(n34898), .I0(n2363), .I1(n88), .CO(n34899));
    SB_LUT4 add_3000_13_lut (.I0(GND_net), .I1(n2364), .I2(n89), .I3(n34897), 
            .O(n6918)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3000_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3000_13 (.CI(n34897), .I0(n2364), .I1(n89), .CO(n34898));
    SB_LUT4 i29985_4_lut (.I0(n44_adj_4080), .I1(n40), .I2(n45), .I3(n44470), 
            .O(n45506));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i29985_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 add_3000_12_lut (.I0(GND_net), .I1(n2365), .I2(n90), .I3(n34896), 
            .O(n6919)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3000_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3000_12 (.CI(n34896), .I0(n2365), .I1(n90), .CO(n34897));
    SB_LUT4 add_3000_11_lut (.I0(GND_net), .I1(n2366), .I2(n91), .I3(n34895), 
            .O(n6920)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3000_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3000_11 (.CI(n34895), .I0(n2366), .I1(n91), .CO(n34896));
    SB_LUT4 add_3000_10_lut (.I0(GND_net), .I1(n2367), .I2(n92), .I3(n34894), 
            .O(n6921)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3000_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3000_10 (.CI(n34894), .I0(n2367), .I1(n92), .CO(n34895));
    SB_LUT4 i1_4_lut_adj_1457 (.I0(n45506), .I1(n22415), .I2(n95), .I3(n914), 
            .O(n938));
    defparam i1_4_lut_adj_1457.LUT_INIT = 16'hceef;
    SB_LUT4 add_3000_9_lut (.I0(GND_net), .I1(n2368), .I2(n93), .I3(n34893), 
            .O(n6922)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3000_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3000_9 (.CI(n34893), .I0(n2368), .I1(n93), .CO(n34894));
    SB_LUT4 i10670_3_lut (.I0(\data_in[1] [4]), .I1(\data_in[2] [4]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n24088));   // verilog/coms.v(126[12] 289[6])
    defparam i10670_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_11_i1717_3_lut_3_lut (.I0(n2558), .I1(n6972), .I2(n2552), 
            .I3(GND_net), .O(n2636));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1717_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_11_i548_4_lut (.I0(n783), .I1(n6_adj_3989), .I2(n806), 
            .I3(n97), .O(n915));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i548_4_lut.LUT_INIT = 16'ha9a6;
    SB_LUT4 div_11_i1716_3_lut_3_lut (.I0(n2558), .I1(n6971), .I2(n2551), 
            .I3(GND_net), .O(n2635));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1716_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_11_i1714_3_lut_3_lut (.I0(n2558), .I1(n6969), .I2(n2549), 
            .I3(GND_net), .O(n2633));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1714_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 add_3000_8_lut (.I0(GND_net), .I1(n2369), .I2(n94), .I3(n34892), 
            .O(n6923)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3000_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3000_8 (.CI(n34892), .I0(n2369), .I1(n94), .CO(n34893));
    SB_LUT4 add_3000_7_lut (.I0(GND_net), .I1(n2370), .I2(n95), .I3(n34891), 
            .O(n6924)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3000_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3000_7 (.CI(n34891), .I0(n2370), .I1(n95), .CO(n34892));
    SB_LUT4 div_11_i1713_3_lut_3_lut (.I0(n2558), .I1(n6968), .I2(n2548), 
            .I3(GND_net), .O(n2632));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1713_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_11_i1769_3_lut_3_lut (.I0(n2642), .I1(n6992), .I2(n2633), 
            .I3(GND_net), .O(n2714));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1769_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 add_3000_6_lut (.I0(GND_net), .I1(n2371), .I2(n96), .I3(n34890), 
            .O(n6925)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3000_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3000_6 (.CI(n34890), .I0(n2371), .I1(n96), .CO(n34891));
    SB_LUT4 add_3000_5_lut (.I0(GND_net), .I1(n2372), .I2(n97), .I3(n34889), 
            .O(n6926)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3000_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3000_5 (.CI(n34889), .I0(n2372), .I1(n97), .CO(n34890));
    SB_LUT4 div_11_i1754_3_lut_3_lut (.I0(n2642), .I1(n6977), .I2(n2618), 
            .I3(GND_net), .O(n2699));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1754_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 add_3000_4_lut (.I0(GND_net), .I1(n2373), .I2(n98), .I3(n34888), 
            .O(n6927)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3000_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3000_4 (.CI(n34888), .I0(n2373), .I1(n98), .CO(n34889));
    SB_LUT4 displacement_23__I_0_add_2_8_lut (.I0(GND_net), .I1(displacement_23__N_93[6]), 
            .I2(n19_adj_3970), .I3(n34245), .O(displacement_23__N_1[6])) /* synthesis syn_instantiated=1 */ ;
    defparam displacement_23__I_0_add_2_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3000_3_lut (.I0(GND_net), .I1(n2374), .I2(n99), .I3(n34887), 
            .O(n6928)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3000_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_11_LessThan_657_i38_4_lut (.I0(n374), .I1(n99), .I2(n1048), 
            .I3(n558), .O(n38));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_657_i38_4_lut.LUT_INIT = 16'h0317;
    SB_LUT4 div_11_LessThan_657_i42_3_lut (.I0(n40_adj_4081), .I1(n96), 
            .I2(n43), .I3(GND_net), .O(n42_adj_4082));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_657_i42_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i30369_4_lut (.I0(n42_adj_4082), .I1(n38), .I2(n43), .I3(n44464), 
            .O(n45890));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i30369_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i30370_3_lut (.I0(n45890), .I1(n95), .I2(n1044), .I3(GND_net), 
            .O(n45891));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i30370_3_lut.LUT_INIT = 16'h2b2b;
    SB_LUT4 i1_4_lut_adj_1458 (.I0(n45891), .I1(n22418), .I2(n94), .I3(n1043), 
            .O(n1067));
    defparam i1_4_lut_adj_1458.LUT_INIT = 16'hceef;
    SB_LUT4 div_11_i635_3_lut (.I0(n915), .I1(n5823), .I2(n938), .I3(GND_net), 
            .O(n1044));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i635_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_11_i1756_3_lut_3_lut (.I0(n2642), .I1(n6979), .I2(n2620), 
            .I3(GND_net), .O(n2701));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1756_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_CARRY displacement_23__I_0_add_2_8 (.CI(n34245), .I0(displacement_23__N_93[6]), 
            .I1(n19_adj_3970), .CO(n34246));
    SB_LUT4 div_11_LessThan_742_i36_4_lut (.I0(n375), .I1(n99), .I2(n1175), 
            .I3(n558), .O(n36));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_742_i36_4_lut.LUT_INIT = 16'h0317;
    SB_LUT4 div_11_i1755_3_lut_3_lut (.I0(n2642), .I1(n6978), .I2(n2619), 
            .I3(GND_net), .O(n2700));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1755_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_11_i1757_3_lut_3_lut (.I0(n2642), .I1(n6980), .I2(n2621), 
            .I3(GND_net), .O(n2702));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1757_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_11_i1758_3_lut_3_lut (.I0(n2642), .I1(n6981), .I2(n2622), 
            .I3(GND_net), .O(n2703));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1758_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_11_LessThan_742_i40_3_lut (.I0(n38_adj_4083), .I1(n96), 
            .I2(n41), .I3(GND_net), .O(n40_adj_4084));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_742_i40_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 div_11_i1761_3_lut_3_lut (.I0(n2642), .I1(n6984), .I2(n2625), 
            .I3(GND_net), .O(n2706));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1761_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i30562_4_lut (.I0(n40_adj_4084), .I1(n36), .I2(n41), .I3(n44430), 
            .O(n46083));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i30562_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i30563_3_lut (.I0(n46083), .I1(n95), .I2(n1171), .I3(GND_net), 
            .O(n46084));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i30563_3_lut.LUT_INIT = 16'h2b2b;
    SB_LUT4 div_11_i1762_3_lut_3_lut (.I0(n2642), .I1(n6985), .I2(n2626), 
            .I3(GND_net), .O(n2707));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1762_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i30510_3_lut (.I0(n46084), .I1(n94), .I2(n1170), .I3(GND_net), 
            .O(n46031));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i30510_3_lut.LUT_INIT = 16'h2b2b;
    SB_LUT4 i1_4_lut_adj_1459 (.I0(n46031), .I1(n22421), .I2(n93), .I3(n1169), 
            .O(n1193));
    defparam i1_4_lut_adj_1459.LUT_INIT = 16'hceef;
    SB_LUT4 div_11_i1759_3_lut_3_lut (.I0(n2642), .I1(n6982), .I2(n2623), 
            .I3(GND_net), .O(n2704));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1759_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_11_i1760_3_lut_3_lut (.I0(n2642), .I1(n6983), .I2(n2624), 
            .I3(GND_net), .O(n2705));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1760_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_11_i1775_3_lut_3_lut (.I0(n2642), .I1(n6998), .I2(n389), 
            .I3(GND_net), .O(n2720));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1775_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 displacement_23__I_0_add_2_7_lut (.I0(GND_net), .I1(displacement_23__N_93[5]), 
            .I2(n20_adj_3969), .I3(n34244), .O(displacement_23__N_1[5])) /* synthesis syn_instantiated=1 */ ;
    defparam displacement_23__I_0_add_2_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i10671_3_lut (.I0(\data_in[1] [3]), .I1(\data_in[2] [3]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n24089));   // verilog/coms.v(126[12] 289[6])
    defparam i10671_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_11_i720_3_lut (.I0(n1044), .I1(n6215), .I2(n1067), .I3(GND_net), 
            .O(n1170));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i720_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY add_3000_3 (.CI(n34887), .I0(n2374), .I1(n99), .CO(n34888));
    SB_LUT4 div_11_i1764_3_lut_3_lut (.I0(n2642), .I1(n6987), .I2(n2628), 
            .I3(GND_net), .O(n2709));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1764_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 add_3000_2_lut (.I0(GND_net), .I1(n386), .I2(n558), .I3(VCC_net), 
            .O(n6929)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3000_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3000_2 (.CI(VCC_net), .I0(n386), .I1(n558), .CO(n34887));
    SB_LUT4 div_11_i1765_3_lut_3_lut (.I0(n2642), .I1(n6988), .I2(n2629), 
            .I3(GND_net), .O(n2710));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1765_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_11_i1766_3_lut_3_lut (.I0(n2642), .I1(n6989), .I2(n2630), 
            .I3(GND_net), .O(n2711));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1766_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_11_i1767_3_lut_3_lut (.I0(n2642), .I1(n6990), .I2(n2631), 
            .I3(GND_net), .O(n2712));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1767_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_11_LessThan_742_i38_3_lut_3_lut (.I0(n1173), .I1(n97), .I2(n98), 
            .I3(GND_net), .O(n38_adj_4083));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_742_i38_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_CARRY displacement_23__I_0_add_2_7 (.CI(n34244), .I0(displacement_23__N_93[5]), 
            .I1(n20_adj_3969), .CO(n34245));
    SB_LUT4 displacement_23__I_0_add_2_6_lut (.I0(GND_net), .I1(displacement_23__N_93[4]), 
            .I2(n21_adj_3968), .I3(n34243), .O(displacement_23__N_1[4])) /* synthesis syn_instantiated=1 */ ;
    defparam displacement_23__I_0_add_2_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY displacement_23__I_0_add_2_6 (.CI(n34243), .I0(displacement_23__N_93[4]), 
            .I1(n21_adj_3968), .CO(n34244));
    SB_LUT4 displacement_23__I_0_add_2_5_lut (.I0(GND_net), .I1(displacement_23__N_93[3]), 
            .I2(n22_adj_3967), .I3(n34242), .O(displacement_23__N_1[3])) /* synthesis syn_instantiated=1 */ ;
    defparam displacement_23__I_0_add_2_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_11_i1773_3_lut_3_lut (.I0(n2642), .I1(n6996), .I2(n2637), 
            .I3(GND_net), .O(n2718));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1773_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_CARRY displacement_23__I_0_add_2_5 (.CI(n34242), .I0(displacement_23__N_93[3]), 
            .I1(n22_adj_3967), .CO(n34243));
    SB_LUT4 div_11_i1774_3_lut_3_lut (.I0(n2642), .I1(n6997), .I2(n2638), 
            .I3(GND_net), .O(n2719));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1774_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_11_LessThan_825_i34_4_lut (.I0(n376), .I1(n99), .I2(n1299), 
            .I3(n558), .O(n34));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_825_i34_4_lut.LUT_INIT = 16'h0317;
    SB_LUT4 i30365_3_lut (.I0(n34), .I1(n95), .I2(n41_adj_4087), .I3(GND_net), 
            .O(n45886));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i30365_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i30366_3_lut (.I0(n45886), .I1(n94), .I2(n43_adj_4088), .I3(GND_net), 
            .O(n45887));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i30366_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 div_11_i1771_3_lut_3_lut (.I0(n2642), .I1(n6994), .I2(n2635), 
            .I3(GND_net), .O(n2716));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1771_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 displacement_23__I_0_add_2_4_lut (.I0(GND_net), .I1(displacement_23__N_93[2]), 
            .I2(n23_adj_3966), .I3(n34241), .O(displacement_23__N_1[2])) /* synthesis syn_instantiated=1 */ ;
    defparam displacement_23__I_0_add_2_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY displacement_23__I_0_add_2_4 (.CI(n34241), .I0(displacement_23__N_93[2]), 
            .I1(n23_adj_3966), .CO(n34242));
    SB_LUT4 i29570_4_lut (.I0(n43_adj_4088), .I1(n41_adj_4087), .I2(n39), 
            .I3(n44422), .O(n45091));
    defparam i29570_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 displacement_23__I_0_add_2_3_lut (.I0(GND_net), .I1(displacement_23__N_93[1]), 
            .I2(n24_adj_3965), .I3(n34240), .O(displacement_23__N_1[1])) /* synthesis syn_instantiated=1 */ ;
    defparam displacement_23__I_0_add_2_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_11_i1763_3_lut_3_lut (.I0(n2642), .I1(n6986), .I2(n2627), 
            .I3(GND_net), .O(n2708));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1763_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_CARRY displacement_23__I_0_add_2_3 (.CI(n34240), .I0(displacement_23__N_93[1]), 
            .I1(n24_adj_3965), .CO(n34241));
    SB_LUT4 displacement_23__I_0_add_2_2_lut (.I0(GND_net), .I1(displacement_23__N_93[0]), 
            .I2(n25_adj_3964), .I3(VCC_net), .O(displacement_23__N_1[0])) /* synthesis syn_instantiated=1 */ ;
    defparam displacement_23__I_0_add_2_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY displacement_23__I_0_add_2_2 (.CI(VCC_net), .I0(displacement_23__N_93[0]), 
            .I1(n25_adj_3964), .CO(n34240));
    SB_LUT4 div_11_LessThan_825_i38_3_lut (.I0(n36_adj_4085), .I1(n96), 
            .I2(n39), .I3(GND_net), .O(n38_adj_4086));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_825_i38_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i30206_3_lut (.I0(n45887), .I1(n93), .I2(n45_adj_4090), .I3(GND_net), 
            .O(n44_adj_4089));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i30206_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i29989_4_lut (.I0(n44_adj_4089), .I1(n38_adj_4086), .I2(n45_adj_4090), 
            .I3(n45091), .O(n45510));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i29989_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i28911_3_lut_4_lut (.I0(n1173), .I1(n97), .I2(n98), .I3(n1174), 
            .O(n44430));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i28911_3_lut_4_lut.LUT_INIT = 16'hf99f;
    SB_LUT4 div_11_LessThan_657_i40_3_lut_3_lut (.I0(n1046), .I1(n97), .I2(n98), 
            .I3(GND_net), .O(n40_adj_4081));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_657_i40_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 div_11_i1772_3_lut_3_lut (.I0(n2642), .I1(n6995), .I2(n2636), 
            .I3(GND_net), .O(n2717));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1772_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i1_4_lut_adj_1460 (.I0(n45510), .I1(n22424), .I2(n92), .I3(n1292), 
            .O(n1316));
    defparam i1_4_lut_adj_1460.LUT_INIT = 16'hceef;
    SB_LUT4 div_11_i803_3_lut (.I0(n1170), .I1(n6576), .I2(n1193), .I3(GND_net), 
            .O(n1293));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i803_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_11_i1768_3_lut_3_lut (.I0(n2642), .I1(n6991), .I2(n2632), 
            .I3(GND_net), .O(n2713));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1768_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_11_i1770_3_lut_3_lut (.I0(n2642), .I1(n6993), .I2(n2634), 
            .I3(GND_net), .O(n2715));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1770_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_11_LessThan_906_i32_4_lut (.I0(n377), .I1(n99), .I2(n1420), 
            .I3(n558), .O(n32));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_906_i32_4_lut.LUT_INIT = 16'h0317;
    SB_LUT4 i30363_3_lut (.I0(n32), .I1(n95), .I2(n39_adj_4092), .I3(GND_net), 
            .O(n45884));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i30363_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i30364_3_lut (.I0(n45884), .I1(n94), .I2(n41_adj_4093), .I3(GND_net), 
            .O(n45885));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i30364_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i29538_4_lut (.I0(n41_adj_4093), .I1(n39_adj_4092), .I2(n37), 
            .I3(n44407), .O(n45059));
    defparam i29538_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i29991_3_lut (.I0(n34_adj_4091), .I1(n96), .I2(n37), .I3(GND_net), 
            .O(n45512));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i29991_3_lut.LUT_INIT = 16'h3a3a;
    GND i1 (.Y(GND_net));
    SB_LUT4 i30208_3_lut (.I0(n45885), .I1(n93), .I2(n43_adj_4094), .I3(GND_net), 
            .O(n45729));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i30208_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i30361_4_lut (.I0(n45729), .I1(n45512), .I2(n43_adj_4094), 
            .I3(n45059), .O(n45882));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i30361_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i30362_3_lut (.I0(n45882), .I1(n92), .I2(n1413), .I3(GND_net), 
            .O(n45883));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i30362_3_lut.LUT_INIT = 16'h2b2b;
    SB_LUT4 i1_4_lut_adj_1461 (.I0(n45883), .I1(n22427), .I2(n91), .I3(n1412), 
            .O(n1436));
    defparam i1_4_lut_adj_1461.LUT_INIT = 16'hceef;
    SB_LUT4 div_11_i884_3_lut (.I0(n1293), .I1(n6647), .I2(n1316), .I3(GND_net), 
            .O(n1413));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i884_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_11_LessThan_985_i31_2_lut (.I0(n1537), .I1(n98), .I2(GND_net), 
            .I3(GND_net), .O(n31));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_985_i31_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i28872_4_lut (.I0(n37_adj_4098), .I1(n35), .I2(n33), .I3(n31), 
            .O(n44391));
    defparam i28872_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 div_11_LessThan_985_i42_3_lut (.I0(n34_adj_4097), .I1(n91), 
            .I2(n45_adj_4103), .I3(GND_net), .O(n42_adj_4101));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_985_i42_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 div_11_LessThan_985_i30_4_lut (.I0(n378), .I1(n99), .I2(n1538), 
            .I3(n558), .O(n30_adj_4095));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_985_i30_4_lut.LUT_INIT = 16'h0317;
    SB_LUT4 i30359_3_lut (.I0(n30_adj_4095), .I1(n95), .I2(n37_adj_4098), 
            .I3(GND_net), .O(n45880));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i30359_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i30360_3_lut (.I0(n45880), .I1(n94), .I2(n39_adj_4099), .I3(GND_net), 
            .O(n45881));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i30360_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i28866_4_lut (.I0(n43_adj_4102), .I1(n41_adj_4100), .I2(n39_adj_4099), 
            .I3(n44391), .O(n44385));
    defparam i28866_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i29993_4_lut (.I0(n42_adj_4101), .I1(n32_adj_4096), .I2(n45_adj_4103), 
            .I3(n44381), .O(n45514));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i29993_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i10672_3_lut (.I0(\data_in[1] [2]), .I1(\data_in[2] [2]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n24090));   // verilog/coms.v(126[12] 289[6])
    defparam i10672_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i30212_3_lut (.I0(n45881), .I1(n93), .I2(n41_adj_4100), .I3(GND_net), 
            .O(n45733));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i30212_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i10707_3_lut (.I0(Kd[5]), .I1(\data_in_frame[4] [5]), .I2(n23399), 
            .I3(GND_net), .O(n24125));   // verilog/coms.v(126[12] 289[6])
    defparam i10707_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i30423_4_lut (.I0(n45733), .I1(n45514), .I2(n45_adj_4103), 
            .I3(n44385), .O(n45944));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i30423_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i1_4_lut_adj_1462 (.I0(n45944), .I1(n22430), .I2(n90), .I3(n1529), 
            .O(n1553));
    defparam i1_4_lut_adj_1462.LUT_INIT = 16'hceef;
    SB_LUT4 div_11_i963_3_lut (.I0(n1413), .I1(n6687), .I2(n1436), .I3(GND_net), 
            .O(n1530));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i963_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_11_LessThan_1062_i29_2_lut (.I0(n1652), .I1(n98), .I2(GND_net), 
            .I3(GND_net), .O(n29));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1062_i29_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i28848_4_lut (.I0(n35_adj_4109), .I1(n33_adj_4108), .I2(n31_adj_4106), 
            .I3(n29), .O(n44367));
    defparam i28848_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i28944_3_lut_4_lut (.I0(n1046), .I1(n97), .I2(n98), .I3(n1047), 
            .O(n44464));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i28944_3_lut_4_lut.LUT_INIT = 16'hf99f;
    SB_LUT4 div_11_LessThan_570_i42_3_lut_3_lut (.I0(n916), .I1(n97), .I2(n98), 
            .I3(GND_net), .O(n42_adj_4079));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_570_i42_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 div_11_LessThan_1062_i40_3_lut (.I0(n32_adj_4107), .I1(n91), 
            .I2(n43_adj_4114), .I3(GND_net), .O(n40_adj_4112));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1062_i40_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 div_11_LessThan_1062_i28_4_lut (.I0(n379), .I1(n99), .I2(n1653), 
            .I3(n558), .O(n28_adj_4104));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1062_i28_4_lut.LUT_INIT = 16'h0317;
    SB_LUT4 i30357_3_lut (.I0(n28_adj_4104), .I1(n95), .I2(n35_adj_4109), 
            .I3(GND_net), .O(n45878));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i30357_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i30358_3_lut (.I0(n45878), .I1(n94), .I2(n37_adj_4110), .I3(GND_net), 
            .O(n45879));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i30358_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i28829_4_lut (.I0(n41_adj_4113), .I1(n39_adj_4111), .I2(n37_adj_4110), 
            .I3(n44367), .O(n44348));
    defparam i28829_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i28950_3_lut_4_lut (.I0(n916), .I1(n97), .I2(n98), .I3(n917), 
            .O(n44470));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i28950_3_lut_4_lut.LUT_INIT = 16'hf99f;
    SB_LUT4 i30355_4_lut (.I0(n40_adj_4112), .I1(n30_adj_4105), .I2(n43_adj_4114), 
            .I3(n44346), .O(n45876));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i30355_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i10708_3_lut (.I0(Kd[4]), .I1(\data_in_frame[4] [4]), .I2(n23399), 
            .I3(GND_net), .O(n24126));   // verilog/coms.v(126[12] 289[6])
    defparam i10708_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i30214_3_lut (.I0(n45879), .I1(n93), .I2(n39_adj_4111), .I3(GND_net), 
            .O(n45735));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i30214_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i30560_4_lut (.I0(n45735), .I1(n45876), .I2(n43_adj_4114), 
            .I3(n44348), .O(n46081));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i30560_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i10709_3_lut (.I0(Kd[3]), .I1(\data_in_frame[4] [3]), .I2(n23399), 
            .I3(GND_net), .O(n24127));   // verilog/coms.v(126[12] 289[6])
    defparam i10709_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i30561_3_lut (.I0(n46081), .I1(n90), .I2(n1644), .I3(GND_net), 
            .O(n46082));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i30561_3_lut.LUT_INIT = 16'h2b2b;
    SB_LUT4 i10710_3_lut (.I0(Kd[2]), .I1(\data_in_frame[4] [2]), .I2(n23399), 
            .I3(GND_net), .O(n24128));   // verilog/coms.v(126[12] 289[6])
    defparam i10710_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_1463 (.I0(n46082), .I1(n22433), .I2(n89), .I3(n1643), 
            .O(n1667));
    defparam i1_4_lut_adj_1463.LUT_INIT = 16'hceef;
    SB_LUT4 i10711_3_lut (.I0(Kd[1]), .I1(\data_in_frame[4] [1]), .I2(n23399), 
            .I3(GND_net), .O(n24129));   // verilog/coms.v(126[12] 289[6])
    defparam i10711_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_11_i1040_3_lut (.I0(n1530), .I1(n6727), .I2(n1553), .I3(GND_net), 
            .O(n1644));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1040_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i10712_3_lut (.I0(Ki[7]), .I1(\data_in_frame[3] [7]), .I2(n23399), 
            .I3(GND_net), .O(n24130));   // verilog/coms.v(126[12] 289[6])
    defparam i10712_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10713_3_lut (.I0(Ki[6]), .I1(\data_in_frame[3] [6]), .I2(n23399), 
            .I3(GND_net), .O(n24131));   // verilog/coms.v(126[12] 289[6])
    defparam i10713_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_11_mux_5_i12_3_lut (.I0(gearBoxRatio[11]), .I1(n64), .I2(gearBoxRatio[23]), 
            .I3(GND_net), .O(n89));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_mux_5_i12_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 div_11_LessThan_1137_i27_2_lut (.I0(n1764), .I1(n98), .I2(GND_net), 
            .I3(GND_net), .O(n27));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1137_i27_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i10714_3_lut (.I0(Ki[5]), .I1(\data_in_frame[3] [5]), .I2(n23399), 
            .I3(GND_net), .O(n24132));   // verilog/coms.v(126[12] 289[6])
    defparam i10714_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i28807_4_lut (.I0(n33_adj_4120), .I1(n31_adj_4119), .I2(n29_adj_4117), 
            .I3(n27), .O(n44326));
    defparam i28807_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 div_11_LessThan_1137_i38_3_lut (.I0(n30_adj_4118), .I1(n91), 
            .I2(n41_adj_4125), .I3(GND_net), .O(n38_adj_4123));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1137_i38_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 div_11_LessThan_1137_i26_4_lut (.I0(n380), .I1(n99), .I2(n1765), 
            .I3(n558), .O(n26_adj_4115));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1137_i26_4_lut.LUT_INIT = 16'h0317;
    SB_LUT4 i30353_3_lut (.I0(n26_adj_4115), .I1(n95), .I2(n33_adj_4120), 
            .I3(GND_net), .O(n45874));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i30353_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i30354_3_lut (.I0(n45874), .I1(n94), .I2(n35_adj_4121), .I3(GND_net), 
            .O(n45875));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i30354_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i10645_4_lut (.I0(\data_out_frame[5] [2]), .I1(control_mode[2]), 
            .I2(n5019), .I3(n22338), .O(n24063));   // verilog/coms.v(126[12] 289[6])
    defparam i10645_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i28795_4_lut (.I0(n39_adj_4124), .I1(n37_adj_4122), .I2(n35_adj_4121), 
            .I3(n44326), .O(n44314));
    defparam i28795_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i30564_4_lut (.I0(n38_adj_4123), .I1(n28_adj_4116), .I2(n41_adj_4125), 
            .I3(n44308), .O(n46085));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i30564_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i30218_3_lut (.I0(n45875), .I1(n93), .I2(n37_adj_4122), .I3(GND_net), 
            .O(n45739));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i30218_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i30663_4_lut (.I0(n45739), .I1(n46085), .I2(n41_adj_4125), 
            .I3(n44314), .O(n46184));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i30663_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i30664_3_lut (.I0(n46184), .I1(n90), .I2(n1756), .I3(GND_net), 
            .O(n46185));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i30664_3_lut.LUT_INIT = 16'h2b2b;
    SB_LUT4 i10648_3_lut (.I0(\data_out_frame[0] [4]), .I1(n5019), .I2(n23458), 
            .I3(GND_net), .O(n24066));   // verilog/coms.v(126[12] 289[6])
    defparam i10648_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i30634_3_lut (.I0(n46185), .I1(n89), .I2(n1755), .I3(GND_net), 
            .O(n46155));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i30634_3_lut.LUT_INIT = 16'h2b2b;
    SB_LUT4 i1_4_lut_adj_1464 (.I0(n46155), .I1(n22436), .I2(n88), .I3(n1754), 
            .O(n1778));
    defparam i1_4_lut_adj_1464.LUT_INIT = 16'hceef;
    SB_LUT4 div_11_i1115_3_lut (.I0(n1644), .I1(n6740), .I2(n1667), .I3(GND_net), 
            .O(n1755));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1115_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i10649_3_lut (.I0(\data_out_frame[0] [3]), .I1(n5019), .I2(n23458), 
            .I3(GND_net), .O(n24067));   // verilog/coms.v(126[12] 289[6])
    defparam i10649_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_11_mux_5_i13_3_lut (.I0(gearBoxRatio[12]), .I1(n63), .I2(gearBoxRatio[23]), 
            .I3(GND_net), .O(n88));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_mux_5_i13_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 div_11_i1188_3_lut (.I0(n1755), .I1(n6781), .I2(n1778), .I3(GND_net), 
            .O(n1863));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1188_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i10650_3_lut (.I0(\data_out_frame[0] [2]), .I1(n5019), .I2(n23458), 
            .I3(GND_net), .O(n24068));   // verilog/coms.v(126[12] 289[6])
    defparam i10650_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_11_LessThan_1210_i45_2_lut (.I0(n1863), .I1(n88), .I2(GND_net), 
            .I3(GND_net), .O(n45_adj_4143));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1210_i45_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i1_2_lut_adj_1465 (.I0(n84), .I1(n22448), .I2(GND_net), .I3(GND_net), 
            .O(n22445));
    defparam i1_2_lut_adj_1465.LUT_INIT = 16'hdddd;
    SB_LUT4 i10651_3_lut (.I0(\data_in[3] [7]), .I1(rx_data[7]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n24069));   // verilog/coms.v(126[12] 289[6])
    defparam i10651_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_11_mux_5_i16_3_lut (.I0(gearBoxRatio[15]), .I1(n60), .I2(gearBoxRatio[23]), 
            .I3(GND_net), .O(n85));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_mux_5_i16_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 i10652_3_lut (.I0(\data_in[3] [6]), .I1(rx_data[6]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n24070));   // verilog/coms.v(126[12] 289[6])
    defparam i10652_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_11_mux_5_i15_3_lut (.I0(gearBoxRatio[14]), .I1(n61), .I2(gearBoxRatio[23]), 
            .I3(GND_net), .O(n86));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_mux_5_i15_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 i10653_3_lut (.I0(\data_in[3] [5]), .I1(rx_data[5]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n24071));   // verilog/coms.v(126[12] 289[6])
    defparam i10653_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_11_i1187_3_lut (.I0(n1754), .I1(n6780), .I2(n1778), .I3(GND_net), 
            .O(n1862));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1187_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i10654_3_lut (.I0(\data_in[3] [4]), .I1(rx_data[4]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n24072));   // verilog/coms.v(126[12] 289[6])
    defparam i10654_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_11_mux_5_i14_3_lut (.I0(gearBoxRatio[13]), .I1(n62), .I2(gearBoxRatio[23]), 
            .I3(GND_net), .O(n87));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_mux_5_i14_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 i10655_3_lut (.I0(\data_in[3] [3]), .I1(rx_data[3]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n24073));   // verilog/coms.v(126[12] 289[6])
    defparam i10655_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_adj_1466 (.I0(n86), .I1(n22442), .I2(GND_net), .I3(GND_net), 
            .O(n22439));
    defparam i1_2_lut_adj_1466.LUT_INIT = 16'hdddd;
    SB_LUT4 i10656_3_lut (.I0(\data_in[3] [2]), .I1(rx_data[2]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n24074));   // verilog/coms.v(126[12] 289[6])
    defparam i10656_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_11_LessThan_1210_i25_2_lut (.I0(n1873), .I1(n98), .I2(GND_net), 
            .I3(GND_net), .O(n25_adj_4127));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1210_i25_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i29006_3_lut_4_lut (.I0(pwm_count[3]), .I1(pwm[3]), .I2(pwm[2]), 
            .I3(pwm_count[2]), .O(n44526));   // verilog/motorControl.v(65[19:32])
    defparam i29006_3_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 i10657_3_lut (.I0(\data_in[3] [1]), .I1(rx_data[1]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n24075));   // verilog/coms.v(126[12] 289[6])
    defparam i10657_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10658_3_lut (.I0(\data_in[3] [0]), .I1(rx_data[0]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n24076));   // verilog/coms.v(126[12] 289[6])
    defparam i10658_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i28777_4_lut (.I0(n31_adj_4133), .I1(n29_adj_4131), .I2(n27_adj_4129), 
            .I3(n25_adj_4127), .O(n44296));
    defparam i28777_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i28766_4_lut (.I0(n37_adj_4138), .I1(n35_adj_4136), .I2(n33_adj_4135), 
            .I3(n44296), .O(n44285));
    defparam i28766_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i10659_3_lut (.I0(\data_in[2] [7]), .I1(\data_in[3] [7]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n24077));   // verilog/coms.v(126[12] 289[6])
    defparam i10659_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10660_3_lut (.I0(\data_in[2] [6]), .I1(\data_in[3] [6]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n24078));   // verilog/coms.v(126[12] 289[6])
    defparam i10660_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_11_LessThan_1210_i24_4_lut (.I0(n381), .I1(n99), .I2(n1874), 
            .I3(n558), .O(n24_adj_4126));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1210_i24_4_lut.LUT_INIT = 16'h0317;
    SB_LUT4 div_11_LessThan_570_i45_2_lut (.I0(n915), .I1(n96), .I2(GND_net), 
            .I3(GND_net), .O(n45));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_570_i45_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_11_LessThan_1210_i32_3_lut (.I0(n30_adj_4132), .I1(n93), 
            .I2(n35_adj_4136), .I3(GND_net), .O(n32_adj_4134));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1210_i32_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i10661_3_lut (.I0(\data_in[2] [5]), .I1(\data_in[3] [5]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n24079));   // verilog/coms.v(126[12] 289[6])
    defparam i10661_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_11_LessThan_657_i43_2_lut (.I0(n1045), .I1(n96), .I2(GND_net), 
            .I3(GND_net), .O(n43));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_657_i43_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 LessThan_539_i6_3_lut_3_lut (.I0(pwm_count[3]), .I1(pwm[3]), 
            .I2(pwm[2]), .I3(GND_net), .O(n6_adj_4020));   // verilog/motorControl.v(65[19:32])
    defparam LessThan_539_i6_3_lut_3_lut.LUT_INIT = 16'hd4d4;
    SB_LUT4 div_11_LessThan_742_i41_2_lut (.I0(n1172), .I1(n96), .I2(GND_net), 
            .I3(GND_net), .O(n41));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_742_i41_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i10748_3_lut (.I0(IntegralLimit[4]), .I1(\data_in_frame[10] [4]), 
            .I2(n23399), .I3(GND_net), .O(n24166));   // verilog/coms.v(126[12] 289[6])
    defparam i10748_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_11_LessThan_825_i41_2_lut (.I0(n1295), .I1(n95), .I2(GND_net), 
            .I3(GND_net), .O(n41_adj_4087));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_825_i41_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_11_LessThan_1210_i36_3_lut (.I0(n28_adj_4130), .I1(n91), 
            .I2(n39_adj_4139), .I3(GND_net), .O(n36_adj_4137));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1210_i36_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 div_11_LessThan_825_i43_2_lut (.I0(n1294), .I1(n94), .I2(GND_net), 
            .I3(GND_net), .O(n43_adj_4088));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_825_i43_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_11_LessThan_825_i39_2_lut (.I0(n1296), .I1(n96), .I2(GND_net), 
            .I3(GND_net), .O(n39));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_825_i39_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i10749_3_lut (.I0(IntegralLimit[3]), .I1(\data_in_frame[10] [3]), 
            .I2(n23399), .I3(GND_net), .O(n24167));   // verilog/coms.v(126[12] 289[6])
    defparam i10749_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i30566_4_lut (.I0(n36_adj_4137), .I1(n26_adj_4128), .I2(n39_adj_4139), 
            .I3(n44281), .O(n46087));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i30566_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i30567_3_lut (.I0(n46087), .I1(n90), .I2(n41_adj_4140), .I3(GND_net), 
            .O(n46088));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i30567_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 div_11_LessThan_825_i45_2_lut (.I0(n1293), .I1(n93), .I2(GND_net), 
            .I3(GND_net), .O(n45_adj_4090));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_825_i45_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i10750_3_lut (.I0(IntegralLimit[2]), .I1(\data_in_frame[10] [2]), 
            .I2(n23399), .I3(GND_net), .O(n24168));   // verilog/coms.v(126[12] 289[6])
    defparam i10750_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i30506_3_lut (.I0(n46088), .I1(n89), .I2(n43_adj_4141), .I3(GND_net), 
            .O(n46027));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i30506_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 div_11_LessThan_906_i39_2_lut (.I0(n1416), .I1(n95), .I2(GND_net), 
            .I3(GND_net), .O(n39_adj_4092));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_906_i39_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i10751_3_lut (.I0(IntegralLimit[1]), .I1(\data_in_frame[10] [1]), 
            .I2(n23399), .I3(GND_net), .O(n24169));   // verilog/coms.v(126[12] 289[6])
    defparam i10751_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_11_LessThan_906_i41_2_lut (.I0(n1415), .I1(n94), .I2(GND_net), 
            .I3(GND_net), .O(n41_adj_4093));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_906_i41_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_11_LessThan_906_i37_2_lut (.I0(n1417), .I1(n96), .I2(GND_net), 
            .I3(GND_net), .O(n37));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_906_i37_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_11_LessThan_906_i43_2_lut (.I0(n1414), .I1(n93), .I2(GND_net), 
            .I3(GND_net), .O(n43_adj_4094));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_906_i43_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_11_LessThan_985_i35_2_lut (.I0(n1535), .I1(n96), .I2(GND_net), 
            .I3(GND_net), .O(n35));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_985_i35_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i30163_4_lut (.I0(n43_adj_4141), .I1(n41_adj_4140), .I2(n39_adj_4139), 
            .I3(n44285), .O(n45684));
    defparam i30163_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i10752_3_lut (.I0(encoder1_position[1]), .I1(n2249), .I2(count_enable_adj_3992), 
            .I3(GND_net), .O(n24170));   // quad.v(35[10] 41[6])
    defparam i10752_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i30223_4_lut (.I0(n32_adj_4134), .I1(n24_adj_4126), .I2(n35_adj_4136), 
            .I3(n44291), .O(n45744));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i30223_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 div_11_LessThan_985_i33_2_lut (.I0(n1536), .I1(n97), .I2(GND_net), 
            .I3(GND_net), .O(n33));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_985_i33_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_11_LessThan_985_i37_2_lut (.I0(n1534), .I1(n95), .I2(GND_net), 
            .I3(GND_net), .O(n37_adj_4098));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_985_i37_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_11_LessThan_985_i39_2_lut (.I0(n1533), .I1(n94), .I2(GND_net), 
            .I3(GND_net), .O(n39_adj_4099));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_985_i39_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_11_LessThan_985_i43_2_lut (.I0(n1531), .I1(n92), .I2(GND_net), 
            .I3(GND_net), .O(n43_adj_4102));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_985_i43_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_11_LessThan_985_i41_2_lut (.I0(n1532), .I1(n93), .I2(GND_net), 
            .I3(GND_net), .O(n41_adj_4100));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_985_i41_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_11_LessThan_985_i45_2_lut (.I0(n1530), .I1(n91), .I2(GND_net), 
            .I3(GND_net), .O(n45_adj_4103));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_985_i45_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i30428_3_lut (.I0(n46027), .I1(n88), .I2(n45_adj_4143), .I3(GND_net), 
            .O(n44_adj_4142));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i30428_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 div_11_LessThan_1062_i33_2_lut (.I0(n1650), .I1(n96), .I2(GND_net), 
            .I3(GND_net), .O(n33_adj_4108));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1062_i33_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_11_LessThan_1062_i31_2_lut (.I0(n1651), .I1(n97), .I2(GND_net), 
            .I3(GND_net), .O(n31_adj_4106));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1062_i31_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_11_LessThan_1062_i35_2_lut (.I0(n1649), .I1(n95), .I2(GND_net), 
            .I3(GND_net), .O(n35_adj_4109));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1062_i35_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i10753_4_lut (.I0(r_Rx_Data), .I1(rx_data[0]), .I2(n4_adj_3984), 
            .I3(n22466), .O(n24171));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i10753_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 div_11_LessThan_1062_i37_2_lut (.I0(n1648), .I1(n94), .I2(GND_net), 
            .I3(GND_net), .O(n37_adj_4110));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1062_i37_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_11_LessThan_1062_i41_2_lut (.I0(n1646), .I1(n92), .I2(GND_net), 
            .I3(GND_net), .O(n41_adj_4113));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1062_i41_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_11_LessThan_1062_i39_2_lut (.I0(n1647), .I1(n93), .I2(GND_net), 
            .I3(GND_net), .O(n39_adj_4111));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1062_i39_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_11_LessThan_1062_i43_2_lut (.I0(n1645), .I1(n91), .I2(GND_net), 
            .I3(GND_net), .O(n43_adj_4114));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1062_i43_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i30225_4_lut (.I0(n44_adj_4142), .I1(n45744), .I2(n45_adj_4143), 
            .I3(n45684), .O(n45746));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i30225_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i1_4_lut_adj_1467 (.I0(n45746), .I1(n22439), .I2(n87), .I3(n1862), 
            .O(n1886));
    defparam i1_4_lut_adj_1467.LUT_INIT = 16'hceef;
    SB_LUT4 i1_2_lut_adj_1468 (.I0(n88), .I1(n22436), .I2(GND_net), .I3(GND_net), 
            .O(n22433));
    defparam i1_2_lut_adj_1468.LUT_INIT = 16'hdddd;
    SB_LUT4 i10754_4_lut (.I0(pwm_23__N_2957), .I1(n471), .I2(PWMLimit[0]), 
            .I3(n387), .O(n24172));   // verilog/motorControl.v(38[14] 59[8])
    defparam i10754_4_lut.LUT_INIT = 16'ha088;
    SB_LUT4 div_11_mux_3_i11_3_lut (.I0(encoder0_position[10]), .I1(n15), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n381));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_mux_3_i11_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_11_LessThan_1137_i31_2_lut (.I0(n1762), .I1(n96), .I2(GND_net), 
            .I3(GND_net), .O(n31_adj_4119));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1137_i31_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_11_LessThan_1137_i29_2_lut (.I0(n1763), .I1(n97), .I2(GND_net), 
            .I3(GND_net), .O(n29_adj_4117));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1137_i29_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i10280_3_lut (.I0(n23560), .I1(r_Bit_Index[0]), .I2(n23471), 
            .I3(GND_net), .O(n23698));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i10280_3_lut.LUT_INIT = 16'h1414;
    SB_LUT4 div_11_LessThan_1137_i33_2_lut (.I0(n1761), .I1(n95), .I2(GND_net), 
            .I3(GND_net), .O(n33_adj_4120));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1137_i33_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_11_LessThan_1137_i35_2_lut (.I0(n1760), .I1(n94), .I2(GND_net), 
            .I3(GND_net), .O(n35_adj_4121));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1137_i35_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_11_LessThan_1137_i39_2_lut (.I0(n1758), .I1(n92), .I2(GND_net), 
            .I3(GND_net), .O(n39_adj_4124));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1137_i39_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_11_LessThan_1137_i37_2_lut (.I0(n1759), .I1(n93), .I2(GND_net), 
            .I3(GND_net), .O(n37_adj_4122));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1137_i37_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_11_mux_5_i1_3_lut (.I0(gearBoxRatio[0]), .I1(n75), .I2(gearBoxRatio[23]), 
            .I3(GND_net), .O(n558));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_mux_5_i1_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 i10277_3_lut (.I0(n23562), .I1(r_Bit_Index_adj_4399[0]), .I2(n23477), 
            .I3(GND_net), .O(n23695));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i10277_3_lut.LUT_INIT = 16'h1414;
    SB_LUT4 div_11_i1271_3_lut (.I0(n381), .I1(n6834), .I2(n1886), .I3(GND_net), 
            .O(n1980));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1271_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_11_LessThan_1137_i41_2_lut (.I0(n1757), .I1(n91), .I2(GND_net), 
            .I3(GND_net), .O(n41_adj_4125));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1137_i41_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_11_LessThan_1210_i31_2_lut (.I0(n1870), .I1(n95), .I2(GND_net), 
            .I3(GND_net), .O(n31_adj_4133));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1210_i31_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_11_LessThan_1210_i33_2_lut (.I0(n1869), .I1(n94), .I2(GND_net), 
            .I3(GND_net), .O(n33_adj_4135));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1210_i33_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_11_LessThan_1210_i29_2_lut (.I0(n1871), .I1(n96), .I2(GND_net), 
            .I3(GND_net), .O(n29_adj_4131));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1210_i29_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_11_LessThan_1210_i37_2_lut (.I0(n1867), .I1(n92), .I2(GND_net), 
            .I3(GND_net), .O(n37_adj_4138));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1210_i37_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_11_mux_5_i2_3_lut (.I0(gearBoxRatio[1]), .I1(n74), .I2(gearBoxRatio[23]), 
            .I3(GND_net), .O(n99));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_mux_5_i2_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 div_11_LessThan_1210_i27_2_lut (.I0(n1872), .I1(n97), .I2(GND_net), 
            .I3(GND_net), .O(n27_adj_4129));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1210_i27_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_11_LessThan_1210_i39_2_lut (.I0(n1866), .I1(n91), .I2(GND_net), 
            .I3(GND_net), .O(n39_adj_4139));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1210_i39_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_11_mux_3_i10_3_lut (.I0(encoder0_position[9]), .I1(n16), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n382));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_mux_3_i10_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_11_LessThan_1210_i41_2_lut (.I0(n1865), .I1(n90), .I2(GND_net), 
            .I3(GND_net), .O(n41_adj_4140));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1210_i41_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_11_LessThan_1210_i43_2_lut (.I0(n1864), .I1(n89), .I2(GND_net), 
            .I3(GND_net), .O(n43_adj_4141));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1210_i43_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_11_LessThan_1210_i35_2_lut (.I0(n1868), .I1(n93), .I2(GND_net), 
            .I3(GND_net), .O(n35_adj_4136));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1210_i35_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i10162_3_lut (.I0(IntegralLimit[0]), .I1(\data_in_frame[10] [0]), 
            .I2(n23399), .I3(GND_net), .O(n23580));   // verilog/coms.v(126[12] 289[6])
    defparam i10162_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10163_3_lut (.I0(Kp[0]), .I1(\data_in_frame[2] [0]), .I2(n23399), 
            .I3(GND_net), .O(n23581));   // verilog/coms.v(126[12] 289[6])
    defparam i10163_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10164_3_lut (.I0(Ki[0]), .I1(\data_in_frame[3] [0]), .I2(n23399), 
            .I3(GND_net), .O(n23582));   // verilog/coms.v(126[12] 289[6])
    defparam i10164_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_11_LessThan_1281_i33_2_lut (.I0(n1974), .I1(n93), .I2(GND_net), 
            .I3(GND_net), .O(n33_adj_4154));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1281_i33_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_11_mux_5_i8_3_lut (.I0(gearBoxRatio[7]), .I1(n68), .I2(gearBoxRatio[23]), 
            .I3(GND_net), .O(n93));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_mux_5_i8_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 i10165_3_lut (.I0(Kd[0]), .I1(\data_in_frame[4] [0]), .I2(n23399), 
            .I3(GND_net), .O(n23583));   // verilog/coms.v(126[12] 289[6])
    defparam i10165_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_11_LessThan_1281_i29_2_lut (.I0(n1976), .I1(n95), .I2(GND_net), 
            .I3(GND_net), .O(n29_adj_4151));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1281_i29_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i10166_3_lut (.I0(gearBoxRatio[0]), .I1(\data_in_frame[19] [0]), 
            .I2(n23399), .I3(GND_net), .O(n23584));   // verilog/coms.v(126[12] 289[6])
    defparam i10166_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10167_3_lut (.I0(\data_in[0] [0]), .I1(\data_in[1] [0]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n23585));   // verilog/coms.v(126[12] 289[6])
    defparam i10167_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_11_LessThan_1281_i31_2_lut (.I0(n1975), .I1(n94), .I2(GND_net), 
            .I3(GND_net), .O(n31_adj_4153));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1281_i31_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_11_LessThan_1281_i23_2_lut (.I0(n1979), .I1(n98), .I2(GND_net), 
            .I3(GND_net), .O(n23_adj_4145));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1281_i23_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i10765_3_lut (.I0(encoder1_position[2]), .I1(n2248), .I2(count_enable_adj_3992), 
            .I3(GND_net), .O(n24183));   // quad.v(35[10] 41[6])
    defparam i10765_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i28738_4_lut (.I0(n29_adj_4151), .I1(n27_adj_4149), .I2(n25_adj_4147), 
            .I3(n23_adj_4145), .O(n44257));
    defparam i28738_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i10169_3_lut (.I0(control_mode[0]), .I1(\data_in_frame[1] [0]), 
            .I2(n23399), .I3(GND_net), .O(n23587));   // verilog/coms.v(126[12] 289[6])
    defparam i10169_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10766_3_lut (.I0(encoder1_position[3]), .I1(n2247), .I2(count_enable_adj_3992), 
            .I3(GND_net), .O(n24184));   // quad.v(35[10] 41[6])
    defparam i10766_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10170_3_lut (.I0(PWMLimit[0]), .I1(\data_in_frame[7] [0]), 
            .I2(n23399), .I3(GND_net), .O(n23588));   // verilog/coms.v(126[12] 289[6])
    defparam i10170_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10171_3_lut (.I0(\PID_CONTROLLER.err_prev [0]), .I1(\PID_CONTROLLER.err [0]), 
            .I2(n41887), .I3(GND_net), .O(n23589));   // verilog/motorControl.v(38[14] 59[8])
    defparam i10171_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i28730_4_lut (.I0(n35_adj_4156), .I1(n33_adj_4154), .I2(n31_adj_4153), 
            .I3(n44257), .O(n44249));
    defparam i28730_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i10767_3_lut (.I0(encoder1_position[4]), .I1(n2246), .I2(count_enable_adj_3992), 
            .I3(GND_net), .O(n24185));   // quad.v(35[10] 41[6])
    defparam i10767_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10768_3_lut (.I0(encoder1_position[5]), .I1(n2245), .I2(count_enable_adj_3992), 
            .I3(GND_net), .O(n24186));   // quad.v(35[10] 41[6])
    defparam i10768_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_11_LessThan_1281_i22_4_lut (.I0(n382), .I1(n99), .I2(n1980), 
            .I3(n558), .O(n22_adj_4144));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1281_i22_4_lut.LUT_INIT = 16'h0317;
    SB_LUT4 i10173_3_lut (.I0(encoder0_position[0]), .I1(n2300), .I2(count_enable), 
            .I3(GND_net), .O(n23591));   // quad.v(35[10] 41[6])
    defparam i10173_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10174_3_lut (.I0(encoder1_position[0]), .I1(n2250), .I2(count_enable_adj_3992), 
            .I3(GND_net), .O(n23592));   // quad.v(35[10] 41[6])
    defparam i10174_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10769_3_lut (.I0(encoder1_position[6]), .I1(n2244), .I2(count_enable_adj_3992), 
            .I3(GND_net), .O(n24187));   // quad.v(35[10] 41[6])
    defparam i10769_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10175_3_lut (.I0(quadB_debounced), .I1(reg_B[0]), .I2(n41998), 
            .I3(GND_net), .O(n23593));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(186[9] 190[16])
    defparam i10175_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_11_LessThan_1281_i30_3_lut (.I0(n28_adj_4150), .I1(n93), 
            .I2(n33_adj_4154), .I3(GND_net), .O(n30_adj_4152));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1281_i30_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i10176_4_lut (.I0(r_SM_Main[2]), .I1(n1_adj_4357), .I2(n28231), 
            .I3(r_SM_Main[1]), .O(n23594));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i10176_4_lut.LUT_INIT = 16'h0544;
    SB_LUT4 i10770_3_lut (.I0(encoder1_position[7]), .I1(n2243), .I2(count_enable_adj_3992), 
            .I3(GND_net), .O(n24188));   // quad.v(35[10] 41[6])
    defparam i10770_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10177_3_lut (.I0(quadB_debounced_adj_3991), .I1(reg_B_adj_4406[0]), 
            .I2(n41767), .I3(GND_net), .O(n23595));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(186[9] 190[16])
    defparam i10177_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i10771_3_lut (.I0(encoder1_position[8]), .I1(n2242), .I2(count_enable_adj_3992), 
            .I3(GND_net), .O(n24189));   // quad.v(35[10] 41[6])
    defparam i10771_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10772_3_lut (.I0(encoder1_position[9]), .I1(n2241), .I2(count_enable_adj_3992), 
            .I3(GND_net), .O(n24190));   // quad.v(35[10] 41[6])
    defparam i10772_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10773_3_lut (.I0(encoder1_position[10]), .I1(n2240), .I2(count_enable_adj_3992), 
            .I3(GND_net), .O(n24191));   // quad.v(35[10] 41[6])
    defparam i10773_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10774_3_lut (.I0(encoder1_position[11]), .I1(n2239), .I2(count_enable_adj_3992), 
            .I3(GND_net), .O(n24192));   // quad.v(35[10] 41[6])
    defparam i10774_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_11_LessThan_1281_i34_3_lut (.I0(n26_adj_4148), .I1(n91), 
            .I2(n37_adj_4157), .I3(GND_net), .O(n34_adj_4155));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1281_i34_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i10775_3_lut (.I0(encoder1_position[12]), .I1(n2238), .I2(count_enable_adj_3992), 
            .I3(GND_net), .O(n24193));   // quad.v(35[10] 41[6])
    defparam i10775_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i30568_4_lut (.I0(n34_adj_4155), .I1(n24_adj_4146), .I2(n37_adj_4157), 
            .I3(n44245), .O(n46089));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i30568_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i10181_3_lut (.I0(setpoint[0]), .I1(n3792), .I2(n23430), .I3(GND_net), 
            .O(n23599));   // verilog/coms.v(126[12] 289[6])
    defparam i10181_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10776_3_lut (.I0(encoder1_position[13]), .I1(n2237), .I2(count_enable_adj_3992), 
            .I3(GND_net), .O(n24194));   // quad.v(35[10] 41[6])
    defparam i10776_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10777_3_lut (.I0(encoder1_position[14]), .I1(n2236), .I2(count_enable_adj_3992), 
            .I3(GND_net), .O(n24195));   // quad.v(35[10] 41[6])
    defparam i10777_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i30569_3_lut (.I0(n46089), .I1(n90), .I2(n39_adj_4158), .I3(GND_net), 
            .O(n46090));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i30569_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i10778_3_lut (.I0(encoder1_position[15]), .I1(n2235), .I2(count_enable_adj_3992), 
            .I3(GND_net), .O(n24196));   // quad.v(35[10] 41[6])
    defparam i10778_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10779_3_lut (.I0(encoder1_position[16]), .I1(n2234), .I2(count_enable_adj_3992), 
            .I3(GND_net), .O(n24197));   // quad.v(35[10] 41[6])
    defparam i10779_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i30504_3_lut (.I0(n46090), .I1(n89), .I2(n41_adj_4159), .I3(GND_net), 
            .O(n46025));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i30504_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i30153_4_lut (.I0(n41_adj_4159), .I1(n39_adj_4158), .I2(n37_adj_4157), 
            .I3(n44249), .O(n45674));
    defparam i30153_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i30345_4_lut (.I0(n30_adj_4152), .I1(n22_adj_4144), .I2(n33_adj_4154), 
            .I3(n44255), .O(n45866));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i30345_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i10780_3_lut (.I0(encoder1_position[17]), .I1(n2233), .I2(count_enable_adj_3992), 
            .I3(GND_net), .O(n24198));   // quad.v(35[10] 41[6])
    defparam i10780_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10781_3_lut (.I0(encoder1_position[18]), .I1(n2232), .I2(count_enable_adj_3992), 
            .I3(GND_net), .O(n24199));   // quad.v(35[10] 41[6])
    defparam i10781_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10782_3_lut (.I0(encoder1_position[19]), .I1(n2231), .I2(count_enable_adj_3992), 
            .I3(GND_net), .O(n24200));   // quad.v(35[10] 41[6])
    defparam i10782_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10783_3_lut (.I0(encoder1_position[20]), .I1(n2230), .I2(count_enable_adj_3992), 
            .I3(GND_net), .O(n24201));   // quad.v(35[10] 41[6])
    defparam i10783_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i30430_3_lut (.I0(n46025), .I1(n88), .I2(n43_adj_4161), .I3(GND_net), 
            .O(n42_adj_4160));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i30430_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i30525_4_lut (.I0(n42_adj_4160), .I1(n45866), .I2(n43_adj_4161), 
            .I3(n45674), .O(n46046));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i30525_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i10784_3_lut (.I0(encoder1_position[21]), .I1(n2229), .I2(count_enable_adj_3992), 
            .I3(GND_net), .O(n24202));   // quad.v(35[10] 41[6])
    defparam i10784_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10785_3_lut (.I0(encoder1_position[22]), .I1(n2228), .I2(count_enable_adj_3992), 
            .I3(GND_net), .O(n24203));   // quad.v(35[10] 41[6])
    defparam i10785_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i30526_3_lut (.I0(n46046), .I1(n87), .I2(n1968), .I3(GND_net), 
            .O(n46047));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i30526_3_lut.LUT_INIT = 16'h2b2b;
    SB_LUT4 mux_22_i17_4_lut (.I0(encoder1_position[16]), .I1(displacement[16]), 
            .I2(n15_adj_3962), .I3(n15_adj_3963), .O(motor_state_23__N_27[16]));   // verilog/TinyFPGA_B.v(138[5] 141[10])
    defparam mux_22_i17_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i10786_3_lut (.I0(encoder1_position[23]), .I1(n2227), .I2(count_enable_adj_3992), 
            .I3(GND_net), .O(n24204));   // quad.v(35[10] 41[6])
    defparam i10786_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_1469 (.I0(n46047), .I1(n22442), .I2(n86), .I3(n1967), 
            .O(n1991));
    defparam i1_4_lut_adj_1469.LUT_INIT = 16'hceef;
    SB_LUT4 mux_21_i17_3_lut (.I0(encoder0_position[16]), .I1(motor_state_23__N_27[16]), 
            .I2(n15_adj_3961), .I3(GND_net), .O(motor_state[16]));   // verilog/TinyFPGA_B.v(137[5] 141[10])
    defparam mux_21_i17_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10182_3_lut (.I0(deadband[0]), .I1(\data_in_frame[13] [0]), 
            .I2(n23399), .I3(GND_net), .O(n23600));   // verilog/coms.v(126[12] 289[6])
    defparam i10182_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_11_i1265_3_lut (.I0(n1869), .I1(n6828), .I2(n1886), .I3(GND_net), 
            .O(n1974));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1265_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_11_mux_5_i9_3_lut (.I0(gearBoxRatio[8]), .I1(n67), .I2(gearBoxRatio[23]), 
            .I3(GND_net), .O(n92));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_mux_5_i9_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 i10787_4_lut (.I0(pwm_23__N_2957), .I1(n470), .I2(PWMLimit[1]), 
            .I3(n387), .O(n24205));   // verilog/motorControl.v(38[14] 59[8])
    defparam i10787_4_lut.LUT_INIT = 16'ha088;
    SB_LUT4 i10700_3_lut (.I0(gearBoxRatio[5]), .I1(\data_in_frame[19] [5]), 
            .I2(n23399), .I3(GND_net), .O(n24118));   // verilog/coms.v(126[12] 289[6])
    defparam i10700_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_11_i1334_3_lut (.I0(n1974), .I1(n6844), .I2(n1991), .I3(GND_net), 
            .O(n2076));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1334_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i10701_3_lut (.I0(gearBoxRatio[4]), .I1(\data_in_frame[19] [4]), 
            .I2(n23399), .I3(GND_net), .O(n24119));   // verilog/coms.v(126[12] 289[6])
    defparam i10701_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10788_4_lut (.I0(pwm_23__N_2957), .I1(n469), .I2(PWMLimit[2]), 
            .I3(n387), .O(n24206));   // verilog/motorControl.v(38[14] 59[8])
    defparam i10788_4_lut.LUT_INIT = 16'ha088;
    SB_LUT4 div_11_mux_5_i7_3_lut (.I0(gearBoxRatio[6]), .I1(n69), .I2(gearBoxRatio[23]), 
            .I3(GND_net), .O(n94));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_mux_5_i7_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 i10702_3_lut (.I0(gearBoxRatio[3]), .I1(\data_in_frame[19] [3]), 
            .I2(n23399), .I3(GND_net), .O(n24120));   // verilog/coms.v(126[12] 289[6])
    defparam i10702_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10789_4_lut (.I0(pwm_23__N_2957), .I1(n468), .I2(PWMLimit[3]), 
            .I3(n387), .O(n24207));   // verilog/motorControl.v(38[14] 59[8])
    defparam i10789_4_lut.LUT_INIT = 16'ha088;
    SB_LUT4 div_11_i1336_3_lut (.I0(n1976), .I1(n6846), .I2(n1991), .I3(GND_net), 
            .O(n2078));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1336_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_11_LessThan_1350_i29_2_lut (.I0(n2078), .I1(n94), .I2(GND_net), 
            .I3(GND_net), .O(n29_adj_4171));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1350_i29_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i10790_4_lut (.I0(pwm_23__N_2957), .I1(n467), .I2(PWMLimit[4]), 
            .I3(n387), .O(n24208));   // verilog/motorControl.v(38[14] 59[8])
    defparam i10790_4_lut.LUT_INIT = 16'ha088;
    SB_LUT4 div_11_LessThan_1350_i31_2_lut (.I0(n2077), .I1(n93), .I2(GND_net), 
            .I3(GND_net), .O(n31_adj_4172));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1350_i31_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 mux_22_i18_4_lut (.I0(encoder1_position[17]), .I1(displacement[17]), 
            .I2(n15_adj_3962), .I3(n15_adj_3963), .O(motor_state_23__N_27[17]));   // verilog/TinyFPGA_B.v(138[5] 141[10])
    defparam mux_22_i18_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i5_3_lut (.I0(\PID_CONTROLLER.result [5]), .I1(n415), .I2(n421), 
            .I3(GND_net), .O(n1));
    defparam i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_21_i18_3_lut (.I0(encoder0_position[17]), .I1(motor_state_23__N_27[17]), 
            .I2(n15_adj_3961), .I3(GND_net), .O(motor_state[17]));   // verilog/TinyFPGA_B.v(137[5] 141[10])
    defparam mux_21_i18_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10703_3_lut (.I0(gearBoxRatio[2]), .I1(\data_in_frame[19] [2]), 
            .I2(n23399), .I3(GND_net), .O(n24121));   // verilog/coms.v(126[12] 289[6])
    defparam i10703_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_11_LessThan_1350_i33_2_lut (.I0(n2076), .I1(n92), .I2(GND_net), 
            .I3(GND_net), .O(n33_adj_4174));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1350_i33_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i13810_3_lut (.I0(\PID_CONTROLLER.result [6]), .I1(n414), .I2(n421), 
            .I3(GND_net), .O(n27212));
    defparam i13810_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_22_i19_4_lut (.I0(encoder1_position[18]), .I1(displacement[18]), 
            .I2(n15_adj_3962), .I3(n15_adj_3963), .O(motor_state_23__N_27[18]));   // verilog/TinyFPGA_B.v(138[5] 141[10])
    defparam mux_22_i19_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_21_i19_3_lut (.I0(encoder0_position[18]), .I1(motor_state_23__N_27[18]), 
            .I2(n15_adj_3961), .I3(GND_net), .O(motor_state[18]));   // verilog/TinyFPGA_B.v(137[5] 141[10])
    defparam mux_21_i19_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_11_mux_5_i3_3_lut (.I0(gearBoxRatio[2]), .I1(n73), .I2(gearBoxRatio[23]), 
            .I3(GND_net), .O(n98));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_mux_5_i3_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 i10793_4_lut (.I0(pwm_23__N_2957), .I1(n464), .I2(PWMLimit[7]), 
            .I3(n387), .O(n24211));   // verilog/motorControl.v(38[14] 59[8])
    defparam i10793_4_lut.LUT_INIT = 16'ha088;
    SB_LUT4 div_11_i1340_3_lut (.I0(n1980), .I1(n6850), .I2(n1991), .I3(GND_net), 
            .O(n2082));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1340_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_11_LessThan_1350_i21_2_lut (.I0(n2082), .I1(n98), .I2(GND_net), 
            .I3(GND_net), .O(n21_adj_4163));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1350_i21_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i10794_4_lut (.I0(pwm_23__N_2957), .I1(n463), .I2(PWMLimit[8]), 
            .I3(n387), .O(n24212));   // verilog/motorControl.v(38[14] 59[8])
    defparam i10794_4_lut.LUT_INIT = 16'ha088;
    SB_LUT4 i28710_4_lut (.I0(n27_adj_4169), .I1(n25_adj_4167), .I2(n23_adj_4165), 
            .I3(n21_adj_4163), .O(n44229));
    defparam i28710_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i10795_4_lut (.I0(pwm_23__N_2957), .I1(n462), .I2(PWMLimit[9]), 
            .I3(n387), .O(n24213));   // verilog/motorControl.v(38[14] 59[8])
    defparam i10795_4_lut.LUT_INIT = 16'ha088;
    SB_LUT4 i28704_4_lut (.I0(n33_adj_4174), .I1(n31_adj_4172), .I2(n29_adj_4171), 
            .I3(n44229), .O(n44223));
    defparam i28704_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 div_11_LessThan_1350_i20_4_lut (.I0(n383), .I1(n99), .I2(n2083), 
            .I3(n558), .O(n20_adj_4162));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1350_i20_4_lut.LUT_INIT = 16'h0317;
    SB_LUT4 i10796_4_lut (.I0(pwm_23__N_2957), .I1(n461), .I2(PWMLimit[9]), 
            .I3(n387), .O(n24214));   // verilog/motorControl.v(38[14] 59[8])
    defparam i10796_4_lut.LUT_INIT = 16'ha088;
    SB_LUT4 div_11_LessThan_1350_i28_3_lut (.I0(n26_adj_4168), .I1(n93), 
            .I2(n31_adj_4172), .I3(GND_net), .O(n28_adj_4170));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1350_i28_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i10797_4_lut (.I0(pwm_23__N_2957), .I1(n460), .I2(PWMLimit[9]), 
            .I3(n387), .O(n24215));   // verilog/motorControl.v(38[14] 59[8])
    defparam i10797_4_lut.LUT_INIT = 16'ha088;
    SB_LUT4 i10798_4_lut (.I0(pwm_23__N_2957), .I1(n459), .I2(PWMLimit[9]), 
            .I3(n387), .O(n24216));   // verilog/motorControl.v(38[14] 59[8])
    defparam i10798_4_lut.LUT_INIT = 16'ha088;
    SB_LUT4 i10799_4_lut (.I0(pwm_23__N_2957), .I1(n458), .I2(PWMLimit[9]), 
            .I3(n387), .O(n24217));   // verilog/motorControl.v(38[14] 59[8])
    defparam i10799_4_lut.LUT_INIT = 16'ha088;
    SB_LUT4 div_11_LessThan_1350_i32_3_lut (.I0(n24_adj_4166), .I1(n91), 
            .I2(n35_adj_4175), .I3(GND_net), .O(n32_adj_4173));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1350_i32_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i30570_4_lut (.I0(n32_adj_4173), .I1(n22_adj_4164), .I2(n35_adj_4175), 
            .I3(n44221), .O(n46091));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i30570_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i10800_4_lut (.I0(pwm_23__N_2957), .I1(n457), .I2(PWMLimit[9]), 
            .I3(n387), .O(n24218));   // verilog/motorControl.v(38[14] 59[8])
    defparam i10800_4_lut.LUT_INIT = 16'ha088;
    SB_LUT4 i30571_3_lut (.I0(n46091), .I1(n90), .I2(n37_adj_4176), .I3(GND_net), 
            .O(n46092));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i30571_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i30502_3_lut (.I0(n46092), .I1(n89), .I2(n39_adj_4177), .I3(GND_net), 
            .O(n46023));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i30502_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i10801_4_lut (.I0(pwm_23__N_2957), .I1(n456), .I2(PWMLimit[9]), 
            .I3(n387), .O(n24219));   // verilog/motorControl.v(38[14] 59[8])
    defparam i10801_4_lut.LUT_INIT = 16'ha088;
    SB_LUT4 i30137_4_lut (.I0(n39_adj_4177), .I1(n37_adj_4176), .I2(n35_adj_4175), 
            .I3(n44223), .O(n45658));
    defparam i30137_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i30572_4_lut (.I0(n28_adj_4170), .I1(n20_adj_4162), .I2(n31_adj_4172), 
            .I3(n44225), .O(n46093));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i30572_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i30434_3_lut (.I0(n46023), .I1(n88), .I2(n41_adj_4178), .I3(GND_net), 
            .O(n45955));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i30434_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i10802_4_lut (.I0(pwm_23__N_2957), .I1(n455), .I2(PWMLimit[9]), 
            .I3(n387), .O(n24220));   // verilog/motorControl.v(38[14] 59[8])
    defparam i10802_4_lut.LUT_INIT = 16'ha088;
    SB_LUT4 i30647_4_lut (.I0(n45955), .I1(n46093), .I2(n41_adj_4178), 
            .I3(n45658), .O(n46168));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i30647_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i30648_3_lut (.I0(n46168), .I1(n87), .I2(n2071), .I3(GND_net), 
            .O(n46169));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i30648_3_lut.LUT_INIT = 16'h2b2b;
    SB_LUT4 i30583_3_lut (.I0(n46169), .I1(n86), .I2(n2070), .I3(GND_net), 
            .O(n46104));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i30583_3_lut.LUT_INIT = 16'h2b2b;
    SB_LUT4 i1_4_lut_adj_1470 (.I0(pwm_23__N_2957), .I1(n44153), .I2(PWMLimit[9]), 
            .I3(n387), .O(n39110));   // verilog/motorControl.v(38[14] 59[8])
    defparam i1_4_lut_adj_1470.LUT_INIT = 16'ha088;
    SB_LUT4 i1_4_lut_adj_1471 (.I0(n46104), .I1(n22445), .I2(n85), .I3(n2069), 
            .O(n2093));
    defparam i1_4_lut_adj_1471.LUT_INIT = 16'hceef;
    SB_LUT4 div_11_i1338_3_lut (.I0(n1978), .I1(n6848), .I2(n1991), .I3(GND_net), 
            .O(n2080));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1338_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_11_mux_5_i6_3_lut (.I0(gearBoxRatio[5]), .I1(n70), .I2(gearBoxRatio[23]), 
            .I3(GND_net), .O(n95));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_mux_5_i6_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 div_11_i1405_3_lut (.I0(n2080), .I1(n6865), .I2(n2093), .I3(GND_net), 
            .O(n2179));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1405_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i10805_4_lut (.I0(pwm_23__N_2957), .I1(n44109), .I2(PWMLimit[9]), 
            .I3(n387), .O(n24223));   // verilog/motorControl.v(38[14] 59[8])
    defparam i10805_4_lut.LUT_INIT = 16'ha088;
    SB_LUT4 LessThan_542_i6_3_lut_3_lut (.I0(pwm_count[3]), .I1(n873), .I2(n874), 
            .I3(GND_net), .O(n6_adj_4027));   // verilog/motorControl.v(86[28:44])
    defparam LessThan_542_i6_3_lut_3_lut.LUT_INIT = 16'hd4d4;
    SB_LUT4 i10806_4_lut (.I0(pwm_23__N_2957), .I1(n44111), .I2(PWMLimit[9]), 
            .I3(n387), .O(n24224));   // verilog/motorControl.v(38[14] 59[8])
    defparam i10806_4_lut.LUT_INIT = 16'ha088;
    SB_LUT4 div_11_LessThan_1417_i25_2_lut (.I0(n2179), .I1(n95), .I2(GND_net), 
            .I3(GND_net), .O(n25_adj_4186));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1417_i25_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_11_LessThan_1417_i27_2_lut (.I0(n2178), .I1(n94), .I2(GND_net), 
            .I3(GND_net), .O(n27_adj_4188));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1417_i27_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_11_LessThan_1417_i19_2_lut (.I0(n2182), .I1(n98), .I2(GND_net), 
            .I3(GND_net), .O(n19_adj_4180));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1417_i19_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i10720_3_lut (.I0(Kp[6]), .I1(\data_in_frame[2] [6]), .I2(n23399), 
            .I3(GND_net), .O(n24138));   // verilog/coms.v(126[12] 289[6])
    defparam i10720_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10807_4_lut (.I0(pwm_23__N_2957), .I1(n44113), .I2(PWMLimit[9]), 
            .I3(n387), .O(n24225));   // verilog/motorControl.v(38[14] 59[8])
    defparam i10807_4_lut.LUT_INIT = 16'ha088;
    SB_LUT4 i10721_3_lut (.I0(Kp[5]), .I1(\data_in_frame[2] [5]), .I2(n23399), 
            .I3(GND_net), .O(n24139));   // verilog/coms.v(126[12] 289[6])
    defparam i10721_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i28684_4_lut (.I0(n25_adj_4186), .I1(n23_adj_4184), .I2(n21_adj_4182), 
            .I3(n19_adj_4180), .O(n44203));
    defparam i28684_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i10722_3_lut (.I0(Kp[4]), .I1(\data_in_frame[2] [4]), .I2(n23399), 
            .I3(GND_net), .O(n24140));   // verilog/coms.v(126[12] 289[6])
    defparam i10722_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10723_3_lut (.I0(Kp[3]), .I1(\data_in_frame[2] [3]), .I2(n23399), 
            .I3(GND_net), .O(n24141));   // verilog/coms.v(126[12] 289[6])
    defparam i10723_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10724_3_lut (.I0(Kp[2]), .I1(\data_in_frame[2] [2]), .I2(n23399), 
            .I3(GND_net), .O(n24142));   // verilog/coms.v(126[12] 289[6])
    defparam i10724_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10725_3_lut (.I0(Kp[1]), .I1(\data_in_frame[2] [1]), .I2(n23399), 
            .I3(GND_net), .O(n24143));   // verilog/coms.v(126[12] 289[6])
    defparam i10725_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10726_3_lut (.I0(IntegralLimit[23]), .I1(\data_in_frame[8] [7]), 
            .I2(n23399), .I3(GND_net), .O(n24144));   // verilog/coms.v(126[12] 289[6])
    defparam i10726_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i28680_4_lut (.I0(n31_adj_4191), .I1(n29_adj_4189), .I2(n27_adj_4188), 
            .I3(n44203), .O(n44199));
    defparam i28680_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i30123_4_lut (.I0(n37_adj_4194), .I1(n35_adj_4193), .I2(n33_adj_4192), 
            .I3(n44199), .O(n45644));
    defparam i30123_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i10808_4_lut (.I0(pwm_23__N_2957), .I1(n44115), .I2(PWMLimit[9]), 
            .I3(n387), .O(n24226));   // verilog/motorControl.v(38[14] 59[8])
    defparam i10808_4_lut.LUT_INIT = 16'ha088;
    SB_LUT4 div_11_LessThan_1417_i18_4_lut (.I0(n384), .I1(n99), .I2(n2183), 
            .I3(n558), .O(n18_adj_4179));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1417_i18_4_lut.LUT_INIT = 16'h0317;
    SB_LUT4 i30131_3_lut (.I0(n18_adj_4179), .I1(n87), .I2(n41_adj_4196), 
            .I3(GND_net), .O(n45652));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i30131_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i30132_3_lut (.I0(n45652), .I1(n86), .I2(n43_adj_4197), .I3(GND_net), 
            .O(n45653));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i30132_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i29856_4_lut (.I0(n43_adj_4197), .I1(n41_adj_4196), .I2(n29_adj_4189), 
            .I3(n44201), .O(n45377));
    defparam i29856_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 div_11_LessThan_1417_i26_3_lut (.I0(n24_adj_4185), .I1(n93), 
            .I2(n29_adj_4189), .I3(GND_net), .O(n26_adj_4187));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1417_i26_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i9_2_lut (.I0(n414), .I1(\PID_CONTROLLER.result [6]), .I2(GND_net), 
            .I3(GND_net), .O(n13_adj_4018));   // verilog/motorControl.v(32[23:29])
    defparam i9_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i29613_3_lut (.I0(n45653), .I1(n85), .I2(n45_adj_4198), .I3(GND_net), 
            .O(n45134));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i29613_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i16_2_lut (.I0(n415), .I1(\PID_CONTROLLER.result [5]), .I2(GND_net), 
            .I3(GND_net), .O(n11_adj_4017));   // verilog/motorControl.v(32[23:29])
    defparam i16_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i10727_3_lut (.I0(IntegralLimit[22]), .I1(\data_in_frame[8] [6]), 
            .I2(n23399), .I3(GND_net), .O(n24145));   // verilog/coms.v(126[12] 289[6])
    defparam i10727_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_11_LessThan_1417_i30_3_lut (.I0(n22_adj_4183), .I1(n91), 
            .I2(n33_adj_4192), .I3(GND_net), .O(n30_adj_4190));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1417_i30_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i30574_4_lut (.I0(n30_adj_4190), .I1(n20_adj_4181), .I2(n33_adj_4192), 
            .I3(n44195), .O(n46095));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i30574_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i30575_3_lut (.I0(n46095), .I1(n90), .I2(n35_adj_4193), .I3(GND_net), 
            .O(n46096));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i30575_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i12039_3_lut (.I0(\data_out_frame[20] [7]), .I1(\data_out_frame[22] [7]), 
            .I2(byte_transmit_counter[1]), .I3(GND_net), .O(n25455));   // verilog/coms.v(100[12:33])
    defparam i12039_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i30498_3_lut (.I0(n46096), .I1(n89), .I2(n37_adj_4194), .I3(GND_net), 
            .O(n46019));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i30498_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i12042_4_lut (.I0(n25455), .I1(\data_out_frame[21] [7]), .I2(byte_transmit_counter[0]), 
            .I3(byte_transmit_counter[1]), .O(n21_adj_4359));   // verilog/coms.v(100[12:33])
    defparam i12042_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i29264_4_lut (.I0(n43_adj_4197), .I1(n41_adj_4196), .I2(n39_adj_4195), 
            .I3(n45644), .O(n44785));
    defparam i29264_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i30241_4_lut (.I0(n45134), .I1(n26_adj_4187), .I2(n45_adj_4198), 
            .I3(n45377), .O(n45762));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i30241_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i30440_3_lut (.I0(n46019), .I1(n88), .I2(n39_adj_4195), .I3(GND_net), 
            .O(n45961));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i30440_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i28966_3_lut_4_lut (.I0(pwm_count[3]), .I1(n873), .I2(n874), 
            .I3(pwm_count[2]), .O(n44486));   // verilog/motorControl.v(86[28:44])
    defparam i28966_3_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 i30545_4_lut (.I0(n45961), .I1(n45762), .I2(n45_adj_4198), 
            .I3(n44785), .O(n46066));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i30545_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i1_4_lut_adj_1472 (.I0(n46066), .I1(n22448), .I2(n84), .I3(n2168), 
            .O(n2192));
    defparam i1_4_lut_adj_1472.LUT_INIT = 16'hceef;
    SB_LUT4 div_11_i1394_3_lut (.I0(n2069), .I1(n6854), .I2(n2093), .I3(GND_net), 
            .O(n2168));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1394_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_11_mux_5_i18_3_lut (.I0(gearBoxRatio[17]), .I1(n58), .I2(gearBoxRatio[23]), 
            .I3(GND_net), .O(n83));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_mux_5_i18_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 div_11_i1459_3_lut (.I0(n2168), .I1(n6872), .I2(n2192), .I3(GND_net), 
            .O(n2264));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1459_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mux_22_i13_4_lut (.I0(encoder1_position[12]), .I1(displacement[12]), 
            .I2(n15_adj_3962), .I3(n15_adj_3963), .O(motor_state_23__N_27[12]));   // verilog/TinyFPGA_B.v(138[5] 141[10])
    defparam mux_22_i13_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_21_i13_3_lut (.I0(encoder0_position[12]), .I1(motor_state_23__N_27[12]), 
            .I2(n15_adj_3961), .I3(GND_net), .O(motor_state[12]));   // verilog/TinyFPGA_B.v(137[5] 141[10])
    defparam mux_21_i13_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i6_2_lut (.I0(pwm_23__N_2960[6]), .I1(\PID_CONTROLLER.result [6]), 
            .I2(GND_net), .I3(GND_net), .O(n13_adj_4014));   // verilog/motorControl.v(32[23:29])
    defparam i6_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mux_22_i14_4_lut (.I0(encoder1_position[13]), .I1(displacement[13]), 
            .I2(n15_adj_3962), .I3(n15_adj_3963), .O(motor_state_23__N_27[13]));   // verilog/TinyFPGA_B.v(138[5] 141[10])
    defparam mux_22_i14_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i20_2_lut (.I0(deadband[5]), .I1(\PID_CONTROLLER.result [5]), 
            .I2(GND_net), .I3(GND_net), .O(n11_adj_4011));   // verilog/motorControl.v(32[23:29])
    defparam i20_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mux_21_i14_3_lut (.I0(encoder0_position[13]), .I1(motor_state_23__N_27[13]), 
            .I2(n15_adj_3961), .I3(GND_net), .O(motor_state[13]));   // verilog/TinyFPGA_B.v(137[5] 141[10])
    defparam mux_21_i14_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i5_2_lut (.I0(deadband[6]), .I1(\PID_CONTROLLER.result [6]), 
            .I2(GND_net), .I3(GND_net), .O(n13_adj_4012));   // verilog/motorControl.v(32[23:29])
    defparam i5_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mux_22_i15_4_lut (.I0(encoder1_position[14]), .I1(displacement[14]), 
            .I2(n15_adj_3962), .I3(n15_adj_3963), .O(motor_state_23__N_27[14]));   // verilog/TinyFPGA_B.v(138[5] 141[10])
    defparam mux_22_i15_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_21_i15_3_lut (.I0(encoder0_position[14]), .I1(motor_state_23__N_27[14]), 
            .I2(n15_adj_3961), .I3(GND_net), .O(motor_state[14]));   // verilog/TinyFPGA_B.v(137[5] 141[10])
    defparam mux_21_i15_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10241_4_lut (.I0(r_Rx_Data), .I1(rx_data[7]), .I2(n27725), 
            .I3(n22471), .O(n23659));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i10241_4_lut.LUT_INIT = 16'hccac;
    SB_LUT4 mux_22_i20_4_lut (.I0(encoder1_position[19]), .I1(displacement[19]), 
            .I2(n15_adj_3962), .I3(n15_adj_3963), .O(motor_state_23__N_27[19]));   // verilog/TinyFPGA_B.v(138[5] 141[10])
    defparam mux_22_i20_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_21_i20_3_lut (.I0(encoder0_position[19]), .I1(motor_state_23__N_27[19]), 
            .I2(n15_adj_3961), .I3(GND_net), .O(motor_state[19]));   // verilog/TinyFPGA_B.v(137[5] 141[10])
    defparam mux_21_i20_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10728_3_lut (.I0(IntegralLimit[21]), .I1(\data_in_frame[8] [5]), 
            .I2(n23399), .I3(GND_net), .O(n24146));   // verilog/coms.v(126[12] 289[6])
    defparam i10728_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10242_4_lut (.I0(r_Rx_Data), .I1(rx_data[6]), .I2(n27725), 
            .I3(n22466), .O(n23660));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i10242_4_lut.LUT_INIT = 16'hccac;
    SB_LUT4 i10704_3_lut (.I0(gearBoxRatio[1]), .I1(\data_in_frame[19] [1]), 
            .I2(n23399), .I3(GND_net), .O(n24122));   // verilog/coms.v(126[12] 289[6])
    defparam i10704_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10662_3_lut (.I0(\data_in[2] [4]), .I1(\data_in[3] [4]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n24080));   // verilog/coms.v(126[12] 289[6])
    defparam i10662_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_22_i21_4_lut (.I0(encoder1_position[20]), .I1(displacement[20]), 
            .I2(n15_adj_3962), .I3(n15_adj_3963), .O(motor_state_23__N_27[20]));   // verilog/TinyFPGA_B.v(138[5] 141[10])
    defparam mux_22_i21_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_21_i21_3_lut (.I0(encoder0_position[20]), .I1(motor_state_23__N_27[20]), 
            .I2(n15_adj_3961), .I3(GND_net), .O(motor_state[20]));   // verilog/TinyFPGA_B.v(137[5] 141[10])
    defparam mux_21_i21_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10663_3_lut (.I0(\data_in[2] [3]), .I1(\data_in[3] [3]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n24081));   // verilog/coms.v(126[12] 289[6])
    defparam i10663_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_22_i22_4_lut (.I0(encoder1_position[21]), .I1(displacement[21]), 
            .I2(n15_adj_3962), .I3(n15_adj_3963), .O(motor_state_23__N_27[21]));   // verilog/TinyFPGA_B.v(138[5] 141[10])
    defparam mux_22_i22_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_21_i22_3_lut (.I0(encoder0_position[21]), .I1(motor_state_23__N_27[21]), 
            .I2(n15_adj_3961), .I3(GND_net), .O(motor_state[21]));   // verilog/TinyFPGA_B.v(137[5] 141[10])
    defparam mux_21_i22_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10243_4_lut (.I0(r_Rx_Data), .I1(rx_data[5]), .I2(n4_adj_3987), 
            .I3(n22471), .O(n23661));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i10243_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i10244_4_lut (.I0(r_Rx_Data), .I1(rx_data[4]), .I2(n4_adj_3987), 
            .I3(n22466), .O(n23662));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i10244_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i10245_4_lut (.I0(r_Rx_Data), .I1(rx_data[3]), .I2(n4_adj_3985), 
            .I3(n22471), .O(n23663));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i10245_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i10705_3_lut (.I0(Kd[7]), .I1(\data_in_frame[4] [7]), .I2(n23399), 
            .I3(GND_net), .O(n24123));   // verilog/coms.v(126[12] 289[6])
    defparam i10705_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10246_4_lut (.I0(r_Rx_Data), .I1(rx_data[2]), .I2(n4_adj_3985), 
            .I3(n22466), .O(n23664));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i10246_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i10247_4_lut (.I0(r_Rx_Data), .I1(rx_data[1]), .I2(n4_adj_3984), 
            .I3(n22471), .O(n23665));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i10247_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i10664_3_lut (.I0(\data_in[2] [2]), .I1(\data_in[3] [2]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n24082));   // verilog/coms.v(126[12] 289[6])
    defparam i10664_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10665_3_lut (.I0(\data_in[2] [1]), .I1(\data_in[3] [1]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n24083));   // verilog/coms.v(126[12] 289[6])
    defparam i10665_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_22_i23_4_lut (.I0(encoder1_position[22]), .I1(displacement[22]), 
            .I2(n15_adj_3962), .I3(n15_adj_3963), .O(motor_state_23__N_27[22]));   // verilog/TinyFPGA_B.v(138[5] 141[10])
    defparam mux_22_i23_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_21_i23_3_lut (.I0(encoder0_position[22]), .I1(motor_state_23__N_27[22]), 
            .I2(n15_adj_3961), .I3(GND_net), .O(motor_state[22]));   // verilog/TinyFPGA_B.v(137[5] 141[10])
    defparam mux_21_i23_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_22_i24_4_lut (.I0(encoder1_position[23]), .I1(displacement[23]), 
            .I2(n15_adj_3962), .I3(n15_adj_3963), .O(motor_state_23__N_27[23]));   // verilog/TinyFPGA_B.v(138[5] 141[10])
    defparam mux_22_i24_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_21_i24_3_lut (.I0(encoder0_position[23]), .I1(motor_state_23__N_27[23]), 
            .I2(n15_adj_3961), .I3(GND_net), .O(motor_state[23]));   // verilog/TinyFPGA_B.v(137[5] 141[10])
    defparam mux_21_i24_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 displacement_23__I_0_inv_0_i1_1_lut (.I0(encoder1_position[3]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n25_adj_3964));   // verilog/TinyFPGA_B.v(162[21:79])
    defparam displacement_23__I_0_inv_0_i1_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 displacement_23__I_0_inv_0_i2_1_lut (.I0(encoder1_position[4]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n24_adj_3965));   // verilog/TinyFPGA_B.v(162[21:79])
    defparam displacement_23__I_0_inv_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 displacement_23__I_0_inv_0_i3_1_lut (.I0(encoder1_position[5]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n23_adj_3966));   // verilog/TinyFPGA_B.v(162[21:79])
    defparam displacement_23__I_0_inv_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i10281_3_lut (.I0(encoder0_position[23]), .I1(n2277), .I2(count_enable), 
            .I3(GND_net), .O(n23699));   // quad.v(35[10] 41[6])
    defparam i10281_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10282_3_lut (.I0(encoder0_position[22]), .I1(n2278), .I2(count_enable), 
            .I3(GND_net), .O(n23700));   // quad.v(35[10] 41[6])
    defparam i10282_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10283_3_lut (.I0(encoder0_position[21]), .I1(n2279), .I2(count_enable), 
            .I3(GND_net), .O(n23701));   // quad.v(35[10] 41[6])
    defparam i10283_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10284_3_lut (.I0(encoder0_position[20]), .I1(n2280), .I2(count_enable), 
            .I3(GND_net), .O(n23702));   // quad.v(35[10] 41[6])
    defparam i10284_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10285_3_lut (.I0(encoder0_position[19]), .I1(n2281), .I2(count_enable), 
            .I3(GND_net), .O(n23703));   // quad.v(35[10] 41[6])
    defparam i10285_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10286_3_lut (.I0(encoder0_position[18]), .I1(n2282), .I2(count_enable), 
            .I3(GND_net), .O(n23704));   // quad.v(35[10] 41[6])
    defparam i10286_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10287_3_lut (.I0(encoder0_position[17]), .I1(n2283), .I2(count_enable), 
            .I3(GND_net), .O(n23705));   // quad.v(35[10] 41[6])
    defparam i10287_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10288_3_lut (.I0(encoder0_position[16]), .I1(n2284), .I2(count_enable), 
            .I3(GND_net), .O(n23706));   // quad.v(35[10] 41[6])
    defparam i10288_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10289_3_lut (.I0(encoder0_position[15]), .I1(n2285), .I2(count_enable), 
            .I3(GND_net), .O(n23707));   // quad.v(35[10] 41[6])
    defparam i10289_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10290_3_lut (.I0(encoder0_position[14]), .I1(n2286), .I2(count_enable), 
            .I3(GND_net), .O(n23708));   // quad.v(35[10] 41[6])
    defparam i10290_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10291_3_lut (.I0(encoder0_position[13]), .I1(n2287), .I2(count_enable), 
            .I3(GND_net), .O(n23709));   // quad.v(35[10] 41[6])
    defparam i10291_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10292_3_lut (.I0(encoder0_position[12]), .I1(n2288), .I2(count_enable), 
            .I3(GND_net), .O(n23710));   // quad.v(35[10] 41[6])
    defparam i10292_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10293_3_lut (.I0(encoder0_position[11]), .I1(n2289), .I2(count_enable), 
            .I3(GND_net), .O(n23711));   // quad.v(35[10] 41[6])
    defparam i10293_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10294_3_lut (.I0(encoder0_position[10]), .I1(n2290), .I2(count_enable), 
            .I3(GND_net), .O(n23712));   // quad.v(35[10] 41[6])
    defparam i10294_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10295_3_lut (.I0(encoder0_position[9]), .I1(n2291), .I2(count_enable), 
            .I3(GND_net), .O(n23713));   // quad.v(35[10] 41[6])
    defparam i10295_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10296_3_lut (.I0(encoder0_position[8]), .I1(n2292), .I2(count_enable), 
            .I3(GND_net), .O(n23714));   // quad.v(35[10] 41[6])
    defparam i10296_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10297_3_lut (.I0(encoder0_position[7]), .I1(n2293), .I2(count_enable), 
            .I3(GND_net), .O(n23715));   // quad.v(35[10] 41[6])
    defparam i10297_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10298_3_lut (.I0(encoder0_position[6]), .I1(n2294), .I2(count_enable), 
            .I3(GND_net), .O(n23716));   // quad.v(35[10] 41[6])
    defparam i10298_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10299_3_lut (.I0(encoder0_position[5]), .I1(n2295), .I2(count_enable), 
            .I3(GND_net), .O(n23717));   // quad.v(35[10] 41[6])
    defparam i10299_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10300_3_lut (.I0(encoder0_position[4]), .I1(n2296), .I2(count_enable), 
            .I3(GND_net), .O(n23718));   // quad.v(35[10] 41[6])
    defparam i10300_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10301_3_lut (.I0(encoder0_position[3]), .I1(n2297), .I2(count_enable), 
            .I3(GND_net), .O(n23719));   // quad.v(35[10] 41[6])
    defparam i10301_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10302_3_lut (.I0(encoder0_position[2]), .I1(n2298), .I2(count_enable), 
            .I3(GND_net), .O(n23720));   // quad.v(35[10] 41[6])
    defparam i10302_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10303_3_lut (.I0(encoder0_position[1]), .I1(n2299), .I2(count_enable), 
            .I3(GND_net), .O(n23721));   // quad.v(35[10] 41[6])
    defparam i10303_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 displacement_23__I_0_inv_0_i4_1_lut (.I0(encoder1_position[6]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n22_adj_3967));   // verilog/TinyFPGA_B.v(162[21:79])
    defparam displacement_23__I_0_inv_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i10305_3_lut (.I0(\PID_CONTROLLER.err_prev [31]), .I1(\PID_CONTROLLER.err [31]), 
            .I2(n41887), .I3(GND_net), .O(n23723));   // verilog/motorControl.v(38[14] 59[8])
    defparam i10305_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i10306_3_lut (.I0(\PID_CONTROLLER.err_prev [23]), .I1(\PID_CONTROLLER.err [23]), 
            .I2(n41887), .I3(GND_net), .O(n23724));   // verilog/motorControl.v(38[14] 59[8])
    defparam i10306_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i10307_3_lut (.I0(\PID_CONTROLLER.err_prev [22]), .I1(\PID_CONTROLLER.err [22]), 
            .I2(n41887), .I3(GND_net), .O(n23725));   // verilog/motorControl.v(38[14] 59[8])
    defparam i10307_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i10308_3_lut (.I0(\PID_CONTROLLER.err_prev [21]), .I1(\PID_CONTROLLER.err [21]), 
            .I2(n41887), .I3(GND_net), .O(n23726));   // verilog/motorControl.v(38[14] 59[8])
    defparam i10308_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i10309_3_lut (.I0(\PID_CONTROLLER.err_prev [20]), .I1(\PID_CONTROLLER.err [20]), 
            .I2(n41887), .I3(GND_net), .O(n23727));   // verilog/motorControl.v(38[14] 59[8])
    defparam i10309_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i10310_3_lut (.I0(\PID_CONTROLLER.err_prev [19]), .I1(\PID_CONTROLLER.err [19]), 
            .I2(n41887), .I3(GND_net), .O(n23728));   // verilog/motorControl.v(38[14] 59[8])
    defparam i10310_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i10311_3_lut (.I0(\PID_CONTROLLER.err_prev [18]), .I1(\PID_CONTROLLER.err [18]), 
            .I2(n41887), .I3(GND_net), .O(n23729));   // verilog/motorControl.v(38[14] 59[8])
    defparam i10311_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i10312_3_lut (.I0(\PID_CONTROLLER.err_prev [17]), .I1(\PID_CONTROLLER.err [17]), 
            .I2(n41887), .I3(GND_net), .O(n23730));   // verilog/motorControl.v(38[14] 59[8])
    defparam i10312_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i10313_3_lut (.I0(\PID_CONTROLLER.err_prev [16]), .I1(\PID_CONTROLLER.err [16]), 
            .I2(n41887), .I3(GND_net), .O(n23731));   // verilog/motorControl.v(38[14] 59[8])
    defparam i10313_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i10314_3_lut (.I0(\PID_CONTROLLER.err_prev [15]), .I1(\PID_CONTROLLER.err [15]), 
            .I2(n41887), .I3(GND_net), .O(n23732));   // verilog/motorControl.v(38[14] 59[8])
    defparam i10314_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i10315_3_lut (.I0(\PID_CONTROLLER.err_prev [14]), .I1(\PID_CONTROLLER.err [14]), 
            .I2(n41887), .I3(GND_net), .O(n23733));   // verilog/motorControl.v(38[14] 59[8])
    defparam i10315_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i10316_3_lut (.I0(\PID_CONTROLLER.err_prev [13]), .I1(\PID_CONTROLLER.err [13]), 
            .I2(n41887), .I3(GND_net), .O(n23734));   // verilog/motorControl.v(38[14] 59[8])
    defparam i10316_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 displacement_23__I_0_inv_0_i5_1_lut (.I0(encoder1_position[7]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n21_adj_3968));   // verilog/TinyFPGA_B.v(162[21:79])
    defparam displacement_23__I_0_inv_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i10317_3_lut (.I0(\PID_CONTROLLER.err_prev [12]), .I1(\PID_CONTROLLER.err [12]), 
            .I2(n41887), .I3(GND_net), .O(n23735));   // verilog/motorControl.v(38[14] 59[8])
    defparam i10317_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14_2_lut (.I0(pwm_23__N_2960[5]), .I1(\PID_CONTROLLER.result [5]), 
            .I2(GND_net), .I3(GND_net), .O(n11_adj_4013));   // verilog/motorControl.v(32[23:29])
    defparam i14_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i10318_3_lut (.I0(\PID_CONTROLLER.err_prev [11]), .I1(\PID_CONTROLLER.err [11]), 
            .I2(n41887), .I3(GND_net), .O(n23736));   // verilog/motorControl.v(38[14] 59[8])
    defparam i10318_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i10319_3_lut (.I0(\PID_CONTROLLER.err_prev [10]), .I1(\PID_CONTROLLER.err [10]), 
            .I2(n41887), .I3(GND_net), .O(n23737));   // verilog/motorControl.v(38[14] 59[8])
    defparam i10319_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i10320_3_lut (.I0(\PID_CONTROLLER.err_prev [9]), .I1(\PID_CONTROLLER.err [9]), 
            .I2(n41887), .I3(GND_net), .O(n23738));   // verilog/motorControl.v(38[14] 59[8])
    defparam i10320_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i10321_3_lut (.I0(\PID_CONTROLLER.err_prev [8]), .I1(\PID_CONTROLLER.err [8]), 
            .I2(n41887), .I3(GND_net), .O(n23739));   // verilog/motorControl.v(38[14] 59[8])
    defparam i10321_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i10322_3_lut (.I0(\PID_CONTROLLER.err_prev [7]), .I1(\PID_CONTROLLER.err [7]), 
            .I2(n41887), .I3(GND_net), .O(n23740));   // verilog/motorControl.v(38[14] 59[8])
    defparam i10322_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i10323_3_lut (.I0(\PID_CONTROLLER.err_prev [6]), .I1(\PID_CONTROLLER.err [6]), 
            .I2(n41887), .I3(GND_net), .O(n23741));   // verilog/motorControl.v(38[14] 59[8])
    defparam i10323_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i10324_3_lut (.I0(\PID_CONTROLLER.err_prev [5]), .I1(\PID_CONTROLLER.err [5]), 
            .I2(n41887), .I3(GND_net), .O(n23742));   // verilog/motorControl.v(38[14] 59[8])
    defparam i10324_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i10325_3_lut (.I0(\PID_CONTROLLER.err_prev [4]), .I1(\PID_CONTROLLER.err [4]), 
            .I2(n41887), .I3(GND_net), .O(n23743));   // verilog/motorControl.v(38[14] 59[8])
    defparam i10325_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i10326_3_lut (.I0(\PID_CONTROLLER.err_prev [3]), .I1(\PID_CONTROLLER.err [3]), 
            .I2(n41887), .I3(GND_net), .O(n23744));   // verilog/motorControl.v(38[14] 59[8])
    defparam i10326_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i10327_3_lut (.I0(\PID_CONTROLLER.err_prev [2]), .I1(\PID_CONTROLLER.err [2]), 
            .I2(n41887), .I3(GND_net), .O(n23745));   // verilog/motorControl.v(38[14] 59[8])
    defparam i10327_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i8_2_lut (.I0(PWMLimit[6]), .I1(\PID_CONTROLLER.result [6]), 
            .I2(GND_net), .I3(GND_net), .O(n13_adj_4016));   // verilog/motorControl.v(32[23:29])
    defparam i8_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i10328_3_lut (.I0(\PID_CONTROLLER.err_prev [1]), .I1(\PID_CONTROLLER.err [1]), 
            .I2(n41887), .I3(GND_net), .O(n23746));   // verilog/motorControl.v(38[14] 59[8])
    defparam i10328_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i17_2_lut (.I0(PWMLimit[5]), .I1(\PID_CONTROLLER.result [5]), 
            .I2(GND_net), .I3(GND_net), .O(n11_adj_4015));   // verilog/motorControl.v(32[23:29])
    defparam i17_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i10329_3_lut (.I0(PWMLimit[9]), .I1(\data_in_frame[6] [1]), 
            .I2(n23399), .I3(GND_net), .O(n23747));   // verilog/coms.v(126[12] 289[6])
    defparam i10329_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10330_3_lut (.I0(PWMLimit[8]), .I1(\data_in_frame[6] [0]), 
            .I2(n23399), .I3(GND_net), .O(n23748));   // verilog/coms.v(126[12] 289[6])
    defparam i10330_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10331_3_lut (.I0(PWMLimit[7]), .I1(\data_in_frame[7] [7]), 
            .I2(n23399), .I3(GND_net), .O(n23749));   // verilog/coms.v(126[12] 289[6])
    defparam i10331_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13818_3_lut (.I0(PWMLimit[6]), .I1(\data_in_frame[7] [6]), 
            .I2(n23399), .I3(GND_net), .O(n27220));
    defparam i13818_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 displacement_23__I_0_inv_0_i6_1_lut (.I0(encoder1_position[8]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n20_adj_3969));   // verilog/TinyFPGA_B.v(162[21:79])
    defparam displacement_23__I_0_inv_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 displacement_23__I_0_inv_0_i7_1_lut (.I0(encoder1_position[9]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n19_adj_3970));   // verilog/TinyFPGA_B.v(162[21:79])
    defparam displacement_23__I_0_inv_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i13763_3_lut (.I0(PWMLimit[5]), .I1(\data_in_frame[7] [5]), 
            .I2(n23399), .I3(GND_net), .O(n23751));
    defparam i13763_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10334_3_lut (.I0(PWMLimit[4]), .I1(\data_in_frame[7] [4]), 
            .I2(n23399), .I3(GND_net), .O(n23752));   // verilog/coms.v(126[12] 289[6])
    defparam i10334_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10335_3_lut (.I0(PWMLimit[3]), .I1(\data_in_frame[7] [3]), 
            .I2(n23399), .I3(GND_net), .O(n23753));   // verilog/coms.v(126[12] 289[6])
    defparam i10335_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10336_3_lut (.I0(PWMLimit[2]), .I1(\data_in_frame[7] [2]), 
            .I2(n23399), .I3(GND_net), .O(n23754));   // verilog/coms.v(126[12] 289[6])
    defparam i10336_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10337_3_lut (.I0(PWMLimit[1]), .I1(\data_in_frame[7] [1]), 
            .I2(n23399), .I3(GND_net), .O(n23755));   // verilog/coms.v(126[12] 289[6])
    defparam i10337_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10338_3_lut (.I0(control_mode[7]), .I1(\data_in_frame[1] [7]), 
            .I2(n23399), .I3(GND_net), .O(n23756));   // verilog/coms.v(126[12] 289[6])
    defparam i10338_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10339_3_lut (.I0(control_mode[6]), .I1(\data_in_frame[1] [6]), 
            .I2(n23399), .I3(GND_net), .O(n23757));   // verilog/coms.v(126[12] 289[6])
    defparam i10339_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10340_3_lut (.I0(control_mode[5]), .I1(\data_in_frame[1] [5]), 
            .I2(n23399), .I3(GND_net), .O(n23758));   // verilog/coms.v(126[12] 289[6])
    defparam i10340_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10341_3_lut (.I0(control_mode[4]), .I1(\data_in_frame[1] [4]), 
            .I2(n23399), .I3(GND_net), .O(n23759));   // verilog/coms.v(126[12] 289[6])
    defparam i10341_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10342_3_lut (.I0(control_mode[3]), .I1(\data_in_frame[1] [3]), 
            .I2(n23399), .I3(GND_net), .O(n23760));   // verilog/coms.v(126[12] 289[6])
    defparam i10342_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10343_3_lut (.I0(control_mode[2]), .I1(\data_in_frame[1] [2]), 
            .I2(n23399), .I3(GND_net), .O(n23761));   // verilog/coms.v(126[12] 289[6])
    defparam i10343_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10344_3_lut (.I0(control_mode[1]), .I1(\data_in_frame[1] [1]), 
            .I2(n23399), .I3(GND_net), .O(n23762));   // verilog/coms.v(126[12] 289[6])
    defparam i10344_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10345_3_lut (.I0(\data_in_frame[21] [7]), .I1(rx_data[7]), 
            .I2(n40207), .I3(GND_net), .O(n23763));   // verilog/coms.v(126[12] 289[6])
    defparam i10345_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i10346_3_lut (.I0(\data_in_frame[21] [6]), .I1(rx_data[6]), 
            .I2(n40207), .I3(GND_net), .O(n23764));   // verilog/coms.v(126[12] 289[6])
    defparam i10346_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i10347_3_lut (.I0(\data_in_frame[21] [5]), .I1(rx_data[5]), 
            .I2(n40207), .I3(GND_net), .O(n23765));   // verilog/coms.v(126[12] 289[6])
    defparam i10347_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i10348_3_lut (.I0(\data_in_frame[21] [4]), .I1(rx_data[4]), 
            .I2(n40207), .I3(GND_net), .O(n23766));   // verilog/coms.v(126[12] 289[6])
    defparam i10348_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_adj_1473 (.I0(\data_in_frame[10] [6]), .I1(\data_in_frame[13] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n22_adj_3988));   // verilog/coms.v(94[12:25])
    defparam i1_2_lut_adj_1473.LUT_INIT = 16'h6666;
    SB_LUT4 i10349_3_lut (.I0(\data_in_frame[21] [3]), .I1(rx_data[3]), 
            .I2(n40207), .I3(GND_net), .O(n23767));   // verilog/coms.v(126[12] 289[6])
    defparam i10349_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i10350_3_lut (.I0(\data_in_frame[21] [2]), .I1(rx_data[2]), 
            .I2(n40207), .I3(GND_net), .O(n23768));   // verilog/coms.v(126[12] 289[6])
    defparam i10350_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i10351_3_lut (.I0(\data_in_frame[21] [1]), .I1(rx_data[1]), 
            .I2(n40207), .I3(GND_net), .O(n23769));   // verilog/coms.v(126[12] 289[6])
    defparam i10351_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i10352_3_lut (.I0(\data_in_frame[21] [0]), .I1(rx_data[0]), 
            .I2(n40207), .I3(GND_net), .O(n23770));   // verilog/coms.v(126[12] 289[6])
    defparam i10352_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 displacement_23__I_0_inv_0_i8_1_lut (.I0(encoder1_position[10]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n18_adj_3971));   // verilog/TinyFPGA_B.v(162[21:79])
    defparam displacement_23__I_0_inv_0_i8_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 displacement_23__I_0_inv_0_i9_1_lut (.I0(encoder1_position[11]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n17_adj_3972));   // verilog/TinyFPGA_B.v(162[21:79])
    defparam displacement_23__I_0_inv_0_i9_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i10361_3_lut (.I0(\data_in_frame[19] [7]), .I1(rx_data[7]), 
            .I2(n40211), .I3(GND_net), .O(n23779));   // verilog/coms.v(126[12] 289[6])
    defparam i10361_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i10362_3_lut (.I0(\data_in_frame[19] [6]), .I1(rx_data[6]), 
            .I2(n40211), .I3(GND_net), .O(n23780));   // verilog/coms.v(126[12] 289[6])
    defparam i10362_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i10715_3_lut (.I0(Ki[4]), .I1(\data_in_frame[3] [4]), .I2(n23399), 
            .I3(GND_net), .O(n24133));   // verilog/coms.v(126[12] 289[6])
    defparam i10715_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10363_3_lut (.I0(\data_in_frame[19] [5]), .I1(rx_data[5]), 
            .I2(n40211), .I3(GND_net), .O(n23781));   // verilog/coms.v(126[12] 289[6])
    defparam i10363_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i10716_3_lut (.I0(Ki[3]), .I1(\data_in_frame[3] [3]), .I2(n23399), 
            .I3(GND_net), .O(n24134));   // verilog/coms.v(126[12] 289[6])
    defparam i10716_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10364_3_lut (.I0(\data_in_frame[19] [4]), .I1(rx_data[4]), 
            .I2(n40211), .I3(GND_net), .O(n23782));   // verilog/coms.v(126[12] 289[6])
    defparam i10364_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i10717_3_lut (.I0(Ki[2]), .I1(\data_in_frame[3] [2]), .I2(n23399), 
            .I3(GND_net), .O(n24135));   // verilog/coms.v(126[12] 289[6])
    defparam i10717_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10365_3_lut (.I0(\data_in_frame[19] [3]), .I1(rx_data[3]), 
            .I2(n40211), .I3(GND_net), .O(n23783));   // verilog/coms.v(126[12] 289[6])
    defparam i10365_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 displacement_23__I_0_inv_0_i10_1_lut (.I0(encoder1_position[12]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n16_adj_3973));   // verilog/TinyFPGA_B.v(162[21:79])
    defparam displacement_23__I_0_inv_0_i10_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 displacement_23__I_0_inv_0_i11_1_lut (.I0(encoder1_position[13]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n15_adj_3974));   // verilog/TinyFPGA_B.v(162[21:79])
    defparam displacement_23__I_0_inv_0_i11_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 displacement_23__I_0_inv_0_i12_1_lut (.I0(encoder1_position[14]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n14_adj_3975));   // verilog/TinyFPGA_B.v(162[21:79])
    defparam displacement_23__I_0_inv_0_i12_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 displacement_23__I_0_inv_0_i13_1_lut (.I0(encoder1_position[15]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n13_adj_3976));   // verilog/TinyFPGA_B.v(162[21:79])
    defparam displacement_23__I_0_inv_0_i13_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i10366_3_lut (.I0(\data_in_frame[19] [2]), .I1(rx_data[2]), 
            .I2(n40211), .I3(GND_net), .O(n23784));   // verilog/coms.v(126[12] 289[6])
    defparam i10366_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i10809_4_lut (.I0(pwm_23__N_2957), .I1(n44117), .I2(PWMLimit[9]), 
            .I3(n387), .O(n24227));   // verilog/motorControl.v(38[14] 59[8])
    defparam i10809_4_lut.LUT_INIT = 16'ha088;
    SB_LUT4 i10811_3_lut (.I0(quadA_debounced), .I1(reg_B[1]), .I2(n41998), 
            .I3(GND_net), .O(n24229));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(186[9] 190[16])
    defparam i10811_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i31359_4_lut (.I0(r_SM_Main[2]), .I1(n44133), .I2(n44134), 
            .I3(r_SM_Main[1]), .O(n28263));
    defparam i31359_4_lut.LUT_INIT = 16'h0511;
    SB_LUT4 i4_4_lut (.I0(control_mode[3]), .I1(control_mode[5]), .I2(control_mode[4]), 
            .I3(control_mode[7]), .O(n10_adj_4356));   // verilog/TinyFPGA_B.v(137[5:22])
    defparam i4_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i10813_3_lut (.I0(quadA_debounced_adj_3990), .I1(reg_B_adj_4406[1]), 
            .I2(n41767), .I3(GND_net), .O(n24231));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(186[9] 190[16])
    defparam i10813_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i5_3_lut_adj_1474 (.I0(control_mode[6]), .I1(n10_adj_4356), 
            .I2(control_mode[2]), .I3(GND_net), .O(n22371));   // verilog/TinyFPGA_B.v(137[5:22])
    defparam i5_3_lut_adj_1474.LUT_INIT = 16'hfefe;
    SB_LUT4 displacement_23__I_0_inv_0_i14_1_lut (.I0(encoder1_position[16]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n12_adj_3977));   // verilog/TinyFPGA_B.v(162[21:79])
    defparam displacement_23__I_0_inv_0_i14_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 displacement_23__I_0_inv_0_i15_1_lut (.I0(encoder1_position[17]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n11_adj_3978));   // verilog/TinyFPGA_B.v(162[21:79])
    defparam displacement_23__I_0_inv_0_i15_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 displacement_23__I_0_inv_0_i16_1_lut (.I0(encoder1_position[18]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n10_adj_3979));   // verilog/TinyFPGA_B.v(162[21:79])
    defparam displacement_23__I_0_inv_0_i16_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 displacement_23__I_0_inv_0_i17_1_lut (.I0(encoder1_position[19]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n9_adj_3980));   // verilog/TinyFPGA_B.v(162[21:79])
    defparam displacement_23__I_0_inv_0_i17_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 displacement_23__I_0_inv_0_i18_1_lut (.I0(encoder1_position[20]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n8_adj_3981));   // verilog/TinyFPGA_B.v(162[21:79])
    defparam displacement_23__I_0_inv_0_i18_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 displacement_23__I_0_inv_0_i19_1_lut (.I0(encoder1_position[21]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n7_adj_3982));   // verilog/TinyFPGA_B.v(162[21:79])
    defparam displacement_23__I_0_inv_0_i19_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i10240_4_lut (.I0(n23560), .I1(r_Bit_Index[1]), .I2(r_Bit_Index[0]), 
            .I3(n23471), .O(n23658));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i10240_4_lut.LUT_INIT = 16'h1444;
    SB_LUT4 displacement_23__I_0_inv_0_i20_1_lut (.I0(encoder1_position[22]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n6_adj_3983));   // verilog/TinyFPGA_B.v(162[21:79])
    defparam displacement_23__I_0_inv_0_i20_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 displacement_23__I_0_inv_0_i24_1_lut (.I0(encoder1_position[23]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n3_adj_4000));   // verilog/TinyFPGA_B.v(162[21:79])
    defparam displacement_23__I_0_inv_0_i24_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i10367_3_lut (.I0(\data_in_frame[19] [1]), .I1(rx_data[1]), 
            .I2(n40211), .I3(GND_net), .O(n23785));   // verilog/coms.v(126[12] 289[6])
    defparam i10367_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i10819_3_lut (.I0(setpoint[1]), .I1(n3793), .I2(n23430), .I3(GND_net), 
            .O(n24237));   // verilog/coms.v(126[12] 289[6])
    defparam i10819_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10820_3_lut (.I0(setpoint[2]), .I1(n3794), .I2(n23430), .I3(GND_net), 
            .O(n24238));   // verilog/coms.v(126[12] 289[6])
    defparam i10820_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10821_3_lut (.I0(setpoint[3]), .I1(n3795), .I2(n23430), .I3(GND_net), 
            .O(n24239));   // verilog/coms.v(126[12] 289[6])
    defparam i10821_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10822_3_lut (.I0(setpoint[4]), .I1(n3796), .I2(n23430), .I3(GND_net), 
            .O(n24240));   // verilog/coms.v(126[12] 289[6])
    defparam i10822_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10823_3_lut (.I0(setpoint[5]), .I1(n3797), .I2(n23430), .I3(GND_net), 
            .O(n24241));   // verilog/coms.v(126[12] 289[6])
    defparam i10823_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10824_3_lut (.I0(setpoint[6]), .I1(n3798), .I2(n23430), .I3(GND_net), 
            .O(n24242));   // verilog/coms.v(126[12] 289[6])
    defparam i10824_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10825_3_lut (.I0(setpoint[7]), .I1(n3799), .I2(n23430), .I3(GND_net), 
            .O(n24243));   // verilog/coms.v(126[12] 289[6])
    defparam i10825_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10826_3_lut (.I0(setpoint[8]), .I1(n3800), .I2(n23430), .I3(GND_net), 
            .O(n24244));   // verilog/coms.v(126[12] 289[6])
    defparam i10826_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10827_3_lut (.I0(setpoint[9]), .I1(n3801), .I2(n23430), .I3(GND_net), 
            .O(n24245));   // verilog/coms.v(126[12] 289[6])
    defparam i10827_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10828_3_lut (.I0(setpoint[10]), .I1(n3802), .I2(n23430), 
            .I3(GND_net), .O(n24246));   // verilog/coms.v(126[12] 289[6])
    defparam i10828_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10829_3_lut (.I0(setpoint[11]), .I1(n3803), .I2(n23430), 
            .I3(GND_net), .O(n24247));   // verilog/coms.v(126[12] 289[6])
    defparam i10829_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10830_3_lut (.I0(setpoint[12]), .I1(n3804), .I2(n23430), 
            .I3(GND_net), .O(n24248));   // verilog/coms.v(126[12] 289[6])
    defparam i10830_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10831_3_lut (.I0(setpoint[13]), .I1(n3805), .I2(n23430), 
            .I3(GND_net), .O(n24249));   // verilog/coms.v(126[12] 289[6])
    defparam i10831_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10832_3_lut (.I0(setpoint[14]), .I1(n3806), .I2(n23430), 
            .I3(GND_net), .O(n24250));   // verilog/coms.v(126[12] 289[6])
    defparam i10832_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10833_3_lut (.I0(setpoint[15]), .I1(n3807), .I2(n23430), 
            .I3(GND_net), .O(n24251));   // verilog/coms.v(126[12] 289[6])
    defparam i10833_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10834_3_lut (.I0(setpoint[16]), .I1(n3808), .I2(n23430), 
            .I3(GND_net), .O(n24252));   // verilog/coms.v(126[12] 289[6])
    defparam i10834_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10835_3_lut (.I0(setpoint[17]), .I1(n3809), .I2(n23430), 
            .I3(GND_net), .O(n24253));   // verilog/coms.v(126[12] 289[6])
    defparam i10835_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10836_3_lut (.I0(setpoint[18]), .I1(n3810), .I2(n23430), 
            .I3(GND_net), .O(n24254));   // verilog/coms.v(126[12] 289[6])
    defparam i10836_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10837_3_lut (.I0(setpoint[19]), .I1(n3811), .I2(n23430), 
            .I3(GND_net), .O(n24255));   // verilog/coms.v(126[12] 289[6])
    defparam i10837_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10838_3_lut (.I0(setpoint[20]), .I1(n3812), .I2(n23430), 
            .I3(GND_net), .O(n24256));   // verilog/coms.v(126[12] 289[6])
    defparam i10838_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2_3_lut (.I0(control_mode[0]), .I1(control_mode[1]), .I2(n22371), 
            .I3(GND_net), .O(n15_adj_3962));   // verilog/TinyFPGA_B.v(138[5:22])
    defparam i2_3_lut.LUT_INIT = 16'hfdfd;
    SB_LUT4 i10839_3_lut (.I0(setpoint[21]), .I1(n3813), .I2(n23430), 
            .I3(GND_net), .O(n24257));   // verilog/coms.v(126[12] 289[6])
    defparam i10839_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10840_3_lut (.I0(setpoint[22]), .I1(n3814), .I2(n23430), 
            .I3(GND_net), .O(n24258));   // verilog/coms.v(126[12] 289[6])
    defparam i10840_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10841_3_lut (.I0(setpoint[23]), .I1(n3815), .I2(n23430), 
            .I3(GND_net), .O(n24259));   // verilog/coms.v(126[12] 289[6])
    defparam i10841_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10842_3_lut (.I0(deadband[1]), .I1(\data_in_frame[13] [1]), 
            .I2(n23399), .I3(GND_net), .O(n24260));   // verilog/coms.v(126[12] 289[6])
    defparam i10842_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10237_4_lut (.I0(n23560), .I1(r_Bit_Index[2]), .I2(n4012), 
            .I3(n23471), .O(n23655));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i10237_4_lut.LUT_INIT = 16'h1444;
    SB_LUT4 i10844_3_lut (.I0(deadband[2]), .I1(\data_in_frame[13] [2]), 
            .I2(n23399), .I3(GND_net), .O(n24262));   // verilog/coms.v(126[12] 289[6])
    defparam i10844_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10845_3_lut (.I0(deadband[3]), .I1(\data_in_frame[13] [3]), 
            .I2(n23399), .I3(GND_net), .O(n24263));   // verilog/coms.v(126[12] 289[6])
    defparam i10845_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10846_3_lut (.I0(deadband[4]), .I1(\data_in_frame[13] [4]), 
            .I2(n23399), .I3(GND_net), .O(n24264));   // verilog/coms.v(126[12] 289[6])
    defparam i10846_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13764_3_lut (.I0(deadband[5]), .I1(\data_in_frame[13] [5]), 
            .I2(n23399), .I3(GND_net), .O(n24265));
    defparam i13764_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13813_3_lut (.I0(deadband[6]), .I1(\data_in_frame[13] [6]), 
            .I2(n23399), .I3(GND_net), .O(n24266));
    defparam i13813_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10849_3_lut (.I0(deadband[7]), .I1(\data_in_frame[13] [7]), 
            .I2(n23399), .I3(GND_net), .O(n24267));   // verilog/coms.v(126[12] 289[6])
    defparam i10849_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10850_3_lut (.I0(deadband[8]), .I1(\data_in_frame[12] [0]), 
            .I2(n23399), .I3(GND_net), .O(n24268));   // verilog/coms.v(126[12] 289[6])
    defparam i10850_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10851_3_lut (.I0(deadband[9]), .I1(\data_in_frame[12] [1]), 
            .I2(n23399), .I3(GND_net), .O(n24269));   // verilog/coms.v(126[12] 289[6])
    defparam i10851_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10234_4_lut (.I0(n23562), .I1(r_Bit_Index_adj_4399[1]), .I2(r_Bit_Index_adj_4399[0]), 
            .I3(n23477), .O(n23652));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i10234_4_lut.LUT_INIT = 16'h1444;
    SB_LUT4 i10231_4_lut (.I0(n23562), .I1(r_Bit_Index_adj_4399[2]), .I2(n4034), 
            .I3(n23477), .O(n23649));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i10231_4_lut.LUT_INIT = 16'h1444;
    SB_LUT4 i10227_4_lut (.I0(n23644), .I1(r_Clock_Count_adj_4398[1]), .I2(n320), 
            .I3(r_SM_Main_adj_4397[2]), .O(n23645));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i10227_4_lut.LUT_INIT = 16'h88a0;
    SB_LUT4 i10224_4_lut (.I0(n23644), .I1(r_Clock_Count_adj_4398[2]), .I2(n319), 
            .I3(r_SM_Main_adj_4397[2]), .O(n23642));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i10224_4_lut.LUT_INIT = 16'h88a0;
    SB_LUT4 i10221_4_lut (.I0(n23644), .I1(r_Clock_Count_adj_4398[3]), .I2(n318), 
            .I3(r_SM_Main_adj_4397[2]), .O(n23639));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i10221_4_lut.LUT_INIT = 16'h88a0;
    SB_LUT4 i10218_4_lut (.I0(n23644), .I1(r_Clock_Count_adj_4398[4]), .I2(n317), 
            .I3(r_SM_Main_adj_4397[2]), .O(n23636));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i10218_4_lut.LUT_INIT = 16'h88a0;
    SB_LUT4 i10215_4_lut (.I0(n23644), .I1(r_Clock_Count_adj_4398[5]), .I2(n316), 
            .I3(r_SM_Main_adj_4397[2]), .O(n23633));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i10215_4_lut.LUT_INIT = 16'h88a0;
    SB_LUT4 i10212_4_lut (.I0(n23644), .I1(r_Clock_Count_adj_4398[6]), .I2(n315), 
            .I3(r_SM_Main_adj_4397[2]), .O(n23630));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i10212_4_lut.LUT_INIT = 16'h88a0;
    SB_LUT4 i10209_4_lut (.I0(n23644), .I1(r_Clock_Count_adj_4398[7]), .I2(n314), 
            .I3(r_SM_Main_adj_4397[2]), .O(n23627));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i10209_4_lut.LUT_INIT = 16'h88a0;
    SB_LUT4 i10206_4_lut (.I0(n23644), .I1(r_Clock_Count_adj_4398[8]), .I2(n313), 
            .I3(r_SM_Main_adj_4397[2]), .O(n23624));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i10206_4_lut.LUT_INIT = 16'h88a0;
    SB_LUT4 i10368_3_lut (.I0(\data_in_frame[19] [0]), .I1(rx_data[0]), 
            .I2(n40211), .I3(GND_net), .O(n23786));   // verilog/coms.v(126[12] 289[6])
    defparam i10368_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i10377_3_lut (.I0(\data_in_frame[17] [7]), .I1(rx_data[7]), 
            .I2(n40209), .I3(GND_net), .O(n23795));   // verilog/coms.v(126[12] 289[6])
    defparam i10377_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i10378_3_lut (.I0(\data_in_frame[17] [6]), .I1(rx_data[6]), 
            .I2(n40209), .I3(GND_net), .O(n23796));   // verilog/coms.v(126[12] 289[6])
    defparam i10378_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i10379_3_lut (.I0(\data_in_frame[17] [5]), .I1(rx_data[5]), 
            .I2(n40209), .I3(GND_net), .O(n23797));   // verilog/coms.v(126[12] 289[6])
    defparam i10379_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i10380_3_lut (.I0(\data_in_frame[17] [4]), .I1(rx_data[4]), 
            .I2(n40209), .I3(GND_net), .O(n23798));   // verilog/coms.v(126[12] 289[6])
    defparam i10380_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i10381_3_lut (.I0(\data_in_frame[17] [3]), .I1(rx_data[3]), 
            .I2(n40209), .I3(GND_net), .O(n23799));   // verilog/coms.v(126[12] 289[6])
    defparam i10381_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i10382_3_lut (.I0(\data_in_frame[17] [2]), .I1(rx_data[2]), 
            .I2(n40209), .I3(GND_net), .O(n23800));   // verilog/coms.v(126[12] 289[6])
    defparam i10382_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i10383_3_lut (.I0(\data_in_frame[17] [1]), .I1(rx_data[1]), 
            .I2(n40209), .I3(GND_net), .O(n23801));   // verilog/coms.v(126[12] 289[6])
    defparam i10383_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i10666_3_lut (.I0(\data_in[2] [0]), .I1(\data_in[3] [0]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n24084));   // verilog/coms.v(126[12] 289[6])
    defparam i10666_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10384_3_lut (.I0(\data_in_frame[17] [0]), .I1(rx_data[0]), 
            .I2(n40209), .I3(GND_net), .O(n23802));   // verilog/coms.v(126[12] 289[6])
    defparam i10384_3_lut.LUT_INIT = 16'hacac;
    pll32MHz pll32MHz_inst (.GND_net(GND_net), .CLK_c(CLK_c), .VCC_net(VCC_net), 
            .clk32MHz(clk32MHz)) /* synthesis lattice_noprune=1, syn_preserve=0, syn_module_defined=1, syn_noprune=0 */ ;   // verilog/TinyFPGA_B.v(35[12] 38[39])
    SB_LUT4 i1_2_lut_3_lut (.I0(control_mode[0]), .I1(n22371), .I2(control_mode[1]), 
            .I3(GND_net), .O(n15_adj_3961));   // verilog/TinyFPGA_B.v(137[5:22])
    defparam i1_2_lut_3_lut.LUT_INIT = 16'hfefe;
    coms setpoint_23__I_0 (.clk32MHz(clk32MHz), .n24165(n24165), .IntegralLimit({IntegralLimit}), 
         .GND_net(GND_net), .n24164(n24164), .n24163(n24163), .n24117(n24117), 
         .gearBoxRatio({gearBoxRatio}), .n24116(n24116), .n24115(n24115), 
         .n24114(n24114), .n24113(n24113), .n24112(n24112), .n24111(n24111), 
         .n24110(n24110), .\data_in_frame[5] ({\data_in_frame[5] }), .\data_in_frame[3] ({\data_in_frame[3] }), 
         .n22338(n22338), .pwm({pwm}), .n24109(n24109), .n24108(n24108), 
         .n24107(n24107), .n24106(n24106), .n24105(n24105), .encoder0_position({encoder0_position}), 
         .n24104(n24104), .n24103(n24103), .n24102(n24102), .n24101(n24101), 
         .n24100(n24100), .n24099(n24099), .\data_in[0] ({\data_in[0] }), 
         .n24098(n24098), .n24097(n24097), .n24096(n24096), .n24095(n24095), 
         .n24094(n24094), .n24093(n24093), .n24092(n24092), .\data_in[1] ({\data_in[1] }), 
         .n24091(n24091), .encoder1_position({encoder1_position}), .n24269(n24269), 
         .\deadband[9] (deadband[9]), .n24268(n24268), .\deadband[8] (deadband[8]), 
         .n24267(n24267), .\deadband[7] (deadband[7]), .n24266(n24266), 
         .\deadband[6] (deadband[6]), .n24265(n24265), .\deadband[5] (deadband[5]), 
         .n24264(n24264), .\deadband[4] (deadband[4]), .n24263(n24263), 
         .\deadband[3] (deadband[3]), .n24262(n24262), .\deadband[2] (deadband[2]), 
         .n24260(n24260), .\deadband[1] (deadband[1]), .n24259(n24259), 
         .setpoint({setpoint}), .n24258(n24258), .n24257(n24257), .n24256(n24256), 
         .n24255(n24255), .n24254(n24254), .n24253(n24253), .n24252(n24252), 
         .n24251(n24251), .n24250(n24250), .n24249(n24249), .n24248(n24248), 
         .n24247(n24247), .n24246(n24246), .n24245(n24245), .n24244(n24244), 
         .n24243(n24243), .n24242(n24242), .n24241(n24241), .n24240(n24240), 
         .n24239(n24239), .n24238(n24238), .n24237(n24237), .VCC_net(VCC_net), 
         .byte_transmit_counter({Open_0, Open_1, Open_2, Open_3, Open_4, 
         Open_5, byte_transmit_counter[1:0]}), .n24169(n24169), .n24168(n24168), 
         .n24167(n24167), .n24166(n24166), .n24079(n24079), .\data_in[2] ({\data_in[2] }), 
         .n24078(n24078), .n24077(n24077), .n24076(n24076), .\data_in[3] ({\data_in[3] }), 
         .n24075(n24075), .n24074(n24074), .n24073(n24073), .n24072(n24072), 
         .n24071(n24071), .n24070(n24070), .n24069(n24069), .n24068(n24068), 
         .\data_out_frame[0][2] (\data_out_frame[0] [2]), .n24067(n24067), 
         .\data_out_frame[0][3] (\data_out_frame[0] [3]), .n24066(n24066), 
         .\data_out_frame[0][4] (\data_out_frame[0] [4]), .n24063(n24063), 
         .\data_out_frame[5][2] (\data_out_frame[5] [2]), .n24132(n24132), 
         .\Ki[5] (Ki[5]), .n24131(n24131), .\Ki[6] (Ki[6]), .n24130(n24130), 
         .\Ki[7] (Ki[7]), .n24129(n24129), .\Kd[1] (Kd[1]), .n24128(n24128), 
         .\Kd[2] (Kd[2]), .n24127(n24127), .\Kd[3] (Kd[3]), .n24126(n24126), 
         .\Kd[4] (Kd[4]), .\data_in_frame[9] ({\data_in_frame[9] }), .\data_in_frame[7] ({\data_in_frame[7] }), 
         .n24125(n24125), .\Kd[5] (Kd[5]), .n24090(n24090), .n24089(n24089), 
         .n24088(n24088), .n24087(n24087), .n40207(n40207), .rx_data_ready(rx_data_ready), 
         .displacement({displacement}), .n24086(n24086), .n24137(n24137), 
         .\Kp[7] (Kp[7]), .n24136(n24136), .\Ki[1] (Ki[1]), .n24124(n24124), 
         .\Kd[6] (Kd[6]), .n24085(n24085), .n24162(n24162), .n24161(n24161), 
         .n24160(n24160), .n24159(n24159), .n24158(n24158), .\data_out_frame[18][3] (\data_out_frame[18] [3]), 
         .\data_in_frame[8] ({\data_in_frame[8] }), .rx_data({rx_data}), 
         .\data_out_frame[19][3] (\data_out_frame[19] [3]), .n24157(n24157), 
         .\data_out_frame[20][7] (\data_out_frame[20] [7]), .n24156(n24156), 
         .n23930(n23930), .\data_in_frame[1] ({\data_in_frame[1] }), .n23929(n23929), 
         .n23928(n23928), .n23927(n23927), .n23926(n23926), .\data_in_frame[6][1] (\data_in_frame[6] [1]), 
         .\data_in_frame[6][0] (\data_in_frame[6] [0]), .n23925(n23925), 
         .n23924(n23924), .n23923(n23923), .\data_in_frame[13] ({\data_in_frame[13] }), 
         .\data_in_frame[2] ({\data_in_frame[2] }), .n23914(n23914), .n24155(n24155), 
         .n23913(n23913), .n23912(n23912), .n23911(n23911), .n23910(n23910), 
         .n23909(n23909), .n23908(n23908), .n23907(n23907), .\data_in_frame[4] ({\data_in_frame[4] }), 
         .n23898(n23898), .n23897(n23897), .n23896(n23896), .\data_in_frame[10] ({\data_in_frame[10] }), 
         .n23895(n23895), .n23894(n23894), .n23893(n23893), .n23892(n23892), 
         .n23891(n23891), .\data_in_frame[12][1] (\data_in_frame[12] [1]), 
         .\data_in_frame[12][0] (\data_in_frame[12] [0]), .n24151(n24151), 
         .n23866(n23866), .n23865(n23865), .n23864(n23864), .n23863(n23863), 
         .n23862(n23862), .n23861(n23861), .n23860(n23860), .n23859(n23859), 
         .n23850(n23850), .\data_in_frame[11] ({\data_in_frame[11] }), .n23849(n23849), 
         .n23848(n23848), .n23847(n23847), .n23846(n23846), .n23845(n23845), 
         .n23844(n23844), .n23843(n23843), .n24150(n24150), .n24149(n24149), 
         .n17(n17_adj_4358), .\data_in_frame[19] ({\data_in_frame[19] }), 
         .n40227(n40227), .n24148(n24148), .n24147(n24147), .n23834(n23834), 
         .\data_in_frame[18] ({\data_in_frame[18] }), .n23833(n23833), .n23832(n23832), 
         .n23831(n23831), .n23830(n23830), .n23829(n23829), .n23828(n23828), 
         .n23827(n23827), .\data_in_frame[21] ({\data_in_frame[21] }), .\data_in_frame[17] ({\data_in_frame[17] }), 
         .n23802(n23802), .n24084(n24084), .n23801(n23801), .n23800(n23800), 
         .n23799(n23799), .n23798(n23798), .n23797(n23797), .n23796(n23796), 
         .n23795(n23795), .n23786(n23786), .\data_out_frame[22][7] (\data_out_frame[22] [7]), 
         .\data_out_frame[21][7] (\data_out_frame[21] [7]), .n23785(n23785), 
         .n23784(n23784), .n23783(n23783), .n24135(n24135), .\Ki[2] (Ki[2]), 
         .n23782(n23782), .n24134(n24134), .\Ki[3] (Ki[3]), .n23781(n23781), 
         .n24133(n24133), .\Ki[4] (Ki[4]), .n23780(n23780), .n23779(n23779), 
         .n23770(n23770), .n23769(n23769), .n23768(n23768), .n23767(n23767), 
         .n23766(n23766), .n23765(n23765), .n23764(n23764), .n23763(n23763), 
         .n23762(n23762), .control_mode({control_mode}), .n23761(n23761), 
         .n23760(n23760), .n23759(n23759), .n23758(n23758), .n23757(n23757), 
         .n23756(n23756), .n23755(n23755), .\PWMLimit[1] (PWMLimit[1]), 
         .n23754(n23754), .\PWMLimit[2] (PWMLimit[2]), .n23753(n23753), 
         .\PWMLimit[3] (PWMLimit[3]), .n23752(n23752), .\PWMLimit[4] (PWMLimit[4]), 
         .n23751(n23751), .\PWMLimit[5] (PWMLimit[5]), .n27220(n27220), 
         .\PWMLimit[6] (PWMLimit[6]), .n23749(n23749), .\PWMLimit[7] (PWMLimit[7]), 
         .n23748(n23748), .\PWMLimit[8] (PWMLimit[8]), .n23747(n23747), 
         .\PWMLimit[9] (PWMLimit[9]), .n24083(n24083), .n24082(n24082), 
         .n24123(n24123), .\Kd[7] (Kd[7]), .n24081(n24081), .n24080(n24080), 
         .n24122(n24122), .n24146(n24146), .n24145(n24145), .n24144(n24144), 
         .n24143(n24143), .\Kp[1] (Kp[1]), .n24142(n24142), .\Kp[2] (Kp[2]), 
         .n24141(n24141), .\Kp[3] (Kp[3]), .n24140(n24140), .\Kp[4] (Kp[4]), 
         .n24139(n24139), .\Kp[5] (Kp[5]), .n24138(n24138), .\Kp[6] (Kp[6]), 
         .LED_c(LED_c), .n24121(n24121), .n24120(n24120), .n24119(n24119), 
         .n24118(n24118), .n23600(n23600), .\deadband[0] (deadband[0]), 
         .n23599(n23599), .n23588(n23588), .\PWMLimit[0] (PWMLimit[0]), 
         .n23587(n23587), .n23585(n23585), .n23584(n23584), .n23583(n23583), 
         .\Kd[0] (Kd[0]), .n23582(n23582), .\Ki[0] (Ki[0]), .n23581(n23581), 
         .\Kp[0] (Kp[0]), .n23580(n23580), .n5019(n5019), .n23458(n23458), 
         .n40218(n40218), .n21(n21_adj_4359), .Kp_23__N_516(Kp_23__N_516), 
         .n22(n22_adj_3988), .n3792(n3792), .n3793(n3793), .n23430(n23430), 
         .n3794(n3794), .n3795(n3795), .n3796(n3796), .n3797(n3797), 
         .n3798(n3798), .n3799(n3799), .n3800(n3800), .n3801(n3801), 
         .n3802(n3802), .n3803(n3803), .n3804(n3804), .n3805(n3805), 
         .n3806(n3806), .n3807(n3807), .n3808(n3808), .n3809(n3809), 
         .n3810(n3810), .n3811(n3811), .n3812(n3812), .n3813(n3813), 
         .n3815(n3815), .n3814(n3814), .n40209(n40209), .n40222(n40222), 
         .n40213(n40213), .n23399(n23399), .n40216(n40216), .n40225(n40225), 
         .n40211(n40211), .n313(n313), .\r_Clock_Count[8] (r_Clock_Count_adj_4398[8]), 
         .n314(n314), .\r_Clock_Count[7] (r_Clock_Count_adj_4398[7]), .n23624(n23624), 
         .n23627(n23627), .n23630(n23630), .\r_Clock_Count[6] (r_Clock_Count_adj_4398[6]), 
         .n23633(n23633), .\r_Clock_Count[5] (r_Clock_Count_adj_4398[5]), 
         .n23636(n23636), .\r_Clock_Count[4] (r_Clock_Count_adj_4398[4]), 
         .n23639(n23639), .\r_Clock_Count[3] (r_Clock_Count_adj_4398[3]), 
         .n23642(n23642), .\r_Clock_Count[2] (r_Clock_Count_adj_4398[2]), 
         .n23645(n23645), .\r_Clock_Count[1] (r_Clock_Count_adj_4398[1]), 
         .n23649(n23649), .r_Bit_Index({r_Bit_Index_adj_4399}), .n23652(n23652), 
         .n23695(n23695), .n315(n315), .n316(n316), .n317(n317), .n318(n318), 
         .n319(n319), .n320(n320), .n23644(n23644), .\r_SM_Main[2] (r_SM_Main_adj_4397[2]), 
         .tx_o(tx_o), .tx_enable(tx_enable), .n23477(n23477), .n23562(n23562), 
         .n4034(n4034), .r_Rx_Data(r_Rx_Data), .\r_SM_Main[2]_adj_3 (r_SM_Main[2]), 
         .\r_SM_Main[1] (r_SM_Main[1]), .n23655(n23655), .r_Bit_Index_adj_9({r_Bit_Index}), 
         .n23658(n23658), .n28263(n28263), .n23698(n23698), .n24171(n24171), 
         .PIN_13_N_26(PIN_13_N_26), .n23665(n23665), .n23664(n23664), 
         .n23663(n23663), .n23662(n23662), .n23661(n23661), .n23660(n23660), 
         .n23659(n23659), .n23594(n23594), .n22466(n22466), .n4(n4_adj_3984), 
         .n28231(n28231), .n1(n1_adj_4357), .n27725(n27725), .n4_adj_7(n4_adj_3987), 
         .n4_adj_8(n4_adj_3985), .n22471(n22471), .n44134(n44134), .n44133(n44133), 
         .n23471(n23471), .n23560(n23560), .n4012(n4012)) /* synthesis lattice_noprune=1, syn_preserve=0, syn_module_defined=1, syn_noprune=0 */ ;   // verilog/TinyFPGA_B.v(68[8] 88[4])
    SB_LUT4 i1_2_lut_3_lut_adj_1475 (.I0(control_mode[0]), .I1(n22371), 
            .I2(control_mode[1]), .I3(GND_net), .O(n15_adj_3963));   // verilog/TinyFPGA_B.v(137[5:22])
    defparam i1_2_lut_3_lut_adj_1475.LUT_INIT = 16'hefef;
    SB_LUT4 i1_2_lut_3_lut_4_lut (.I0(n90), .I1(n89), .I2(n88), .I3(n22436), 
            .O(n22427));
    defparam i1_2_lut_3_lut_4_lut.LUT_INIT = 16'hff7f;
    SB_LUT4 div_11_i107_1_lut_4_lut (.I0(n558), .I1(n99), .I2(n224), .I3(n22403), 
            .O(n249));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i107_1_lut_4_lut.LUT_INIT = 16'h00c8;
    SB_LUT4 div_11_LessThan_1482_i18_3_lut_3_lut (.I0(n98), .I1(n97), .I2(n2278_adj_4003), 
            .I3(GND_net), .O(n18_adj_4201));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1482_i18_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 i29240_2_lut_4_lut (.I0(n2273), .I1(n92), .I2(n2277_adj_4002), 
            .I3(n96), .O(n44761));
    defparam i29240_2_lut_4_lut.LUT_INIT = 16'hf99f;
    SB_LUT4 mux_22_i16_4_lut (.I0(encoder1_position[15]), .I1(displacement[15]), 
            .I2(n15_adj_3962), .I3(n15_adj_3963), .O(motor_state_23__N_27[15]));   // verilog/TinyFPGA_B.v(138[5] 141[10])
    defparam mux_22_i16_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 div_11_LessThan_1482_i20_3_lut_3_lut (.I0(n96), .I1(n92), .I2(n2273), 
            .I3(GND_net), .O(n20_adj_4203));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1482_i20_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 div_11_LessThan_1482_i22_3_lut_3_lut (.I0(n95), .I1(n94), .I2(n2275), 
            .I3(GND_net), .O(n22_adj_4205));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1482_i22_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 i29248_2_lut_4_lut (.I0(n2275), .I1(n94), .I2(n2276), .I3(n95), 
            .O(n44769));
    defparam i29248_2_lut_4_lut.LUT_INIT = 16'hf99f;
    SB_LUT4 div_11_LessThan_1545_i16_3_lut_3_lut (.I0(n98), .I1(n97), .I2(n2372), 
            .I3(GND_net), .O(n16_adj_4219));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1545_i16_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 i29200_2_lut_4_lut (.I0(n2367), .I1(n92), .I2(n2371), .I3(n96), 
            .O(n44721));
    defparam i29200_2_lut_4_lut.LUT_INIT = 16'hf99f;
    SB_LUT4 div_11_LessThan_1545_i18_3_lut_3_lut (.I0(n96), .I1(n92), .I2(n2367), 
            .I3(GND_net), .O(n18_adj_4221));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1545_i18_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 div_11_LessThan_1545_i20_3_lut_3_lut (.I0(n95), .I1(n94), .I2(n2369), 
            .I3(GND_net), .O(n20_adj_4223));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1545_i20_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 i29173_2_lut_4_lut (.I0(n2359), .I1(n84), .I2(n2368), .I3(n93), 
            .O(n44694));
    defparam i29173_2_lut_4_lut.LUT_INIT = 16'hf99f;
    SB_LUT4 div_11_LessThan_1545_i22_3_lut_3_lut (.I0(n93), .I1(n84), .I2(n2359), 
            .I3(GND_net), .O(n22_adj_4225));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1545_i22_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 div_11_LessThan_1606_i14_3_lut_3_lut (.I0(n98), .I1(n97), .I2(n2463), 
            .I3(GND_net), .O(n14_adj_4241));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1606_i14_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 i29157_2_lut_4_lut (.I0(n2458), .I1(n92), .I2(n2462), .I3(n96), 
            .O(n44678));
    defparam i29157_2_lut_4_lut.LUT_INIT = 16'hf99f;
    SB_LUT4 div_11_LessThan_1606_i16_3_lut_3_lut (.I0(n96), .I1(n92), .I2(n2458), 
            .I3(GND_net), .O(n16_adj_4243));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1606_i16_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 div_11_LessThan_1606_i18_3_lut_3_lut (.I0(n95), .I1(n94), .I2(n2460), 
            .I3(GND_net), .O(n18_adj_4245));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1606_i18_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 i29133_2_lut_4_lut (.I0(n2450), .I1(n84), .I2(n2459), .I3(n93), 
            .O(n44654));
    defparam i29133_2_lut_4_lut.LUT_INIT = 16'hf99f;
    SB_LUT4 div_11_LessThan_1606_i20_3_lut_3_lut (.I0(n93), .I1(n84), .I2(n2450), 
            .I3(GND_net), .O(n20_adj_4247));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1606_i20_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 div_11_LessThan_1665_i12_3_lut_3_lut (.I0(n98), .I1(n97), .I2(n2551), 
            .I3(GND_net), .O(n12_adj_4263));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1665_i12_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 i29113_2_lut_4_lut (.I0(n2546), .I1(n92), .I2(n2550), .I3(n96), 
            .O(n44634));
    defparam i29113_2_lut_4_lut.LUT_INIT = 16'hf99f;
    SB_LUT4 div_11_LessThan_1665_i14_3_lut_3_lut (.I0(n96), .I1(n92), .I2(n2546), 
            .I3(GND_net), .O(n14_adj_4265));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1665_i14_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 div_11_LessThan_1665_i16_3_lut_3_lut (.I0(n95), .I1(n94), .I2(n2548), 
            .I3(GND_net), .O(n16_adj_4267));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1665_i16_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 i29095_2_lut_4_lut (.I0(n2538), .I1(n84), .I2(n2547), .I3(n93), 
            .O(n44616));
    defparam i29095_2_lut_4_lut.LUT_INIT = 16'hf99f;
    SB_LUT4 i10409_3_lut (.I0(\data_in_frame[13] [7]), .I1(rx_data[7]), 
            .I2(n40227), .I3(GND_net), .O(n23827));   // verilog/coms.v(126[12] 289[6])
    defparam i10409_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i10410_3_lut (.I0(\data_in_frame[13] [6]), .I1(rx_data[6]), 
            .I2(n40227), .I3(GND_net), .O(n23828));   // verilog/coms.v(126[12] 289[6])
    defparam i10410_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i10411_3_lut (.I0(\data_in_frame[13] [5]), .I1(rx_data[5]), 
            .I2(n40227), .I3(GND_net), .O(n23829));   // verilog/coms.v(126[12] 289[6])
    defparam i10411_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i10412_3_lut (.I0(\data_in_frame[13] [4]), .I1(rx_data[4]), 
            .I2(n40227), .I3(GND_net), .O(n23830));   // verilog/coms.v(126[12] 289[6])
    defparam i10412_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i10413_3_lut (.I0(\data_in_frame[13] [3]), .I1(rx_data[3]), 
            .I2(n40227), .I3(GND_net), .O(n23831));   // verilog/coms.v(126[12] 289[6])
    defparam i10413_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i10414_3_lut (.I0(\data_in_frame[13] [2]), .I1(rx_data[2]), 
            .I2(n40227), .I3(GND_net), .O(n23832));   // verilog/coms.v(126[12] 289[6])
    defparam i10414_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i10415_3_lut (.I0(\data_in_frame[13] [1]), .I1(rx_data[1]), 
            .I2(n40227), .I3(GND_net), .O(n23833));   // verilog/coms.v(126[12] 289[6])
    defparam i10415_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_11_LessThan_1665_i18_3_lut_3_lut (.I0(n93), .I1(n84), .I2(n2538), 
            .I3(GND_net), .O(n18_adj_4269));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1665_i18_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 i10416_3_lut (.I0(\data_in_frame[13] [0]), .I1(rx_data[0]), 
            .I2(n40227), .I3(GND_net), .O(n23834));   // verilog/coms.v(126[12] 289[6])
    defparam i10416_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_11_LessThan_1722_i10_3_lut_3_lut (.I0(n98), .I1(n97), .I2(n2636), 
            .I3(GND_net), .O(n10_adj_4285));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1722_i10_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 div_11_LessThan_1722_i14_3_lut_3_lut (.I0(n95), .I1(n94), .I2(n2633), 
            .I3(GND_net), .O(n14_adj_4289));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1722_i14_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 i28942_2_lut_4_lut (.I0(n2623), .I1(n84), .I2(n2632), .I3(n93), 
            .O(n44462));
    defparam i28942_2_lut_4_lut.LUT_INIT = 16'hf99f;
    SB_LUT4 div_11_LessThan_1722_i16_3_lut_3_lut (.I0(n93), .I1(n84), .I2(n2623), 
            .I3(GND_net), .O(n16_adj_4291));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1722_i16_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 div_11_LessThan_1722_i12_3_lut_3_lut (.I0(n96), .I1(n92), .I2(n2631), 
            .I3(GND_net), .O(n12_adj_4287));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1722_i12_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 i10729_3_lut (.I0(IntegralLimit[20]), .I1(\data_in_frame[8] [4]), 
            .I2(n23399), .I3(GND_net), .O(n24147));   // verilog/coms.v(126[12] 289[6])
    defparam i10729_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10730_3_lut (.I0(IntegralLimit[19]), .I1(\data_in_frame[8] [3]), 
            .I2(n23399), .I3(GND_net), .O(n24148));   // verilog/coms.v(126[12] 289[6])
    defparam i10730_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_11_LessThan_1830_i41_4_lut (.I0(n2702), .I1(n80), .I2(n7004), 
            .I3(n2724), .O(n41_adj_4353));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1830_i41_4_lut.LUT_INIT = 16'hc399;
    SB_LUT4 div_11_LessThan_1830_i39_4_lut (.I0(n2703), .I1(n81), .I2(n7005), 
            .I3(n2724), .O(n39_adj_4351));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1830_i39_4_lut.LUT_INIT = 16'hc399;
    SB_LUT4 div_11_mux_3_i1_3_lut (.I0(encoder0_position[0]), .I1(n25), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n391));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_mux_3_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_11_LessThan_1830_i45_4_lut (.I0(n2700), .I1(n78), .I2(n7002), 
            .I3(n2724), .O(n45_adj_4355));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1830_i45_4_lut.LUT_INIT = 16'hc399;
    SB_LUT4 div_11_LessThan_1830_i43_4_lut (.I0(n2701), .I1(n79), .I2(n7003), 
            .I3(n2724), .O(n43_adj_4354));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1830_i43_4_lut.LUT_INIT = 16'hc399;
    SB_LUT4 div_11_LessThan_1830_i37_4_lut (.I0(n2704), .I1(n82), .I2(n7006), 
            .I3(n2724), .O(n37_adj_4350));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1830_i37_4_lut.LUT_INIT = 16'hc399;
    SB_LUT4 div_11_LessThan_1830_i29_4_lut (.I0(n2708), .I1(n86), .I2(n7010), 
            .I3(n2724), .O(n29_adj_4345));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1830_i29_4_lut.LUT_INIT = 16'hc399;
    SB_LUT4 div_11_LessThan_1830_i31_4_lut (.I0(n2707), .I1(n85), .I2(n7009), 
            .I3(n2724), .O(n31_adj_4347));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1830_i31_4_lut.LUT_INIT = 16'hc399;
    SB_LUT4 div_11_LessThan_1830_i9_4_lut (.I0(n2718), .I1(n96), .I2(n7020), 
            .I3(n2724), .O(n9_adj_4331));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1830_i9_4_lut.LUT_INIT = 16'hc399;
    SB_LUT4 div_11_LessThan_1830_i21_4_lut (.I0(n2712), .I1(n90), .I2(n7014), 
            .I3(n2724), .O(n21_adj_4340));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1830_i21_4_lut.LUT_INIT = 16'hc399;
    SB_LUT4 div_11_LessThan_1830_i23_4_lut (.I0(n2711), .I1(n89), .I2(n7013), 
            .I3(n2724), .O(n23_adj_4341));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1830_i23_4_lut.LUT_INIT = 16'hc399;
    SB_LUT4 div_11_LessThan_1830_i25_4_lut (.I0(n2710), .I1(n88), .I2(n7012), 
            .I3(n2724), .O(n25_adj_4343));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1830_i25_4_lut.LUT_INIT = 16'hc399;
    SB_LUT4 div_11_LessThan_1830_i7_4_lut (.I0(n2719), .I1(n97), .I2(n7021), 
            .I3(n2724), .O(n7_adj_4329));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1830_i7_4_lut.LUT_INIT = 16'hc399;
    SB_LUT4 div_11_LessThan_1830_i35_4_lut (.I0(n2705), .I1(n83), .I2(n7007), 
            .I3(n2724), .O(n35_adj_4349));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1830_i35_4_lut.LUT_INIT = 16'hc399;
    SB_LUT4 div_11_LessThan_1830_i17_4_lut (.I0(n2714), .I1(n92), .I2(n7016), 
            .I3(n2724), .O(n17_adj_4338));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1830_i17_4_lut.LUT_INIT = 16'hc399;
    SB_LUT4 div_11_LessThan_1830_i19_4_lut (.I0(n2713), .I1(n91), .I2(n7015), 
            .I3(n2724), .O(n19_adj_4339));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1830_i19_4_lut.LUT_INIT = 16'hc399;
    SB_LUT4 div_11_LessThan_1830_i11_4_lut (.I0(n2717), .I1(n95), .I2(n7019), 
            .I3(n2724), .O(n11_adj_4333));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1830_i11_4_lut.LUT_INIT = 16'hc399;
    SB_LUT4 div_11_LessThan_1830_i13_4_lut (.I0(n2716), .I1(n94), .I2(n7018), 
            .I3(n2724), .O(n13_adj_4335));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1830_i13_4_lut.LUT_INIT = 16'hc399;
    SB_LUT4 div_11_LessThan_1830_i27_4_lut (.I0(n2709), .I1(n87), .I2(n7011), 
            .I3(n2724), .O(n27_adj_4344));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1830_i27_4_lut.LUT_INIT = 16'hc399;
    SB_LUT4 div_11_LessThan_1830_i15_4_lut (.I0(n2715), .I1(n93), .I2(n7017), 
            .I3(n2724), .O(n15_adj_4336));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1830_i15_4_lut.LUT_INIT = 16'hc399;
    SB_LUT4 div_11_LessThan_1830_i33_4_lut (.I0(n2706), .I1(n84), .I2(n7008), 
            .I3(n2724), .O(n33_adj_4348));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1830_i33_4_lut.LUT_INIT = 16'hc399;
    SB_LUT4 div_11_i1832_1_lut (.I0(n2801), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n2802));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1832_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i28734_4_lut (.I0(n27_adj_4344), .I1(n15_adj_4336), .I2(n13_adj_4335), 
            .I3(n11_adj_4333), .O(n44253));
    defparam i28734_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 div_11_LessThan_1830_i12_3_lut (.I0(n93), .I1(n84), .I2(n33_adj_4348), 
            .I3(GND_net), .O(n12_adj_4334));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1830_i12_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 i28724_2_lut (.I0(n33_adj_4348), .I1(n15_adj_4336), .I2(GND_net), 
            .I3(GND_net), .O(n44243));
    defparam i28724_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 div_11_LessThan_1830_i10_3_lut (.I0(n95), .I1(n94), .I2(n13_adj_4335), 
            .I3(GND_net), .O(n10_adj_4332));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1830_i10_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 div_11_LessThan_1830_i30_3_lut (.I0(n12_adj_4334), .I1(n83), 
            .I2(n35_adj_4349), .I3(GND_net), .O(n30_adj_4346));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1830_i30_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 div_11_i1828_3_lut (.I0(n2720), .I1(n7022), .I2(n2724), .I3(GND_net), 
            .O(n2798));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1828_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i28768_3_lut (.I0(n7_adj_4329), .I1(n2798), .I2(n98), .I3(GND_net), 
            .O(n44287));
    defparam i28768_3_lut.LUT_INIT = 16'hebeb;
    SB_LUT4 i29452_4_lut (.I0(n13_adj_4335), .I1(n11_adj_4333), .I2(n9_adj_4331), 
            .I3(n44287), .O(n44973));
    defparam i29452_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i29443_4_lut (.I0(n19_adj_4339), .I1(n17_adj_4338), .I2(n15_adj_4336), 
            .I3(n44973), .O(n44964));
    defparam i29443_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i30399_4_lut (.I0(n25_adj_4343), .I1(n23_adj_4341), .I2(n21_adj_4340), 
            .I3(n44964), .O(n45920));
    defparam i30399_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i29923_4_lut (.I0(n31_adj_4347), .I1(n29_adj_4345), .I2(n27_adj_4344), 
            .I3(n45920), .O(n45444));
    defparam i29923_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i30529_4_lut (.I0(n37_adj_4350), .I1(n35_adj_4349), .I2(n33_adj_4348), 
            .I3(n45444), .O(n46050));
    defparam i30529_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 div_11_LessThan_1830_i16_3_lut (.I0(n91), .I1(n79), .I2(n43_adj_4354), 
            .I3(GND_net), .O(n16_adj_4337));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1830_i16_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 div_11_LessThan_1830_i6_3_lut (.I0(n98), .I1(n97), .I2(n7_adj_4329), 
            .I3(GND_net), .O(n6_adj_4328));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1830_i6_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 i30327_3_lut (.I0(n6_adj_4328), .I1(n90), .I2(n21_adj_4340), 
            .I3(GND_net), .O(n45848));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i30327_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i30328_3_lut (.I0(n45848), .I1(n89), .I2(n23_adj_4341), .I3(GND_net), 
            .O(n45849));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i30328_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i28749_4_lut (.I0(n21_adj_4340), .I1(n19_adj_4339), .I2(n17_adj_4338), 
            .I3(n9_adj_4331), .O(n44268));
    defparam i28749_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i28678_2_lut (.I0(n43_adj_4354), .I1(n19_adj_4339), .I2(GND_net), 
            .I3(GND_net), .O(n44197));
    defparam i28678_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 div_11_LessThan_1830_i8_3_lut (.I0(n96), .I1(n92), .I2(n17_adj_4338), 
            .I3(GND_net), .O(n8_adj_4330));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1830_i8_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 div_11_LessThan_1830_i24_3_lut (.I0(n16_adj_4337), .I1(n78), 
            .I2(n45_adj_4355), .I3(GND_net), .O(n24_adj_4342));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1830_i24_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i28692_4_lut (.I0(n43_adj_4354), .I1(n25_adj_4343), .I2(n23_adj_4341), 
            .I3(n44268), .O(n44211));
    defparam i28692_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i30275_4_lut (.I0(n24_adj_4342), .I1(n8_adj_4330), .I2(n45_adj_4355), 
            .I3(n44197), .O(n45796));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i30275_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i30270_3_lut (.I0(n45849), .I1(n88), .I2(n25_adj_4343), .I3(GND_net), 
            .O(n45791));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i30270_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 div_11_i1829_3_lut (.I0(n390), .I1(n7023), .I2(n2724), .I3(GND_net), 
            .O(n2799));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1829_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_11_LessThan_1830_i4_4_lut (.I0(n391), .I1(n99), .I2(n2799), 
            .I3(n558), .O(n4_adj_4327));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1830_i4_4_lut.LUT_INIT = 16'h0317;
    SB_LUT4 i30325_3_lut (.I0(n4_adj_4327), .I1(n87), .I2(n27_adj_4344), 
            .I3(GND_net), .O(n45846));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i30325_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i30326_3_lut (.I0(n45846), .I1(n86), .I2(n29_adj_4345), .I3(GND_net), 
            .O(n45847));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i30326_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i28728_4_lut (.I0(n33_adj_4348), .I1(n31_adj_4347), .I2(n29_adj_4345), 
            .I3(n44253), .O(n44247));
    defparam i28728_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i30580_4_lut (.I0(n30_adj_4346), .I1(n10_adj_4332), .I2(n35_adj_4349), 
            .I3(n44243), .O(n46101));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i30580_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i30272_3_lut (.I0(n45847), .I1(n85), .I2(n31_adj_4347), .I3(GND_net), 
            .O(n45793));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i30272_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i30669_4_lut (.I0(n45793), .I1(n46101), .I2(n35_adj_4349), 
            .I3(n44247), .O(n46190));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i30669_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i30670_3_lut (.I0(n46190), .I1(n82), .I2(n37_adj_4350), .I3(GND_net), 
            .O(n46191));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i30670_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i30626_3_lut (.I0(n46191), .I1(n81), .I2(n39_adj_4351), .I3(GND_net), 
            .O(n46147));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i30626_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i28698_4_lut (.I0(n43_adj_4354), .I1(n41_adj_4353), .I2(n39_adj_4351), 
            .I3(n46050), .O(n44217));
    defparam i28698_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i30449_4_lut (.I0(n45791), .I1(n45796), .I2(n45_adj_4355), 
            .I3(n44211), .O(n45970));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i30449_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i30616_3_lut (.I0(n46147), .I1(n80), .I2(n41_adj_4353), .I3(GND_net), 
            .O(n40_adj_4352));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i30616_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 div_11_i1807_3_lut (.I0(n2699), .I1(n7001), .I2(n2724), .I3(GND_net), 
            .O(n2777));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1807_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i30451_4_lut (.I0(n40_adj_4352), .I1(n45970), .I2(n45_adj_4355), 
            .I3(n44217), .O(n45972));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i30451_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i30452_3_lut (.I0(n45972), .I1(n77), .I2(n2777), .I3(GND_net), 
            .O(n2801));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i30452_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i29030_2_lut_4_lut (.I0(n2631), .I1(n92), .I2(n2635), .I3(n96), 
            .O(n44550));
    defparam i29030_2_lut_4_lut.LUT_INIT = 16'hf99f;
    SB_LUT4 div_11_LessThan_1777_i8_3_lut_3_lut (.I0(n98), .I1(n97), .I2(n2718), 
            .I3(GND_net), .O(n8_adj_4307));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1777_i8_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 div_11_LessThan_1777_i12_3_lut_3_lut (.I0(n95), .I1(n94), .I2(n2715), 
            .I3(GND_net), .O(n12_adj_4311));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1777_i12_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 i28793_2_lut_4_lut (.I0(n2705), .I1(n84), .I2(n2714), .I3(n93), 
            .O(n44312));
    defparam i28793_2_lut_4_lut.LUT_INIT = 16'hf99f;
    SB_LUT4 div_11_LessThan_1777_i14_3_lut_3_lut (.I0(n93), .I1(n84), .I2(n2705), 
            .I3(GND_net), .O(n14_adj_4313));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1777_i14_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 div_11_LessThan_1777_i10_3_lut_3_lut (.I0(n96), .I1(n92), .I2(n2713), 
            .I3(GND_net), .O(n10_adj_4309));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1777_i10_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 i28846_2_lut_4_lut (.I0(n2713), .I1(n92), .I2(n2717), .I3(n96), 
            .O(n44365));
    defparam i28846_2_lut_4_lut.LUT_INIT = 16'hf99f;
    SB_LUT4 div_11_LessThan_1777_i33_2_lut (.I0(n2706), .I1(n85), .I2(GND_net), 
            .I3(GND_net), .O(n33_adj_4324));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1777_i33_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_11_LessThan_1777_i31_2_lut (.I0(n2707), .I1(n86), .I2(GND_net), 
            .I3(GND_net), .O(n31_adj_4322));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1777_i31_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_11_LessThan_1777_i37_2_lut (.I0(n2704), .I1(n83), .I2(GND_net), 
            .I3(GND_net), .O(n37_adj_4326));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1777_i37_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_11_LessThan_1777_i35_2_lut (.I0(n2705), .I1(n84), .I2(GND_net), 
            .I3(GND_net), .O(n35_adj_4325));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1777_i35_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_11_mux_3_i2_3_lut (.I0(encoder0_position[1]), .I1(n24), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n390));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_mux_3_i2_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_11_LessThan_1777_i25_2_lut (.I0(n2710), .I1(n89), .I2(GND_net), 
            .I3(GND_net), .O(n25_adj_4319));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1777_i25_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_11_LessThan_1777_i27_2_lut (.I0(n2709), .I1(n88), .I2(GND_net), 
            .I3(GND_net), .O(n27_adj_4320));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1777_i27_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_11_LessThan_1777_i21_2_lut (.I0(n2712), .I1(n91), .I2(GND_net), 
            .I3(GND_net), .O(n21_adj_4317));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1777_i21_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_11_LessThan_1777_i23_2_lut (.I0(n2711), .I1(n90), .I2(GND_net), 
            .I3(GND_net), .O(n23_adj_4318));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1777_i23_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_11_LessThan_1777_i9_2_lut (.I0(n2718), .I1(n97), .I2(GND_net), 
            .I3(GND_net), .O(n9_adj_4308));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1777_i9_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_11_LessThan_1777_i11_2_lut (.I0(n2717), .I1(n96), .I2(GND_net), 
            .I3(GND_net), .O(n11_adj_4310));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1777_i11_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_11_LessThan_1777_i19_2_lut (.I0(n2713), .I1(n92), .I2(GND_net), 
            .I3(GND_net), .O(n19_adj_4316));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1777_i19_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_11_LessThan_1777_i13_2_lut (.I0(n2716), .I1(n95), .I2(GND_net), 
            .I3(GND_net), .O(n13_adj_4312));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1777_i13_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_11_LessThan_1777_i15_2_lut (.I0(n2715), .I1(n94), .I2(GND_net), 
            .I3(GND_net), .O(n15_adj_4314));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1777_i15_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_11_LessThan_1777_i17_2_lut (.I0(n2714), .I1(n93), .I2(GND_net), 
            .I3(GND_net), .O(n17_adj_4315));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1777_i17_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_11_LessThan_1777_i29_2_lut (.I0(n2708), .I1(n87), .I2(GND_net), 
            .I3(GND_net), .O(n29_adj_4321));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1777_i29_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_11_i1779_1_lut (.I0(n2723), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n2724));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1779_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i28813_4_lut (.I0(n29_adj_4321), .I1(n17_adj_4315), .I2(n15_adj_4314), 
            .I3(n13_adj_4312), .O(n44332));
    defparam i28813_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i29520_4_lut (.I0(n11_adj_4310), .I1(n9_adj_4308), .I2(n2719), 
            .I3(n98), .O(n45041));
    defparam i29520_4_lut.LUT_INIT = 16'hfeef;
    SB_LUT4 i29959_4_lut (.I0(n17_adj_4315), .I1(n15_adj_4314), .I2(n13_adj_4312), 
            .I3(n45041), .O(n45480));
    defparam i29959_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i29957_4_lut (.I0(n23_adj_4318), .I1(n21_adj_4317), .I2(n19_adj_4316), 
            .I3(n45480), .O(n45478));
    defparam i29957_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i28821_4_lut (.I0(n29_adj_4321), .I1(n27_adj_4320), .I2(n25_adj_4319), 
            .I3(n45478), .O(n44340));
    defparam i28821_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 div_11_LessThan_1777_i6_4_lut (.I0(n390), .I1(n99), .I2(n2720), 
            .I3(n558), .O(n6_adj_4306));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1777_i6_4_lut.LUT_INIT = 16'h0317;
    SB_LUT4 i30333_3_lut (.I0(n6_adj_4306), .I1(n87), .I2(n29_adj_4321), 
            .I3(GND_net), .O(n45854));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i30333_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 div_11_LessThan_1777_i32_3_lut (.I0(n14_adj_4313), .I1(n83), 
            .I2(n37_adj_4326), .I3(GND_net), .O(n32_adj_4323));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1777_i32_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i30334_3_lut (.I0(n45854), .I1(n86), .I2(n31_adj_4322), .I3(GND_net), 
            .O(n45855));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i30334_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i28799_4_lut (.I0(n35_adj_4325), .I1(n33_adj_4324), .I2(n31_adj_4322), 
            .I3(n44332), .O(n44318));
    defparam i28799_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i30578_4_lut (.I0(n32_adj_4323), .I1(n12_adj_4311), .I2(n37_adj_4326), 
            .I3(n44312), .O(n46099));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i30578_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i30262_3_lut (.I0(n45855), .I1(n85), .I2(n33_adj_4324), .I3(GND_net), 
            .O(n45783));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i30262_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i30335_3_lut (.I0(n8_adj_4307), .I1(n90), .I2(n23_adj_4318), 
            .I3(GND_net), .O(n45856));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i30335_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i30336_3_lut (.I0(n45856), .I1(n89), .I2(n25_adj_4319), .I3(GND_net), 
            .O(n45857));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i30336_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i29500_4_lut (.I0(n25_adj_4319), .I1(n23_adj_4318), .I2(n21_adj_4317), 
            .I3(n44365), .O(n45021));
    defparam i29500_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i30259_3_lut (.I0(n10_adj_4309), .I1(n91), .I2(n21_adj_4317), 
            .I3(GND_net), .O(n45780));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i30259_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i30258_3_lut (.I0(n45857), .I1(n88), .I2(n27_adj_4320), .I3(GND_net), 
            .O(n45779));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i30258_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i30169_4_lut (.I0(n35_adj_4325), .I1(n33_adj_4324), .I2(n31_adj_4322), 
            .I3(n44340), .O(n45690));
    defparam i30169_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i30667_4_lut (.I0(n45783), .I1(n46099), .I2(n37_adj_4326), 
            .I3(n44318), .O(n46188));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i30667_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i30329_4_lut (.I0(n45779), .I1(n45780), .I2(n27_adj_4320), 
            .I3(n45021), .O(n45850));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i30329_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i30681_4_lut (.I0(n45850), .I1(n46188), .I2(n37_adj_4326), 
            .I3(n45690), .O(n46202));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i30681_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i30682_3_lut (.I0(n46202), .I1(n82), .I2(n2703), .I3(GND_net), 
            .O(n46203));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i30682_3_lut.LUT_INIT = 16'h2b2b;
    SB_LUT4 i30676_3_lut (.I0(n46203), .I1(n81), .I2(n2702), .I3(GND_net), 
            .O(n46197));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i30676_3_lut.LUT_INIT = 16'h2b2b;
    SB_LUT4 i30523_3_lut (.I0(n46197), .I1(n80), .I2(n2701), .I3(GND_net), 
            .O(n46044));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i30523_3_lut.LUT_INIT = 16'h2b2b;
    SB_LUT4 i30524_3_lut (.I0(n46044), .I1(n79), .I2(n2700), .I3(GND_net), 
            .O(n46045));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i30524_3_lut.LUT_INIT = 16'h2b2b;
    SB_LUT4 i1806_4_lut (.I0(n46045), .I1(n77), .I2(n78), .I3(n2699), 
            .O(n2723));
    defparam i1806_4_lut.LUT_INIT = 16'hceef;
    SB_LUT4 div_11_LessThan_1722_i35_2_lut (.I0(n2624), .I1(n85), .I2(GND_net), 
            .I3(GND_net), .O(n35_adj_4303));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1722_i35_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_11_LessThan_1722_i39_2_lut (.I0(n2622), .I1(n83), .I2(GND_net), 
            .I3(GND_net), .O(n39_adj_4305));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1722_i39_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_11_LessThan_1722_i33_2_lut (.I0(n2625), .I1(n86), .I2(GND_net), 
            .I3(GND_net), .O(n33_adj_4301));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1722_i33_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_11_mux_3_i3_3_lut (.I0(encoder0_position[2]), .I1(n23), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n389));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_mux_3_i3_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_11_LessThan_1722_i37_2_lut (.I0(n2623), .I1(n84), .I2(GND_net), 
            .I3(GND_net), .O(n37_adj_4304));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1722_i37_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_11_LessThan_1722_i27_2_lut (.I0(n2628), .I1(n89), .I2(GND_net), 
            .I3(GND_net), .O(n27_adj_4298));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1722_i27_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_11_LessThan_1722_i29_2_lut (.I0(n2627), .I1(n88), .I2(GND_net), 
            .I3(GND_net), .O(n29_adj_4299));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1722_i29_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_11_LessThan_1722_i23_2_lut (.I0(n2630), .I1(n91), .I2(GND_net), 
            .I3(GND_net), .O(n23_adj_4296));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1722_i23_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_11_LessThan_1722_i25_2_lut (.I0(n2629), .I1(n90), .I2(GND_net), 
            .I3(GND_net), .O(n25_adj_4297));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1722_i25_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_11_LessThan_1722_i11_2_lut (.I0(n2636), .I1(n97), .I2(GND_net), 
            .I3(GND_net), .O(n11_adj_4286));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1722_i11_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_11_LessThan_1722_i13_2_lut (.I0(n2635), .I1(n96), .I2(GND_net), 
            .I3(GND_net), .O(n13_adj_4288));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1722_i13_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_11_LessThan_1722_i21_2_lut (.I0(n2631), .I1(n92), .I2(GND_net), 
            .I3(GND_net), .O(n21_adj_4295));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1722_i21_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_11_LessThan_1722_i15_2_lut (.I0(n2634), .I1(n95), .I2(GND_net), 
            .I3(GND_net), .O(n15_adj_4290));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1722_i15_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_11_LessThan_1722_i17_2_lut (.I0(n2633), .I1(n94), .I2(GND_net), 
            .I3(GND_net), .O(n17_adj_4292));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1722_i17_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_11_LessThan_1722_i19_2_lut (.I0(n2632), .I1(n93), .I2(GND_net), 
            .I3(GND_net), .O(n19_adj_4293));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1722_i19_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_11_LessThan_1722_i31_2_lut (.I0(n2626), .I1(n87), .I2(GND_net), 
            .I3(GND_net), .O(n31_adj_4300));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1722_i31_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_11_i1724_1_lut (.I0(n2642), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n2643));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1724_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i28973_4_lut (.I0(n31_adj_4300), .I1(n19_adj_4293), .I2(n17_adj_4292), 
            .I3(n15_adj_4290), .O(n44493));
    defparam i28973_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i29694_4_lut (.I0(n13_adj_4288), .I1(n11_adj_4286), .I2(n2637), 
            .I3(n98), .O(n45215));
    defparam i29694_4_lut.LUT_INIT = 16'hfeef;
    SB_LUT4 i30009_4_lut (.I0(n19_adj_4293), .I1(n17_adj_4292), .I2(n15_adj_4290), 
            .I3(n45215), .O(n45530));
    defparam i30009_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i30005_4_lut (.I0(n25_adj_4297), .I1(n23_adj_4296), .I2(n21_adj_4295), 
            .I3(n45530), .O(n45526));
    defparam i30005_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i28997_4_lut (.I0(n31_adj_4300), .I1(n29_adj_4299), .I2(n27_adj_4298), 
            .I3(n45526), .O(n44517));
    defparam i28997_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 div_11_LessThan_1722_i8_4_lut (.I0(n389), .I1(n99), .I2(n2638), 
            .I3(n558), .O(n8_adj_4284));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1722_i8_4_lut.LUT_INIT = 16'h0317;
    SB_LUT4 i30339_3_lut (.I0(n8_adj_4284), .I1(n87), .I2(n31_adj_4300), 
            .I3(GND_net), .O(n45860));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i30339_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i30340_3_lut (.I0(n45860), .I1(n86), .I2(n33_adj_4301), .I3(GND_net), 
            .O(n45861));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i30340_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 div_11_LessThan_1722_i34_3_lut (.I0(n16_adj_4291), .I1(n83), 
            .I2(n39_adj_4305), .I3(GND_net), .O(n34_adj_4302));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1722_i34_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i28948_4_lut (.I0(n37_adj_4304), .I1(n35_adj_4303), .I2(n33_adj_4301), 
            .I3(n44493), .O(n44468));
    defparam i28948_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i30576_4_lut (.I0(n34_adj_4302), .I1(n14_adj_4289), .I2(n39_adj_4305), 
            .I3(n44462), .O(n46097));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i30576_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i30250_3_lut (.I0(n45861), .I1(n85), .I2(n35_adj_4303), .I3(GND_net), 
            .O(n45771));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i30250_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i30107_3_lut (.I0(n10_adj_4285), .I1(n90), .I2(n25_adj_4297), 
            .I3(GND_net), .O(n45628));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i30107_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i30108_3_lut (.I0(n45628), .I1(n89), .I2(n27_adj_4298), .I3(GND_net), 
            .O(n45629));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i30108_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i29660_4_lut (.I0(n27_adj_4298), .I1(n25_adj_4297), .I2(n23_adj_4296), 
            .I3(n44550), .O(n45181));
    defparam i29660_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 div_11_LessThan_1722_i20_3_lut (.I0(n12_adj_4287), .I1(n91), 
            .I2(n23_adj_4296), .I3(GND_net), .O(n20_adj_4294));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1722_i20_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i29651_3_lut (.I0(n45629), .I1(n88), .I2(n29_adj_4299), .I3(GND_net), 
            .O(n45172));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i29651_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i30195_4_lut (.I0(n37_adj_4304), .I1(n35_adj_4303), .I2(n33_adj_4301), 
            .I3(n44517), .O(n45716));
    defparam i30195_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i30665_4_lut (.I0(n45771), .I1(n46097), .I2(n39_adj_4305), 
            .I3(n44468), .O(n46186));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i30665_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i30253_4_lut (.I0(n45172), .I1(n20_adj_4294), .I2(n29_adj_4299), 
            .I3(n45181), .O(n45774));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i30253_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i30683_4_lut (.I0(n45774), .I1(n46186), .I2(n39_adj_4305), 
            .I3(n45716), .O(n46204));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i30683_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i30684_3_lut (.I0(n46204), .I1(n82), .I2(n2621), .I3(GND_net), 
            .O(n46205));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i30684_3_lut.LUT_INIT = 16'h2b2b;
    SB_LUT4 i30674_3_lut (.I0(n46205), .I1(n81), .I2(n2620), .I3(GND_net), 
            .O(n46195));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i30674_3_lut.LUT_INIT = 16'h2b2b;
    SB_LUT4 i30255_3_lut (.I0(n46195), .I1(n80), .I2(n2619), .I3(GND_net), 
            .O(n45776));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i30255_3_lut.LUT_INIT = 16'h2b2b;
    SB_LUT4 i1_4_lut_adj_1476 (.I0(n45776), .I1(n22463), .I2(n79), .I3(n2618), 
            .O(n2642));
    defparam i1_4_lut_adj_1476.LUT_INIT = 16'hceef;
    SB_LUT4 div_11_LessThan_1665_i37_2_lut (.I0(n2539), .I1(n85), .I2(GND_net), 
            .I3(GND_net), .O(n37_adj_4281));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1665_i37_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_11_LessThan_1665_i41_2_lut (.I0(n2537), .I1(n83), .I2(GND_net), 
            .I3(GND_net), .O(n41_adj_4283));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1665_i41_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_11_LessThan_1665_i35_2_lut (.I0(n2540), .I1(n86), .I2(GND_net), 
            .I3(GND_net), .O(n35_adj_4279));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1665_i35_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_11_mux_3_i4_3_lut (.I0(encoder0_position[3]), .I1(n22), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n388));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_mux_3_i4_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_11_LessThan_1665_i39_2_lut (.I0(n2538), .I1(n84), .I2(GND_net), 
            .I3(GND_net), .O(n39_adj_4282));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1665_i39_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_11_LessThan_1665_i29_2_lut (.I0(n2543), .I1(n89), .I2(GND_net), 
            .I3(GND_net), .O(n29_adj_4276));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1665_i29_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_11_LessThan_1665_i31_2_lut (.I0(n2542), .I1(n88), .I2(GND_net), 
            .I3(GND_net), .O(n31_adj_4277));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1665_i31_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_11_LessThan_1665_i23_2_lut (.I0(n2546), .I1(n92), .I2(GND_net), 
            .I3(GND_net), .O(n23_adj_4273));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1665_i23_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_11_LessThan_1665_i25_2_lut (.I0(n2545), .I1(n91), .I2(GND_net), 
            .I3(GND_net), .O(n25_adj_4274));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1665_i25_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_11_LessThan_1665_i27_2_lut (.I0(n2544), .I1(n90), .I2(GND_net), 
            .I3(GND_net), .O(n27_adj_4275));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1665_i27_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_11_LessThan_1665_i33_2_lut (.I0(n2541), .I1(n87), .I2(GND_net), 
            .I3(GND_net), .O(n33_adj_4278));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1665_i33_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_11_LessThan_1665_i17_2_lut (.I0(n2549), .I1(n95), .I2(GND_net), 
            .I3(GND_net), .O(n17_adj_4268));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1665_i17_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_11_LessThan_1665_i19_2_lut (.I0(n2548), .I1(n94), .I2(GND_net), 
            .I3(GND_net), .O(n19_adj_4270));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1665_i19_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_11_LessThan_1665_i21_2_lut (.I0(n2547), .I1(n93), .I2(GND_net), 
            .I3(GND_net), .O(n21_adj_4271));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1665_i21_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_11_LessThan_1665_i13_2_lut (.I0(n2551), .I1(n97), .I2(GND_net), 
            .I3(GND_net), .O(n13_adj_4264));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1665_i13_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_11_LessThan_1665_i15_2_lut (.I0(n2550), .I1(n96), .I2(GND_net), 
            .I3(GND_net), .O(n15_adj_4266));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1665_i15_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_11_i1667_1_lut (.I0(n2558), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n2559));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1667_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i29101_4_lut (.I0(n33_adj_4278), .I1(n21_adj_4271), .I2(n19_adj_4270), 
            .I3(n17_adj_4268), .O(n44622));
    defparam i29101_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i29738_4_lut (.I0(n15_adj_4266), .I1(n13_adj_4264), .I2(n2552), 
            .I3(n98), .O(n45259));
    defparam i29738_4_lut.LUT_INIT = 16'hfeef;
    SB_LUT4 i30029_4_lut (.I0(n21_adj_4271), .I1(n19_adj_4270), .I2(n17_adj_4268), 
            .I3(n45259), .O(n45550));
    defparam i30029_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i30027_4_lut (.I0(n27_adj_4275), .I1(n25_adj_4274), .I2(n23_adj_4273), 
            .I3(n45550), .O(n45548));
    defparam i30027_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i29105_4_lut (.I0(n33_adj_4278), .I1(n31_adj_4277), .I2(n29_adj_4276), 
            .I3(n45548), .O(n44626));
    defparam i29105_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 div_11_LessThan_1665_i10_4_lut (.I0(n388), .I1(n99), .I2(n2553), 
            .I3(n558), .O(n10_adj_4262));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1665_i10_4_lut.LUT_INIT = 16'h0317;
    SB_LUT4 i30113_3_lut (.I0(n10_adj_4262), .I1(n87), .I2(n33_adj_4278), 
            .I3(GND_net), .O(n45634));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i30113_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i30114_3_lut (.I0(n45634), .I1(n86), .I2(n35_adj_4279), .I3(GND_net), 
            .O(n45635));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i30114_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 div_11_LessThan_1665_i36_3_lut (.I0(n18_adj_4269), .I1(n83), 
            .I2(n41_adj_4283), .I3(GND_net), .O(n36_adj_4280));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1665_i36_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i29097_4_lut (.I0(n39_adj_4282), .I1(n37_adj_4281), .I2(n35_adj_4279), 
            .I3(n44622), .O(n44618));
    defparam i29097_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i30521_4_lut (.I0(n36_adj_4280), .I1(n16_adj_4267), .I2(n41_adj_4283), 
            .I3(n44616), .O(n46042));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i30521_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i29641_3_lut (.I0(n45635), .I1(n85), .I2(n37_adj_4281), .I3(GND_net), 
            .O(n45162));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i29641_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 div_11_LessThan_1665_i22_3_lut (.I0(n14_adj_4265), .I1(n91), 
            .I2(n25_adj_4274), .I3(GND_net), .O(n22_adj_4272));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1665_i22_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i30527_4_lut (.I0(n22_adj_4272), .I1(n12_adj_4263), .I2(n25_adj_4274), 
            .I3(n44634), .O(n46048));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i30527_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i30528_3_lut (.I0(n46048), .I1(n90), .I2(n27_adj_4275), .I3(GND_net), 
            .O(n46049));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i30528_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i30376_3_lut (.I0(n46049), .I1(n89), .I2(n29_adj_4276), .I3(GND_net), 
            .O(n45897));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i30376_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i30291_4_lut (.I0(n39_adj_4282), .I1(n37_adj_4281), .I2(n35_adj_4279), 
            .I3(n44626), .O(n45812));
    defparam i30291_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i30645_4_lut (.I0(n45162), .I1(n46042), .I2(n41_adj_4283), 
            .I3(n44618), .O(n46166));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i30645_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i29639_3_lut (.I0(n45897), .I1(n88), .I2(n31_adj_4277), .I3(GND_net), 
            .O(n45160));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i29639_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i30679_4_lut (.I0(n45160), .I1(n46166), .I2(n41_adj_4283), 
            .I3(n45812), .O(n46200));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i30679_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i30680_3_lut (.I0(n46200), .I1(n82), .I2(n2536), .I3(GND_net), 
            .O(n46201));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i30680_3_lut.LUT_INIT = 16'h2b2b;
    SB_LUT4 i30678_3_lut (.I0(n46201), .I1(n81), .I2(n2535), .I3(GND_net), 
            .O(n46199));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i30678_3_lut.LUT_INIT = 16'h2b2b;
    SB_LUT4 i1_4_lut_adj_1477 (.I0(n46199), .I1(n22460), .I2(n80), .I3(n2534), 
            .O(n2558));
    defparam i1_4_lut_adj_1477.LUT_INIT = 16'hceef;
    SB_LUT4 div_11_LessThan_1606_i39_2_lut (.I0(n2451), .I1(n85), .I2(GND_net), 
            .I3(GND_net), .O(n39_adj_4259));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1606_i39_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_11_LessThan_1606_i37_2_lut (.I0(n2452), .I1(n86), .I2(GND_net), 
            .I3(GND_net), .O(n37_adj_4257));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1606_i37_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_11_LessThan_1606_i43_2_lut (.I0(n2449), .I1(n83), .I2(GND_net), 
            .I3(GND_net), .O(n43_adj_4261));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1606_i43_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_11_LessThan_1606_i41_2_lut (.I0(n2450), .I1(n84), .I2(GND_net), 
            .I3(GND_net), .O(n41_adj_4260));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1606_i41_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_11_mux_3_i5_3_lut (.I0(encoder0_position[4]), .I1(n21), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n387_adj_4001));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_mux_3_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_11_LessThan_1606_i31_2_lut (.I0(n2455), .I1(n89), .I2(GND_net), 
            .I3(GND_net), .O(n31_adj_4254));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1606_i31_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_11_LessThan_1606_i33_2_lut (.I0(n2454), .I1(n88), .I2(GND_net), 
            .I3(GND_net), .O(n33_adj_4255));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1606_i33_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_11_LessThan_1606_i25_2_lut (.I0(n2458), .I1(n92), .I2(GND_net), 
            .I3(GND_net), .O(n25_adj_4251));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1606_i25_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_11_LessThan_1606_i27_2_lut (.I0(n2457), .I1(n91), .I2(GND_net), 
            .I3(GND_net), .O(n27_adj_4252));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1606_i27_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_11_LessThan_1606_i29_2_lut (.I0(n2456), .I1(n90), .I2(GND_net), 
            .I3(GND_net), .O(n29_adj_4253));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1606_i29_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_11_LessThan_1606_i15_2_lut (.I0(n2463), .I1(n97), .I2(GND_net), 
            .I3(GND_net), .O(n15_adj_4242));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1606_i15_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_11_LessThan_1606_i17_2_lut (.I0(n2462), .I1(n96), .I2(GND_net), 
            .I3(GND_net), .O(n17_adj_4244));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1606_i17_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_11_LessThan_1606_i19_2_lut (.I0(n2461), .I1(n95), .I2(GND_net), 
            .I3(GND_net), .O(n19_adj_4246));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1606_i19_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_11_LessThan_1606_i21_2_lut (.I0(n2460), .I1(n94), .I2(GND_net), 
            .I3(GND_net), .O(n21_adj_4248));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1606_i21_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_11_LessThan_1606_i23_2_lut (.I0(n2459), .I1(n93), .I2(GND_net), 
            .I3(GND_net), .O(n23_adj_4249));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1606_i23_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_11_LessThan_1606_i35_2_lut (.I0(n2453), .I1(n87), .I2(GND_net), 
            .I3(GND_net), .O(n35_adj_4256));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1606_i35_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_11_i1608_1_lut (.I0(n2471), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n2472));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1608_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i29141_4_lut (.I0(n35_adj_4256), .I1(n23_adj_4249), .I2(n21_adj_4248), 
            .I3(n19_adj_4246), .O(n44662));
    defparam i29141_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i29776_4_lut (.I0(n17_adj_4244), .I1(n15_adj_4242), .I2(n2464), 
            .I3(n98), .O(n45297));
    defparam i29776_4_lut.LUT_INIT = 16'hfeef;
    SB_LUT4 i30051_4_lut (.I0(n23_adj_4249), .I1(n21_adj_4248), .I2(n19_adj_4246), 
            .I3(n45297), .O(n45572));
    defparam i30051_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i30047_4_lut (.I0(n29_adj_4253), .I1(n27_adj_4252), .I2(n25_adj_4251), 
            .I3(n45572), .O(n45568));
    defparam i30047_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i29145_4_lut (.I0(n35_adj_4256), .I1(n33_adj_4255), .I2(n31_adj_4254), 
            .I3(n45568), .O(n44666));
    defparam i29145_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 div_11_LessThan_1606_i12_4_lut (.I0(n387_adj_4001), .I1(n99), 
            .I2(n2465), .I3(n558), .O(n12_adj_4240));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1606_i12_4_lut.LUT_INIT = 16'h0317;
    SB_LUT4 i30117_3_lut (.I0(n12_adj_4240), .I1(n87), .I2(n35_adj_4256), 
            .I3(GND_net), .O(n45638));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i30117_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 div_11_LessThan_1606_i38_3_lut (.I0(n20_adj_4247), .I1(n83), 
            .I2(n43_adj_4261), .I3(GND_net), .O(n38_adj_4258));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1606_i38_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i30118_3_lut (.I0(n45638), .I1(n86), .I2(n37_adj_4257), .I3(GND_net), 
            .O(n45639));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i30118_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i29135_4_lut (.I0(n41_adj_4260), .I1(n39_adj_4259), .I2(n37_adj_4257), 
            .I3(n44662), .O(n44656));
    defparam i29135_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i30495_4_lut (.I0(n38_adj_4258), .I1(n18_adj_4245), .I2(n43_adj_4261), 
            .I3(n44654), .O(n46016));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i30495_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i29635_3_lut (.I0(n45639), .I1(n85), .I2(n39_adj_4259), .I3(GND_net), 
            .O(n45156));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i29635_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 div_11_LessThan_1606_i24_3_lut (.I0(n16_adj_4243), .I1(n91), 
            .I2(n27_adj_4252), .I3(GND_net), .O(n24_adj_4250));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1606_i24_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i30519_4_lut (.I0(n24_adj_4250), .I1(n14_adj_4241), .I2(n27_adj_4252), 
            .I3(n44678), .O(n46040));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i30519_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i30520_3_lut (.I0(n46040), .I1(n90), .I2(n29_adj_4253), .I3(GND_net), 
            .O(n46041));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i30520_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i30380_3_lut (.I0(n46041), .I1(n89), .I2(n31_adj_4254), .I3(GND_net), 
            .O(n45901));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i30380_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i30301_4_lut (.I0(n41_adj_4260), .I1(n39_adj_4259), .I2(n37_adj_4257), 
            .I3(n44666), .O(n45822));
    defparam i30301_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i30631_4_lut (.I0(n45156), .I1(n46016), .I2(n43_adj_4261), 
            .I3(n44656), .O(n46152));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i30631_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i29633_3_lut (.I0(n45901), .I1(n88), .I2(n33_adj_4255), .I3(GND_net), 
            .O(n45154));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i29633_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i30671_4_lut (.I0(n45154), .I1(n46152), .I2(n43_adj_4261), 
            .I3(n45822), .O(n46192));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i30671_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i30672_3_lut (.I0(n46192), .I1(n82), .I2(n2448), .I3(GND_net), 
            .O(n46193));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i30672_3_lut.LUT_INIT = 16'h2b2b;
    SB_LUT4 i1_4_lut_adj_1478 (.I0(n46193), .I1(n22457), .I2(n81), .I3(n2447), 
            .O(n2471));
    defparam i1_4_lut_adj_1478.LUT_INIT = 16'hceef;
    SB_LUT4 div_11_LessThan_1417_i20_3_lut_3_lut (.I0(n98), .I1(n97), .I2(n2181), 
            .I3(GND_net), .O(n20_adj_4181));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1417_i20_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 i28676_2_lut_4_lut (.I0(n2176), .I1(n92), .I2(n2180), .I3(n96), 
            .O(n44195));
    defparam i28676_2_lut_4_lut.LUT_INIT = 16'hf99f;
    SB_LUT4 div_11_LessThan_1417_i22_3_lut_3_lut (.I0(n96), .I1(n92), .I2(n2176), 
            .I3(GND_net), .O(n22_adj_4183));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1417_i22_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 div_11_LessThan_1545_i41_2_lut (.I0(n2360), .I1(n85), .I2(GND_net), 
            .I3(GND_net), .O(n41_adj_4237));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1545_i41_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_11_LessThan_1417_i24_3_lut_3_lut (.I0(n95), .I1(n94), .I2(n2178), 
            .I3(GND_net), .O(n24_adj_4185));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1417_i24_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 div_11_LessThan_1545_i45_2_lut (.I0(n2358), .I1(n83), .I2(GND_net), 
            .I3(GND_net), .O(n45_adj_4239));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1545_i45_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_11_LessThan_1545_i39_2_lut (.I0(n2361), .I1(n86), .I2(GND_net), 
            .I3(GND_net), .O(n39_adj_4235));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1545_i39_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i28682_2_lut_4_lut (.I0(n2178), .I1(n94), .I2(n2179), .I3(n95), 
            .O(n44201));
    defparam i28682_2_lut_4_lut.LUT_INIT = 16'hf99f;
    SB_LUT4 div_11_mux_3_i6_3_lut (.I0(encoder0_position[5]), .I1(n20), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n386));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_mux_3_i6_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_11_LessThan_1545_i43_2_lut (.I0(n2359), .I1(n84), .I2(GND_net), 
            .I3(GND_net), .O(n43_adj_4238));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1545_i43_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_11_LessThan_1350_i22_3_lut_3_lut (.I0(n98), .I1(n97), .I2(n2081), 
            .I3(GND_net), .O(n22_adj_4164));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1350_i22_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 div_11_LessThan_1545_i27_2_lut (.I0(n2367), .I1(n92), .I2(GND_net), 
            .I3(GND_net), .O(n27_adj_4229));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1545_i27_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_11_LessThan_1545_i29_2_lut (.I0(n2366), .I1(n91), .I2(GND_net), 
            .I3(GND_net), .O(n29_adj_4230));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1545_i29_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_11_LessThan_1545_i31_2_lut (.I0(n2365), .I1(n90), .I2(GND_net), 
            .I3(GND_net), .O(n31_adj_4231));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1545_i31_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i28702_2_lut_4_lut (.I0(n2076), .I1(n92), .I2(n2080), .I3(n96), 
            .O(n44221));
    defparam i28702_2_lut_4_lut.LUT_INIT = 16'hf99f;
    SB_LUT4 div_11_LessThan_1350_i24_3_lut_3_lut (.I0(n96), .I1(n92), .I2(n2076), 
            .I3(GND_net), .O(n24_adj_4166));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1350_i24_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 div_11_LessThan_1545_i17_2_lut (.I0(n2372), .I1(n97), .I2(GND_net), 
            .I3(GND_net), .O(n17_adj_4220));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1545_i17_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_11_LessThan_1545_i19_2_lut (.I0(n2371), .I1(n96), .I2(GND_net), 
            .I3(GND_net), .O(n19_adj_4222));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1545_i19_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i28706_2_lut_4_lut (.I0(n2078), .I1(n94), .I2(n2079), .I3(n95), 
            .O(n44225));
    defparam i28706_2_lut_4_lut.LUT_INIT = 16'hf99f;
    SB_LUT4 div_11_LessThan_1545_i33_2_lut (.I0(n2364), .I1(n89), .I2(GND_net), 
            .I3(GND_net), .O(n33_adj_4232));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1545_i33_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_11_LessThan_1545_i35_2_lut (.I0(n2363), .I1(n88), .I2(GND_net), 
            .I3(GND_net), .O(n35_adj_4233));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1545_i35_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_11_LessThan_1545_i37_2_lut (.I0(n2362), .I1(n87), .I2(GND_net), 
            .I3(GND_net), .O(n37_adj_4234));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1545_i37_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_11_LessThan_1350_i26_3_lut_3_lut (.I0(n95), .I1(n94), .I2(n2078), 
            .I3(GND_net), .O(n26_adj_4168));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1350_i26_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 div_11_LessThan_1545_i21_2_lut (.I0(n2370), .I1(n95), .I2(GND_net), 
            .I3(GND_net), .O(n21_adj_4224));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1545_i21_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_11_LessThan_1545_i23_2_lut (.I0(n2369), .I1(n94), .I2(GND_net), 
            .I3(GND_net), .O(n23_adj_4226));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1545_i23_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_11_LessThan_1545_i25_2_lut (.I0(n2368), .I1(n93), .I2(GND_net), 
            .I3(GND_net), .O(n25_adj_4227));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1545_i25_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_11_i1547_1_lut (.I0(n2381), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n2382));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1547_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i29184_4_lut (.I0(n37_adj_4234), .I1(n25_adj_4227), .I2(n23_adj_4226), 
            .I3(n21_adj_4224), .O(n44705));
    defparam i29184_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i29814_4_lut (.I0(n19_adj_4222), .I1(n17_adj_4220), .I2(n2373), 
            .I3(n98), .O(n45335));
    defparam i29814_4_lut.LUT_INIT = 16'hfeef;
    SB_LUT4 i30067_4_lut (.I0(n25_adj_4227), .I1(n23_adj_4226), .I2(n21_adj_4224), 
            .I3(n45335), .O(n45588));
    defparam i30067_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i30065_4_lut (.I0(n31_adj_4231), .I1(n29_adj_4230), .I2(n27_adj_4229), 
            .I3(n45588), .O(n45586));
    defparam i30065_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i29189_4_lut (.I0(n37_adj_4234), .I1(n35_adj_4233), .I2(n33_adj_4232), 
            .I3(n45586), .O(n44710));
    defparam i29189_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 div_11_LessThan_1545_i14_4_lut (.I0(n386), .I1(n99), .I2(n2374), 
            .I3(n558), .O(n14_adj_4218));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1545_i14_4_lut.LUT_INIT = 16'h0317;
    SB_LUT4 i30121_3_lut (.I0(n14_adj_4218), .I1(n87), .I2(n37_adj_4234), 
            .I3(GND_net), .O(n45642));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i30121_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i30122_3_lut (.I0(n45642), .I1(n86), .I2(n39_adj_4235), .I3(GND_net), 
            .O(n45643));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i30122_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 div_11_LessThan_1545_i40_3_lut (.I0(n22_adj_4225), .I1(n83), 
            .I2(n45_adj_4239), .I3(GND_net), .O(n40_adj_4236));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1545_i40_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i29175_4_lut (.I0(n43_adj_4238), .I1(n41_adj_4237), .I2(n39_adj_4235), 
            .I3(n44705), .O(n44696));
    defparam i29175_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i30245_4_lut (.I0(n40_adj_4236), .I1(n20_adj_4223), .I2(n45_adj_4239), 
            .I3(n44694), .O(n45766));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i30245_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i29629_3_lut (.I0(n45643), .I1(n85), .I2(n41_adj_4237), .I3(GND_net), 
            .O(n45150));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i29629_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 div_11_LessThan_1281_i24_3_lut_3_lut (.I0(n98), .I1(n97), .I2(n1978), 
            .I3(GND_net), .O(n24_adj_4146));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1281_i24_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 div_11_LessThan_1545_i26_3_lut (.I0(n18_adj_4221), .I1(n91), 
            .I2(n29_adj_4230), .I3(GND_net), .O(n26_adj_4228));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1545_i26_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i30517_4_lut (.I0(n26_adj_4228), .I1(n16_adj_4219), .I2(n29_adj_4230), 
            .I3(n44721), .O(n46038));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i30517_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i30518_3_lut (.I0(n46038), .I1(n90), .I2(n31_adj_4231), .I3(GND_net), 
            .O(n46039));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i30518_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i30382_3_lut (.I0(n46039), .I1(n89), .I2(n33_adj_4232), .I3(GND_net), 
            .O(n45903));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i30382_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i30309_4_lut (.I0(n43_adj_4238), .I1(n41_adj_4237), .I2(n39_adj_4235), 
            .I3(n44710), .O(n45830));
    defparam i30309_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i28726_2_lut_4_lut (.I0(n1973), .I1(n92), .I2(n1977), .I3(n96), 
            .O(n44245));
    defparam i28726_2_lut_4_lut.LUT_INIT = 16'hf99f;
    SB_LUT4 i30547_4_lut (.I0(n45150), .I1(n45766), .I2(n45_adj_4239), 
            .I3(n44696), .O(n46068));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i30547_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i29627_3_lut (.I0(n45903), .I1(n88), .I2(n35_adj_4233), .I3(GND_net), 
            .O(n45148));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i29627_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i30549_4_lut (.I0(n45148), .I1(n46068), .I2(n45_adj_4239), 
            .I3(n45830), .O(n46070));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i30549_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i1_4_lut_adj_1479 (.I0(n46070), .I1(n22454), .I2(n82), .I3(n2357), 
            .O(n2381));
    defparam i1_4_lut_adj_1479.LUT_INIT = 16'hceef;
    SB_LUT4 div_11_LessThan_1281_i26_3_lut_3_lut (.I0(n96), .I1(n92), .I2(n1973), 
            .I3(GND_net), .O(n26_adj_4148));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1281_i26_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 i12052_3_lut (.I0(\data_out_frame[18] [3]), .I1(\data_out_frame[19] [3]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n17_adj_4358));   // verilog/coms.v(100[12:33])
    defparam i12052_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_11_LessThan_1482_i37_2_lut (.I0(n2269), .I1(n88), .I2(GND_net), 
            .I3(GND_net), .O(n37_adj_4214));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1482_i37_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_11_LessThan_1482_i43_2_lut (.I0(n2266), .I1(n85), .I2(GND_net), 
            .I3(GND_net), .O(n43_adj_4217));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1482_i43_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_11_LessThan_1482_i41_2_lut (.I0(n2267), .I1(n86), .I2(GND_net), 
            .I3(GND_net), .O(n41_adj_4216));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1482_i41_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_11_LessThan_1482_i39_2_lut (.I0(n2268), .I1(n87), .I2(GND_net), 
            .I3(GND_net), .O(n39_adj_4215));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1482_i39_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_11_LessThan_1482_i31_2_lut (.I0(n2272), .I1(n91), .I2(GND_net), 
            .I3(GND_net), .O(n31_adj_4211));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1482_i31_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_11_LessThan_1482_i33_2_lut (.I0(n2271), .I1(n90), .I2(GND_net), 
            .I3(GND_net), .O(n33_adj_4212));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1482_i33_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_11_LessThan_1482_i35_2_lut (.I0(n2270), .I1(n89), .I2(GND_net), 
            .I3(GND_net), .O(n35_adj_4213));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1482_i35_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_11_LessThan_1482_i27_2_lut (.I0(n2274), .I1(n93), .I2(GND_net), 
            .I3(GND_net), .O(n27_adj_4208));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1482_i27_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_11_LessThan_1482_i29_2_lut (.I0(n2273), .I1(n92), .I2(GND_net), 
            .I3(GND_net), .O(n29_adj_4210));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1482_i29_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_11_LessThan_1482_i19_2_lut (.I0(n2278_adj_4003), .I1(n97), 
            .I2(GND_net), .I3(GND_net), .O(n19_adj_4202));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1482_i19_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_11_LessThan_1482_i21_2_lut (.I0(n2277_adj_4002), .I1(n96), 
            .I2(GND_net), .I3(GND_net), .O(n21_adj_4204));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1482_i21_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_11_LessThan_1482_i23_2_lut (.I0(n2276), .I1(n95), .I2(GND_net), 
            .I3(GND_net), .O(n23_adj_4206));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1482_i23_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_11_LessThan_1482_i25_2_lut (.I0(n2275), .I1(n94), .I2(GND_net), 
            .I3(GND_net), .O(n25_adj_4207));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1482_i25_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_11_i1484_1_lut (.I0(n2288_adj_4006), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n2289_adj_4007));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1484_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_11_LessThan_1482_i17_2_lut (.I0(n2279_adj_4004), .I1(n98), 
            .I2(GND_net), .I3(GND_net), .O(n17_adj_4200));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1482_i17_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i29250_4_lut (.I0(n23_adj_4206), .I1(n21_adj_4204), .I2(n19_adj_4202), 
            .I3(n17_adj_4200), .O(n44771));
    defparam i29250_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i29244_4_lut (.I0(n29_adj_4210), .I1(n27_adj_4208), .I2(n25_adj_4207), 
            .I3(n44771), .O(n44765));
    defparam i29244_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i30315_4_lut (.I0(n35_adj_4213), .I1(n33_adj_4212), .I2(n31_adj_4211), 
            .I3(n44765), .O(n45836));
    defparam i30315_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 div_11_LessThan_1482_i16_4_lut (.I0(n385), .I1(n99), .I2(n2280_adj_4005), 
            .I3(n558), .O(n16_adj_4199));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1482_i16_4_lut.LUT_INIT = 16'h0317;
    SB_LUT4 i30127_3_lut (.I0(n16_adj_4199), .I1(n87), .I2(n39_adj_4215), 
            .I3(GND_net), .O(n45648));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i30127_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i30128_3_lut (.I0(n45648), .I1(n86), .I2(n41_adj_4216), .I3(GND_net), 
            .O(n45649));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i30128_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i29826_4_lut (.I0(n41_adj_4216), .I1(n39_adj_4215), .I2(n27_adj_4208), 
            .I3(n44769), .O(n45347));
    defparam i29826_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i30243_3_lut (.I0(n22_adj_4205), .I1(n93), .I2(n27_adj_4208), 
            .I3(GND_net), .O(n45764));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i30243_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i29619_3_lut (.I0(n45649), .I1(n85), .I2(n43_adj_4217), .I3(GND_net), 
            .O(n45140));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i29619_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 div_11_LessThan_1482_i28_3_lut (.I0(n20_adj_4203), .I1(n91), 
            .I2(n31_adj_4211), .I3(GND_net), .O(n28_adj_4209));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1482_i28_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i30515_4_lut (.I0(n28_adj_4209), .I1(n18_adj_4201), .I2(n31_adj_4211), 
            .I3(n44761), .O(n46036));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i30515_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i30516_3_lut (.I0(n46036), .I1(n90), .I2(n33_adj_4212), .I3(GND_net), 
            .O(n46037));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i30516_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i30386_3_lut (.I0(n46037), .I1(n89), .I2(n35_adj_4213), .I3(GND_net), 
            .O(n45907));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i30386_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i29830_4_lut (.I0(n41_adj_4216), .I1(n39_adj_4215), .I2(n37_adj_4214), 
            .I3(n45836), .O(n45351));
    defparam i29830_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i30383_4_lut (.I0(n45140), .I1(n45764), .I2(n43_adj_4217), 
            .I3(n45347), .O(n45904));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i30383_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i29617_3_lut (.I0(n45907), .I1(n88), .I2(n37_adj_4214), .I3(GND_net), 
            .O(n45138));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i29617_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i30588_4_lut (.I0(n45138), .I1(n45904), .I2(n43_adj_4217), 
            .I3(n45351), .O(n46109));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i30588_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i30589_3_lut (.I0(n46109), .I1(n84), .I2(n2265), .I3(GND_net), 
            .O(n46110));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i30589_3_lut.LUT_INIT = 16'h2b2b;
    SB_LUT4 i1_4_lut_adj_1480 (.I0(n46110), .I1(n22451), .I2(n83), .I3(n2264), 
            .O(n2288_adj_4006));
    defparam i1_4_lut_adj_1480.LUT_INIT = 16'hceef;
    SB_LUT4 div_11_i1419_1_lut (.I0(n2192), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n2193));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1419_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_11_i1352_1_lut (.I0(n2093), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n2094));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1352_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_11_i1283_1_lut (.I0(n1991), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n1992));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1283_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_11_i1212_1_lut (.I0(n1886), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n1887));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1212_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_11_i1139_1_lut (.I0(n1778), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n1779));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1139_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_11_i1064_1_lut (.I0(n1667), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n1668));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1064_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_11_i987_1_lut (.I0(n1553), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n1554));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i987_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_11_i908_1_lut (.I0(n1436), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n1437));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i908_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_11_i827_1_lut (.I0(n1316), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n1317));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i827_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_11_i744_1_lut (.I0(n1193), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n1194));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i744_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i10731_3_lut (.I0(IntegralLimit[18]), .I1(\data_in_frame[8] [2]), 
            .I2(n23399), .I3(GND_net), .O(n24149));   // verilog/coms.v(126[12] 289[6])
    defparam i10731_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_11_i659_1_lut (.I0(n1067), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n1068));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i659_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_11_i572_1_lut (.I0(n938), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n939));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i572_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_11_i483_1_lut (.I0(n806), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n807));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i483_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_11_i392_1_lut (.I0(n671), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n672));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i392_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_11_i299_1_lut (.I0(n533), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n534));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i299_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i10747_3_lut (.I0(IntegralLimit[5]), .I1(\data_in_frame[10] [5]), 
            .I2(n23399), .I3(GND_net), .O(n24165));   // verilog/coms.v(126[12] 289[6])
    defparam i10747_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_11_i204_1_lut (.I0(n392), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n393));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i204_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i2_4_lut (.I0(n558), .I1(n99), .I2(n224), .I3(n22403), .O(n248));
    defparam i2_4_lut.LUT_INIT = 16'hff37;
    SB_LUT4 i31368_2_lut (.I0(encoder0_position[23]), .I1(gearBoxRatio[23]), 
            .I2(GND_net), .I3(GND_net), .O(n46887));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i31368_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i28736_2_lut_4_lut (.I0(n1975), .I1(n94), .I2(n1976), .I3(n95), 
            .O(n44255));
    defparam i28736_2_lut_4_lut.LUT_INIT = 16'hf99f;
    SB_LUT4 i10732_3_lut (.I0(IntegralLimit[17]), .I1(\data_in_frame[8] [1]), 
            .I2(n23399), .I3(GND_net), .O(n24150));   // verilog/coms.v(126[12] 289[6])
    defparam i10732_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_11_LessThan_1281_i28_3_lut_3_lut (.I0(n95), .I1(n94), .I2(n1975), 
            .I3(GND_net), .O(n28_adj_4150));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1281_i28_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 i1_2_lut_3_lut_adj_1481 (.I0(n89), .I1(n88), .I2(n22436), 
            .I3(GND_net), .O(n22430));
    defparam i1_2_lut_3_lut_adj_1481.LUT_INIT = 16'hf7f7;
    SB_LUT4 div_11_LessThan_1210_i26_3_lut_3_lut (.I0(n98), .I1(n97), .I2(n1872), 
            .I3(GND_net), .O(n26_adj_4128));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1210_i26_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 i28762_2_lut_4_lut (.I0(n1867), .I1(n92), .I2(n1871), .I3(n96), 
            .O(n44281));
    defparam i28762_2_lut_4_lut.LUT_INIT = 16'hf99f;
    SB_LUT4 div_11_LessThan_1210_i28_3_lut_3_lut (.I0(n96), .I1(n92), .I2(n1867), 
            .I3(GND_net), .O(n28_adj_4130));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1210_i28_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 i10425_3_lut (.I0(\data_in_frame[11] [7]), .I1(rx_data[7]), 
            .I2(n40225), .I3(GND_net), .O(n23843));   // verilog/coms.v(126[12] 289[6])
    defparam i10425_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i10426_3_lut (.I0(\data_in_frame[11] [6]), .I1(rx_data[6]), 
            .I2(n40225), .I3(GND_net), .O(n23844));   // verilog/coms.v(126[12] 289[6])
    defparam i10426_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i10427_3_lut (.I0(\data_in_frame[11] [5]), .I1(rx_data[5]), 
            .I2(n40225), .I3(GND_net), .O(n23845));   // verilog/coms.v(126[12] 289[6])
    defparam i10427_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i10428_3_lut (.I0(\data_in_frame[11] [4]), .I1(rx_data[4]), 
            .I2(n40225), .I3(GND_net), .O(n23846));   // verilog/coms.v(126[12] 289[6])
    defparam i10428_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i10429_3_lut (.I0(\data_in_frame[11] [3]), .I1(rx_data[3]), 
            .I2(n40225), .I3(GND_net), .O(n23847));   // verilog/coms.v(126[12] 289[6])
    defparam i10429_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i10430_3_lut (.I0(\data_in_frame[11] [2]), .I1(rx_data[2]), 
            .I2(n40225), .I3(GND_net), .O(n23848));   // verilog/coms.v(126[12] 289[6])
    defparam i10430_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i10431_3_lut (.I0(\data_in_frame[11] [1]), .I1(rx_data[1]), 
            .I2(n40225), .I3(GND_net), .O(n23849));   // verilog/coms.v(126[12] 289[6])
    defparam i10431_3_lut.LUT_INIT = 16'hacac;
    \quad(DEBOUNCE_TICKS=100)_U1  quad_counter0 (.n2276({n2277, n2278, n2279, 
            n2280, n2281, n2282, n2283, n2284, n2285, n2286, n2287, 
            n2288, n2289, n2290, n2291, n2292, n2293, n2294, n2295, 
            n2296, n2297, n2298, n2299, n2300}), .encoder0_position({encoder0_position}), 
            .GND_net(GND_net), .data_o({quadA_debounced, quadB_debounced}), 
            .clk32MHz(clk32MHz), .n23721(n23721), .n23720(n23720), .n23719(n23719), 
            .n23718(n23718), .n23717(n23717), .n23716(n23716), .n23715(n23715), 
            .n23714(n23714), .n23713(n23713), .n23712(n23712), .n23711(n23711), 
            .n23710(n23710), .n23709(n23709), .n23708(n23708), .n23707(n23707), 
            .n23706(n23706), .n23705(n23705), .n23704(n23704), .n23703(n23703), 
            .n23702(n23702), .n23701(n23701), .n23700(n23700), .n23699(n23699), 
            .n23591(n23591), .count_enable(count_enable), .n24229(n24229), 
            .reg_B({reg_B}), .PIN_23_c_1(PIN_23_c_1), .PIN_24_c_0(PIN_24_c_0), 
            .n23593(n23593), .n41998(n41998)) /* synthesis lattice_noprune=1, syn_preserve=0, syn_module_defined=1, syn_noprune=0 */ ;   // verilog/TinyFPGA_B.v(166[15] 171[4])
    SB_LUT4 i28772_2_lut_4_lut (.I0(n1869), .I1(n94), .I2(n1870), .I3(n95), 
            .O(n44291));
    defparam i28772_2_lut_4_lut.LUT_INIT = 16'hf99f;
    SB_LUT4 i10432_3_lut (.I0(\data_in_frame[11] [0]), .I1(rx_data[0]), 
            .I2(n40225), .I3(GND_net), .O(n23850));   // verilog/coms.v(126[12] 289[6])
    defparam i10432_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_11_LessThan_1210_i30_3_lut_3_lut (.I0(n95), .I1(n94), .I2(n1869), 
            .I3(GND_net), .O(n30_adj_4132));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1210_i30_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 i1_2_lut_3_lut_adj_1482 (.I0(n85), .I1(n84), .I2(n22448), 
            .I3(GND_net), .O(n22442));
    defparam i1_2_lut_3_lut_adj_1482.LUT_INIT = 16'hf7f7;
    SB_LUT4 div_11_LessThan_1137_i28_3_lut_3_lut (.I0(n98), .I1(n97), .I2(n1763), 
            .I3(GND_net), .O(n28_adj_4116));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1137_i28_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 i28789_2_lut_4_lut (.I0(n1758), .I1(n92), .I2(n1762), .I3(n96), 
            .O(n44308));
    defparam i28789_2_lut_4_lut.LUT_INIT = 16'hf99f;
    SB_LUT4 div_11_LessThan_1137_i30_3_lut_3_lut (.I0(n96), .I1(n92), .I2(n1758), 
            .I3(GND_net), .O(n30_adj_4118));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1137_i30_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 div_11_LessThan_1062_i30_3_lut_3_lut (.I0(n98), .I1(n97), .I2(n1651), 
            .I3(GND_net), .O(n30_adj_4105));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1062_i30_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 i28827_2_lut_4_lut (.I0(n1646), .I1(n92), .I2(n1650), .I3(n96), 
            .O(n44346));
    defparam i28827_2_lut_4_lut.LUT_INIT = 16'hf99f;
    SB_LUT4 div_11_LessThan_1062_i32_3_lut_3_lut (.I0(n96), .I1(n92), .I2(n1646), 
            .I3(GND_net), .O(n32_adj_4107));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1062_i32_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 i10441_3_lut (.I0(\data_in_frame[9] [7]), .I1(rx_data[7]), .I2(n40222), 
            .I3(GND_net), .O(n23859));   // verilog/coms.v(126[12] 289[6])
    defparam i10441_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i10442_3_lut (.I0(\data_in_frame[9] [6]), .I1(rx_data[6]), .I2(n40222), 
            .I3(GND_net), .O(n23860));   // verilog/coms.v(126[12] 289[6])
    defparam i10442_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_11_LessThan_985_i32_3_lut_3_lut (.I0(n98), .I1(n97), .I2(n1536), 
            .I3(GND_net), .O(n32_adj_4096));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_985_i32_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 mux_21_i16_3_lut (.I0(encoder0_position[15]), .I1(motor_state_23__N_27[15]), 
            .I2(n15_adj_3961), .I3(GND_net), .O(motor_state[15]));   // verilog/TinyFPGA_B.v(137[5] 141[10])
    defparam mux_21_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10443_3_lut (.I0(\data_in_frame[9] [5]), .I1(rx_data[5]), .I2(n40222), 
            .I3(GND_net), .O(n23861));   // verilog/coms.v(126[12] 289[6])
    defparam i10443_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i10444_3_lut (.I0(\data_in_frame[9] [4]), .I1(rx_data[4]), .I2(n40222), 
            .I3(GND_net), .O(n23862));   // verilog/coms.v(126[12] 289[6])
    defparam i10444_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i10445_3_lut (.I0(\data_in_frame[9] [3]), .I1(rx_data[3]), .I2(n40222), 
            .I3(GND_net), .O(n23863));   // verilog/coms.v(126[12] 289[6])
    defparam i10445_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i10446_3_lut (.I0(\data_in_frame[9] [2]), .I1(rx_data[2]), .I2(n40222), 
            .I3(GND_net), .O(n23864));   // verilog/coms.v(126[12] 289[6])
    defparam i10446_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i10447_3_lut (.I0(\data_in_frame[9] [1]), .I1(rx_data[1]), .I2(n40222), 
            .I3(GND_net), .O(n23865));   // verilog/coms.v(126[12] 289[6])
    defparam i10447_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i28862_2_lut_4_lut (.I0(n1531), .I1(n92), .I2(n1535), .I3(n96), 
            .O(n44381));
    defparam i28862_2_lut_4_lut.LUT_INIT = 16'hf99f;
    SB_LUT4 i10448_3_lut (.I0(\data_in_frame[9] [0]), .I1(rx_data[0]), .I2(n40222), 
            .I3(GND_net), .O(n23866));   // verilog/coms.v(126[12] 289[6])
    defparam i10448_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_11_LessThan_985_i34_3_lut_3_lut (.I0(n96), .I1(n92), .I2(n1531), 
            .I3(GND_net), .O(n34_adj_4097));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_985_i34_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 i10733_3_lut (.I0(IntegralLimit[16]), .I1(\data_in_frame[8] [0]), 
            .I2(n23399), .I3(GND_net), .O(n24151));   // verilog/coms.v(126[12] 289[6])
    defparam i10733_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i20165_3_lut_4_lut (.I0(n649), .I1(n99), .I2(n371), .I3(n558), 
            .O(n4));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i20165_3_lut_4_lut.LUT_INIT = 16'heee8;
    SB_LUT4 i1_2_lut_3_lut_adj_1483 (.I0(n87), .I1(n86), .I2(n22442), 
            .I3(GND_net), .O(n22436));
    defparam i1_2_lut_3_lut_adj_1483.LUT_INIT = 16'hf7f7;
    SB_LUT4 i20141_3_lut_4_lut (.I0(n510), .I1(n99), .I2(n370), .I3(n558), 
            .O(n4_adj_3956));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i20141_3_lut_4_lut.LUT_INIT = 16'heee8;
    SB_LUT4 i1_2_lut_4_lut (.I0(n97), .I1(n96), .I2(n95), .I3(n22415), 
            .O(n22406));
    defparam i1_2_lut_4_lut.LUT_INIT = 16'hff7f;
    SB_LUT4 i1_2_lut_3_lut_adj_1484 (.I0(n96), .I1(n95), .I2(n22415), 
            .I3(GND_net), .O(n22409));
    defparam i1_2_lut_3_lut_adj_1484.LUT_INIT = 16'hf7f7;
    SB_LUT4 i1_2_lut_4_lut_adj_1485 (.I0(n94), .I1(n93), .I2(n92), .I3(n22424), 
            .O(n22415));
    defparam i1_2_lut_4_lut_adj_1485.LUT_INIT = 16'hff7f;
    SB_LUT4 i1_2_lut_3_lut_adj_1486 (.I0(n93), .I1(n92), .I2(n22424), 
            .I3(GND_net), .O(n22418));
    defparam i1_2_lut_3_lut_adj_1486.LUT_INIT = 16'hf7f7;
    SB_LUT4 i1_2_lut_4_lut_adj_1487 (.I0(n91), .I1(n90), .I2(n89), .I3(n22433), 
            .O(n22424));
    defparam i1_2_lut_4_lut_adj_1487.LUT_INIT = 16'hff7f;
    SB_LUT4 i20197_3_lut_4_lut (.I0(n785), .I1(n99), .I2(n372), .I3(n558), 
            .O(n4_adj_3993));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i20197_3_lut_4_lut.LUT_INIT = 16'heee8;
    \quad(DEBOUNCE_TICKS=100)  quad_counter1 (.n24204(n24204), .encoder1_position({encoder1_position}), 
            .clk32MHz(clk32MHz), .n24203(n24203), .n24202(n24202), .n24201(n24201), 
            .n24200(n24200), .n24199(n24199), .n24198(n24198), .n24197(n24197), 
            .n24196(n24196), .n24195(n24195), .n24194(n24194), .n24193(n24193), 
            .n24192(n24192), .n24191(n24191), .n24190(n24190), .n24189(n24189), 
            .n24188(n24188), .n24187(n24187), .n24186(n24186), .n24185(n24185), 
            .n24184(n24184), .n24183(n24183), .n24170(n24170), .data_o({quadA_debounced_adj_3990, 
            quadB_debounced_adj_3991}), .n2226({n2227, n2228, n2229, 
            n2230, n2231, n2232, n2233, n2234, n2235, n2236, n2237, 
            n2238, n2239, n2240, n2241, n2242, n2243, n2244, n2245, 
            n2246, n2247, n2248, n2249, n2250}), .GND_net(GND_net), 
            .n23592(n23592), .count_enable(count_enable_adj_3992), .n24231(n24231), 
            .reg_B({reg_B_adj_4406}), .PIN_18_c_1(PIN_18_c_1), .PIN_19_c_0(PIN_19_c_0), 
            .n23595(n23595), .n41767(n41767)) /* synthesis lattice_noprune=1, syn_preserve=0, syn_module_defined=1, syn_noprune=0 */ ;   // verilog/TinyFPGA_B.v(174[15] 179[4])
    SB_LUT4 i1_2_lut_4_lut_adj_1488 (.I0(n83), .I1(n82), .I2(n81), .I3(n22457), 
            .O(n22448));
    defparam i1_2_lut_4_lut_adj_1488.LUT_INIT = 16'hff7f;
    SB_LUT4 i1_2_lut_3_lut_adj_1489 (.I0(n82), .I1(n81), .I2(n22457), 
            .I3(GND_net), .O(n22451));
    defparam i1_2_lut_3_lut_adj_1489.LUT_INIT = 16'hf7f7;
    SB_LUT4 i1_2_lut_4_lut_adj_1490 (.I0(n80), .I1(n79), .I2(n78), .I3(n77), 
            .O(n22457));
    defparam i1_2_lut_4_lut_adj_1490.LUT_INIT = 16'hff7f;
    SB_LUT4 i1_2_lut_3_lut_adj_1491 (.I0(n79), .I1(n78), .I2(n77), .I3(GND_net), 
            .O(n22460));
    defparam i1_2_lut_3_lut_adj_1491.LUT_INIT = 16'hf7f7;
    SB_LUT4 i10473_3_lut (.I0(\data_in_frame[5] [7]), .I1(rx_data[7]), .I2(n40218), 
            .I3(GND_net), .O(n23891));   // verilog/coms.v(126[12] 289[6])
    defparam i10473_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i10474_3_lut (.I0(\data_in_frame[5] [6]), .I1(rx_data[6]), .I2(n40218), 
            .I3(GND_net), .O(n23892));   // verilog/coms.v(126[12] 289[6])
    defparam i10474_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i10475_3_lut (.I0(\data_in_frame[5] [5]), .I1(rx_data[5]), .I2(n40218), 
            .I3(GND_net), .O(n23893));   // verilog/coms.v(126[12] 289[6])
    defparam i10475_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i10476_3_lut (.I0(\data_in_frame[5] [4]), .I1(rx_data[4]), .I2(n40218), 
            .I3(GND_net), .O(n23894));   // verilog/coms.v(126[12] 289[6])
    defparam i10476_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i10477_3_lut (.I0(\data_in_frame[5] [3]), .I1(rx_data[3]), .I2(n40218), 
            .I3(GND_net), .O(n23895));   // verilog/coms.v(126[12] 289[6])
    defparam i10477_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i10478_3_lut (.I0(\data_in_frame[5] [2]), .I1(rx_data[2]), .I2(n40218), 
            .I3(GND_net), .O(n23896));   // verilog/coms.v(126[12] 289[6])
    defparam i10478_3_lut.LUT_INIT = 16'hacac;
    
endmodule
//
// Verilog Description of module motorControl
//

module motorControl (\Kd[3] , GND_net, \motor_state[15] , \Kp[6] , \PID_CONTROLLER.err[18] , 
            \Kd[4] , \motor_state[14] , \motor_state[13] , \motor_state[12] , 
            \motor_state[11] , \motor_state[10] , \motor_state[9] , \motor_state[8] , 
            \Kd[5] , \motor_state[7] , \Kd[6] , \motor_state[6] , \Kd[1] , 
            \motor_state[5] , \Kd[0] , \motor_state[4] , \motor_state[3] , 
            \Kd[7] , \motor_state[2] , \Kd[2] , \motor_state[1] , \Kp[7] , 
            \motor_state[0] , VCC_net, \PID_CONTROLLER.err_prev[31] , 
            \PID_CONTROLLER.err_prev[23] , \PID_CONTROLLER.err_prev[22] , 
            \PID_CONTROLLER.err_prev[21] , \Kp[1] , \PID_CONTROLLER.err[6] , 
            \PID_CONTROLLER.err_prev[20] , \PID_CONTROLLER.err_prev[19] , 
            \Kp[0] , \PID_CONTROLLER.err[7] , \Kp[2] , \Kp[3] , \Kp[4] , 
            \PID_CONTROLLER.err_prev[18] , \PID_CONTROLLER.err_prev[17] , 
            \Kp[5] , \PID_CONTROLLER.err_prev[16] , \PID_CONTROLLER.err[9] , 
            \PID_CONTROLLER.err[8] , \PID_CONTROLLER.err[5] , \PID_CONTROLLER.err[4] , 
            \PID_CONTROLLER.err[3] , \PID_CONTROLLER.err[2] , \PID_CONTROLLER.err[1] , 
            \PID_CONTROLLER.err[0] , pwm_count, \PID_CONTROLLER.err[31] , 
            n24227, pwm, clk32MHz, n24226, n24225, n24224, n24223, 
            n39110, n24220, n24219, n24218, n24217, n24216, n24215, 
            n24214, n24213, n24212, n24211, n24208, n24207, n24206, 
            n24205, n24172, \PID_CONTROLLER.err[16] , \PID_CONTROLLER.err_prev[15] , 
            \PID_CONTROLLER.err[17] , \PID_CONTROLLER.err[21] , \Ki[5] , 
            \Ki[6] , \Ki[7] , \PID_CONTROLLER.err_prev[14] , \PID_CONTROLLER.err_prev[13] , 
            \PID_CONTROLLER.err_prev[12] , \PID_CONTROLLER.err[19] , \PID_CONTROLLER.err_prev[11] , 
            \PID_CONTROLLER.err[20] , \PID_CONTROLLER.err[22] , \PID_CONTROLLER.err[23] , 
            PIN_7_c_1, setpoint, \PID_CONTROLLER.err[10] , PIN_6_c_0, 
            \PID_CONTROLLER.err_prev[10] , \PID_CONTROLLER.err[11] , \PID_CONTROLLER.err_prev[9] , 
            \PID_CONTROLLER.err_prev[8] , \PID_CONTROLLER.err_prev[7] , 
            \PID_CONTROLLER.err_prev[6] , \PID_CONTROLLER.err_prev[5] , 
            \PWMLimit[3] , \PWMLimit[2] , \Ki[0] , \PID_CONTROLLER.err_prev[4] , 
            \Ki[1] , \Ki[2] , \PID_CONTROLLER.err_prev[3] , \Ki[3] , 
            hall1, hall2, \Ki[4] , \PID_CONTROLLER.err_prev[2] , \PID_CONTROLLER.err_prev[1] , 
            n421, n44153, \PID_CONTROLLER.err_prev[0] , hall3, n44109, 
            n44111, n44117, n44113, n44115, n25, n30, n26, n853, 
            n21, n855, n856, n857, n859, n860, n861, n862, n863, 
            n864, n865, n866, n867, n868, n869, n870, n871, 
            n872, n873, n874, n875, n44074, n414, n415, n45714, 
            \pwm_23__N_2960[6] , \pwm_23__N_2960[5] , \PID_CONTROLLER.err[12] , 
            \PID_CONTROLLER.err[13] , \PID_CONTROLLER.err[14] , n23746, 
            n23745, n23744, n23743, n23742, n23741, n23740, n23739, 
            n23738, n23737, n23736, n23735, n23734, n23733, n23732, 
            n23731, n23730, n23729, n23728, n23727, n23726, n23725, 
            n23724, n23723, \motor_state[23] , \PID_CONTROLLER.result[5] , 
            \PID_CONTROLLER.result[6] , PIN_8_c_2, PIN_9_c_3, PIN_10_c_4, 
            PIN_11_c_5, \motor_state[22] , \PID_CONTROLLER.err[15] , \motor_state[21] , 
            \motor_state[20] , \motor_state[19] , \motor_state[18] , \motor_state[17] , 
            \motor_state[16] , n23589, n471, n470, n469, n468, n467, 
            pwm_23__N_2957, n1, \PWMLimit[5] , n387, n27212, \PWMLimit[6] , 
            n464, n463, n462, n461, n460, n459, n458, n457, 
            n456, n455, \PWMLimit[9] , n11, n13, \deadband[3] , 
            \deadband[7] , \deadband[4] , \deadband[8] , \deadband[9] , 
            n13_adj_10, n11_adj_11, \deadband[2] , \deadband[0] , \deadband[1] , 
            n16, \PWMLimit[7] , \PWMLimit[4] , n41887, \PWMLimit[0] , 
            \PWMLimit[1] , n11_adj_12, n13_adj_13, \PWMLimit[8] , n11_adj_14, 
            n13_adj_15, \deadband[5] , \deadband[6] , IntegralLimit) /* synthesis lattice_noprune=1, syn_preserve=0, syn_module_defined=1, syn_noprune=0 */ ;
    input \Kd[3] ;
    input GND_net;
    input \motor_state[15] ;
    input \Kp[6] ;
    output \PID_CONTROLLER.err[18] ;
    input \Kd[4] ;
    input \motor_state[14] ;
    input \motor_state[13] ;
    input \motor_state[12] ;
    input \motor_state[11] ;
    input \motor_state[10] ;
    input \motor_state[9] ;
    input \motor_state[8] ;
    input \Kd[5] ;
    input \motor_state[7] ;
    input \Kd[6] ;
    input \motor_state[6] ;
    input \Kd[1] ;
    input \motor_state[5] ;
    input \Kd[0] ;
    input \motor_state[4] ;
    input \motor_state[3] ;
    input \Kd[7] ;
    input \motor_state[2] ;
    input \Kd[2] ;
    input \motor_state[1] ;
    input \Kp[7] ;
    input \motor_state[0] ;
    input VCC_net;
    output \PID_CONTROLLER.err_prev[31] ;
    output \PID_CONTROLLER.err_prev[23] ;
    output \PID_CONTROLLER.err_prev[22] ;
    output \PID_CONTROLLER.err_prev[21] ;
    input \Kp[1] ;
    output \PID_CONTROLLER.err[6] ;
    output \PID_CONTROLLER.err_prev[20] ;
    output \PID_CONTROLLER.err_prev[19] ;
    input \Kp[0] ;
    output \PID_CONTROLLER.err[7] ;
    input \Kp[2] ;
    input \Kp[3] ;
    input \Kp[4] ;
    output \PID_CONTROLLER.err_prev[18] ;
    output \PID_CONTROLLER.err_prev[17] ;
    input \Kp[5] ;
    output \PID_CONTROLLER.err_prev[16] ;
    output \PID_CONTROLLER.err[9] ;
    output \PID_CONTROLLER.err[8] ;
    output \PID_CONTROLLER.err[5] ;
    output \PID_CONTROLLER.err[4] ;
    output \PID_CONTROLLER.err[3] ;
    output \PID_CONTROLLER.err[2] ;
    output \PID_CONTROLLER.err[1] ;
    output \PID_CONTROLLER.err[0] ;
    output [8:0]pwm_count;
    output \PID_CONTROLLER.err[31] ;
    input n24227;
    output [23:0]pwm;
    input clk32MHz;
    input n24226;
    input n24225;
    input n24224;
    input n24223;
    input n39110;
    input n24220;
    input n24219;
    input n24218;
    input n24217;
    input n24216;
    input n24215;
    input n24214;
    input n24213;
    input n24212;
    input n24211;
    input n24208;
    input n24207;
    input n24206;
    input n24205;
    input n24172;
    output \PID_CONTROLLER.err[16] ;
    output \PID_CONTROLLER.err_prev[15] ;
    output \PID_CONTROLLER.err[17] ;
    output \PID_CONTROLLER.err[21] ;
    input \Ki[5] ;
    input \Ki[6] ;
    input \Ki[7] ;
    output \PID_CONTROLLER.err_prev[14] ;
    output \PID_CONTROLLER.err_prev[13] ;
    output \PID_CONTROLLER.err_prev[12] ;
    output \PID_CONTROLLER.err[19] ;
    output \PID_CONTROLLER.err_prev[11] ;
    output \PID_CONTROLLER.err[20] ;
    output \PID_CONTROLLER.err[22] ;
    output \PID_CONTROLLER.err[23] ;
    output PIN_7_c_1;
    input [23:0]setpoint;
    output \PID_CONTROLLER.err[10] ;
    output PIN_6_c_0;
    output \PID_CONTROLLER.err_prev[10] ;
    output \PID_CONTROLLER.err[11] ;
    output \PID_CONTROLLER.err_prev[9] ;
    output \PID_CONTROLLER.err_prev[8] ;
    output \PID_CONTROLLER.err_prev[7] ;
    output \PID_CONTROLLER.err_prev[6] ;
    output \PID_CONTROLLER.err_prev[5] ;
    input \PWMLimit[3] ;
    input \PWMLimit[2] ;
    input \Ki[0] ;
    output \PID_CONTROLLER.err_prev[4] ;
    input \Ki[1] ;
    input \Ki[2] ;
    output \PID_CONTROLLER.err_prev[3] ;
    input \Ki[3] ;
    input hall1;
    input hall2;
    input \Ki[4] ;
    output \PID_CONTROLLER.err_prev[2] ;
    output \PID_CONTROLLER.err_prev[1] ;
    output n421;
    output n44153;
    output \PID_CONTROLLER.err_prev[0] ;
    input hall3;
    output n44109;
    output n44111;
    output n44117;
    output n44113;
    output n44115;
    input n25;
    input n30;
    input n26;
    output n853;
    output n21;
    output n855;
    output n856;
    output n857;
    output n859;
    output n860;
    output n861;
    output n862;
    output n863;
    output n864;
    output n865;
    output n866;
    output n867;
    output n868;
    output n869;
    output n870;
    output n871;
    output n872;
    output n873;
    output n874;
    output n875;
    output n44074;
    output n414;
    output n415;
    input n45714;
    output \pwm_23__N_2960[6] ;
    output \pwm_23__N_2960[5] ;
    output \PID_CONTROLLER.err[12] ;
    output \PID_CONTROLLER.err[13] ;
    output \PID_CONTROLLER.err[14] ;
    input n23746;
    input n23745;
    input n23744;
    input n23743;
    input n23742;
    input n23741;
    input n23740;
    input n23739;
    input n23738;
    input n23737;
    input n23736;
    input n23735;
    input n23734;
    input n23733;
    input n23732;
    input n23731;
    input n23730;
    input n23729;
    input n23728;
    input n23727;
    input n23726;
    input n23725;
    input n23724;
    input n23723;
    input \motor_state[23] ;
    output \PID_CONTROLLER.result[5] ;
    output \PID_CONTROLLER.result[6] ;
    output PIN_8_c_2;
    output PIN_9_c_3;
    output PIN_10_c_4;
    output PIN_11_c_5;
    input \motor_state[22] ;
    output \PID_CONTROLLER.err[15] ;
    input \motor_state[21] ;
    input \motor_state[20] ;
    input \motor_state[19] ;
    input \motor_state[18] ;
    input \motor_state[17] ;
    input \motor_state[16] ;
    input n23589;
    output n471;
    output n470;
    output n469;
    output n468;
    output n467;
    output pwm_23__N_2957;
    input n1;
    input \PWMLimit[5] ;
    output n387;
    input n27212;
    input \PWMLimit[6] ;
    output n464;
    output n463;
    output n462;
    output n461;
    output n460;
    output n459;
    output n458;
    output n457;
    output n456;
    output n455;
    input \PWMLimit[9] ;
    input n11;
    input n13;
    input \deadband[3] ;
    input \deadband[7] ;
    input \deadband[4] ;
    input \deadband[8] ;
    input \deadband[9] ;
    input n13_adj_10;
    input n11_adj_11;
    input \deadband[2] ;
    input \deadband[0] ;
    input \deadband[1] ;
    input n16;
    input \PWMLimit[7] ;
    input \PWMLimit[4] ;
    output n41887;
    input \PWMLimit[0] ;
    input \PWMLimit[1] ;
    input n11_adj_12;
    input n13_adj_13;
    input \PWMLimit[8] ;
    input n11_adj_14;
    input n13_adj_15;
    input \deadband[5] ;
    input \deadband[6] ;
    input [23:0]IntegralLimit;
    
    wire clk32MHz /* synthesis SET_AS_NETWORK=clk32MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(34[8:16])
    wire [31:0]n57;
    
    wire n298;
    wire [20:0]n13594;
    wire [19:0]n14035;
    
    wire n34385, n34230;
    wire [24:0]n58;
    
    wire n34231, n34864;
    wire [33:0]n282;
    wire [55:0]n61;
    
    wire n34865, n637;
    wire [31:0]n63;
    
    wire n34863, n395;
    wire [26:0]n8049;
    wire [25:0]n8078;
    
    wire n304, n35299, n34862, n35396;
    wire [21:0]n8184;
    
    wire n219, n35397, n35300, n34861, n207, n35298, n34860, n35448;
    wire [19:0]n8231;
    
    wire n35449;
    wire [22:0]n8159;
    
    wire n29, n122, n34859, n17, n110, n34858, n34386;
    wire [15:0]n12157;
    wire [14:0]n12732;
    
    wire n326, n35125;
    wire [24:0]\PID_CONTROLLER.err_31__N_2825 ;
    
    wire n34229, n34857, n34576;
    wire [25:0]n10671;
    
    wire n34577;
    wire [27:0]n8019;
    
    wire n35297, n34384, n35296, n34228, n34227;
    wire [23:0]n8133;
    
    wire n35395;
    wire [20:0]n8208;
    
    wire n35447, n35487;
    wire [17:0]n8274;
    
    wire n35488;
    wire [16:0]n8294;
    wire [15:0]n8313;
    
    wire n35528;
    wire [26:0]n9929;
    
    wire n34575, n34856, n35126, n34574, n253, n35124, n34573, 
        n34572, n180, n35123, n35295, n35394, n34571, n34570, 
        n35, n107, n34569, n34568, n35294, n34567, n34566, n34565, 
        n692, n34564, n35293, n35393, n595, n34563, n498, n34562, 
        n35292, n34383, n34226, n34225, n34382, n34381, n34224, 
        n35446, n35392, n35291, n401, n34561, n34223, n507;
    wire [18:0]n8253;
    
    wire n35486, n34380, n34222, n35290, n34379, n34378, n604, 
        n35289, n34377, n304_adj_3378, n34560, n207_adj_3379, n34559, 
        n34221, n35445, n128, n34376, n34220, n35_adj_3381, n35391, 
        n710, n34375, n613, n34374, n516, n34373, n35288, n34219, 
        n419, n34372, n34218, n701, n322, n34371, n35390, n34217, 
        n225, n34370, n225_adj_3382, n34216, n35287, n35_adj_3383, 
        n128_adj_3384, n734;
    wire [9:0]n16420;
    wire [8:0]n16505;
    
    wire n34369;
    wire [31:0]n64;
    
    wire n34215, n34214, n34368, n34213, n34212, n35286, n34367, 
        n716, n34211, n743, n34366, n116, n34210, n646, n34365, 
        n34209, n23_adj_3389, n213, n310_adj_3390, n407, n492, n34208;
    wire [12:0]n16031;
    wire [11:0]n16185;
    
    wire n35677, n35676, n35585;
    wire [10:0]n8393;
    
    wire n446, n35586, n35527, n710_adj_3392, n35444, n35389, n35285, 
        n17_adj_3393, n110_adj_3394;
    wire [11:0]n14168;
    wire [10:0]n14560;
    
    wire n34558, n34557, n34556, n34555, n35284, n34554, n545, 
        n34553, n472, n34552, n399, n34551, n35388, n35283, n549, 
        n34364, n34550, n34207;
    wire [11:0]n8379;
    
    wire n349, n35584, n34549, n34548, n35282;
    wire [24:0]n11358;
    
    wire n34547, n34546, n34545, n35485, n613_adj_3396, n35443, 
        n35387, n35281, n34544, n34543, n34542, n504, n34541, 
        n35280, n34540, n34539, n34538, n34537, n35386, n35279, 
        n34536, n601, n34535, n34534, n34533, n35278, n34532, 
        n34531, n34530, n698, n34529, n516_adj_3397, n35442, n35385, 
        n35277, n695, n34528, n34206, n598, n34527, n501, n34526, 
        n404, n34525, n689, n35276, n307_adj_3399, n34524, n210, 
        n34523, n20_adj_3400, n113;
    wire [9:0]n14912;
    
    wire n34522, n34521, n35384, n592, n35275, n34520, n34519, 
        n34518, n322_adj_3401, n34517, n495, n35274, n34516, n34515, 
        n34514, n34513, n35484, n419_adj_3402, n35441, n35383, n107_adj_3403, 
        n398, n35273, n14_adj_3404;
    wire [23:0]n11992;
    
    wire n34512, n204, n34511, n34510, n301, n35272, n34509, n34508, 
        n34507, n34506, n35382, n35271, n34505, n34504, n34503, 
        n34502, n34501, n34500;
    wire [9:0]n66;
    wire [9:0]\PID_CONTROLLER.integral ;   // verilog/motorControl.v(33[22:30])
    
    wire n35076, n34499, n35075, n34498, n35526, n35440, n35381;
    wire [28:0]n7988;
    
    wire n35270, n34497, n35074, n34496, n35269, n34495, n35073, 
        n34494, n34493, n35072, n34492, n35268, n34491, n35071, 
        n34490, n35380, n34489, n35070, n35267;
    wire [8:0]n15226;
    
    wire n34488, n34487, n35069, n34486, n34485, n35068, n34484, 
        n35266, n589, n34483, n34482, n35483, n35439, n35379, 
        n34481;
    wire [8:0]n67;
    
    wire n35067, n34480, n35265, n35066, n35065, n134, n35264, 
        n35064, n35378, n35063, n35263, n35062;
    wire [22:0]n12575;
    
    wire n34473, n34472, n34471, n35061, n34470, n41, n34469, 
        n35262, n35060, n34468, n34467, n35377, n34466, n34465, 
        n35261;
    wire [29:0]n7956;
    
    wire n35059, n34464, n35058, n34463, n34462, n35057, n34461, 
        n35260, n34460, n686, n35056, n34459;
    wire [0:0]n5786;
    wire [29:0]n6542;
    
    wire n34730, n35376, n34729, n34458, n35055, n34728, n39108, 
        n24210, n24209, n34457, n34727, n35259, n231, n328, n34726, 
        n34205, n701_adj_3413, n34456, n452, n34363, n425, n252, 
        n35583, n98, n5, n35675, n62, n155_adj_3414, n35525, n35524, 
        n35674, n35054, n34725, n35438, n34204, n35258, n34203, 
        n35053, n34724, n355, n34362, n258, n34361, n604_adj_3417, 
        n34455, n35052, n34202, n34723, n34722, n34201, n410, 
        n35375, n35257, n195, n507_adj_3421, n34454, n34721, n35051, 
        n34720;
    wire [31:0]\PID_CONTROLLER.result_31__N_3003 ;
    wire [31:0]\PID_CONTROLLER.result ;   // verilog/motorControl.v(32[23:29])
    
    wire n68, n161, n410_adj_3422, n34453;
    wire [5:0]GATES_5__N_2788;
    
    wire n313_adj_3423, n34452, n619, n35482, n34719;
    wire [18:0]n14434;
    
    wire n34360, n35050, n34359, n35256, n216, n34451, n35049, 
        n34718, n34200, n26_adj_3425, n119, n34717, n35437, n313_adj_3426, 
        n35374, n35255, n522, n292, n34716, n34450, n583, n34449, 
        n510, n34448, n34715, n437, n34447, n389, n35254, n35048, 
        n34714, n364, n34446, n34713, n291, n34445, n35047, n34712, 
        n218, n34444, n486, n145, n34443, n34711, n216_adj_3429, 
        n35373, n35046, n34358, n72, n34710, n35673;
    wire [12:0]n8364;
    
    wire n35582, n35253, n35581, n34709, n34199;
    wire [21:0]n13109;
    
    wire n34442, n35045, n35252, n34708, n34441, n34198, n34707, 
        n34440, n35044, n26_adj_3432, n119_adj_3433, n680, n34706, 
        n34439, n35436, n35251, n35043, n583_adj_3434, n34705, n34438, 
        n35042, n34704, n34703, n34357, n34437, n34197, n34356, 
        n35250, n34702, n35481, n34196, n35041, n34436, n34355, 
        n34354, n34701, n35040, n34435, n34195;
    wire [24:0]n8106;
    
    wire n35372, n35371, n35249, n35480, n35370, n35435, n35434, 
        n35479, n35523, n34434, n35478, n35580, n35369, n35522, 
        n35248, n44552, n35672, n35579, n35039, n35038, n35521, 
        n35247, n34433, n34194, n35368, n6, n34432, n35578, n35037, 
        n35246, n35671, n35433, n34431, n34353, n35245, n34430, 
        n35670, n35244, n540, n35669, n443, n35668, n34429, n346, 
        n35667, n34193, n683, n35036, n35520, n34352, n249, n35666, 
        n35577, n586, n35035, n59, n152_adj_3435, n35367, n34428, 
        n201, n35243, n35366, n489, n35034;
    wire [28:0]n7760;
    
    wire n34693, n34692, n35365, n392, n35033, n734_adj_3436, n35576, 
        n35519, n35432, n637_adj_3437, n35575;
    wire [10:0]n16314;
    
    wire n35665, n34427, n35364, n34691, n35477, n11_adj_3438, n104, 
        n35664, n722, n35518, n35363, n35431, n704, n34426;
    wire [6:0]n69;
    wire [6:0]Kd_delay_counter;   // verilog/motorControl.v(27[13:29])
    
    wire n34690;
    wire [0:0]n7061;
    
    wire n35242, n35362, n295, n35032, n35663, n540_adj_3439, n35574, 
        n625, n35517;
    wire [55:0]n191;
    
    wire n35241, n35476, n35475, n198, n35031, n35240, n35662, 
        n607, n34425, n34689;
    wire [5:0]GATES_5__N_3048;
    
    wire n5_adj_3441, n35661, n510_adj_3442, n34424, n34688, n528, 
        n35516, n35430, n443_adj_3443, n35573, n35361, n34687, n737, 
        n35660, n34351, n413, n34423, n35239, n8, n101, n431, 
        n35515, n346_adj_3445, n35572, n35238, n640, n35659, n34350, 
        n543, n35658, n334, n35514, n34192, n35360, n446_adj_3446, 
        n35657, n35429, n35359, n35237;
    wire [13:0]n13256;
    
    wire n35030, n34686, n316_adj_3447, n34422, n219_adj_3448, n34421, 
        n35236, n34685, n35029, n29_adj_3449, n122_adj_3450, n34684, 
        n34420, n34419, n34683, n34418, n35474, n35428, n34417, 
        n35028, n34682, n34681, n34349, n35235, n35027, n740, 
        n34416, n35358, n34680, n34679, n35026, n643, n34415, 
        n34678, n546, n34414, n34677, n35234, n449, n34413, n34191, 
        n35233, n35025, n34676, n34675, n352, n34412, n255, n34411, 
        n35024;
    wire [31:0]n70;
    
    wire n34674, n34348, n65, n158, n35232, n35023, n35022, n35357, 
        n34673, n35473, n349_adj_3453, n35656, n713, n34347, n35427, 
        n34672, n35231, n34671, n616, n34346, n683_adj_3454, n34670, 
        n586_adj_3455, n34669, n35230, n878, n17_adj_3456, n35356, 
        n489_adj_3457, n34668, n35021, n35229, n519, n34345, n44151, 
        n392_adj_3458, n34667, n35020, n249_adj_3459, n35571, n35426, 
        n252_adj_3460, n35655, n422, n34344, n325, n34343, n295_adj_3461, 
        n34666, n35228, n228_adj_3462, n34342, n35019, n35355, n237, 
        n35513, n38, n131_adj_3463, n35227, n35018, n59_adj_3465, 
        n152_adj_3466;
    wire [17:0]n14793;
    
    wire n34341, n34340, n35017, n62_adj_3467, n155_adj_3468, n198_adj_3469, 
        n34665, n35226, n34339, n34410, n8_adj_3470, n101_adj_3471, 
        n34338, n698_adj_3472, n35354, n35225, n34337, n35472;
    wire [13:0]n8348;
    
    wire n35570, n47_adj_3473, n140_adj_3474, n35471;
    wire [27:0]n9125;
    
    wire n34664, n34336, n34663, n34335, n35470, n35569, n34334;
    wire [21:0]n8448;
    wire [20:0]n8472;
    
    wire n35654, n35469, n35568, n35512, n35511, n35567, n35653, 
        n35468, n35510, n35016, n35015, n35652, n35467, n34333, 
        n35566, n34662, n35651, n35565, n35650, n35564, n731, 
        n35563, n35649, n34332, n35014, n35648, n35509, n35647, 
        n35646, n35425, n35645, n35644, n34331, n35643, n35224, 
        n34661, n35642, n35424, n34660, n35641, n34330, n35013, 
        n601_adj_3476, n35353, n35223, n716_adj_3477, n34329;
    wire [4:0]n16637;
    
    wire n35466, n35990, n35012, n34659, n35640, n707, n35423, 
        n35508, n634, n35562, n35639, n537, n35561, n440, n35560, 
        n35638, n35637, n343, n35559, n246, n35558, n35636, n35635, 
        n34658, n35222, n34657, n504_adj_3479, n35352, n34656, n619_adj_3480, 
        n34328, n35221, n34655, n34409, n35634, n407_adj_3482, n35351, 
        n56, n149_adj_3483, n35011;
    wire [14:0]n8331;
    
    wire n35557, n522_adj_3484, n34327, n34408;
    wire [6:0]n8439;
    wire [5:0]n9319;
    
    wire n752, n35633, n34654, n34653, n425_adj_3485, n34326, n35556, 
        n328_adj_3486, n34325, n610, n35422, n34407, n231_adj_3487, 
        n34324, n655, n35632, n35220, n41_adj_3488, n134_adj_3489, 
        n35507, n35555, n34652;
    wire [7:0]n16571;
    
    wire n34323, n34322, n746, n34321, n35465, n513, n35421, n40121, 
        n34651, n35219, n34650, n649, n34320, GATES_5__N_3055, n34166;
    wire [23:0]n73;
    
    wire n34165;
    wire [23:0]n852;
    
    wire n552, n34319, n310_adj_3494, n35350, n680_adj_3495, n35218, 
        n455_c, n34318, n358, n34317, n34649, n261, n34316, n583_adj_3496, 
        n35217, n34648, n71, n164, n34164, n34647, n486_adj_3497, 
        n35216, n34646, n34163, n558, n35631, n461_c, n35630, 
        n34162, n34161, n34160, n34645, n213_adj_3502, n35349, n34159, 
        n34310, n34309, n34644, n34308, n34307, n34158, n416, 
        n35420, n389_adj_3504, n35215, n34643, n34306, n34157, n686_adj_3506, 
        n34642, n364_adj_3507, n35629, n267, n35628, n34156, n34305, 
        n34155, n23_adj_3510, n116_adj_3511, n34304, n292_adj_3512, 
        n35214, n589_adj_3513, n34641, n34303, n34154, n492_adj_3515, 
        n34640, n34302, n34301, n34153, n34152, n34300, n34151, 
        n40176, n34150, n395_adj_3520, n34639, n86, n170_adj_3521, 
        n34299;
    wire [7:0]n8429;
    
    wire n35627, n749, n35626, n34149, n34298, n34148, n34147, 
        n195_adj_3525, n35213, n298_adj_3526, n34638, n34297, n34146, 
        n34145, n35554, n652, n35625, n35506, n713_adj_3529, n35464, 
        n35348, n5_adj_3531, n98_adj_3532, n34296, n201_adj_3533, 
        n34637, n34144, n34295, n25474, n6_adj_3536, n34143, n11_adj_3537, 
        n104_adj_3538, n34294, n34293, n34142;
    wire [31:0]n75;
    
    wire n34141, n555, n35624, n458_c, n35623, n35347;
    wire [19:0]n9327;
    wire [18:0]n10118;
    
    wire n35212;
    wire [8:0]n7065;
    wire [22:0]n1804;
    
    wire n1711, n35987;
    wire [22:0]n1803;
    
    wire n1707, n35986;
    wire [22:0]n1802;
    
    wire n1703, n35985;
    wire [22:0]n1801;
    
    wire n1699, n35984;
    wire [22:0]n1800;
    
    wire n1695, n35983;
    wire [22:0]n1799;
    
    wire n1691, n35982;
    wire [22:0]n1798;
    
    wire n1687, n35981, n35553, n35552;
    wire [22:0]n1797;
    
    wire n1683, n35980;
    wire [22:0]n1796;
    
    wire n35979, n34292, n34140, n35978, n35211, n35977, n35976, 
        n35975, n35974, n35505, n35551, n361, n35622, n35504, 
        n264, n35621, n35503, n35550, n74, n167_adj_3542, n35210;
    wire [8:0]n8418;
    
    wire n35620, n35619, n746_adj_3543, n35618, n319, n35419, n35346, 
        n649_adj_3544, n35617, n35209, n35973, n35972, n35971, n35970, 
        n35969, n35208, n34139, n35968, n34138, n35967, n35966, 
        n35965, n616_adj_3547, n35463, n35964, n35963, n35962, n552_adj_3548, 
        n35616, n35502, n35961, n35960, n35345, n728, n35549, 
        n455_adj_3549, n35615, n35959, n35207, n358_adj_3550, n35614, 
        n35958, n719, n35501;
    wire [12:0]n13734;
    
    wire n34636, n34635, n519_adj_3551, n35462, n34291, n34137, 
        n20_adj_3554, n34136, n34290, n35957, n261_adj_3556, n35613, 
        n35956, n34135, n631, n35548, n222_adj_3558, n35418, n35955, 
        n34289, n34634, n35954, n35953, n35952, n35951, n35950, 
        n35949, n35948, n35947, n35344, n35946, n26_adj_3559, n34134, 
        n32_adj_3562, n125, n35945, n35343, n35206, n35944, n536, 
        n35943, n463_c, n35942, n390, n35941, n35342, n534, n35547, 
        n422_adj_3566, n35461, n71_adj_3567, n164_adj_3568, n317, 
        n35940, n34288, n244_adj_3571, n35939;
    wire [23:0]n76;
    wire [23:0]n79;
    
    wire n34133, n35205, n34633, n34287, n45_adj_3573, n34132, n43_adj_3575, 
        n34131, n35341, n35417, n35204, n35203;
    wire [9:0]n8406;
    
    wire n35612, n35611, n35610, n24_adj_3577, n171_adj_3579, n35938, 
        n98_adj_3580, n35936, n35935, n35934, n35933, n35932, n35931, 
        n437_adj_3581, n35546, n743_adj_3582, n35609, n646_adj_3583, 
        n35608, n549_adj_3584, n35607, n452_adj_3585, n35606, n355_adj_3586, 
        n35605, n258_adj_3587, n35604, n68_adj_3588, n161_adj_3589, 
        n622, n35500, n35930, n35929, n35928, n35927, n35926, 
        n35925, n35924, n35923, n340, n35545, n243_adj_3590, n35544, 
        n28_adj_3591, n34286, n41_adj_3592, n34130, n55_adj_3594, 
        n35922, n23_adj_3596, n39_adj_3597, n34129, n35340, n35202, 
        n53_adj_3599, n146_adj_3600, n35416, n525, n35499, n35201, 
        n40975, n34632, n35339, n44158, n37_adj_3601, n34128, n34285, 
        n18_adj_3603, n35200, n34284, n35415, n35338, n35_adj_3604, 
        n34127, n35199, n34631, n35921, n34283, n533, n35920, 
        n34282, n33_adj_3608, n34126, n35198, n35197, n34630, n460_c, 
        n35919, n31_adj_3611, n34125, n34281, n387_c, n35918, n35196, 
        n428, n35498, n325_adj_3613, n35460, n314_adj_3615, n35917, 
        n35337, n241_adj_3617, n35916, n35195, n35194, n168_adj_3619, 
        n35915, n26_adj_3620, n95, n35603, n35602, n35913, n35601, 
        n34629, n34280, n35600, n35912, n29_adj_3621, n34124, n35543, 
        n35542, n35414, n34628, n27_adj_3623, n34123;
    wire [16:0]n15114;
    
    wire n34279, n34278, n35336, n41372, n658, n35193, n34277, 
        n331, n35497, n35335;
    wire [4:0]n10111;
    
    wire n564, n35192, n740_adj_3625, n35599, n35911, n228_adj_3626, 
        n35459, n643_adj_3627, n35598, n464_adj_3628, n35191, n25_adj_3629, 
        n34122, n23_adj_3631, n34121, n34276, n34627, n35541, n21_adj_3633, 
        n34120, n35334, n370, n35190, n546_adj_3635, n35597, n34275, 
        n19_adj_3636, n34119, n276, n35189, n35413, n17_adj_3638, 
        n34118, n35333, n182_adj_3640, n38_adj_3641, n131_adj_3642;
    wire [17:0]n10852;
    
    wire n35188, n35187, n35332, n35186, n35910, n234_adj_3643, 
        n35496, n35909, n35908, n35907, n34626, n34274, n15_adj_3644, 
        n34117, n35185, n13_adj_3646, n34116, n35906, n34273, n11_adj_3648, 
        n34115, n35905, n34625, n34272, n9_adj_3650, n34114, n7_adj_3652, 
        n34113, n34271, n5_adj_3654, n34112, n44_adj_3656, n137_adj_3657, 
        n35904, n35412, n35331, n35184, n35903, n34270, n3_adj_3658, 
        n34111, n35902, n35901, n35458, n34624, n35900, n34269, 
        n719_adj_3660, n34268, n35183, n622_adj_3661, n34267, n35899, 
        n525_adj_3664, n34266, n35898, n34623;
    wire [31:0]pwm_23__N_2960;
    wire [31:0]n82;
    
    wire n34110, n34109, n34108, n35330, n34622, n428_adj_3668, 
        n34265, n331_adj_3669, n34264, n35495, n35457, n35411, n35182, 
        n234_adj_3670, n34263, n34621, n44_adj_3671, n137_adj_3672, 
        n34107, n530, n35897, n34620, n35181, n34106, n34105, 
        n34619, n34104, n695_adj_3677, n35329, n34618, n457_c, n35896, 
        n35180, n35540, n35410, n384, n35895, n34103, n35179, 
        n34617, n311_adj_3681, n35894, n35178, n598_adj_3682, n35328, 
        n35177, n35456, n501_adj_3683, n35327, n238_adj_3685, n35893, 
        n35494, n165_adj_3687, n35892, n35539, n35176, n23_adj_3688, 
        n92, n449_adj_3689, n35596, n34616, n35890, n35889, n35888, 
        n352_adj_3690, n35595, n35887, n35886, n34102, n35175, n34615, 
        n35885, n34614, n34613, n35538, n35493, n35409, n404_adj_3692, 
        n35326, n35174, n35173, n35172, n35455, n307_adj_3693, n35325, 
        n35171, n35884, n35883, n35408, n210_adj_3694, n35324, n35537, 
        n35882, n255_adj_3695, n35594, n35881, n35536, n34101, n35880, 
        n35879;
    wire [16:0]n11531;
    
    wire n35170, n35169, n35454, n20_adj_3697, n113_adj_3698, n35168, 
        n35167, n35535, n35407, n35323, n35492, n35166, n35322, 
        n35165, n35321, n35164, n65_adj_3699, n158_adj_3700, n35163, 
        n44044, n28200, n35406, n35878, n35877, n35876, n35453, 
        n35875, n35593, n35592, n527, n35874, n35491, n454, n35873, 
        n381, n35872, n308_adj_3706, n35871, n235_adj_3708, n35870, 
        n725, n35534, n162, n35869, n20_adj_3709, n89, n35867, 
        n35591, n35866, n34612, n35865, n35320, n35864, n35590, 
        n35863, n35490, n35862, n35861, n35162, n35860, n35859, 
        n35858, n35857, n35405, n35161, n34611, n35856, n35319, 
        n35855, n35160, n35854, n34610, n34609, n34608, n35159, 
        n34607, n35318, n34606, n35158, n34605, n35452, n35404, 
        n35157, n35317, n35156, n34604, n35155, n35853, n34603, 
        n35316, n689_adj_3710, n34602, n35154, n592_adj_3711, n34601, 
        n495_adj_3712, n34600, n398_adj_3713, n34599, n35315, n35451, 
        n35852, n35403, n524, n35851, n35153, n35152, n35314, 
        n35151, n35402, n451, n35850, n378, n35849, n35150, n35313, 
        n305, n35848, n35149, n35312, n232_adj_3718, n35847, n35148, 
        n159, n35846, n17_adj_3719, n86_adj_3720, n35311, n35147, 
        n35844, n704_adj_3721, n35401, n301_adj_3722, n34598, n35843, 
        n628, n35533, n35146, n204_adj_3723, n34597, n35842, n35841, 
        n35145, n35310, n34886, n34885, n35144, n34884, n14_adj_3724, 
        n107_adj_3725, n35840, n35489, n34883, n35450, n35143, n35839, 
        n35838, n35837, n35836, n35835, n35834, n35309, n35833, 
        n35832, n35142, n35831, n35830, n531_adj_3726, n35532, n35829, 
        n607_adj_3728, n35400, n521, n35828, n35141, n34882, n34596, 
        n35140, n35308, n34881, n448, n35827, n35139, n34880, 
        n35307, n34879, n34595, n510_adj_3731, n35399, n375, n35826, 
        n302, n35825, n34594, n35138, n35589, n229_adj_3733, n35824, 
        n156_adj_3735, n35823, n34239, n34238, n34878, n34877, n34593, 
        n34876, n14_adj_3738, n83, n35821, n35820, n35819, n35818, 
        n34237, n35306, n35137, n35817, n35305, n35136, n413_adj_3740, 
        n35398, n35135, n34875, n35134, n34874, n35816, n35304, 
        n35815, n34873, n35133, n34872, n434, n35531, n34871, 
        n316_adj_3742, n692_adj_3743, n35303, n35132, n34592, n35814, 
        n34236, n35813, n35812, n35811, n34870, n34235, n34591, 
        n34406, n35810, n34234, n35809, n34405, n34590, n34404, 
        n34403, n35131, n34589, n34402, n34401, n337, n35530, 
        n240_adj_3748, n35529, n50_adj_3749, n143_adj_3750, n35808, 
        n35807, n35806, n518, n35805, n445, n35804, n372, n35803, 
        n299_adj_3755, n35802, n226_adj_3757, n35801, n153_adj_3759, 
        n35800, n11_adj_3760, n80, n35798, n35797, n34588, n34400, 
        n35796, n35795, n35794, n35793, n35792, n35791, n35790, 
        n35789, n35788, n35787, n35786, n35785, n35784, n35783, 
        n515, n35782, n442, n35781, n369, n35780, n296_adj_3766, 
        n35779, n223_adj_3768, n35778, n150_adj_3770, n35777, n8_adj_3771, 
        n77, n35775, n35774, n35773, n35772, n35771, n35770, n35769, 
        n35768, n35767, n35766, n35765, n35764, n35763, n35762, 
        n35761, n35760, n512, n35759, n439, n35758, n366, n35757, 
        n293, n35756, n220_adj_3777, n35755, n147_adj_3778, n35754, 
        n5_adj_3779, n74_adj_3780;
    wire [15:0]n15399;
    
    wire n35753, n35752, n35751, n35750, n35749, n35748, n35747, 
        n35746, n35745, n35744, n722_adj_3781, n35743, n625_adj_3782, 
        n35742, n528_adj_3783, n35741, n431_adj_3784, n35740, n334_adj_3785, 
        n35739, n237_adj_3786, n35738, n47_adj_3787, n140_adj_3788;
    wire [6:0]n16620;
    
    wire n35737, n749_adj_3789, n35736, n652_adj_3790, n35735, n595_adj_3791, 
        n35302, n34399, n35130, n34587, n34398, n555_adj_3792, n35734, 
        n458_adj_3793, n35733, n361_adj_3794, n35732, n264_adj_3795, 
        n35731, n86_adj_3796, n167_adj_3797;
    wire [14:0]n15640;
    
    wire n35730, n35729, n35728, n35727, n35726, n35725, n35724, 
        n35723, n35722, n725_adj_3798, n35721, n628_adj_3799, n35720, 
        n531_adj_3800, n35719, n434_adj_3801, n35718, n337_adj_3802, 
        n35717, n240_adj_3803, n35716, n50_adj_3804, n143_adj_3805;
    wire [5:0]n16629;
    
    wire n41719, n658_adj_3806, n35715, n558_adj_3807, n35714, n464_adj_3808, 
        n35713;
    wire [3:0]n16644;
    
    wire n370_adj_3809, n35712, n276_adj_3810, n35711, n182_adj_3811;
    wire [13:0]n15850;
    
    wire n35710, n35709, n35708, n35707, n35706, n35705, n35704, 
        n35703, n728_adj_3812, n35702, n631_adj_3813, n35701, n534_adj_3814, 
        n35700, n437_adj_3815, n35699, n340_adj_3816, n35698, n243_adj_3817, 
        n35697, n53_adj_3818, n146_adj_3819, n752_adj_3820, n35696, 
        n35695, n35694, n34233, n34869, n35693, n34397, n34586, 
        n34396, n35129, n34585, n707_adj_3822, n34395, n35692, n35691, 
        n35690, n35689, n35688, n35687, n35686, n35685, n610_adj_3823, 
        n34394, n35684, n34232, n498_adj_3825, n35301, n513_adj_3826, 
        n34393, n35128, n34584, n416_adj_3827, n34392, n34583, n34868, 
        n34582, n319_adj_3828, n34391, n34581, n222_adj_3829, n34390, 
        n35127, n34867, n34580, n731_adj_3830, n35683, n737_adj_3831, 
        n35588, n634_adj_3832, n35682, n537_adj_3833, n35681, n32_adj_3834, 
        n125_adj_3835, n640_adj_3836, n35587, n440_adj_3837, n35680, 
        n34579, n343_adj_3839, n35679, n34389, n246_adj_3840, n35678, 
        n401_adj_3841, n543_adj_3842, n34866, n34578, n34388, n56_adj_3843, 
        n149_adj_3844, n34387, n33546, n7_adj_3851, n8_adj_3852, n8_adj_3853, 
        n33872, n4_adj_3856, n7_adj_3857, n19_adj_3858, n15_adj_3859, 
        n17_adj_3860, n7_adj_3861, n9_adj_3862, n18_adj_3863, n24_adj_3864, 
        n5_adj_3865, n44539, n4_adj_3867, n45656, n45657, n10_adj_3869, 
        n49_adj_3870, n22_adj_3871, n12_adj_3872, n16_adj_3873, n62_adj_3874, 
        n26_adj_3875, n40200, n40124, n44166, n25_adj_3876, n6_adj_3877, 
        n45808, n45809, n44530, n45098, n45627, n20_adj_3878, n45712, 
        n7_adj_3879, n15_adj_3880, n9_adj_3881, n17_adj_3882, n45305, 
        n45299, n45313, n45283, n45263, n30_adj_3885, n45325, n45582, 
        n45309, n45828, n44676, n45566, n45988, n46140, n6_adj_3886, 
        n45670, n45229, n24_adj_3887, n44632, n47290, n8_adj_3888, 
        n45924, n45076, n4_adj_3889, n45668, n44664, n47267, n10_adj_3890, 
        n46034, n45078, n46162, n46163, n44638, n46117, n45084, 
        n46158, n50_adj_3891, n19_adj_3893, n42185, n42181, n42183, 
        n29_adj_3894, n6_adj_3895, n44119, n17_adj_3896, n7_adj_3897, 
        n9_adj_3898, n15_adj_3899, n19_adj_3900, n14_adj_3901, n15_adj_3902, 
        n15_adj_3903, n9_adj_3904, n6_adj_3905, n4_adj_3906, n45660, 
        n45661, n45197, n8_adj_3909, n45088, n45710, n18_adj_3910, 
        n41755, n41486, n26_adj_3911, n6_adj_3912, n41766, n41485, 
        n34_adj_3913, n41915, n41828, n56_adj_3914, n41769, n40126, 
        n4_adj_3915, n13_adj_3916, n18_adj_3917, n16_adj_3918, n17_adj_3919, 
        n15_adj_3920, n41951, n5_adj_3921, n44602, n8_adj_3923, n6_adj_3924, 
        n16_adj_3925, n44041, n4_adj_3926, n45662, n45663, n14_adj_3928, 
        n12_adj_3929, n13_adj_3930, n11_adj_3931, n44592, n44590, 
        n46008, n45086, n41904, n46156, n45227, n56_adj_3932, n60, 
        pwm_23__N_2959, n45706, n33897, n8_adj_3933, n8_adj_3934, 
        n18_adj_3935, n24_adj_3936, n22_adj_3937, n26_adj_3938, n41724, 
        n11_adj_3939, n9_adj_3940, n17_adj_3941, n45395, n45393, n44745, 
        n47477, n45399, n45387, n44787, n47465, n10_adj_3942, n30_adj_3943, 
        n5_adj_3944, n45403, n45401, n44811, n45620, n46006, n45389, 
        n45840, n46079, n46182, n6_adj_3945, n44888, n24_adj_3946, 
        n45698, n44763, n47430, n8_adj_3947, n45700, n45064, n4_adj_3948, 
        n45672, n45673, n8_adj_3949, n44735, n6_adj_3950, n16_adj_3951, 
        n44739, n45798, n45074, n46056, n4_adj_3952, n45678, n44789, 
        n46032, n45066, n46160, n46161, n45365, n45936, n45072, 
        n46057, n46054, n6_adj_3953, n6_adj_3954, n4_adj_3955;
    
    SB_LUT4 mult_12_i201_2_lut (.I0(\Kd[3] ), .I1(n57[2]), .I2(GND_net), 
            .I3(GND_net), .O(n298));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i201_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_3294_18_lut (.I0(GND_net), .I1(n14035[15]), .I2(GND_net), 
            .I3(n34385), .O(n13594[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3294_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY state_23__I_0_add_2_17 (.CI(n34230), .I0(\motor_state[15] ), 
            .I1(n58[15]), .CO(n34231));
    SB_CARRY add_13_add_1_20061_add_1_11 (.CI(n34864), .I0(n282[9]), .I1(n61[9]), 
            .CO(n34865));
    SB_LUT4 mult_10_i428_2_lut (.I0(\Kp[6] ), .I1(\PID_CONTROLLER.err[18] ), 
            .I2(GND_net), .I3(GND_net), .O(n637));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i428_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_13_add_1_20061_add_1_10_lut (.I0(GND_net), .I1(n282[8]), 
            .I2(n61[8]), .I3(n34863), .O(n63[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_13_add_1_20061_add_1_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_12_i266_2_lut (.I0(\Kd[4] ), .I1(n57[2]), .I2(GND_net), 
            .I3(GND_net), .O(n395));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i266_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_3059_4_lut (.I0(GND_net), .I1(n8078[1]), .I2(n304), .I3(n35299), 
            .O(n8049[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3059_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_13_add_1_20061_add_1_10 (.CI(n34863), .I0(n282[8]), .I1(n61[8]), 
            .CO(n34864));
    SB_LUT4 add_13_add_1_20061_add_1_9_lut (.I0(GND_net), .I1(n282[7]), 
            .I2(n61[7]), .I3(n34862), .O(n63[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_13_add_1_20061_add_1_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3063_3 (.CI(n35396), .I0(n8184[0]), .I1(n219), .CO(n35397));
    SB_CARRY add_3059_4 (.CI(n35299), .I0(n8078[1]), .I1(n304), .CO(n35300));
    SB_CARRY add_13_add_1_20061_add_1_9 (.CI(n34862), .I0(n282[7]), .I1(n61[7]), 
            .CO(n34863));
    SB_LUT4 add_13_add_1_20061_add_1_8_lut (.I0(GND_net), .I1(n282[6]), 
            .I2(n61[6]), .I3(n34861), .O(n63[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_13_add_1_20061_add_1_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3059_3_lut (.I0(GND_net), .I1(n8078[0]), .I2(n207), .I3(n35298), 
            .O(n8049[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3059_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_13_add_1_20061_add_1_8 (.CI(n34861), .I0(n282[6]), .I1(n61[6]), 
            .CO(n34862));
    SB_LUT4 add_13_add_1_20061_add_1_7_lut (.I0(GND_net), .I1(n282[5]), 
            .I2(n61[5]), .I3(n34860), .O(n63[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_13_add_1_20061_add_1_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3065_12 (.CI(n35448), .I0(n8231[9]), .I1(GND_net), .CO(n35449));
    SB_LUT4 add_3063_2_lut (.I0(GND_net), .I1(n29), .I2(n122), .I3(GND_net), 
            .O(n8159[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3063_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3059_3 (.CI(n35298), .I0(n8078[0]), .I1(n207), .CO(n35299));
    SB_CARRY add_13_add_1_20061_add_1_7 (.CI(n34860), .I0(n282[5]), .I1(n61[5]), 
            .CO(n34861));
    SB_LUT4 add_13_add_1_20061_add_1_6_lut (.I0(GND_net), .I1(n282[4]), 
            .I2(n61[4]), .I3(n34859), .O(n63[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_13_add_1_20061_add_1_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3059_2_lut (.I0(GND_net), .I1(n17), .I2(n110), .I3(GND_net), 
            .O(n8049[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3059_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_13_add_1_20061_add_1_6 (.CI(n34859), .I0(n282[4]), .I1(n61[4]), 
            .CO(n34860));
    SB_LUT4 add_13_add_1_20061_add_1_5_lut (.I0(GND_net), .I1(n282[3]), 
            .I2(n61[3]), .I3(n34858), .O(n63[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_13_add_1_20061_add_1_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3294_18 (.CI(n34385), .I0(n14035[15]), .I1(GND_net), 
            .CO(n34386));
    SB_CARRY add_3059_2 (.CI(GND_net), .I0(n17), .I1(n110), .CO(n35298));
    SB_LUT4 add_3231_5_lut (.I0(GND_net), .I1(n12732[2]), .I2(n326), .I3(n35125), 
            .O(n12157[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3231_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 state_23__I_0_add_2_16_lut (.I0(GND_net), .I1(\motor_state[14] ), 
            .I2(n58[14]), .I3(n34229), .O(\PID_CONTROLLER.err_31__N_2825 [14])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_13_add_1_20061_add_1_5 (.CI(n34858), .I0(n282[3]), .I1(n61[3]), 
            .CO(n34859));
    SB_LUT4 add_13_add_1_20061_add_1_4_lut (.I0(GND_net), .I1(n282[2]), 
            .I2(n61[2]), .I3(n34857), .O(n63[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_13_add_1_20061_add_1_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3142_20 (.CI(n34576), .I0(n10671[17]), .I1(GND_net), 
            .CO(n34577));
    SB_LUT4 add_3058_29_lut (.I0(GND_net), .I1(n8049[26]), .I2(GND_net), 
            .I3(n35297), .O(n8019[27])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3058_29_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3294_17_lut (.I0(GND_net), .I1(n14035[14]), .I2(GND_net), 
            .I3(n34384), .O(n13594[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3294_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3063_2 (.CI(GND_net), .I0(n29), .I1(n122), .CO(n35396));
    SB_CARRY state_23__I_0_add_2_16 (.CI(n34229), .I0(\motor_state[14] ), 
            .I1(n58[14]), .CO(n34230));
    SB_LUT4 add_3058_28_lut (.I0(GND_net), .I1(n8049[25]), .I2(GND_net), 
            .I3(n35296), .O(n8019[26])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3058_28_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 state_23__I_0_add_2_15_lut (.I0(GND_net), .I1(\motor_state[13] ), 
            .I2(n58[13]), .I3(n34228), .O(\PID_CONTROLLER.err_31__N_2825 [13])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY state_23__I_0_add_2_15 (.CI(n34228), .I0(\motor_state[13] ), 
            .I1(n58[13]), .CO(n34229));
    SB_LUT4 state_23__I_0_add_2_14_lut (.I0(GND_net), .I1(\motor_state[12] ), 
            .I2(n58[12]), .I3(n34227), .O(\PID_CONTROLLER.err_31__N_2825 [12])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3062_25_lut (.I0(GND_net), .I1(n8159[22]), .I2(GND_net), 
            .I3(n35395), .O(n8133[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3062_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3065_11_lut (.I0(GND_net), .I1(n8231[8]), .I2(GND_net), 
            .I3(n35447), .O(n8208[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3065_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3067_12 (.CI(n35487), .I0(n8274[9]), .I1(GND_net), .CO(n35488));
    SB_LUT4 add_3069_18_lut (.I0(GND_net), .I1(n8313[15]), .I2(GND_net), 
            .I3(n35528), .O(n8294[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3069_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3142_19_lut (.I0(GND_net), .I1(n10671[16]), .I2(GND_net), 
            .I3(n34575), .O(n9929[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3142_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3142_19 (.CI(n34575), .I0(n10671[16]), .I1(GND_net), 
            .CO(n34576));
    SB_CARRY add_13_add_1_20061_add_1_4 (.CI(n34857), .I0(n282[2]), .I1(n61[2]), 
            .CO(n34858));
    SB_LUT4 add_13_add_1_20061_add_1_3_lut (.I0(GND_net), .I1(n282[1]), 
            .I2(n61[1]), .I3(n34856), .O(n63[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_13_add_1_20061_add_1_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3231_5 (.CI(n35125), .I0(n12732[2]), .I1(n326), .CO(n35126));
    SB_LUT4 add_3142_18_lut (.I0(GND_net), .I1(n10671[15]), .I2(GND_net), 
            .I3(n34574), .O(n9929[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3142_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3142_18 (.CI(n34574), .I0(n10671[15]), .I1(GND_net), 
            .CO(n34575));
    SB_CARRY add_13_add_1_20061_add_1_3 (.CI(n34856), .I0(n282[1]), .I1(n61[1]), 
            .CO(n34857));
    SB_LUT4 add_13_add_1_20061_add_1_2_lut (.I0(GND_net), .I1(n282[0]), 
            .I2(n61[0]), .I3(GND_net), .O(n63[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_13_add_1_20061_add_1_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3231_4_lut (.I0(GND_net), .I1(n12732[1]), .I2(n253), .I3(n35124), 
            .O(n12157[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3231_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3058_28 (.CI(n35296), .I0(n8049[25]), .I1(GND_net), .CO(n35297));
    SB_LUT4 add_3142_17_lut (.I0(GND_net), .I1(n10671[14]), .I2(GND_net), 
            .I3(n34573), .O(n9929[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3142_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3142_17 (.CI(n34573), .I0(n10671[14]), .I1(GND_net), 
            .CO(n34574));
    SB_CARRY add_13_add_1_20061_add_1_2 (.CI(GND_net), .I0(n282[0]), .I1(n61[0]), 
            .CO(n34856));
    SB_CARRY add_3231_4 (.CI(n35124), .I0(n12732[1]), .I1(n253), .CO(n35125));
    SB_LUT4 add_3142_16_lut (.I0(GND_net), .I1(n10671[13]), .I2(GND_net), 
            .I3(n34572), .O(n9929[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3142_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3142_16 (.CI(n34572), .I0(n10671[13]), .I1(GND_net), 
            .CO(n34573));
    SB_LUT4 add_3231_3_lut (.I0(GND_net), .I1(n12732[0]), .I2(n180), .I3(n35123), 
            .O(n12157[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3231_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3058_27_lut (.I0(GND_net), .I1(n8049[24]), .I2(GND_net), 
            .I3(n35295), .O(n8019[25])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3058_27_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3062_24_lut (.I0(GND_net), .I1(n8159[21]), .I2(GND_net), 
            .I3(n35394), .O(n8133[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3062_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3142_15_lut (.I0(GND_net), .I1(n10671[12]), .I2(GND_net), 
            .I3(n34571), .O(n9929[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3142_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3142_15 (.CI(n34571), .I0(n10671[12]), .I1(GND_net), 
            .CO(n34572));
    SB_CARRY add_3231_3 (.CI(n35123), .I0(n12732[0]), .I1(n180), .CO(n35124));
    SB_LUT4 add_3142_14_lut (.I0(GND_net), .I1(n10671[11]), .I2(GND_net), 
            .I3(n34570), .O(n9929[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3142_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3142_14 (.CI(n34570), .I0(n10671[11]), .I1(GND_net), 
            .CO(n34571));
    SB_LUT4 add_3231_2_lut (.I0(GND_net), .I1(n35), .I2(n107), .I3(GND_net), 
            .O(n12157[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3231_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3058_27 (.CI(n35295), .I0(n8049[24]), .I1(GND_net), .CO(n35296));
    SB_LUT4 add_3142_13_lut (.I0(GND_net), .I1(n10671[10]), .I2(GND_net), 
            .I3(n34569), .O(n9929[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3142_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3142_13 (.CI(n34569), .I0(n10671[10]), .I1(GND_net), 
            .CO(n34570));
    SB_CARRY add_3231_2 (.CI(GND_net), .I0(n35), .I1(n107), .CO(n35123));
    SB_LUT4 add_3142_12_lut (.I0(GND_net), .I1(n10671[9]), .I2(GND_net), 
            .I3(n34568), .O(n9929[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3142_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3142_12 (.CI(n34568), .I0(n10671[9]), .I1(GND_net), .CO(n34569));
    SB_LUT4 add_3058_26_lut (.I0(GND_net), .I1(n8049[23]), .I2(GND_net), 
            .I3(n35294), .O(n8019[24])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3058_26_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3062_24 (.CI(n35394), .I0(n8159[21]), .I1(GND_net), .CO(n35395));
    SB_CARRY add_3065_11 (.CI(n35447), .I0(n8231[8]), .I1(GND_net), .CO(n35448));
    SB_LUT4 add_3142_11_lut (.I0(GND_net), .I1(n10671[8]), .I2(GND_net), 
            .I3(n34567), .O(n9929[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3142_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3142_11 (.CI(n34567), .I0(n10671[8]), .I1(GND_net), .CO(n34568));
    SB_LUT4 add_3142_10_lut (.I0(GND_net), .I1(n10671[7]), .I2(GND_net), 
            .I3(n34566), .O(n9929[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3142_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3142_10 (.CI(n34566), .I0(n10671[7]), .I1(GND_net), .CO(n34567));
    SB_CARRY add_3058_26 (.CI(n35294), .I0(n8049[23]), .I1(GND_net), .CO(n35295));
    SB_LUT4 add_3142_9_lut (.I0(GND_net), .I1(n10671[6]), .I2(GND_net), 
            .I3(n34565), .O(n9929[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3142_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3142_9 (.CI(n34565), .I0(n10671[6]), .I1(GND_net), .CO(n34566));
    SB_LUT4 add_3142_8_lut (.I0(GND_net), .I1(n10671[5]), .I2(n692), .I3(n34564), 
            .O(n9929[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3142_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3142_8 (.CI(n34564), .I0(n10671[5]), .I1(n692), .CO(n34565));
    SB_LUT4 add_3058_25_lut (.I0(GND_net), .I1(n8049[22]), .I2(GND_net), 
            .I3(n35293), .O(n8019[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3058_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3062_23_lut (.I0(GND_net), .I1(n8159[20]), .I2(GND_net), 
            .I3(n35393), .O(n8133[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3062_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3142_7_lut (.I0(GND_net), .I1(n10671[4]), .I2(n595), .I3(n34563), 
            .O(n9929[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3142_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3142_7 (.CI(n34563), .I0(n10671[4]), .I1(n595), .CO(n34564));
    SB_LUT4 add_3142_6_lut (.I0(GND_net), .I1(n10671[3]), .I2(n498), .I3(n34562), 
            .O(n9929[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3142_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3062_23 (.CI(n35393), .I0(n8159[20]), .I1(GND_net), .CO(n35394));
    SB_CARRY add_3058_25 (.CI(n35293), .I0(n8049[22]), .I1(GND_net), .CO(n35294));
    SB_CARRY add_3294_17 (.CI(n34384), .I0(n14035[14]), .I1(GND_net), 
            .CO(n34385));
    SB_CARRY state_23__I_0_add_2_14 (.CI(n34227), .I0(\motor_state[12] ), 
            .I1(n58[12]), .CO(n34228));
    SB_LUT4 add_3058_24_lut (.I0(GND_net), .I1(n8049[21]), .I2(GND_net), 
            .I3(n35292), .O(n8019[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3058_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3294_16_lut (.I0(GND_net), .I1(n14035[13]), .I2(GND_net), 
            .I3(n34383), .O(n13594[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3294_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 state_23__I_0_add_2_13_lut (.I0(GND_net), .I1(\motor_state[11] ), 
            .I2(n58[11]), .I3(n34226), .O(\PID_CONTROLLER.err_31__N_2825 [11])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY state_23__I_0_add_2_13 (.CI(n34226), .I0(\motor_state[11] ), 
            .I1(n58[11]), .CO(n34227));
    SB_LUT4 state_23__I_0_add_2_12_lut (.I0(GND_net), .I1(\motor_state[10] ), 
            .I2(n58[10]), .I3(n34225), .O(\PID_CONTROLLER.err_31__N_2825 [10])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3294_16 (.CI(n34383), .I0(n14035[13]), .I1(GND_net), 
            .CO(n34384));
    SB_LUT4 add_3294_15_lut (.I0(GND_net), .I1(n14035[12]), .I2(GND_net), 
            .I3(n34382), .O(n13594[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3294_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3294_15 (.CI(n34382), .I0(n14035[12]), .I1(GND_net), 
            .CO(n34383));
    SB_CARRY state_23__I_0_add_2_12 (.CI(n34225), .I0(\motor_state[10] ), 
            .I1(n58[10]), .CO(n34226));
    SB_CARRY add_3142_6 (.CI(n34562), .I0(n10671[3]), .I1(n498), .CO(n34563));
    SB_LUT4 add_3294_14_lut (.I0(GND_net), .I1(n14035[11]), .I2(GND_net), 
            .I3(n34381), .O(n13594[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3294_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 state_23__I_0_add_2_11_lut (.I0(GND_net), .I1(\motor_state[9] ), 
            .I2(n58[9]), .I3(n34224), .O(\PID_CONTROLLER.err_31__N_2825 [9])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3294_14 (.CI(n34381), .I0(n14035[11]), .I1(GND_net), 
            .CO(n34382));
    SB_LUT4 add_3065_10_lut (.I0(GND_net), .I1(n8231[7]), .I2(GND_net), 
            .I3(n35446), .O(n8208[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3065_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3062_22_lut (.I0(GND_net), .I1(n8159[19]), .I2(GND_net), 
            .I3(n35392), .O(n8133[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3062_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3058_24 (.CI(n35292), .I0(n8049[21]), .I1(GND_net), .CO(n35293));
    SB_LUT4 add_3058_23_lut (.I0(GND_net), .I1(n8049[20]), .I2(GND_net), 
            .I3(n35291), .O(n8019[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3058_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY state_23__I_0_add_2_11 (.CI(n34224), .I0(\motor_state[9] ), 
            .I1(n58[9]), .CO(n34225));
    SB_LUT4 add_3142_5_lut (.I0(GND_net), .I1(n10671[2]), .I2(n401), .I3(n34561), 
            .O(n9929[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3142_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 state_23__I_0_add_2_10_lut (.I0(GND_net), .I1(\motor_state[8] ), 
            .I2(n58[8]), .I3(n34223), .O(\PID_CONTROLLER.err_31__N_2825 [8])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY state_23__I_0_add_2_10 (.CI(n34223), .I0(\motor_state[8] ), 
            .I1(n58[8]), .CO(n34224));
    SB_LUT4 mult_12_i341_2_lut (.I0(\Kd[5] ), .I1(n57[7]), .I2(GND_net), 
            .I3(GND_net), .O(n507));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i341_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_3142_5 (.CI(n34561), .I0(n10671[2]), .I1(n401), .CO(n34562));
    SB_LUT4 add_3067_11_lut (.I0(GND_net), .I1(n8274[8]), .I2(GND_net), 
            .I3(n35486), .O(n8253[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3067_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3065_10 (.CI(n35446), .I0(n8231[7]), .I1(GND_net), .CO(n35447));
    SB_CARRY add_3062_22 (.CI(n35392), .I0(n8159[19]), .I1(GND_net), .CO(n35393));
    SB_CARRY add_3058_23 (.CI(n35291), .I0(n8049[20]), .I1(GND_net), .CO(n35292));
    SB_LUT4 add_3294_13_lut (.I0(GND_net), .I1(n14035[10]), .I2(GND_net), 
            .I3(n34380), .O(n13594[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3294_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3294_13 (.CI(n34380), .I0(n14035[10]), .I1(GND_net), 
            .CO(n34381));
    SB_LUT4 state_23__I_0_add_2_9_lut (.I0(GND_net), .I1(\motor_state[7] ), 
            .I2(n58[7]), .I3(n34222), .O(\PID_CONTROLLER.err_31__N_2825 [7])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3058_22_lut (.I0(GND_net), .I1(n8049[19]), .I2(GND_net), 
            .I3(n35290), .O(n8019[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3058_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3294_12_lut (.I0(GND_net), .I1(n14035[9]), .I2(GND_net), 
            .I3(n34379), .O(n13594[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3294_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3294_12 (.CI(n34379), .I0(n14035[9]), .I1(GND_net), .CO(n34380));
    SB_LUT4 add_3294_11_lut (.I0(GND_net), .I1(n14035[8]), .I2(GND_net), 
            .I3(n34378), .O(n13594[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3294_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3058_22 (.CI(n35290), .I0(n8049[19]), .I1(GND_net), .CO(n35291));
    SB_LUT4 mult_12_i406_2_lut (.I0(\Kd[6] ), .I1(n57[7]), .I2(GND_net), 
            .I3(GND_net), .O(n604));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i406_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_3058_21_lut (.I0(GND_net), .I1(n8049[18]), .I2(GND_net), 
            .I3(n35289), .O(n8019[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3058_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3294_11 (.CI(n34378), .I0(n14035[8]), .I1(GND_net), .CO(n34379));
    SB_CARRY state_23__I_0_add_2_9 (.CI(n34222), .I0(\motor_state[7] ), 
            .I1(n58[7]), .CO(n34223));
    SB_LUT4 add_3294_10_lut (.I0(GND_net), .I1(n14035[7]), .I2(GND_net), 
            .I3(n34377), .O(n13594[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3294_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3142_4_lut (.I0(GND_net), .I1(n10671[1]), .I2(n304_adj_3378), 
            .I3(n34560), .O(n9929[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3142_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3142_4 (.CI(n34560), .I0(n10671[1]), .I1(n304_adj_3378), 
            .CO(n34561));
    SB_LUT4 add_3142_3_lut (.I0(GND_net), .I1(n10671[0]), .I2(n207_adj_3379), 
            .I3(n34559), .O(n9929[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3142_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 state_23__I_0_add_2_8_lut (.I0(GND_net), .I1(\motor_state[6] ), 
            .I2(n58[6]), .I3(n34221), .O(\PID_CONTROLLER.err_31__N_2825 [6])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3065_9_lut (.I0(GND_net), .I1(n8231[6]), .I2(GND_net), 
            .I3(n35445), .O(n8208[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3065_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY state_23__I_0_add_2_8 (.CI(n34221), .I0(\motor_state[6] ), 
            .I1(n58[6]), .CO(n34222));
    SB_CARRY add_3142_3 (.CI(n34559), .I0(n10671[0]), .I1(n207_adj_3379), 
            .CO(n34560));
    SB_CARRY add_3294_10 (.CI(n34377), .I0(n14035[7]), .I1(GND_net), .CO(n34378));
    SB_LUT4 mult_12_i87_2_lut (.I0(\Kd[1] ), .I1(n57[10]), .I2(GND_net), 
            .I3(GND_net), .O(n128));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i87_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_3294_9_lut (.I0(GND_net), .I1(n14035[6]), .I2(GND_net), 
            .I3(n34376), .O(n13594[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3294_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 state_23__I_0_add_2_7_lut (.I0(GND_net), .I1(\motor_state[5] ), 
            .I2(n58[5]), .I3(n34220), .O(\PID_CONTROLLER.err_31__N_2825 [5])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3294_9 (.CI(n34376), .I0(n14035[6]), .I1(GND_net), .CO(n34377));
    SB_CARRY state_23__I_0_add_2_7 (.CI(n34220), .I0(\motor_state[5] ), 
            .I1(n58[5]), .CO(n34221));
    SB_LUT4 mult_12_i24_2_lut (.I0(\Kd[0] ), .I1(n57[11]), .I2(GND_net), 
            .I3(GND_net), .O(n35_adj_3381));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i24_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_3062_21_lut (.I0(GND_net), .I1(n8159[18]), .I2(GND_net), 
            .I3(n35391), .O(n8133[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3062_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3058_21 (.CI(n35289), .I0(n8049[18]), .I1(GND_net), .CO(n35290));
    SB_LUT4 add_3294_8_lut (.I0(GND_net), .I1(n14035[5]), .I2(n710), .I3(n34375), 
            .O(n13594[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3294_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3294_8 (.CI(n34375), .I0(n14035[5]), .I1(n710), .CO(n34376));
    SB_LUT4 add_3294_7_lut (.I0(GND_net), .I1(n14035[4]), .I2(n613), .I3(n34374), 
            .O(n13594[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3294_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3294_7 (.CI(n34374), .I0(n14035[4]), .I1(n613), .CO(n34375));
    SB_CARRY add_3062_21 (.CI(n35391), .I0(n8159[18]), .I1(GND_net), .CO(n35392));
    SB_LUT4 add_3294_6_lut (.I0(GND_net), .I1(n14035[3]), .I2(n516), .I3(n34373), 
            .O(n13594[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3294_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3058_20_lut (.I0(GND_net), .I1(n8049[17]), .I2(GND_net), 
            .I3(n35288), .O(n8019[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3058_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3294_6 (.CI(n34373), .I0(n14035[3]), .I1(n516), .CO(n34374));
    SB_LUT4 state_23__I_0_add_2_6_lut (.I0(GND_net), .I1(\motor_state[4] ), 
            .I2(n58[4]), .I3(n34219), .O(\PID_CONTROLLER.err_31__N_2825 [4])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3294_5_lut (.I0(GND_net), .I1(n14035[2]), .I2(n419), .I3(n34372), 
            .O(n13594[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3294_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY state_23__I_0_add_2_6 (.CI(n34219), .I0(\motor_state[4] ), 
            .I1(n58[4]), .CO(n34220));
    SB_CARRY add_3294_5 (.CI(n34372), .I0(n14035[2]), .I1(n419), .CO(n34373));
    SB_LUT4 state_23__I_0_add_2_5_lut (.I0(GND_net), .I1(\motor_state[3] ), 
            .I2(n58[3]), .I3(n34218), .O(\PID_CONTROLLER.err_31__N_2825 [3])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_12_i471_2_lut (.I0(\Kd[7] ), .I1(n57[7]), .I2(GND_net), 
            .I3(GND_net), .O(n701));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i471_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_3294_4_lut (.I0(GND_net), .I1(n14035[1]), .I2(n322), .I3(n34371), 
            .O(n13594[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3294_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY state_23__I_0_add_2_5 (.CI(n34218), .I0(\motor_state[3] ), 
            .I1(n58[3]), .CO(n34219));
    SB_CARRY add_3065_9 (.CI(n35445), .I0(n8231[6]), .I1(GND_net), .CO(n35446));
    SB_LUT4 add_3062_20_lut (.I0(GND_net), .I1(n8159[17]), .I2(GND_net), 
            .I3(n35390), .O(n8133[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3062_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3058_20 (.CI(n35288), .I0(n8049[17]), .I1(GND_net), .CO(n35289));
    SB_CARRY add_3294_4 (.CI(n34371), .I0(n14035[1]), .I1(n322), .CO(n34372));
    SB_LUT4 state_23__I_0_add_2_4_lut (.I0(GND_net), .I1(\motor_state[2] ), 
            .I2(n58[2]), .I3(n34217), .O(\PID_CONTROLLER.err_31__N_2825 [2])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3294_3_lut (.I0(GND_net), .I1(n14035[0]), .I2(n225), .I3(n34370), 
            .O(n13594[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3294_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY state_23__I_0_add_2_4 (.CI(n34217), .I0(\motor_state[2] ), 
            .I1(n58[2]), .CO(n34218));
    SB_CARRY add_3294_3 (.CI(n34370), .I0(n14035[0]), .I1(n225), .CO(n34371));
    SB_LUT4 mult_12_i152_2_lut (.I0(\Kd[2] ), .I1(n57[10]), .I2(GND_net), 
            .I3(GND_net), .O(n225_adj_3382));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i152_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 state_23__I_0_add_2_3_lut (.I0(GND_net), .I1(\motor_state[1] ), 
            .I2(n58[1]), .I3(n34216), .O(\PID_CONTROLLER.err_31__N_2825 [1])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3058_19_lut (.I0(GND_net), .I1(n8049[16]), .I2(GND_net), 
            .I3(n35287), .O(n8019[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3058_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3294_2_lut (.I0(GND_net), .I1(n35_adj_3383), .I2(n128_adj_3384), 
            .I3(GND_net), .O(n13594[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3294_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i493_2_lut (.I0(\Kp[7] ), .I1(\PID_CONTROLLER.err[18] ), 
            .I2(GND_net), .I3(GND_net), .O(n734));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i493_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY state_23__I_0_add_2_3 (.CI(n34216), .I0(\motor_state[1] ), 
            .I1(n58[1]), .CO(n34217));
    SB_CARRY add_3058_19 (.CI(n35287), .I0(n8049[16]), .I1(GND_net), .CO(n35288));
    SB_CARRY add_3294_2 (.CI(GND_net), .I0(n35_adj_3383), .I1(n128_adj_3384), 
            .CO(n34370));
    SB_LUT4 state_23__I_0_add_2_2_lut (.I0(GND_net), .I1(\motor_state[0] ), 
            .I2(n58[0]), .I3(VCC_net), .O(\PID_CONTROLLER.err_31__N_2825 [0])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY state_23__I_0_add_2_2 (.CI(VCC_net), .I0(\motor_state[0] ), 
            .I1(n58[0]), .CO(n34216));
    SB_LUT4 add_3464_11_lut (.I0(GND_net), .I1(n16505[8]), .I2(GND_net), 
            .I3(n34369), .O(n16420[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3464_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_11_add_2_27_lut (.I0(GND_net), .I1(\PID_CONTROLLER.err_prev[31] ), 
            .I2(n64[26]), .I3(n34215), .O(n57[25])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_11_add_2_27_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_11_add_2_26_lut (.I0(GND_net), .I1(\PID_CONTROLLER.err_prev[31] ), 
            .I2(n64[26]), .I3(n34214), .O(n57[24])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_11_add_2_26_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3464_10_lut (.I0(GND_net), .I1(n16505[7]), .I2(GND_net), 
            .I3(n34368), .O(n16420[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3464_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_11_add_2_26 (.CI(n34214), .I0(\PID_CONTROLLER.err_prev[31] ), 
            .I1(n64[26]), .CO(n34215));
    SB_LUT4 sub_11_add_2_25_lut (.I0(GND_net), .I1(\PID_CONTROLLER.err_prev[23] ), 
            .I2(n64[23]), .I3(n34213), .O(n57[23])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_11_add_2_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3464_10 (.CI(n34368), .I0(n16505[7]), .I1(GND_net), .CO(n34369));
    SB_CARRY sub_11_add_2_25 (.CI(n34213), .I0(\PID_CONTROLLER.err_prev[23] ), 
            .I1(n64[23]), .CO(n34214));
    SB_LUT4 sub_11_add_2_24_lut (.I0(GND_net), .I1(\PID_CONTROLLER.err_prev[22] ), 
            .I2(n64[22]), .I3(n34212), .O(n57[22])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_11_add_2_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3062_20 (.CI(n35390), .I0(n8159[17]), .I1(GND_net), .CO(n35391));
    SB_LUT4 add_3058_18_lut (.I0(GND_net), .I1(n8049[15]), .I2(GND_net), 
            .I3(n35286), .O(n8019[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3058_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3464_9_lut (.I0(GND_net), .I1(n16505[6]), .I2(GND_net), 
            .I3(n34367), .O(n16420[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3464_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_11_add_2_24 (.CI(n34212), .I0(\PID_CONTROLLER.err_prev[22] ), 
            .I1(n64[22]), .CO(n34213));
    SB_CARRY add_3464_9 (.CI(n34367), .I0(n16505[6]), .I1(GND_net), .CO(n34368));
    SB_LUT4 mult_12_i481_2_lut (.I0(\Kd[7] ), .I1(n57[12]), .I2(GND_net), 
            .I3(GND_net), .O(n716));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i481_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 sub_11_add_2_23_lut (.I0(GND_net), .I1(\PID_CONTROLLER.err_prev[21] ), 
            .I2(n64[21]), .I3(n34211), .O(n57[21])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_11_add_2_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3464_8_lut (.I0(GND_net), .I1(n16505[5]), .I2(n743), .I3(n34366), 
            .O(n16420[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3464_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_11_add_2_23 (.CI(n34211), .I0(\PID_CONTROLLER.err_prev[21] ), 
            .I1(n64[21]), .CO(n34212));
    SB_LUT4 mult_10_i79_2_lut (.I0(\Kp[1] ), .I1(\PID_CONTROLLER.err[6] ), 
            .I2(GND_net), .I3(GND_net), .O(n116));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i79_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_3058_18 (.CI(n35286), .I0(n8049[15]), .I1(GND_net), .CO(n35287));
    SB_CARRY add_3464_8 (.CI(n34366), .I0(n16505[5]), .I1(n743), .CO(n34367));
    SB_LUT4 sub_11_add_2_22_lut (.I0(GND_net), .I1(\PID_CONTROLLER.err_prev[20] ), 
            .I2(n64[20]), .I3(n34210), .O(n57[20])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_11_add_2_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_11_add_2_22 (.CI(n34210), .I0(\PID_CONTROLLER.err_prev[20] ), 
            .I1(n64[20]), .CO(n34211));
    SB_LUT4 add_3464_7_lut (.I0(GND_net), .I1(n16505[4]), .I2(n646), .I3(n34365), 
            .O(n16420[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3464_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_11_add_2_21_lut (.I0(GND_net), .I1(\PID_CONTROLLER.err_prev[19] ), 
            .I2(n64[19]), .I3(n34209), .O(n57[19])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_11_add_2_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_11_add_2_21 (.CI(n34209), .I0(\PID_CONTROLLER.err_prev[19] ), 
            .I1(n64[19]), .CO(n34210));
    SB_LUT4 mult_10_i16_2_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err[7] ), 
            .I2(GND_net), .I3(GND_net), .O(n23_adj_3389));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i16_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i144_2_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err[6] ), 
            .I2(GND_net), .I3(GND_net), .O(n213));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i144_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i209_2_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err[6] ), 
            .I2(GND_net), .I3(GND_net), .O(n310_adj_3390));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i209_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i274_2_lut (.I0(\Kp[4] ), .I1(\PID_CONTROLLER.err[6] ), 
            .I2(GND_net), .I3(GND_net), .O(n407));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i274_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i331_2_lut (.I0(\Kd[5] ), .I1(n57[2]), .I2(GND_net), 
            .I3(GND_net), .O(n492));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i331_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 sub_11_add_2_20_lut (.I0(GND_net), .I1(\PID_CONTROLLER.err_prev[18] ), 
            .I2(n64[18]), .I3(n34208), .O(n57[18])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_11_add_2_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_11_add_2_20 (.CI(n34208), .I0(\PID_CONTROLLER.err_prev[18] ), 
            .I1(n64[18]), .CO(n34209));
    SB_CARRY add_3464_7 (.CI(n34365), .I0(n16505[4]), .I1(n646), .CO(n34366));
    SB_LUT4 add_3431_14_lut (.I0(GND_net), .I1(n16185[11]), .I2(GND_net), 
            .I3(n35677), .O(n16031[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3431_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3431_13_lut (.I0(GND_net), .I1(n16185[10]), .I2(GND_net), 
            .I3(n35676), .O(n16031[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3431_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3431_13 (.CI(n35676), .I0(n16185[10]), .I1(GND_net), 
            .CO(n35677));
    SB_CARRY add_3074_5 (.CI(n35585), .I0(n8393[2]), .I1(n446), .CO(n35586));
    SB_LUT4 add_3069_17_lut (.I0(GND_net), .I1(n8313[14]), .I2(GND_net), 
            .I3(n35527), .O(n8294[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3069_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3067_11 (.CI(n35486), .I0(n8274[8]), .I1(GND_net), .CO(n35487));
    SB_LUT4 add_3065_8_lut (.I0(GND_net), .I1(n8231[5]), .I2(n710_adj_3392), 
            .I3(n35444), .O(n8208[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3065_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3062_19_lut (.I0(GND_net), .I1(n8159[16]), .I2(GND_net), 
            .I3(n35389), .O(n8133[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3062_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3058_17_lut (.I0(GND_net), .I1(n8049[14]), .I2(GND_net), 
            .I3(n35285), .O(n8019[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3058_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3142_2_lut (.I0(GND_net), .I1(n17_adj_3393), .I2(n110_adj_3394), 
            .I3(GND_net), .O(n9929[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3142_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3142_2 (.CI(GND_net), .I0(n17_adj_3393), .I1(n110_adj_3394), 
            .CO(n34559));
    SB_LUT4 add_3322_13_lut (.I0(GND_net), .I1(n14560[10]), .I2(GND_net), 
            .I3(n34558), .O(n14168[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3322_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3322_12_lut (.I0(GND_net), .I1(n14560[9]), .I2(GND_net), 
            .I3(n34557), .O(n14168[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3322_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3058_17 (.CI(n35285), .I0(n8049[14]), .I1(GND_net), .CO(n35286));
    SB_CARRY add_3322_12 (.CI(n34557), .I0(n14560[9]), .I1(GND_net), .CO(n34558));
    SB_LUT4 add_3322_11_lut (.I0(GND_net), .I1(n14560[8]), .I2(GND_net), 
            .I3(n34556), .O(n14168[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3322_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3322_11 (.CI(n34556), .I0(n14560[8]), .I1(GND_net), .CO(n34557));
    SB_LUT4 add_3322_10_lut (.I0(GND_net), .I1(n14560[7]), .I2(GND_net), 
            .I3(n34555), .O(n14168[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3322_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3062_19 (.CI(n35389), .I0(n8159[16]), .I1(GND_net), .CO(n35390));
    SB_LUT4 add_3058_16_lut (.I0(GND_net), .I1(n8049[13]), .I2(GND_net), 
            .I3(n35284), .O(n8019[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3058_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3322_10 (.CI(n34555), .I0(n14560[7]), .I1(GND_net), .CO(n34556));
    SB_LUT4 add_3322_9_lut (.I0(GND_net), .I1(n14560[6]), .I2(GND_net), 
            .I3(n34554), .O(n14168[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3322_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3322_9 (.CI(n34554), .I0(n14560[6]), .I1(GND_net), .CO(n34555));
    SB_LUT4 add_3322_8_lut (.I0(GND_net), .I1(n14560[5]), .I2(n545), .I3(n34553), 
            .O(n14168[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3322_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3058_16 (.CI(n35284), .I0(n8049[13]), .I1(GND_net), .CO(n35285));
    SB_CARRY add_3322_8 (.CI(n34553), .I0(n14560[5]), .I1(n545), .CO(n34554));
    SB_LUT4 add_3322_7_lut (.I0(GND_net), .I1(n14560[4]), .I2(n472), .I3(n34552), 
            .O(n14168[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3322_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3322_7 (.CI(n34552), .I0(n14560[4]), .I1(n472), .CO(n34553));
    SB_LUT4 add_3322_6_lut (.I0(GND_net), .I1(n14560[3]), .I2(n399), .I3(n34551), 
            .O(n14168[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3322_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3065_8 (.CI(n35444), .I0(n8231[5]), .I1(n710_adj_3392), 
            .CO(n35445));
    SB_LUT4 add_3062_18_lut (.I0(GND_net), .I1(n8159[15]), .I2(GND_net), 
            .I3(n35388), .O(n8133[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3062_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3058_15_lut (.I0(GND_net), .I1(n8049[12]), .I2(GND_net), 
            .I3(n35283), .O(n8019[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3058_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3322_6 (.CI(n34551), .I0(n14560[3]), .I1(n399), .CO(n34552));
    SB_LUT4 add_3464_6_lut (.I0(GND_net), .I1(n16505[3]), .I2(n549), .I3(n34364), 
            .O(n16420[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3464_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3322_5_lut (.I0(GND_net), .I1(n14560[2]), .I2(n326), .I3(n34550), 
            .O(n14168[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3322_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3322_5 (.CI(n34550), .I0(n14560[2]), .I1(n326), .CO(n34551));
    SB_LUT4 sub_11_add_2_19_lut (.I0(GND_net), .I1(\PID_CONTROLLER.err_prev[17] ), 
            .I2(n64[17]), .I3(n34207), .O(n57[17])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_11_add_2_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3074_4_lut (.I0(GND_net), .I1(n8393[1]), .I2(n349), .I3(n35584), 
            .O(n8379[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3074_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3464_6 (.CI(n34364), .I0(n16505[3]), .I1(n549), .CO(n34365));
    SB_CARRY add_3058_15 (.CI(n35283), .I0(n8049[12]), .I1(GND_net), .CO(n35284));
    SB_LUT4 add_3322_4_lut (.I0(GND_net), .I1(n14560[1]), .I2(n253), .I3(n34549), 
            .O(n14168[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3322_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3322_4 (.CI(n34549), .I0(n14560[1]), .I1(n253), .CO(n34550));
    SB_LUT4 add_3322_3_lut (.I0(GND_net), .I1(n14560[0]), .I2(n180), .I3(n34548), 
            .O(n14168[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3322_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3062_18 (.CI(n35388), .I0(n8159[15]), .I1(GND_net), .CO(n35389));
    SB_LUT4 add_3058_14_lut (.I0(GND_net), .I1(n8049[11]), .I2(GND_net), 
            .I3(n35282), .O(n8019[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3058_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3322_3 (.CI(n34548), .I0(n14560[0]), .I1(n180), .CO(n34549));
    SB_LUT4 add_3322_2_lut (.I0(GND_net), .I1(n35), .I2(n107), .I3(GND_net), 
            .O(n14168[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3322_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3322_2 (.CI(GND_net), .I0(n35), .I1(n107), .CO(n34548));
    SB_LUT4 add_3170_27_lut (.I0(GND_net), .I1(n11358[24]), .I2(GND_net), 
            .I3(n34547), .O(n10671[25])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3170_27_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3058_14 (.CI(n35282), .I0(n8049[11]), .I1(GND_net), .CO(n35283));
    SB_LUT4 add_3170_26_lut (.I0(GND_net), .I1(n11358[23]), .I2(GND_net), 
            .I3(n34546), .O(n10671[24])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3170_26_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3170_26 (.CI(n34546), .I0(n11358[23]), .I1(GND_net), 
            .CO(n34547));
    SB_CARRY sub_11_add_2_19 (.CI(n34207), .I0(\PID_CONTROLLER.err_prev[17] ), 
            .I1(n64[17]), .CO(n34208));
    SB_LUT4 add_3170_25_lut (.I0(GND_net), .I1(n11358[22]), .I2(GND_net), 
            .I3(n34545), .O(n10671[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3170_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3170_25 (.CI(n34545), .I0(n11358[22]), .I1(GND_net), 
            .CO(n34546));
    SB_LUT4 add_3067_10_lut (.I0(GND_net), .I1(n8274[7]), .I2(GND_net), 
            .I3(n35485), .O(n8253[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3067_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3065_7_lut (.I0(GND_net), .I1(n8231[4]), .I2(n613_adj_3396), 
            .I3(n35443), .O(n8208[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3065_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3062_17_lut (.I0(GND_net), .I1(n8159[14]), .I2(GND_net), 
            .I3(n35387), .O(n8133[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3062_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3058_13_lut (.I0(GND_net), .I1(n8049[10]), .I2(GND_net), 
            .I3(n35281), .O(n8019[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3058_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3170_24_lut (.I0(GND_net), .I1(n11358[21]), .I2(GND_net), 
            .I3(n34544), .O(n10671[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3170_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3170_24 (.CI(n34544), .I0(n11358[21]), .I1(GND_net), 
            .CO(n34545));
    SB_LUT4 add_3170_23_lut (.I0(GND_net), .I1(n11358[20]), .I2(GND_net), 
            .I3(n34543), .O(n10671[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3170_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3170_23 (.CI(n34543), .I0(n11358[20]), .I1(GND_net), 
            .CO(n34544));
    SB_CARRY add_3058_13 (.CI(n35281), .I0(n8049[10]), .I1(GND_net), .CO(n35282));
    SB_LUT4 add_3170_22_lut (.I0(GND_net), .I1(n11358[19]), .I2(GND_net), 
            .I3(n34542), .O(n10671[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3170_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i339_2_lut (.I0(\Kp[5] ), .I1(\PID_CONTROLLER.err[6] ), 
            .I2(GND_net), .I3(GND_net), .O(n504));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i339_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_3170_22 (.CI(n34542), .I0(n11358[19]), .I1(GND_net), 
            .CO(n34543));
    SB_LUT4 add_3170_21_lut (.I0(GND_net), .I1(n11358[18]), .I2(GND_net), 
            .I3(n34541), .O(n10671[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3170_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3170_21 (.CI(n34541), .I0(n11358[18]), .I1(GND_net), 
            .CO(n34542));
    SB_CARRY add_3062_17 (.CI(n35387), .I0(n8159[14]), .I1(GND_net), .CO(n35388));
    SB_LUT4 add_3058_12_lut (.I0(GND_net), .I1(n8049[9]), .I2(GND_net), 
            .I3(n35280), .O(n8019[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3058_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3170_20_lut (.I0(GND_net), .I1(n11358[17]), .I2(GND_net), 
            .I3(n34540), .O(n10671[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3170_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3170_20 (.CI(n34540), .I0(n11358[17]), .I1(GND_net), 
            .CO(n34541));
    SB_LUT4 add_3170_19_lut (.I0(GND_net), .I1(n11358[16]), .I2(GND_net), 
            .I3(n34539), .O(n10671[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3170_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3170_19 (.CI(n34539), .I0(n11358[16]), .I1(GND_net), 
            .CO(n34540));
    SB_CARRY add_3058_12 (.CI(n35280), .I0(n8049[9]), .I1(GND_net), .CO(n35281));
    SB_LUT4 add_3170_18_lut (.I0(GND_net), .I1(n11358[15]), .I2(GND_net), 
            .I3(n34538), .O(n10671[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3170_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3170_18 (.CI(n34538), .I0(n11358[15]), .I1(GND_net), 
            .CO(n34539));
    SB_LUT4 add_3170_17_lut (.I0(GND_net), .I1(n11358[14]), .I2(GND_net), 
            .I3(n34537), .O(n10671[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3170_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3170_17 (.CI(n34537), .I0(n11358[14]), .I1(GND_net), 
            .CO(n34538));
    SB_CARRY add_3065_7 (.CI(n35443), .I0(n8231[4]), .I1(n613_adj_3396), 
            .CO(n35444));
    SB_LUT4 add_3062_16_lut (.I0(GND_net), .I1(n8159[13]), .I2(GND_net), 
            .I3(n35386), .O(n8133[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3062_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3058_11_lut (.I0(GND_net), .I1(n8049[8]), .I2(GND_net), 
            .I3(n35279), .O(n8019[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3058_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3170_16_lut (.I0(GND_net), .I1(n11358[13]), .I2(GND_net), 
            .I3(n34536), .O(n10671[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3170_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3170_16 (.CI(n34536), .I0(n11358[13]), .I1(GND_net), 
            .CO(n34537));
    SB_LUT4 mult_10_i404_2_lut (.I0(\Kp[6] ), .I1(\PID_CONTROLLER.err[6] ), 
            .I2(GND_net), .I3(GND_net), .O(n601));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i404_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_3170_15_lut (.I0(GND_net), .I1(n11358[12]), .I2(GND_net), 
            .I3(n34535), .O(n10671[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3170_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3170_15 (.CI(n34535), .I0(n11358[12]), .I1(GND_net), 
            .CO(n34536));
    SB_CARRY add_3058_11 (.CI(n35279), .I0(n8049[8]), .I1(GND_net), .CO(n35280));
    SB_LUT4 add_3170_14_lut (.I0(GND_net), .I1(n11358[11]), .I2(GND_net), 
            .I3(n34534), .O(n10671[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3170_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3170_14 (.CI(n34534), .I0(n11358[11]), .I1(GND_net), 
            .CO(n34535));
    SB_LUT4 add_3170_13_lut (.I0(GND_net), .I1(n11358[10]), .I2(GND_net), 
            .I3(n34533), .O(n10671[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3170_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3170_13 (.CI(n34533), .I0(n11358[10]), .I1(GND_net), 
            .CO(n34534));
    SB_CARRY add_3062_16 (.CI(n35386), .I0(n8159[13]), .I1(GND_net), .CO(n35387));
    SB_LUT4 add_3058_10_lut (.I0(GND_net), .I1(n8049[7]), .I2(GND_net), 
            .I3(n35278), .O(n8019[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3058_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3170_12_lut (.I0(GND_net), .I1(n11358[9]), .I2(GND_net), 
            .I3(n34532), .O(n10671[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3170_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3170_12 (.CI(n34532), .I0(n11358[9]), .I1(GND_net), .CO(n34533));
    SB_LUT4 add_3170_11_lut (.I0(GND_net), .I1(n11358[8]), .I2(GND_net), 
            .I3(n34531), .O(n10671[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3170_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3170_11 (.CI(n34531), .I0(n11358[8]), .I1(GND_net), .CO(n34532));
    SB_CARRY add_3058_10 (.CI(n35278), .I0(n8049[7]), .I1(GND_net), .CO(n35279));
    SB_LUT4 add_3170_10_lut (.I0(GND_net), .I1(n11358[7]), .I2(GND_net), 
            .I3(n34530), .O(n10671[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3170_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i469_2_lut (.I0(\Kp[7] ), .I1(\PID_CONTROLLER.err[6] ), 
            .I2(GND_net), .I3(GND_net), .O(n698));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i469_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_3170_10 (.CI(n34530), .I0(n11358[7]), .I1(GND_net), .CO(n34531));
    SB_LUT4 add_3170_9_lut (.I0(GND_net), .I1(n11358[6]), .I2(GND_net), 
            .I3(n34529), .O(n10671[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3170_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3170_9 (.CI(n34529), .I0(n11358[6]), .I1(GND_net), .CO(n34530));
    SB_CARRY add_3069_17 (.CI(n35527), .I0(n8313[14]), .I1(GND_net), .CO(n35528));
    SB_CARRY add_3067_10 (.CI(n35485), .I0(n8274[7]), .I1(GND_net), .CO(n35486));
    SB_LUT4 add_3065_6_lut (.I0(GND_net), .I1(n8231[3]), .I2(n516_adj_3397), 
            .I3(n35442), .O(n8208[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3065_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3062_15_lut (.I0(GND_net), .I1(n8159[12]), .I2(GND_net), 
            .I3(n35385), .O(n8133[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3062_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3058_9_lut (.I0(GND_net), .I1(n8049[6]), .I2(GND_net), 
            .I3(n35277), .O(n8019[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3058_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3170_8_lut (.I0(GND_net), .I1(n11358[5]), .I2(n695), .I3(n34528), 
            .O(n10671[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3170_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3170_8 (.CI(n34528), .I0(n11358[5]), .I1(n695), .CO(n34529));
    SB_LUT4 sub_11_add_2_18_lut (.I0(GND_net), .I1(\PID_CONTROLLER.err_prev[16] ), 
            .I2(n64[16]), .I3(n34206), .O(n57[16])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_11_add_2_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3170_7_lut (.I0(GND_net), .I1(n11358[4]), .I2(n598), .I3(n34527), 
            .O(n10671[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3170_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3170_7 (.CI(n34527), .I0(n11358[4]), .I1(n598), .CO(n34528));
    SB_CARRY add_3058_9 (.CI(n35277), .I0(n8049[6]), .I1(GND_net), .CO(n35278));
    SB_LUT4 add_3170_6_lut (.I0(GND_net), .I1(n11358[3]), .I2(n501), .I3(n34526), 
            .O(n10671[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3170_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3170_6 (.CI(n34526), .I0(n11358[3]), .I1(n501), .CO(n34527));
    SB_LUT4 add_3170_5_lut (.I0(GND_net), .I1(n11358[2]), .I2(n404), .I3(n34525), 
            .O(n10671[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3170_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3170_5 (.CI(n34525), .I0(n11358[2]), .I1(n404), .CO(n34526));
    SB_CARRY add_3062_15 (.CI(n35385), .I0(n8159[12]), .I1(GND_net), .CO(n35386));
    SB_LUT4 add_3058_8_lut (.I0(GND_net), .I1(n8049[5]), .I2(n689), .I3(n35276), 
            .O(n8019[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3058_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3170_4_lut (.I0(GND_net), .I1(n11358[1]), .I2(n307_adj_3399), 
            .I3(n34524), .O(n10671[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3170_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3170_4 (.CI(n34524), .I0(n11358[1]), .I1(n307_adj_3399), 
            .CO(n34525));
    SB_LUT4 add_3170_3_lut (.I0(GND_net), .I1(n11358[0]), .I2(n210), .I3(n34523), 
            .O(n10671[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3170_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3170_3 (.CI(n34523), .I0(n11358[0]), .I1(n210), .CO(n34524));
    SB_CARRY add_3058_8 (.CI(n35276), .I0(n8049[5]), .I1(n689), .CO(n35277));
    SB_LUT4 add_3170_2_lut (.I0(GND_net), .I1(n20_adj_3400), .I2(n113), 
            .I3(GND_net), .O(n10671[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3170_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3170_2 (.CI(GND_net), .I0(n20_adj_3400), .I1(n113), .CO(n34523));
    SB_LUT4 add_3342_12_lut (.I0(GND_net), .I1(n14912[9]), .I2(GND_net), 
            .I3(n34522), .O(n14560[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3342_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3342_11_lut (.I0(GND_net), .I1(n14912[8]), .I2(GND_net), 
            .I3(n34521), .O(n14560[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3342_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3065_6 (.CI(n35442), .I0(n8231[3]), .I1(n516_adj_3397), 
            .CO(n35443));
    SB_LUT4 add_3062_14_lut (.I0(GND_net), .I1(n8159[11]), .I2(GND_net), 
            .I3(n35384), .O(n8133[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3062_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3058_7_lut (.I0(GND_net), .I1(n8049[4]), .I2(n592), .I3(n35275), 
            .O(n8019[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3058_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3342_11 (.CI(n34521), .I0(n14912[8]), .I1(GND_net), .CO(n34522));
    SB_LUT4 add_3342_10_lut (.I0(GND_net), .I1(n14912[7]), .I2(GND_net), 
            .I3(n34520), .O(n14560[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3342_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3342_10 (.CI(n34520), .I0(n14912[7]), .I1(GND_net), .CO(n34521));
    SB_LUT4 add_3342_9_lut (.I0(GND_net), .I1(n14912[6]), .I2(GND_net), 
            .I3(n34519), .O(n14560[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3342_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3058_7 (.CI(n35275), .I0(n8049[4]), .I1(n592), .CO(n35276));
    SB_CARRY add_3342_9 (.CI(n34519), .I0(n14912[6]), .I1(GND_net), .CO(n34520));
    SB_LUT4 add_3342_8_lut (.I0(GND_net), .I1(n14912[5]), .I2(n545), .I3(n34518), 
            .O(n14560[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3342_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3342_8 (.CI(n34518), .I0(n14912[5]), .I1(n545), .CO(n34519));
    SB_LUT4 mult_12_i217_2_lut (.I0(\Kd[3] ), .I1(n57[10]), .I2(GND_net), 
            .I3(GND_net), .O(n322_adj_3401));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i217_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_3342_7_lut (.I0(GND_net), .I1(n14912[4]), .I2(n472), .I3(n34517), 
            .O(n14560[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3342_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3062_14 (.CI(n35384), .I0(n8159[11]), .I1(GND_net), .CO(n35385));
    SB_LUT4 add_3058_6_lut (.I0(GND_net), .I1(n8049[3]), .I2(n495), .I3(n35274), 
            .O(n8019[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3058_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3342_7 (.CI(n34517), .I0(n14912[4]), .I1(n472), .CO(n34518));
    SB_LUT4 add_3342_6_lut (.I0(GND_net), .I1(n14912[3]), .I2(n399), .I3(n34516), 
            .O(n14560[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3342_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3342_6 (.CI(n34516), .I0(n14912[3]), .I1(n399), .CO(n34517));
    SB_LUT4 add_3342_5_lut (.I0(GND_net), .I1(n14912[2]), .I2(n326), .I3(n34515), 
            .O(n14560[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3342_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3058_6 (.CI(n35274), .I0(n8049[3]), .I1(n495), .CO(n35275));
    SB_CARRY add_3342_5 (.CI(n34515), .I0(n14912[2]), .I1(n326), .CO(n34516));
    SB_LUT4 add_3342_4_lut (.I0(GND_net), .I1(n14912[1]), .I2(n253), .I3(n34514), 
            .O(n14560[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3342_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3342_4 (.CI(n34514), .I0(n14912[1]), .I1(n253), .CO(n34515));
    SB_LUT4 add_3342_3_lut (.I0(GND_net), .I1(n14912[0]), .I2(n180), .I3(n34513), 
            .O(n14560[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3342_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3067_9_lut (.I0(GND_net), .I1(n8274[6]), .I2(GND_net), 
            .I3(n35484), .O(n8253[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3067_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3065_5_lut (.I0(GND_net), .I1(n8231[2]), .I2(n419_adj_3402), 
            .I3(n35441), .O(n8208[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3065_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3062_13_lut (.I0(GND_net), .I1(n8159[10]), .I2(GND_net), 
            .I3(n35383), .O(n8133[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3062_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_12_i73_2_lut (.I0(\Kd[1] ), .I1(n57[3]), .I2(GND_net), 
            .I3(GND_net), .O(n107_adj_3403));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i73_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_3058_5_lut (.I0(GND_net), .I1(n8049[2]), .I2(n398), .I3(n35273), 
            .O(n8019[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3058_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3342_3 (.CI(n34513), .I0(n14912[0]), .I1(n180), .CO(n34514));
    SB_LUT4 add_3342_2_lut (.I0(GND_net), .I1(n35), .I2(n107), .I3(GND_net), 
            .O(n14560[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3342_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_12_i10_2_lut (.I0(\Kd[0] ), .I1(n57[4]), .I2(GND_net), 
            .I3(GND_net), .O(n14_adj_3404));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i10_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_3342_2 (.CI(GND_net), .I0(n35), .I1(n107), .CO(n34513));
    SB_LUT4 add_3197_26_lut (.I0(GND_net), .I1(n11992[23]), .I2(GND_net), 
            .I3(n34512), .O(n11358[24])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3197_26_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3058_5 (.CI(n35273), .I0(n8049[2]), .I1(n398), .CO(n35274));
    SB_LUT4 mult_12_i138_2_lut (.I0(\Kd[2] ), .I1(n57[3]), .I2(GND_net), 
            .I3(GND_net), .O(n204));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i138_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_3197_25_lut (.I0(GND_net), .I1(n11992[22]), .I2(GND_net), 
            .I3(n34511), .O(n11358[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3197_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3197_25 (.CI(n34511), .I0(n11992[22]), .I1(GND_net), 
            .CO(n34512));
    SB_LUT4 add_3197_24_lut (.I0(GND_net), .I1(n11992[21]), .I2(GND_net), 
            .I3(n34510), .O(n11358[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3197_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3197_24 (.CI(n34510), .I0(n11992[21]), .I1(GND_net), 
            .CO(n34511));
    SB_CARRY add_3062_13 (.CI(n35383), .I0(n8159[10]), .I1(GND_net), .CO(n35384));
    SB_LUT4 add_3058_4_lut (.I0(GND_net), .I1(n8049[1]), .I2(n301), .I3(n35272), 
            .O(n8019[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3058_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3197_23_lut (.I0(GND_net), .I1(n11992[20]), .I2(GND_net), 
            .I3(n34509), .O(n11358[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3197_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3197_23 (.CI(n34509), .I0(n11992[20]), .I1(GND_net), 
            .CO(n34510));
    SB_LUT4 add_3197_22_lut (.I0(GND_net), .I1(n11992[19]), .I2(GND_net), 
            .I3(n34508), .O(n11358[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3197_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3197_22 (.CI(n34508), .I0(n11992[19]), .I1(GND_net), 
            .CO(n34509));
    SB_CARRY add_3058_4 (.CI(n35272), .I0(n8049[1]), .I1(n301), .CO(n35273));
    SB_LUT4 add_3197_21_lut (.I0(GND_net), .I1(n11992[18]), .I2(GND_net), 
            .I3(n34507), .O(n11358[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3197_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3197_21 (.CI(n34507), .I0(n11992[18]), .I1(GND_net), 
            .CO(n34508));
    SB_LUT4 add_3197_20_lut (.I0(GND_net), .I1(n11992[17]), .I2(GND_net), 
            .I3(n34506), .O(n11358[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3197_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3197_20 (.CI(n34506), .I0(n11992[17]), .I1(GND_net), 
            .CO(n34507));
    SB_CARRY add_3065_5 (.CI(n35441), .I0(n8231[2]), .I1(n419_adj_3402), 
            .CO(n35442));
    SB_LUT4 add_3062_12_lut (.I0(GND_net), .I1(n8159[9]), .I2(GND_net), 
            .I3(n35382), .O(n8133[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3062_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3058_3_lut (.I0(GND_net), .I1(n8049[0]), .I2(n204), .I3(n35271), 
            .O(n8019[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3058_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3197_19_lut (.I0(GND_net), .I1(n11992[16]), .I2(GND_net), 
            .I3(n34505), .O(n11358[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3197_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3197_19 (.CI(n34505), .I0(n11992[16]), .I1(GND_net), 
            .CO(n34506));
    SB_LUT4 add_3197_18_lut (.I0(GND_net), .I1(n11992[15]), .I2(GND_net), 
            .I3(n34504), .O(n11358[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3197_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3197_18 (.CI(n34504), .I0(n11992[15]), .I1(GND_net), 
            .CO(n34505));
    SB_CARRY add_3058_3 (.CI(n35271), .I0(n8049[0]), .I1(n204), .CO(n35272));
    SB_LUT4 add_3197_17_lut (.I0(GND_net), .I1(n11992[14]), .I2(GND_net), 
            .I3(n34503), .O(n11358[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3197_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3197_17 (.CI(n34503), .I0(n11992[14]), .I1(GND_net), 
            .CO(n34504));
    SB_LUT4 add_3197_16_lut (.I0(GND_net), .I1(n11992[13]), .I2(GND_net), 
            .I3(n34502), .O(n11358[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3197_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3197_16 (.CI(n34502), .I0(n11992[13]), .I1(GND_net), 
            .CO(n34503));
    SB_CARRY add_3062_12 (.CI(n35382), .I0(n8159[9]), .I1(GND_net), .CO(n35383));
    SB_LUT4 add_3058_2_lut (.I0(GND_net), .I1(n14_adj_3404), .I2(n107_adj_3403), 
            .I3(GND_net), .O(n8019[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3058_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3197_15_lut (.I0(GND_net), .I1(n11992[12]), .I2(GND_net), 
            .I3(n34501), .O(n11358[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3197_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3197_15 (.CI(n34501), .I0(n11992[12]), .I1(GND_net), 
            .CO(n34502));
    SB_LUT4 add_3197_14_lut (.I0(GND_net), .I1(n11992[11]), .I2(GND_net), 
            .I3(n34500), .O(n11358[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3197_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3197_14 (.CI(n34500), .I0(n11992[11]), .I1(GND_net), 
            .CO(n34501));
    SB_CARRY add_3058_2 (.CI(GND_net), .I0(n14_adj_3404), .I1(n107_adj_3403), 
            .CO(n35271));
    SB_LUT4 \PID_CONTROLLER.integral_1017_add_4_11_lut  (.I0(GND_net), .I1(\PID_CONTROLLER.err[9] ), 
            .I2(\PID_CONTROLLER.integral [9]), .I3(n35076), .O(n66[9])) /* synthesis syn_instantiated=1 */ ;
    defparam \PID_CONTROLLER.integral_1017_add_4_11_lut .LUT_INIT = 16'hC33C;
    SB_LUT4 add_3197_13_lut (.I0(GND_net), .I1(n11992[10]), .I2(GND_net), 
            .I3(n34499), .O(n11358[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3197_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3197_13 (.CI(n34499), .I0(n11992[10]), .I1(GND_net), 
            .CO(n34500));
    SB_LUT4 \PID_CONTROLLER.integral_1017_add_4_10_lut  (.I0(GND_net), .I1(\PID_CONTROLLER.err[8] ), 
            .I2(\PID_CONTROLLER.integral [8]), .I3(n35075), .O(n66[8])) /* synthesis syn_instantiated=1 */ ;
    defparam \PID_CONTROLLER.integral_1017_add_4_10_lut .LUT_INIT = 16'hC33C;
    SB_LUT4 add_3197_12_lut (.I0(GND_net), .I1(n11992[9]), .I2(GND_net), 
            .I3(n34498), .O(n11358[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3197_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_12_i203_2_lut (.I0(\Kd[3] ), .I1(n57[3]), .I2(GND_net), 
            .I3(GND_net), .O(n301));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i203_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_3197_12 (.CI(n34498), .I0(n11992[9]), .I1(GND_net), .CO(n34499));
    SB_CARRY add_3074_4 (.CI(n35584), .I0(n8393[1]), .I1(n349), .CO(n35585));
    SB_LUT4 add_3069_16_lut (.I0(GND_net), .I1(n8313[13]), .I2(GND_net), 
            .I3(n35526), .O(n8294[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3069_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3067_9 (.CI(n35484), .I0(n8274[6]), .I1(GND_net), .CO(n35485));
    SB_LUT4 add_3065_4_lut (.I0(GND_net), .I1(n8231[1]), .I2(n322_adj_3401), 
            .I3(n35440), .O(n8208[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3065_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3062_11_lut (.I0(GND_net), .I1(n8159[8]), .I2(GND_net), 
            .I3(n35381), .O(n8133[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3062_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3057_30_lut (.I0(GND_net), .I1(n8019[27]), .I2(GND_net), 
            .I3(n35270), .O(n7988[28])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3057_30_lut.LUT_INIT = 16'hC33C;
    SB_CARRY \PID_CONTROLLER.integral_1017_add_4_10  (.CI(n35075), .I0(\PID_CONTROLLER.err[8] ), 
            .I1(\PID_CONTROLLER.integral [8]), .CO(n35076));
    SB_LUT4 add_3197_11_lut (.I0(GND_net), .I1(n11992[8]), .I2(GND_net), 
            .I3(n34497), .O(n11358[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3197_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3197_11 (.CI(n34497), .I0(n11992[8]), .I1(GND_net), .CO(n34498));
    SB_LUT4 \PID_CONTROLLER.integral_1017_add_4_9_lut  (.I0(GND_net), .I1(\PID_CONTROLLER.err[7] ), 
            .I2(\PID_CONTROLLER.integral [7]), .I3(n35074), .O(n66[7])) /* synthesis syn_instantiated=1 */ ;
    defparam \PID_CONTROLLER.integral_1017_add_4_9_lut .LUT_INIT = 16'hC33C;
    SB_LUT4 add_3197_10_lut (.I0(GND_net), .I1(n11992[7]), .I2(GND_net), 
            .I3(n34496), .O(n11358[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3197_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3197_10 (.CI(n34496), .I0(n11992[7]), .I1(GND_net), .CO(n34497));
    SB_LUT4 add_3057_29_lut (.I0(GND_net), .I1(n8019[26]), .I2(GND_net), 
            .I3(n35269), .O(n7988[27])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3057_29_lut.LUT_INIT = 16'hC33C;
    SB_CARRY \PID_CONTROLLER.integral_1017_add_4_9  (.CI(n35074), .I0(\PID_CONTROLLER.err[7] ), 
            .I1(\PID_CONTROLLER.integral [7]), .CO(n35075));
    SB_LUT4 add_3197_9_lut (.I0(GND_net), .I1(n11992[6]), .I2(GND_net), 
            .I3(n34495), .O(n11358[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3197_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3197_9 (.CI(n34495), .I0(n11992[6]), .I1(GND_net), .CO(n34496));
    SB_LUT4 \PID_CONTROLLER.integral_1017_add_4_8_lut  (.I0(GND_net), .I1(\PID_CONTROLLER.err[6] ), 
            .I2(\PID_CONTROLLER.integral [6]), .I3(n35073), .O(n66[6])) /* synthesis syn_instantiated=1 */ ;
    defparam \PID_CONTROLLER.integral_1017_add_4_8_lut .LUT_INIT = 16'hC33C;
    SB_LUT4 add_3197_8_lut (.I0(GND_net), .I1(n11992[5]), .I2(n698), .I3(n34494), 
            .O(n11358[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3197_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3197_8 (.CI(n34494), .I0(n11992[5]), .I1(n698), .CO(n34495));
    SB_CARRY add_3062_11 (.CI(n35381), .I0(n8159[8]), .I1(GND_net), .CO(n35382));
    SB_CARRY add_3057_29 (.CI(n35269), .I0(n8019[26]), .I1(GND_net), .CO(n35270));
    SB_CARRY \PID_CONTROLLER.integral_1017_add_4_8  (.CI(n35073), .I0(\PID_CONTROLLER.err[6] ), 
            .I1(\PID_CONTROLLER.integral [6]), .CO(n35074));
    SB_LUT4 add_3197_7_lut (.I0(GND_net), .I1(n11992[4]), .I2(n601), .I3(n34493), 
            .O(n11358[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3197_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3197_7 (.CI(n34493), .I0(n11992[4]), .I1(n601), .CO(n34494));
    SB_LUT4 \PID_CONTROLLER.integral_1017_add_4_7_lut  (.I0(GND_net), .I1(\PID_CONTROLLER.err[5] ), 
            .I2(\PID_CONTROLLER.integral [5]), .I3(n35072), .O(n66[5])) /* synthesis syn_instantiated=1 */ ;
    defparam \PID_CONTROLLER.integral_1017_add_4_7_lut .LUT_INIT = 16'hC33C;
    SB_LUT4 add_3197_6_lut (.I0(GND_net), .I1(n11992[3]), .I2(n504), .I3(n34492), 
            .O(n11358[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3197_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3197_6 (.CI(n34492), .I0(n11992[3]), .I1(n504), .CO(n34493));
    SB_LUT4 add_3057_28_lut (.I0(GND_net), .I1(n8019[25]), .I2(GND_net), 
            .I3(n35268), .O(n7988[26])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3057_28_lut.LUT_INIT = 16'hC33C;
    SB_CARRY \PID_CONTROLLER.integral_1017_add_4_7  (.CI(n35072), .I0(\PID_CONTROLLER.err[5] ), 
            .I1(\PID_CONTROLLER.integral [5]), .CO(n35073));
    SB_LUT4 add_3197_5_lut (.I0(GND_net), .I1(n11992[2]), .I2(n407), .I3(n34491), 
            .O(n11358[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3197_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3197_5 (.CI(n34491), .I0(n11992[2]), .I1(n407), .CO(n34492));
    SB_LUT4 sub_11_inv_0_i5_1_lut (.I0(\PID_CONTROLLER.err[4] ), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n64[4]));   // verilog/motorControl.v(43[31:45])
    defparam sub_11_inv_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 \PID_CONTROLLER.integral_1017_add_4_6_lut  (.I0(GND_net), .I1(\PID_CONTROLLER.err[4] ), 
            .I2(\PID_CONTROLLER.integral [4]), .I3(n35071), .O(n66[4])) /* synthesis syn_instantiated=1 */ ;
    defparam \PID_CONTROLLER.integral_1017_add_4_6_lut .LUT_INIT = 16'hC33C;
    SB_LUT4 add_3197_4_lut (.I0(GND_net), .I1(n11992[1]), .I2(n310_adj_3390), 
            .I3(n34490), .O(n11358[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3197_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3197_4 (.CI(n34490), .I0(n11992[1]), .I1(n310_adj_3390), 
            .CO(n34491));
    SB_CARRY add_3065_4 (.CI(n35440), .I0(n8231[1]), .I1(n322_adj_3401), 
            .CO(n35441));
    SB_LUT4 add_3062_10_lut (.I0(GND_net), .I1(n8159[7]), .I2(GND_net), 
            .I3(n35380), .O(n8133[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3062_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3057_28 (.CI(n35268), .I0(n8019[25]), .I1(GND_net), .CO(n35269));
    SB_CARRY \PID_CONTROLLER.integral_1017_add_4_6  (.CI(n35071), .I0(\PID_CONTROLLER.err[4] ), 
            .I1(\PID_CONTROLLER.integral [4]), .CO(n35072));
    SB_LUT4 add_3197_3_lut (.I0(GND_net), .I1(n11992[0]), .I2(n213), .I3(n34489), 
            .O(n11358[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3197_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3197_3 (.CI(n34489), .I0(n11992[0]), .I1(n213), .CO(n34490));
    SB_LUT4 \PID_CONTROLLER.integral_1017_add_4_5_lut  (.I0(GND_net), .I1(\PID_CONTROLLER.err[3] ), 
            .I2(\PID_CONTROLLER.integral [3]), .I3(n35070), .O(n66[3])) /* synthesis syn_instantiated=1 */ ;
    defparam \PID_CONTROLLER.integral_1017_add_4_5_lut .LUT_INIT = 16'hC33C;
    SB_LUT4 add_3197_2_lut (.I0(GND_net), .I1(n23_adj_3389), .I2(n116), 
            .I3(GND_net), .O(n11358[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3197_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3197_2 (.CI(GND_net), .I0(n23_adj_3389), .I1(n116), .CO(n34489));
    SB_LUT4 add_3057_27_lut (.I0(GND_net), .I1(n8019[24]), .I2(GND_net), 
            .I3(n35267), .O(n7988[25])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3057_27_lut.LUT_INIT = 16'hC33C;
    SB_CARRY \PID_CONTROLLER.integral_1017_add_4_5  (.CI(n35070), .I0(\PID_CONTROLLER.err[3] ), 
            .I1(\PID_CONTROLLER.integral [3]), .CO(n35071));
    SB_LUT4 add_3361_11_lut (.I0(GND_net), .I1(n15226[8]), .I2(GND_net), 
            .I3(n34488), .O(n14912[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3361_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3361_10_lut (.I0(GND_net), .I1(n15226[7]), .I2(GND_net), 
            .I3(n34487), .O(n14912[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3361_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 \PID_CONTROLLER.integral_1017_add_4_4_lut  (.I0(GND_net), .I1(\PID_CONTROLLER.err[2] ), 
            .I2(\PID_CONTROLLER.integral [2]), .I3(n35069), .O(n66[2])) /* synthesis syn_instantiated=1 */ ;
    defparam \PID_CONTROLLER.integral_1017_add_4_4_lut .LUT_INIT = 16'hC33C;
    SB_CARRY add_3361_10 (.CI(n34487), .I0(n15226[7]), .I1(GND_net), .CO(n34488));
    SB_LUT4 add_3361_9_lut (.I0(GND_net), .I1(n15226[6]), .I2(GND_net), 
            .I3(n34486), .O(n14912[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3361_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3062_10 (.CI(n35380), .I0(n8159[7]), .I1(GND_net), .CO(n35381));
    SB_CARRY add_3057_27 (.CI(n35267), .I0(n8019[24]), .I1(GND_net), .CO(n35268));
    SB_CARRY \PID_CONTROLLER.integral_1017_add_4_4  (.CI(n35069), .I0(\PID_CONTROLLER.err[2] ), 
            .I1(\PID_CONTROLLER.integral [2]), .CO(n35070));
    SB_CARRY add_3361_9 (.CI(n34486), .I0(n15226[6]), .I1(GND_net), .CO(n34487));
    SB_LUT4 add_3361_8_lut (.I0(GND_net), .I1(n15226[5]), .I2(n545), .I3(n34485), 
            .O(n14912[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3361_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 \PID_CONTROLLER.integral_1017_add_4_3_lut  (.I0(GND_net), .I1(\PID_CONTROLLER.err[1] ), 
            .I2(\PID_CONTROLLER.integral [1]), .I3(n35068), .O(n66[1])) /* synthesis syn_instantiated=1 */ ;
    defparam \PID_CONTROLLER.integral_1017_add_4_3_lut .LUT_INIT = 16'hC33C;
    SB_CARRY add_3361_8 (.CI(n34485), .I0(n15226[5]), .I1(n545), .CO(n34486));
    SB_LUT4 add_3361_7_lut (.I0(GND_net), .I1(n15226[4]), .I2(n472), .I3(n34484), 
            .O(n14912[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3361_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3057_26_lut (.I0(GND_net), .I1(n8019[23]), .I2(GND_net), 
            .I3(n35266), .O(n7988[24])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3057_26_lut.LUT_INIT = 16'hC33C;
    SB_CARRY \PID_CONTROLLER.integral_1017_add_4_3  (.CI(n35068), .I0(\PID_CONTROLLER.err[1] ), 
            .I1(\PID_CONTROLLER.integral [1]), .CO(n35069));
    SB_CARRY add_3361_7 (.CI(n34484), .I0(n15226[4]), .I1(n472), .CO(n34485));
    SB_LUT4 mult_12_i396_2_lut (.I0(\Kd[6] ), .I1(n57[2]), .I2(GND_net), 
            .I3(GND_net), .O(n589));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i396_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_3361_6_lut (.I0(GND_net), .I1(n15226[3]), .I2(n399), .I3(n34483), 
            .O(n14912[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3361_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 \PID_CONTROLLER.integral_1017_add_4_2_lut  (.I0(GND_net), .I1(\PID_CONTROLLER.err[0] ), 
            .I2(\PID_CONTROLLER.integral [0]), .I3(GND_net), .O(n66[0])) /* synthesis syn_instantiated=1 */ ;
    defparam \PID_CONTROLLER.integral_1017_add_4_2_lut .LUT_INIT = 16'hC33C;
    SB_CARRY add_3361_6 (.CI(n34483), .I0(n15226[3]), .I1(n399), .CO(n34484));
    SB_LUT4 add_3361_5_lut (.I0(GND_net), .I1(n15226[2]), .I2(n326), .I3(n34482), 
            .O(n14912[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3361_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3067_8_lut (.I0(GND_net), .I1(n8274[5]), .I2(n716), .I3(n35483), 
            .O(n8253[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3067_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3065_3_lut (.I0(GND_net), .I1(n8231[0]), .I2(n225_adj_3382), 
            .I3(n35439), .O(n8208[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3065_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3062_9_lut (.I0(GND_net), .I1(n8159[6]), .I2(GND_net), 
            .I3(n35379), .O(n8133[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3062_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3057_26 (.CI(n35266), .I0(n8019[23]), .I1(GND_net), .CO(n35267));
    SB_CARRY \PID_CONTROLLER.integral_1017_add_4_2  (.CI(GND_net), .I0(\PID_CONTROLLER.err[0] ), 
            .I1(\PID_CONTROLLER.integral [0]), .CO(n35068));
    SB_CARRY add_3361_5 (.CI(n34482), .I0(n15226[2]), .I1(n326), .CO(n34483));
    SB_LUT4 add_3361_4_lut (.I0(GND_net), .I1(n15226[1]), .I2(n253), .I3(n34481), 
            .O(n14912[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3361_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 pwm_count_1016_add_4_10_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_count[8]), 
            .I3(n35067), .O(n67[8])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_count_1016_add_4_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3361_4 (.CI(n34481), .I0(n15226[1]), .I1(n253), .CO(n34482));
    SB_LUT4 add_3361_3_lut (.I0(GND_net), .I1(n15226[0]), .I2(n180), .I3(n34480), 
            .O(n14912[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3361_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3057_25_lut (.I0(GND_net), .I1(n8019[22]), .I2(GND_net), 
            .I3(n35265), .O(n7988[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3057_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 pwm_count_1016_add_4_9_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_count[7]), 
            .I3(n35066), .O(n67[7])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_count_1016_add_4_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3361_3 (.CI(n34480), .I0(n15226[0]), .I1(n180), .CO(n34481));
    SB_LUT4 add_3361_2_lut (.I0(GND_net), .I1(n35), .I2(n107), .I3(GND_net), 
            .O(n14912[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3361_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_count_1016_add_4_9 (.CI(n35066), .I0(GND_net), .I1(pwm_count[7]), 
            .CO(n35067));
    SB_CARRY add_3361_2 (.CI(GND_net), .I0(n35), .I1(n107), .CO(n34480));
    SB_CARRY add_3062_9 (.CI(n35379), .I0(n8159[6]), .I1(GND_net), .CO(n35380));
    SB_CARRY add_3057_25 (.CI(n35265), .I0(n8019[22]), .I1(GND_net), .CO(n35266));
    SB_LUT4 pwm_count_1016_add_4_8_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_count[6]), 
            .I3(n35065), .O(n67[6])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_count_1016_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_count_1016_add_4_8 (.CI(n35065), .I0(GND_net), .I1(pwm_count[6]), 
            .CO(n35066));
    SB_LUT4 mult_12_i91_2_lut (.I0(\Kd[1] ), .I1(n57[12]), .I2(GND_net), 
            .I3(GND_net), .O(n134));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i91_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_3057_24_lut (.I0(GND_net), .I1(n8019[21]), .I2(GND_net), 
            .I3(n35264), .O(n7988[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3057_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 pwm_count_1016_add_4_7_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_count[5]), 
            .I3(n35064), .O(n67[5])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_count_1016_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_count_1016_add_4_7 (.CI(n35064), .I0(GND_net), .I1(pwm_count[5]), 
            .CO(n35065));
    SB_CARRY add_3065_3 (.CI(n35439), .I0(n8231[0]), .I1(n225_adj_3382), 
            .CO(n35440));
    SB_LUT4 add_3062_8_lut (.I0(GND_net), .I1(n8159[5]), .I2(n701), .I3(n35378), 
            .O(n8133[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3062_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3057_24 (.CI(n35264), .I0(n8019[21]), .I1(GND_net), .CO(n35265));
    SB_LUT4 pwm_count_1016_add_4_6_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_count[4]), 
            .I3(n35063), .O(n67[4])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_count_1016_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_count_1016_add_4_6 (.CI(n35063), .I0(GND_net), .I1(pwm_count[4]), 
            .CO(n35064));
    SB_LUT4 add_3057_23_lut (.I0(GND_net), .I1(n8019[20]), .I2(GND_net), 
            .I3(n35263), .O(n7988[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3057_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 pwm_count_1016_add_4_5_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_count[3]), 
            .I3(n35062), .O(n67[3])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_count_1016_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3223_25_lut (.I0(GND_net), .I1(n12575[22]), .I2(GND_net), 
            .I3(n34473), .O(n11992[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3223_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3223_24_lut (.I0(GND_net), .I1(n12575[21]), .I2(GND_net), 
            .I3(n34472), .O(n11992[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3223_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_count_1016_add_4_5 (.CI(n35062), .I0(GND_net), .I1(pwm_count[3]), 
            .CO(n35063));
    SB_CARRY add_3223_24 (.CI(n34472), .I0(n12575[21]), .I1(GND_net), 
            .CO(n34473));
    SB_LUT4 add_3223_23_lut (.I0(GND_net), .I1(n12575[20]), .I2(GND_net), 
            .I3(n34471), .O(n11992[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3223_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3062_8 (.CI(n35378), .I0(n8159[5]), .I1(n701), .CO(n35379));
    SB_CARRY add_3057_23 (.CI(n35263), .I0(n8019[20]), .I1(GND_net), .CO(n35264));
    SB_LUT4 pwm_count_1016_add_4_4_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_count[2]), 
            .I3(n35061), .O(n67[2])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_count_1016_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3223_23 (.CI(n34471), .I0(n12575[20]), .I1(GND_net), 
            .CO(n34472));
    SB_LUT4 add_3223_22_lut (.I0(GND_net), .I1(n12575[19]), .I2(GND_net), 
            .I3(n34470), .O(n11992[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3223_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_count_1016_add_4_4 (.CI(n35061), .I0(GND_net), .I1(pwm_count[2]), 
            .CO(n35062));
    SB_LUT4 mult_12_i28_2_lut (.I0(\Kd[0] ), .I1(n57[13]), .I2(GND_net), 
            .I3(GND_net), .O(n41));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i28_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_3223_22 (.CI(n34470), .I0(n12575[19]), .I1(GND_net), 
            .CO(n34471));
    SB_LUT4 add_3223_21_lut (.I0(GND_net), .I1(n12575[18]), .I2(GND_net), 
            .I3(n34469), .O(n11992[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3223_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3057_22_lut (.I0(GND_net), .I1(n8019[19]), .I2(GND_net), 
            .I3(n35262), .O(n7988[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3057_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 pwm_count_1016_add_4_3_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_count[1]), 
            .I3(n35060), .O(n67[1])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_count_1016_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_11_add_2_18 (.CI(n34206), .I0(\PID_CONTROLLER.err_prev[16] ), 
            .I1(n64[16]), .CO(n34207));
    SB_CARRY add_3223_21 (.CI(n34469), .I0(n12575[18]), .I1(GND_net), 
            .CO(n34470));
    SB_LUT4 add_3223_20_lut (.I0(GND_net), .I1(n12575[17]), .I2(GND_net), 
            .I3(n34468), .O(n11992[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3223_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_count_1016_add_4_3 (.CI(n35060), .I0(GND_net), .I1(pwm_count[1]), 
            .CO(n35061));
    SB_CARRY add_3223_20 (.CI(n34468), .I0(n12575[17]), .I1(GND_net), 
            .CO(n34469));
    SB_LUT4 mult_12_i268_2_lut (.I0(\Kd[4] ), .I1(n57[3]), .I2(GND_net), 
            .I3(GND_net), .O(n398));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i268_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_3223_19_lut (.I0(GND_net), .I1(n12575[16]), .I2(GND_net), 
            .I3(n34467), .O(n11992[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3223_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3069_16 (.CI(n35526), .I0(n8313[13]), .I1(GND_net), .CO(n35527));
    SB_CARRY add_3067_8 (.CI(n35483), .I0(n8274[5]), .I1(n716), .CO(n35484));
    SB_LUT4 add_3065_2_lut (.I0(GND_net), .I1(n35_adj_3381), .I2(n128), 
            .I3(GND_net), .O(n8208[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3065_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3062_7_lut (.I0(GND_net), .I1(n8159[4]), .I2(n604), .I3(n35377), 
            .O(n8133[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3062_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3057_22 (.CI(n35262), .I0(n8019[19]), .I1(GND_net), .CO(n35263));
    SB_LUT4 pwm_count_1016_add_4_2_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_count[0]), 
            .I3(VCC_net), .O(n67[0])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_count_1016_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3223_19 (.CI(n34467), .I0(n12575[16]), .I1(GND_net), 
            .CO(n34468));
    SB_LUT4 add_3223_18_lut (.I0(GND_net), .I1(n12575[15]), .I2(GND_net), 
            .I3(n34466), .O(n11992[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3223_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_count_1016_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(pwm_count[0]), 
            .CO(n35060));
    SB_CARRY add_3223_18 (.CI(n34466), .I0(n12575[15]), .I1(GND_net), 
            .CO(n34467));
    SB_LUT4 add_3223_17_lut (.I0(GND_net), .I1(n12575[14]), .I2(GND_net), 
            .I3(n34465), .O(n11992[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3223_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3057_21_lut (.I0(GND_net), .I1(n8019[18]), .I2(GND_net), 
            .I3(n35261), .O(n7988[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3057_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3056_31_lut (.I0(GND_net), .I1(n7988[28]), .I2(GND_net), 
            .I3(n35059), .O(n7956[29])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3056_31_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3223_17 (.CI(n34465), .I0(n12575[14]), .I1(GND_net), 
            .CO(n34466));
    SB_LUT4 mult_12_i282_2_lut (.I0(\Kd[4] ), .I1(n57[10]), .I2(GND_net), 
            .I3(GND_net), .O(n419_adj_3402));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i282_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_3223_16_lut (.I0(GND_net), .I1(n12575[13]), .I2(GND_net), 
            .I3(n34464), .O(n11992[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3223_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3056_30_lut (.I0(GND_net), .I1(n7988[27]), .I2(GND_net), 
            .I3(n35058), .O(n7956[28])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3056_30_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3223_16 (.CI(n34464), .I0(n12575[13]), .I1(GND_net), 
            .CO(n34465));
    SB_LUT4 add_3223_15_lut (.I0(GND_net), .I1(n12575[12]), .I2(GND_net), 
            .I3(n34463), .O(n11992[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3223_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3062_7 (.CI(n35377), .I0(n8159[4]), .I1(n604), .CO(n35378));
    SB_CARRY add_3057_21 (.CI(n35261), .I0(n8019[18]), .I1(GND_net), .CO(n35262));
    SB_CARRY add_3056_30 (.CI(n35058), .I0(n7988[27]), .I1(GND_net), .CO(n35059));
    SB_CARRY add_3223_15 (.CI(n34463), .I0(n12575[12]), .I1(GND_net), 
            .CO(n34464));
    SB_LUT4 add_3223_14_lut (.I0(GND_net), .I1(n12575[11]), .I2(GND_net), 
            .I3(n34462), .O(n11992[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3223_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3056_29_lut (.I0(GND_net), .I1(n7988[26]), .I2(GND_net), 
            .I3(n35057), .O(n7956[27])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3056_29_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3223_14 (.CI(n34462), .I0(n12575[11]), .I1(GND_net), 
            .CO(n34463));
    SB_LUT4 add_3223_13_lut (.I0(GND_net), .I1(n12575[10]), .I2(GND_net), 
            .I3(n34461), .O(n11992[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3223_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3057_20_lut (.I0(GND_net), .I1(n8019[17]), .I2(GND_net), 
            .I3(n35260), .O(n7988[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3057_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3056_29 (.CI(n35057), .I0(n7988[26]), .I1(GND_net), .CO(n35058));
    SB_CARRY add_3223_13 (.CI(n34461), .I0(n12575[10]), .I1(GND_net), 
            .CO(n34462));
    SB_LUT4 add_3223_12_lut (.I0(GND_net), .I1(n12575[9]), .I2(GND_net), 
            .I3(n34460), .O(n11992[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3223_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_12_i461_2_lut (.I0(\Kd[7] ), .I1(n57[2]), .I2(GND_net), 
            .I3(GND_net), .O(n686));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i461_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_3056_28_lut (.I0(GND_net), .I1(n7988[25]), .I2(GND_net), 
            .I3(n35056), .O(n7956[26])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3056_28_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3223_12 (.CI(n34460), .I0(n12575[9]), .I1(GND_net), .CO(n34461));
    SB_LUT4 add_3223_11_lut (.I0(GND_net), .I1(n12575[8]), .I2(GND_net), 
            .I3(n34459), .O(n11992[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3223_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_add_2137_32_lut (.I0(\PID_CONTROLLER.err[31] ), .I1(n6542[29]), 
            .I2(GND_net), .I3(n34730), .O(n5786[0])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_2137_32_lut.LUT_INIT = 16'h6996;
    SB_CARRY add_3065_2 (.CI(GND_net), .I0(n35_adj_3381), .I1(n128), .CO(n35439));
    SB_LUT4 add_3062_6_lut (.I0(GND_net), .I1(n8159[3]), .I2(n507), .I3(n35376), 
            .O(n8133[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3062_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3057_20 (.CI(n35260), .I0(n8019[17]), .I1(GND_net), .CO(n35261));
    SB_CARRY add_3056_28 (.CI(n35056), .I0(n7988[25]), .I1(GND_net), .CO(n35057));
    SB_LUT4 mult_10_add_2137_31_lut (.I0(GND_net), .I1(n6542[28]), .I2(GND_net), 
            .I3(n34729), .O(n61[30])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_2137_31_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3223_11 (.CI(n34459), .I0(n12575[8]), .I1(GND_net), .CO(n34460));
    SB_LUT4 add_3223_10_lut (.I0(GND_net), .I1(n12575[7]), .I2(GND_net), 
            .I3(n34458), .O(n11992[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3223_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_2137_31 (.CI(n34729), .I0(n6542[28]), .I1(GND_net), 
            .CO(n34730));
    SB_LUT4 add_3056_27_lut (.I0(GND_net), .I1(n7988[24]), .I2(GND_net), 
            .I3(n35055), .O(n7956[25])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3056_27_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_add_2137_30_lut (.I0(GND_net), .I1(n6542[27]), .I2(GND_net), 
            .I3(n34728), .O(n61[29])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_2137_30_lut.LUT_INIT = 16'hC33C;
    SB_DFF pwm__i23 (.Q(pwm[23]), .C(clk32MHz), .D(n24227));   // verilog/motorControl.v(38[14] 59[8])
    SB_DFF pwm__i22 (.Q(pwm[22]), .C(clk32MHz), .D(n24226));   // verilog/motorControl.v(38[14] 59[8])
    SB_DFF pwm__i21 (.Q(pwm[21]), .C(clk32MHz), .D(n24225));   // verilog/motorControl.v(38[14] 59[8])
    SB_DFF pwm__i20 (.Q(pwm[20]), .C(clk32MHz), .D(n24224));   // verilog/motorControl.v(38[14] 59[8])
    SB_DFF pwm__i19 (.Q(pwm[19]), .C(clk32MHz), .D(n24223));   // verilog/motorControl.v(38[14] 59[8])
    SB_DFF pwm__i18 (.Q(pwm[18]), .C(clk32MHz), .D(n39108));   // verilog/motorControl.v(38[14] 59[8])
    SB_DFF pwm__i17 (.Q(pwm[17]), .C(clk32MHz), .D(n39110));   // verilog/motorControl.v(38[14] 59[8])
    SB_DFF pwm__i16 (.Q(pwm[16]), .C(clk32MHz), .D(n24220));   // verilog/motorControl.v(38[14] 59[8])
    SB_DFF pwm__i15 (.Q(pwm[15]), .C(clk32MHz), .D(n24219));   // verilog/motorControl.v(38[14] 59[8])
    SB_DFF pwm__i14 (.Q(pwm[14]), .C(clk32MHz), .D(n24218));   // verilog/motorControl.v(38[14] 59[8])
    SB_DFF pwm__i13 (.Q(pwm[13]), .C(clk32MHz), .D(n24217));   // verilog/motorControl.v(38[14] 59[8])
    SB_DFF pwm__i12 (.Q(pwm[12]), .C(clk32MHz), .D(n24216));   // verilog/motorControl.v(38[14] 59[8])
    SB_DFF pwm__i11 (.Q(pwm[11]), .C(clk32MHz), .D(n24215));   // verilog/motorControl.v(38[14] 59[8])
    SB_DFF pwm__i10 (.Q(pwm[10]), .C(clk32MHz), .D(n24214));   // verilog/motorControl.v(38[14] 59[8])
    SB_DFF pwm__i9 (.Q(pwm[9]), .C(clk32MHz), .D(n24213));   // verilog/motorControl.v(38[14] 59[8])
    SB_DFF pwm__i8 (.Q(pwm[8]), .C(clk32MHz), .D(n24212));   // verilog/motorControl.v(38[14] 59[8])
    SB_DFF pwm__i7 (.Q(pwm[7]), .C(clk32MHz), .D(n24211));   // verilog/motorControl.v(38[14] 59[8])
    SB_DFF pwm__i6 (.Q(pwm[6]), .C(clk32MHz), .D(n24210));   // verilog/motorControl.v(38[14] 59[8])
    SB_DFF pwm__i5 (.Q(pwm[5]), .C(clk32MHz), .D(n24209));   // verilog/motorControl.v(38[14] 59[8])
    SB_DFF pwm__i4 (.Q(pwm[4]), .C(clk32MHz), .D(n24208));   // verilog/motorControl.v(38[14] 59[8])
    SB_DFF pwm__i3 (.Q(pwm[3]), .C(clk32MHz), .D(n24207));   // verilog/motorControl.v(38[14] 59[8])
    SB_DFF pwm__i2 (.Q(pwm[2]), .C(clk32MHz), .D(n24206));   // verilog/motorControl.v(38[14] 59[8])
    SB_DFF pwm__i1 (.Q(pwm[1]), .C(clk32MHz), .D(n24205));   // verilog/motorControl.v(38[14] 59[8])
    SB_DFF pwm__i0 (.Q(pwm[0]), .C(clk32MHz), .D(n24172));   // verilog/motorControl.v(38[14] 59[8])
    SB_LUT4 mult_12_i333_2_lut (.I0(\Kd[5] ), .I1(n57[3]), .I2(GND_net), 
            .I3(GND_net), .O(n495));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i333_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_3223_10 (.CI(n34458), .I0(n12575[7]), .I1(GND_net), .CO(n34459));
    SB_CARRY mult_10_add_2137_30 (.CI(n34728), .I0(n6542[27]), .I1(GND_net), 
            .CO(n34729));
    SB_LUT4 mult_12_i398_2_lut (.I0(\Kd[6] ), .I1(n57[3]), .I2(GND_net), 
            .I3(GND_net), .O(n592));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i398_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_3223_9_lut (.I0(GND_net), .I1(n12575[6]), .I2(GND_net), 
            .I3(n34457), .O(n11992[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3223_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i77_2_lut (.I0(\Kp[1] ), .I1(\PID_CONTROLLER.err[5] ), 
            .I2(GND_net), .I3(GND_net), .O(n113));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i77_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_add_2137_29_lut (.I0(GND_net), .I1(n6542[26]), .I2(GND_net), 
            .I3(n34727), .O(n61[28])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_2137_29_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3057_19_lut (.I0(GND_net), .I1(n8019[16]), .I2(GND_net), 
            .I3(n35259), .O(n7988[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3057_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i14_2_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err[6] ), 
            .I2(GND_net), .I3(GND_net), .O(n20_adj_3400));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i14_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i156_2_lut (.I0(\Kd[2] ), .I1(n57[12]), .I2(GND_net), 
            .I3(GND_net), .O(n231));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i156_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_3056_27 (.CI(n35055), .I0(n7988[24]), .I1(GND_net), .CO(n35056));
    SB_LUT4 mult_10_i142_2_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err[5] ), 
            .I2(GND_net), .I3(GND_net), .O(n210));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i142_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY mult_10_add_2137_29 (.CI(n34727), .I0(n6542[26]), .I1(GND_net), 
            .CO(n34728));
    SB_LUT4 mult_10_i207_2_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err[5] ), 
            .I2(GND_net), .I3(GND_net), .O(n307_adj_3399));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i207_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i463_2_lut (.I0(\Kd[7] ), .I1(n57[3]), .I2(GND_net), 
            .I3(GND_net), .O(n689));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i463_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i221_2_lut (.I0(\Kd[3] ), .I1(n57[12]), .I2(GND_net), 
            .I3(GND_net), .O(n328));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i221_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i272_2_lut (.I0(\Kp[4] ), .I1(\PID_CONTROLLER.err[5] ), 
            .I2(GND_net), .I3(GND_net), .O(n404));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i272_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i337_2_lut (.I0(\Kp[5] ), .I1(\PID_CONTROLLER.err[5] ), 
            .I2(GND_net), .I3(GND_net), .O(n501));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i337_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i402_2_lut (.I0(\Kp[6] ), .I1(\PID_CONTROLLER.err[5] ), 
            .I2(GND_net), .I3(GND_net), .O(n598));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i402_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 sub_11_inv_0_i17_1_lut (.I0(\PID_CONTROLLER.err[16] ), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n64[16]));   // verilog/motorControl.v(43[31:45])
    defparam sub_11_inv_0_i17_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_add_2137_28_lut (.I0(GND_net), .I1(n6542[25]), .I2(GND_net), 
            .I3(n34726), .O(n61[27])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_2137_28_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i467_2_lut (.I0(\Kp[7] ), .I1(\PID_CONTROLLER.err[5] ), 
            .I2(GND_net), .I3(GND_net), .O(n695));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i467_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_3223_9 (.CI(n34457), .I0(n12575[6]), .I1(GND_net), .CO(n34458));
    SB_LUT4 mult_12_i347_2_lut (.I0(\Kd[5] ), .I1(n57[10]), .I2(GND_net), 
            .I3(GND_net), .O(n516_adj_3397));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i347_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 sub_11_add_2_17_lut (.I0(GND_net), .I1(\PID_CONTROLLER.err_prev[15] ), 
            .I2(n64[15]), .I3(n34205), .O(n57[15])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_11_add_2_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3223_8_lut (.I0(GND_net), .I1(n12575[5]), .I2(n701_adj_3413), 
            .I3(n34456), .O(n11992[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3223_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3464_5_lut (.I0(GND_net), .I1(n16505[2]), .I2(n452), .I3(n34363), 
            .O(n16420[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3464_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_12_i286_2_lut (.I0(\Kd[4] ), .I1(n57[12]), .I2(GND_net), 
            .I3(GND_net), .O(n425));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i286_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i412_2_lut (.I0(\Kd[6] ), .I1(n57[10]), .I2(GND_net), 
            .I3(GND_net), .O(n613_adj_3396));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i412_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY sub_11_add_2_17 (.CI(n34205), .I0(\PID_CONTROLLER.err_prev[15] ), 
            .I1(n64[15]), .CO(n34206));
    SB_CARRY add_3464_5 (.CI(n34363), .I0(n16505[2]), .I1(n452), .CO(n34364));
    SB_LUT4 add_3074_3_lut (.I0(GND_net), .I1(n8393[0]), .I2(n252), .I3(n35583), 
            .O(n8379[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3074_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_12_i235_2_lut (.I0(\Kd[3] ), .I1(n57[19]), .I2(GND_net), 
            .I3(GND_net), .O(n349));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i235_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 sub_11_inv_0_i18_1_lut (.I0(\PID_CONTROLLER.err[17] ), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n64[17]));   // verilog/motorControl.v(43[31:45])
    defparam sub_11_inv_0_i18_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i369_2_lut (.I0(\Kp[5] ), .I1(\PID_CONTROLLER.err[21] ), 
            .I2(GND_net), .I3(GND_net), .O(n549));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i369_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i67_2_lut (.I0(\Kp[1] ), .I1(\PID_CONTROLLER.err[0] ), 
            .I2(GND_net), .I3(GND_net), .O(n98));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i67_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i4_2_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err[1] ), 
            .I2(GND_net), .I3(GND_net), .O(n5));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i4_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_14_i291_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral [9]), 
            .I2(GND_net), .I3(GND_net), .O(n399));   // verilog/motorControl.v(43[48:59])
    defparam mult_14_i291_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_14_i340_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral [9]), 
            .I2(GND_net), .I3(GND_net), .O(n472));   // verilog/motorControl.v(43[48:59])
    defparam mult_14_i340_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_3431_12_lut (.I0(GND_net), .I1(n16185[9]), .I2(GND_net), 
            .I3(n35675), .O(n16031[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3431_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3074_3 (.CI(n35583), .I0(n8393[0]), .I1(n252), .CO(n35584));
    SB_LUT4 add_3074_2_lut (.I0(GND_net), .I1(n62), .I2(n155_adj_3414), 
            .I3(GND_net), .O(n8379[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3074_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_i389_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral [9]), 
            .I2(GND_net), .I3(GND_net), .O(n545));   // verilog/motorControl.v(43[48:59])
    defparam mult_14_i389_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 sub_11_inv_0_i6_1_lut (.I0(\PID_CONTROLLER.err[5] ), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n64[5]));   // verilog/motorControl.v(43[31:45])
    defparam sub_11_inv_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_3069_15_lut (.I0(GND_net), .I1(n8313[12]), .I2(GND_net), 
            .I3(n35525), .O(n8294[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3069_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3069_15 (.CI(n35525), .I0(n8313[12]), .I1(GND_net), .CO(n35526));
    SB_CARRY mult_10_add_2137_28 (.CI(n34726), .I0(n6542[25]), .I1(GND_net), 
            .CO(n34727));
    SB_LUT4 add_3069_14_lut (.I0(GND_net), .I1(n8313[11]), .I2(GND_net), 
            .I3(n35524), .O(n8294[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3069_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3431_12 (.CI(n35675), .I0(n16185[9]), .I1(GND_net), .CO(n35676));
    SB_LUT4 add_3431_11_lut (.I0(GND_net), .I1(n16185[8]), .I2(GND_net), 
            .I3(n35674), .O(n16031[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3431_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3056_26_lut (.I0(GND_net), .I1(n7988[23]), .I2(GND_net), 
            .I3(n35054), .O(n7956[24])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3056_26_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i75_2_lut (.I0(\Kp[1] ), .I1(\PID_CONTROLLER.err[4] ), 
            .I2(GND_net), .I3(GND_net), .O(n110_adj_3394));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i75_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i12_2_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err[5] ), 
            .I2(GND_net), .I3(GND_net), .O(n17_adj_3393));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i12_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i477_2_lut (.I0(\Kd[7] ), .I1(n57[10]), .I2(GND_net), 
            .I3(GND_net), .O(n710_adj_3392));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i477_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_add_2137_27_lut (.I0(GND_net), .I1(n6542[24]), .I2(GND_net), 
            .I3(n34725), .O(n61[26])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_2137_27_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_12_i300_2_lut (.I0(\Kd[4] ), .I1(n57[19]), .I2(GND_net), 
            .I3(GND_net), .O(n446));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i300_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_3064_23_lut (.I0(GND_net), .I1(n8208[20]), .I2(GND_net), 
            .I3(n35438), .O(n8184[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3064_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_11_add_2_16_lut (.I0(GND_net), .I1(\PID_CONTROLLER.err_prev[14] ), 
            .I2(n64[14]), .I3(n34204), .O(n57[14])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_11_add_2_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3062_6 (.CI(n35376), .I0(n8159[3]), .I1(n507), .CO(n35377));
    SB_CARRY add_3057_19 (.CI(n35259), .I0(n8019[16]), .I1(GND_net), .CO(n35260));
    SB_LUT4 add_3057_18_lut (.I0(GND_net), .I1(n8019[15]), .I2(GND_net), 
            .I3(n35258), .O(n7988[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3057_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3223_8 (.CI(n34456), .I0(n12575[5]), .I1(n701_adj_3413), 
            .CO(n34457));
    SB_CARRY add_3057_18 (.CI(n35258), .I0(n8019[15]), .I1(GND_net), .CO(n35259));
    SB_CARRY sub_11_add_2_16 (.CI(n34204), .I0(\PID_CONTROLLER.err_prev[14] ), 
            .I1(n64[14]), .CO(n34205));
    SB_LUT4 sub_11_add_2_15_lut (.I0(GND_net), .I1(\PID_CONTROLLER.err_prev[13] ), 
            .I2(n64[13]), .I3(n34203), .O(n57[13])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_11_add_2_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3056_26 (.CI(n35054), .I0(n7988[23]), .I1(GND_net), .CO(n35055));
    SB_LUT4 add_3056_25_lut (.I0(GND_net), .I1(n7988[22]), .I2(GND_net), 
            .I3(n35053), .O(n7956[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3056_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_2137_27 (.CI(n34725), .I0(n6542[24]), .I1(GND_net), 
            .CO(n34726));
    SB_LUT4 mult_10_add_2137_26_lut (.I0(GND_net), .I1(n6542[23]), .I2(GND_net), 
            .I3(n34724), .O(n61[25])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_2137_26_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_11_inv_0_i19_1_lut (.I0(\PID_CONTROLLER.err[18] ), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n64[18]));   // verilog/motorControl.v(43[31:45])
    defparam sub_11_inv_0_i19_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_3464_4_lut (.I0(GND_net), .I1(n16505[1]), .I2(n355), .I3(n34362), 
            .O(n16420[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3464_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3464_4 (.CI(n34362), .I0(n16505[1]), .I1(n355), .CO(n34363));
    SB_LUT4 add_3464_3_lut (.I0(GND_net), .I1(n16505[0]), .I2(n258), .I3(n34361), 
            .O(n16420[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3464_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_11_add_2_15 (.CI(n34203), .I0(\PID_CONTROLLER.err_prev[13] ), 
            .I1(n64[13]), .CO(n34204));
    SB_LUT4 add_3223_7_lut (.I0(GND_net), .I1(n12575[4]), .I2(n604_adj_3417), 
            .I3(n34455), .O(n11992[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3223_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3056_25 (.CI(n35053), .I0(n7988[22]), .I1(GND_net), .CO(n35054));
    SB_LUT4 add_3056_24_lut (.I0(GND_net), .I1(n7988[21]), .I2(GND_net), 
            .I3(n35052), .O(n7956[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3056_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_11_add_2_14_lut (.I0(GND_net), .I1(\PID_CONTROLLER.err_prev[12] ), 
            .I2(n64[12]), .I3(n34202), .O(n57[12])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_11_add_2_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_11_inv_0_i20_1_lut (.I0(\PID_CONTROLLER.err[19] ), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n64[19]));   // verilog/motorControl.v(43[31:45])
    defparam sub_11_inv_0_i20_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY mult_10_add_2137_26 (.CI(n34724), .I0(n6542[23]), .I1(GND_net), 
            .CO(n34725));
    SB_CARRY add_3464_3 (.CI(n34361), .I0(n16505[0]), .I1(n258), .CO(n34362));
    SB_LUT4 mult_10_i434_2_lut (.I0(\Kp[6] ), .I1(\PID_CONTROLLER.err[21] ), 
            .I2(GND_net), .I3(GND_net), .O(n646));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i434_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_add_2137_25_lut (.I0(GND_net), .I1(n6542[22]), .I2(GND_net), 
            .I3(n34723), .O(n61[24])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_2137_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_11_add_2_14 (.CI(n34202), .I0(\PID_CONTROLLER.err_prev[12] ), 
            .I1(n64[12]), .CO(n34203));
    SB_CARRY mult_10_add_2137_25 (.CI(n34723), .I0(n6542[22]), .I1(GND_net), 
            .CO(n34724));
    SB_LUT4 mult_10_add_2137_24_lut (.I0(GND_net), .I1(n6542[21]), .I2(GND_net), 
            .I3(n34722), .O(n61[23])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_2137_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_11_add_2_13_lut (.I0(GND_net), .I1(\PID_CONTROLLER.err_prev[11] ), 
            .I2(n64[11]), .I3(n34201), .O(n57[11])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_11_add_2_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3062_5_lut (.I0(GND_net), .I1(n8159[2]), .I2(n410), .I3(n35375), 
            .O(n8133[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3062_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3057_17_lut (.I0(GND_net), .I1(n8019[14]), .I2(GND_net), 
            .I3(n35257), .O(n7988[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3057_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3431_11 (.CI(n35674), .I0(n16185[8]), .I1(GND_net), .CO(n35675));
    SB_LUT4 sub_11_inv_0_i21_1_lut (.I0(\PID_CONTROLLER.err[20] ), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n64[20]));   // verilog/motorControl.v(43[31:45])
    defparam sub_11_inv_0_i21_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i499_2_lut (.I0(\Kp[7] ), .I1(\PID_CONTROLLER.err[21] ), 
            .I2(GND_net), .I3(GND_net), .O(n743));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i499_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_3056_24 (.CI(n35052), .I0(n7988[21]), .I1(GND_net), .CO(n35053));
    SB_CARRY mult_10_add_2137_24 (.CI(n34722), .I0(n6542[21]), .I1(GND_net), 
            .CO(n34723));
    SB_LUT4 mult_10_i132_2_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err[0] ), 
            .I2(GND_net), .I3(GND_net), .O(n195));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i132_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_3223_7 (.CI(n34455), .I0(n12575[4]), .I1(n604_adj_3417), 
            .CO(n34456));
    SB_LUT4 add_3223_6_lut (.I0(GND_net), .I1(n12575[3]), .I2(n507_adj_3421), 
            .I3(n34454), .O(n11992[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3223_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_add_2137_23_lut (.I0(GND_net), .I1(n6542[20]), .I2(GND_net), 
            .I3(n34721), .O(n61[22])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_2137_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_2137_23 (.CI(n34721), .I0(n6542[20]), .I1(GND_net), 
            .CO(n34722));
    SB_LUT4 add_3056_23_lut (.I0(GND_net), .I1(n7988[20]), .I2(GND_net), 
            .I3(n35051), .O(n7956[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3056_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_add_2137_22_lut (.I0(GND_net), .I1(n6542[19]), .I2(GND_net), 
            .I3(n34720), .O(n61[21])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_2137_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_11_inv_0_i22_1_lut (.I0(\PID_CONTROLLER.err[21] ), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n64[21]));   // verilog/motorControl.v(43[31:45])
    defparam sub_11_inv_0_i22_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_11_inv_0_i23_1_lut (.I0(\PID_CONTROLLER.err[22] ), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n64[22]));   // verilog/motorControl.v(43[31:45])
    defparam sub_11_inv_0_i23_1_lut.LUT_INIT = 16'h5555;
    SB_DFF \PID_CONTROLLER.result_i0  (.Q(\PID_CONTROLLER.result [0]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.result_31__N_3003 [0]));   // verilog/motorControl.v(38[14] 59[8])
    SB_LUT4 sub_11_inv_0_i24_1_lut (.I0(\PID_CONTROLLER.err[23] ), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n64[23]));   // verilog/motorControl.v(43[31:45])
    defparam sub_11_inv_0_i24_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_3223_6 (.CI(n34454), .I0(n12575[3]), .I1(n507_adj_3421), 
            .CO(n34455));
    SB_LUT4 add_3464_2_lut (.I0(GND_net), .I1(n68), .I2(n161), .I3(GND_net), 
            .O(n16420[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3464_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3223_5_lut (.I0(GND_net), .I1(n12575[2]), .I2(n410_adj_3422), 
            .I3(n34453), .O(n11992[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3223_5_lut.LUT_INIT = 16'hC33C;
    SB_DFF \PID_CONTROLLER.err_i1  (.Q(\PID_CONTROLLER.err[0] ), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_31__N_2825 [0]));   // verilog/motorControl.v(38[14] 59[8])
    SB_DFF GATES_i2 (.Q(PIN_7_c_1), .C(clk32MHz), .D(GATES_5__N_2788[1]));   // verilog/motorControl.v(64[10] 111[6])
    SB_CARRY add_3223_5 (.CI(n34453), .I0(n12575[2]), .I1(n410_adj_3422), 
            .CO(n34454));
    SB_CARRY add_3464_2 (.CI(GND_net), .I0(n68), .I1(n161), .CO(n34361));
    SB_LUT4 sub_11_inv_0_i32_1_lut (.I0(\PID_CONTROLLER.err[31] ), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n64[26]));   // verilog/motorControl.v(43[31:45])
    defparam sub_11_inv_0_i32_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_3223_4_lut (.I0(GND_net), .I1(n12575[1]), .I2(n313_adj_3423), 
            .I3(n34452), .O(n11992[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3223_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3067_7_lut (.I0(GND_net), .I1(n8274[4]), .I2(n619), .I3(n35482), 
            .O(n8253[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3067_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 state_23__I_0_inv_0_i1_1_lut (.I0(setpoint[0]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n58[0]));   // verilog/motorControl.v(39[14:30])
    defparam state_23__I_0_inv_0_i1_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY mult_10_add_2137_22 (.CI(n34720), .I0(n6542[19]), .I1(GND_net), 
            .CO(n34721));
    SB_CARRY add_3057_17 (.CI(n35257), .I0(n8019[14]), .I1(GND_net), .CO(n35258));
    SB_CARRY add_3056_23 (.CI(n35051), .I0(n7988[20]), .I1(GND_net), .CO(n35052));
    SB_LUT4 mult_10_i87_2_lut (.I0(\Kp[1] ), .I1(\PID_CONTROLLER.err[10] ), 
            .I2(GND_net), .I3(GND_net), .O(n128_adj_3384));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i87_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_add_2137_21_lut (.I0(GND_net), .I1(n6542[18]), .I2(GND_net), 
            .I3(n34719), .O(n61[20])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_2137_21_lut.LUT_INIT = 16'hC33C;
    SB_DFF GATES_i1 (.Q(PIN_6_c_0), .C(clk32MHz), .D(GATES_5__N_2788[0]));   // verilog/motorControl.v(64[10] 111[6])
    SB_LUT4 add_3315_21_lut (.I0(GND_net), .I1(n14434[18]), .I2(GND_net), 
            .I3(n34360), .O(n14035[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3315_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3056_22_lut (.I0(GND_net), .I1(n7988[19]), .I2(GND_net), 
            .I3(n35050), .O(n7956[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3056_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3062_5 (.CI(n35375), .I0(n8159[2]), .I1(n410), .CO(n35376));
    SB_CARRY sub_11_add_2_13 (.CI(n34201), .I0(\PID_CONTROLLER.err_prev[11] ), 
            .I1(n64[11]), .CO(n34202));
    SB_LUT4 add_3315_20_lut (.I0(GND_net), .I1(n14434[17]), .I2(GND_net), 
            .I3(n34359), .O(n14035[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3315_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3056_22 (.CI(n35050), .I0(n7988[19]), .I1(GND_net), .CO(n35051));
    SB_LUT4 add_3057_16_lut (.I0(GND_net), .I1(n8019[13]), .I2(GND_net), 
            .I3(n35256), .O(n7988[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3057_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_2137_21 (.CI(n34719), .I0(n6542[18]), .I1(GND_net), 
            .CO(n34720));
    SB_CARRY add_3223_4 (.CI(n34452), .I0(n12575[1]), .I1(n313_adj_3423), 
            .CO(n34453));
    SB_CARRY add_3057_16 (.CI(n35256), .I0(n8019[13]), .I1(GND_net), .CO(n35257));
    SB_LUT4 add_3223_3_lut (.I0(GND_net), .I1(n12575[0]), .I2(n216), .I3(n34451), 
            .O(n11992[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3223_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3223_3 (.CI(n34451), .I0(n12575[0]), .I1(n216), .CO(n34452));
    SB_LUT4 add_3056_21_lut (.I0(GND_net), .I1(n7988[18]), .I2(GND_net), 
            .I3(n35049), .O(n7956[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3056_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3315_20 (.CI(n34359), .I0(n14434[17]), .I1(GND_net), 
            .CO(n34360));
    SB_LUT4 mult_10_add_2137_20_lut (.I0(GND_net), .I1(n6542[17]), .I2(GND_net), 
            .I3(n34718), .O(n61[19])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_2137_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_11_add_2_12_lut (.I0(GND_net), .I1(\PID_CONTROLLER.err_prev[10] ), 
            .I2(n64[10]), .I3(n34200), .O(n57[10])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_11_add_2_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3056_21 (.CI(n35049), .I0(n7988[18]), .I1(GND_net), .CO(n35050));
    SB_CARRY mult_10_add_2137_20 (.CI(n34718), .I0(n6542[17]), .I1(GND_net), 
            .CO(n34719));
    SB_LUT4 add_3223_2_lut (.I0(GND_net), .I1(n26_adj_3425), .I2(n119), 
            .I3(GND_net), .O(n11992[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3223_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3223_2 (.CI(GND_net), .I0(n26_adj_3425), .I1(n119), .CO(n34451));
    SB_LUT4 mult_10_add_2137_19_lut (.I0(GND_net), .I1(n6542[16]), .I2(GND_net), 
            .I3(n34717), .O(n61[18])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_2137_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i24_2_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err[11] ), 
            .I2(GND_net), .I3(GND_net), .O(n35_adj_3383));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i24_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 state_23__I_0_inv_0_i2_1_lut (.I0(setpoint[1]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n58[1]));   // verilog/motorControl.v(39[14:30])
    defparam state_23__I_0_inv_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_11_inv_0_i7_1_lut (.I0(\PID_CONTROLLER.err[6] ), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n64[6]));   // verilog/motorControl.v(43[31:45])
    defparam sub_11_inv_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_3064_22_lut (.I0(GND_net), .I1(n8208[19]), .I2(GND_net), 
            .I3(n35437), .O(n8184[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3064_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_2137_19 (.CI(n34717), .I0(n6542[16]), .I1(GND_net), 
            .CO(n34718));
    SB_LUT4 add_3062_4_lut (.I0(GND_net), .I1(n8159[1]), .I2(n313_adj_3426), 
            .I3(n35374), .O(n8133[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3062_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3067_7 (.CI(n35482), .I0(n8274[4]), .I1(n619), .CO(n35483));
    SB_LUT4 add_3057_15_lut (.I0(GND_net), .I1(n8019[12]), .I2(GND_net), 
            .I3(n35255), .O(n7988[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3057_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_12_i351_2_lut (.I0(\Kd[5] ), .I1(n57[12]), .I2(GND_net), 
            .I3(GND_net), .O(n522));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i351_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_3064_22 (.CI(n35437), .I0(n8208[19]), .I1(GND_net), .CO(n35438));
    SB_LUT4 mult_10_i197_2_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err[0] ), 
            .I2(GND_net), .I3(GND_net), .O(n292));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i197_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_3062_4 (.CI(n35374), .I0(n8159[1]), .I1(n313_adj_3426), 
            .CO(n35375));
    SB_LUT4 mult_10_add_2137_18_lut (.I0(GND_net), .I1(n6542[15]), .I2(GND_net), 
            .I3(n34716), .O(n61[17])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_2137_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i152_2_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err[10] ), 
            .I2(GND_net), .I3(GND_net), .O(n225));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i152_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 state_23__I_0_inv_0_i3_1_lut (.I0(setpoint[2]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n58[2]));   // verilog/motorControl.v(39[14:30])
    defparam state_23__I_0_inv_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_3379_10_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [9]), 
            .I2(GND_net), .I3(n34450), .O(n15226[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3379_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3379_9_lut (.I0(GND_net), .I1(n583), .I2(GND_net), .I3(n34449), 
            .O(n15226[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3379_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i217_2_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err[10] ), 
            .I2(GND_net), .I3(GND_net), .O(n322));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i217_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY mult_10_add_2137_18 (.CI(n34716), .I0(n6542[15]), .I1(GND_net), 
            .CO(n34717));
    SB_CARRY add_3379_9 (.CI(n34449), .I0(n583), .I1(GND_net), .CO(n34450));
    SB_LUT4 state_23__I_0_inv_0_i4_1_lut (.I0(setpoint[3]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n58[3]));   // verilog/motorControl.v(39[14:30])
    defparam state_23__I_0_inv_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_3379_8_lut (.I0(GND_net), .I1(n510), .I2(n545), .I3(n34448), 
            .O(n15226[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3379_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3057_15 (.CI(n35255), .I0(n8019[12]), .I1(GND_net), .CO(n35256));
    SB_LUT4 mult_10_i282_2_lut (.I0(\Kp[4] ), .I1(\PID_CONTROLLER.err[10] ), 
            .I2(GND_net), .I3(GND_net), .O(n419));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i282_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_add_2137_17_lut (.I0(GND_net), .I1(n6542[14]), .I2(GND_net), 
            .I3(n34715), .O(n61[16])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_2137_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3379_8 (.CI(n34448), .I0(n510), .I1(n545), .CO(n34449));
    SB_LUT4 state_23__I_0_inv_0_i5_1_lut (.I0(setpoint[4]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n58[4]));   // verilog/motorControl.v(39[14:30])
    defparam state_23__I_0_inv_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_3379_7_lut (.I0(GND_net), .I1(n437), .I2(n472), .I3(n34447), 
            .O(n15226[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3379_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_11_inv_0_i8_1_lut (.I0(\PID_CONTROLLER.err[7] ), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n64[7]));   // verilog/motorControl.v(43[31:45])
    defparam sub_11_inv_0_i8_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY mult_10_add_2137_17 (.CI(n34715), .I0(n6542[14]), .I1(GND_net), 
            .CO(n34716));
    SB_CARRY add_3379_7 (.CI(n34447), .I0(n437), .I1(n472), .CO(n34448));
    SB_LUT4 mult_10_i347_2_lut (.I0(\Kp[5] ), .I1(\PID_CONTROLLER.err[10] ), 
            .I2(GND_net), .I3(GND_net), .O(n516));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i347_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i262_2_lut (.I0(\Kp[4] ), .I1(\PID_CONTROLLER.err[0] ), 
            .I2(GND_net), .I3(GND_net), .O(n389));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i262_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_3057_14_lut (.I0(GND_net), .I1(n8019[11]), .I2(GND_net), 
            .I3(n35254), .O(n7988[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3057_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3056_20_lut (.I0(GND_net), .I1(n7988[17]), .I2(GND_net), 
            .I3(n35048), .O(n7956[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3056_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_add_2137_16_lut (.I0(GND_net), .I1(n6542[13]), .I2(GND_net), 
            .I3(n34714), .O(n61[15])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_2137_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3379_6_lut (.I0(GND_net), .I1(n364), .I2(n399), .I3(n34446), 
            .O(n15226[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3379_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3379_6 (.CI(n34446), .I0(n364), .I1(n399), .CO(n34447));
    SB_CARRY mult_10_add_2137_16 (.CI(n34714), .I0(n6542[13]), .I1(GND_net), 
            .CO(n34715));
    SB_CARRY add_3056_20 (.CI(n35048), .I0(n7988[17]), .I1(GND_net), .CO(n35049));
    SB_LUT4 mult_10_add_2137_15_lut (.I0(GND_net), .I1(n6542[12]), .I2(GND_net), 
            .I3(n34713), .O(n61[14])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_2137_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3379_5_lut (.I0(GND_net), .I1(n291), .I2(n326), .I3(n34445), 
            .O(n15226[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3379_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3379_5 (.CI(n34445), .I0(n291), .I1(n326), .CO(n34446));
    SB_CARRY mult_10_add_2137_15 (.CI(n34713), .I0(n6542[12]), .I1(GND_net), 
            .CO(n34714));
    SB_CARRY add_3057_14 (.CI(n35254), .I0(n8019[11]), .I1(GND_net), .CO(n35255));
    SB_LUT4 add_3056_19_lut (.I0(GND_net), .I1(n7988[16]), .I2(GND_net), 
            .I3(n35047), .O(n7956[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3056_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_add_2137_14_lut (.I0(GND_net), .I1(n6542[11]), .I2(GND_net), 
            .I3(n34712), .O(n61[13])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_2137_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i412_2_lut (.I0(\Kp[6] ), .I1(\PID_CONTROLLER.err[10] ), 
            .I2(GND_net), .I3(GND_net), .O(n613));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i412_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i477_2_lut (.I0(\Kp[7] ), .I1(\PID_CONTROLLER.err[10] ), 
            .I2(GND_net), .I3(GND_net), .O(n710));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i477_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_3379_4_lut (.I0(GND_net), .I1(n218), .I2(n253), .I3(n34444), 
            .O(n15226[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3379_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 state_23__I_0_inv_0_i6_1_lut (.I0(setpoint[5]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n58[5]));   // verilog/motorControl.v(39[14:30])
    defparam state_23__I_0_inv_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_3056_19 (.CI(n35047), .I0(n7988[16]), .I1(GND_net), .CO(n35048));
    SB_CARRY add_3379_4 (.CI(n34444), .I0(n218), .I1(n253), .CO(n34445));
    SB_LUT4 mult_10_i327_2_lut (.I0(\Kp[5] ), .I1(\PID_CONTROLLER.err[0] ), 
            .I2(GND_net), .I3(GND_net), .O(n486));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i327_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 state_23__I_0_inv_0_i7_1_lut (.I0(setpoint[6]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n58[6]));   // verilog/motorControl.v(39[14:30])
    defparam state_23__I_0_inv_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_3379_3_lut (.I0(GND_net), .I1(n145), .I2(n180), .I3(n34443), 
            .O(n15226[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3379_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_2137_14 (.CI(n34712), .I0(n6542[11]), .I1(GND_net), 
            .CO(n34713));
    SB_CARRY sub_11_add_2_12 (.CI(n34200), .I0(\PID_CONTROLLER.err_prev[10] ), 
            .I1(n64[10]), .CO(n34201));
    SB_LUT4 mult_10_add_2137_13_lut (.I0(GND_net), .I1(n6542[10]), .I2(GND_net), 
            .I3(n34711), .O(n61[12])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_2137_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3062_3_lut (.I0(GND_net), .I1(n8159[0]), .I2(n216_adj_3429), 
            .I3(n35373), .O(n8133[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3062_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3056_18_lut (.I0(GND_net), .I1(n7988[15]), .I2(GND_net), 
            .I3(n35046), .O(n7956[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3056_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3074_2 (.CI(GND_net), .I0(n62), .I1(n155_adj_3414), .CO(n35583));
    SB_LUT4 add_3315_19_lut (.I0(GND_net), .I1(n14434[16]), .I2(GND_net), 
            .I3(n34358), .O(n14035[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3315_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_2137_13 (.CI(n34711), .I0(n6542[10]), .I1(GND_net), 
            .CO(n34712));
    SB_CARRY add_3379_3 (.CI(n34443), .I0(n145), .I1(n180), .CO(n34444));
    SB_LUT4 add_3379_2_lut (.I0(GND_net), .I1(n72), .I2(n107), .I3(GND_net), 
            .O(n15226[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3379_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_add_2137_12_lut (.I0(GND_net), .I1(n6542[9]), .I2(GND_net), 
            .I3(n34710), .O(n61[11])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_2137_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3062_3 (.CI(n35373), .I0(n8159[0]), .I1(n216_adj_3429), 
            .CO(n35374));
    SB_LUT4 add_3431_10_lut (.I0(GND_net), .I1(n16185[7]), .I2(GND_net), 
            .I3(n35673), .O(n16031[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3431_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i140_2_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err[4] ), 
            .I2(GND_net), .I3(GND_net), .O(n207_adj_3379));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i140_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_3073_14_lut (.I0(GND_net), .I1(n8379[11]), .I2(GND_net), 
            .I3(n35582), .O(n8364[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3073_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3057_13_lut (.I0(GND_net), .I1(n8019[10]), .I2(GND_net), 
            .I3(n35253), .O(n7988[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3057_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3056_18 (.CI(n35046), .I0(n7988[15]), .I1(GND_net), .CO(n35047));
    SB_LUT4 add_3073_13_lut (.I0(GND_net), .I1(n8379[10]), .I2(GND_net), 
            .I3(n35581), .O(n8364[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3073_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_2137_12 (.CI(n34710), .I0(n6542[9]), .I1(GND_net), 
            .CO(n34711));
    SB_LUT4 mult_10_add_2137_11_lut (.I0(GND_net), .I1(n6542[8]), .I2(GND_net), 
            .I3(n34709), .O(n61[10])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_2137_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3379_2 (.CI(GND_net), .I0(n72), .I1(n107), .CO(n34443));
    SB_LUT4 sub_11_add_2_11_lut (.I0(GND_net), .I1(\PID_CONTROLLER.err_prev[9] ), 
            .I2(n64[9]), .I3(n34199), .O(n57[9])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_11_add_2_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3248_24_lut (.I0(GND_net), .I1(n13109[21]), .I2(GND_net), 
            .I3(n34442), .O(n12575[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3248_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3073_13 (.CI(n35581), .I0(n8379[10]), .I1(GND_net), .CO(n35582));
    SB_CARRY mult_10_add_2137_11 (.CI(n34709), .I0(n6542[8]), .I1(GND_net), 
            .CO(n34710));
    SB_LUT4 add_3056_17_lut (.I0(GND_net), .I1(n7988[14]), .I2(GND_net), 
            .I3(n35045), .O(n7956[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3056_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3315_19 (.CI(n34358), .I0(n14434[16]), .I1(GND_net), 
            .CO(n34359));
    SB_LUT4 mult_10_i205_2_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err[4] ), 
            .I2(GND_net), .I3(GND_net), .O(n304_adj_3378));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i205_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY sub_11_add_2_11 (.CI(n34199), .I0(\PID_CONTROLLER.err_prev[9] ), 
            .I1(n64[9]), .CO(n34200));
    SB_CARRY add_3057_13 (.CI(n35253), .I0(n8019[10]), .I1(GND_net), .CO(n35254));
    SB_LUT4 add_3057_12_lut (.I0(GND_net), .I1(n8019[9]), .I2(GND_net), 
            .I3(n35252), .O(n7988[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3057_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_add_2137_10_lut (.I0(GND_net), .I1(n6542[7]), .I2(GND_net), 
            .I3(n34708), .O(n61[9])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_2137_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3248_23_lut (.I0(GND_net), .I1(n13109[20]), .I2(GND_net), 
            .I3(n34441), .O(n12575[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3248_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3069_14 (.CI(n35524), .I0(n8313[11]), .I1(GND_net), .CO(n35525));
    SB_CARRY add_3248_23 (.CI(n34441), .I0(n13109[20]), .I1(GND_net), 
            .CO(n34442));
    SB_CARRY mult_10_add_2137_10 (.CI(n34708), .I0(n6542[7]), .I1(GND_net), 
            .CO(n34709));
    SB_LUT4 sub_11_add_2_10_lut (.I0(GND_net), .I1(\PID_CONTROLLER.err_prev[8] ), 
            .I2(n64[8]), .I3(n34198), .O(n57[8])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_11_add_2_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3057_12 (.CI(n35252), .I0(n8019[9]), .I1(GND_net), .CO(n35253));
    SB_CARRY add_3056_17 (.CI(n35045), .I0(n7988[14]), .I1(GND_net), .CO(n35046));
    SB_LUT4 mult_10_add_2137_9_lut (.I0(GND_net), .I1(n6542[6]), .I2(GND_net), 
            .I3(n34707), .O(n61[8])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_2137_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_11_add_2_10 (.CI(n34198), .I0(\PID_CONTROLLER.err_prev[8] ), 
            .I1(n64[8]), .CO(n34199));
    SB_LUT4 add_3248_22_lut (.I0(GND_net), .I1(n13109[19]), .I2(GND_net), 
            .I3(n34440), .O(n12575[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3248_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3248_22 (.CI(n34440), .I0(n13109[19]), .I1(GND_net), 
            .CO(n34441));
    SB_CARRY mult_10_add_2137_9 (.CI(n34707), .I0(n6542[6]), .I1(GND_net), 
            .CO(n34708));
    SB_LUT4 add_3056_16_lut (.I0(GND_net), .I1(n7988[13]), .I2(GND_net), 
            .I3(n35044), .O(n7956[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3056_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3062_2_lut (.I0(GND_net), .I1(n26_adj_3432), .I2(n119_adj_3433), 
            .I3(GND_net), .O(n8133[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3062_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_add_2137_8_lut (.I0(GND_net), .I1(n6542[5]), .I2(n680), 
            .I3(n34706), .O(n61[7])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_2137_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3248_21_lut (.I0(GND_net), .I1(n13109[18]), .I2(GND_net), 
            .I3(n34439), .O(n12575[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3248_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3248_21 (.CI(n34439), .I0(n13109[18]), .I1(GND_net), 
            .CO(n34440));
    SB_CARRY mult_10_add_2137_8 (.CI(n34706), .I0(n6542[5]), .I1(n680), 
            .CO(n34707));
    SB_LUT4 add_3064_21_lut (.I0(GND_net), .I1(n8208[18]), .I2(GND_net), 
            .I3(n35436), .O(n8184[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3064_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3431_10 (.CI(n35673), .I0(n16185[7]), .I1(GND_net), .CO(n35674));
    SB_CARRY add_3062_2 (.CI(GND_net), .I0(n26_adj_3432), .I1(n119_adj_3433), 
            .CO(n35373));
    SB_LUT4 add_3057_11_lut (.I0(GND_net), .I1(n8019[8]), .I2(GND_net), 
            .I3(n35251), .O(n7988[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3057_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3056_16 (.CI(n35044), .I0(n7988[13]), .I1(GND_net), .CO(n35045));
    SB_LUT4 add_3056_15_lut (.I0(GND_net), .I1(n7988[12]), .I2(GND_net), 
            .I3(n35043), .O(n7956[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3056_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_add_2137_7_lut (.I0(GND_net), .I1(n6542[4]), .I2(n583_adj_3434), 
            .I3(n34705), .O(n61[6])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_2137_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3248_20_lut (.I0(GND_net), .I1(n13109[17]), .I2(GND_net), 
            .I3(n34438), .O(n12575[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3248_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3248_20 (.CI(n34438), .I0(n13109[17]), .I1(GND_net), 
            .CO(n34439));
    SB_CARRY mult_10_add_2137_7 (.CI(n34705), .I0(n6542[4]), .I1(n583_adj_3434), 
            .CO(n34706));
    SB_CARRY add_3057_11 (.CI(n35251), .I0(n8019[8]), .I1(GND_net), .CO(n35252));
    SB_CARRY add_3056_15 (.CI(n35043), .I0(n7988[12]), .I1(GND_net), .CO(n35044));
    SB_LUT4 add_3056_14_lut (.I0(GND_net), .I1(n7988[11]), .I2(GND_net), 
            .I3(n35042), .O(n7956[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3056_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_add_2137_6_lut (.I0(GND_net), .I1(n6542[3]), .I2(n486), 
            .I3(n34704), .O(n61[5])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_2137_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_2137_6 (.CI(n34704), .I0(n6542[3]), .I1(n486), 
            .CO(n34705));
    SB_LUT4 mult_10_add_2137_5_lut (.I0(GND_net), .I1(n6542[2]), .I2(n389), 
            .I3(n34703), .O(n61[4])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_2137_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3315_18_lut (.I0(GND_net), .I1(n14434[15]), .I2(GND_net), 
            .I3(n34357), .O(n14035[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3315_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3248_19_lut (.I0(GND_net), .I1(n13109[16]), .I2(GND_net), 
            .I3(n34437), .O(n12575[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3248_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_11_add_2_9_lut (.I0(GND_net), .I1(\PID_CONTROLLER.err_prev[7] ), 
            .I2(n64[7]), .I3(n34197), .O(n57[7])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_11_add_2_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 state_23__I_0_inv_0_i8_1_lut (.I0(setpoint[7]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n58[7]));   // verilog/motorControl.v(39[14:30])
    defparam state_23__I_0_inv_0_i8_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_3248_19 (.CI(n34437), .I0(n13109[16]), .I1(GND_net), 
            .CO(n34438));
    SB_CARRY add_3315_18 (.CI(n34357), .I0(n14434[15]), .I1(GND_net), 
            .CO(n34358));
    SB_CARRY mult_10_add_2137_5 (.CI(n34703), .I0(n6542[2]), .I1(n389), 
            .CO(n34704));
    SB_LUT4 add_3315_17_lut (.I0(GND_net), .I1(n14434[14]), .I2(GND_net), 
            .I3(n34356), .O(n14035[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3315_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3315_17 (.CI(n34356), .I0(n14434[14]), .I1(GND_net), 
            .CO(n34357));
    SB_LUT4 add_3057_10_lut (.I0(GND_net), .I1(n8019[7]), .I2(GND_net), 
            .I3(n35250), .O(n7988[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3057_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3056_14 (.CI(n35042), .I0(n7988[11]), .I1(GND_net), .CO(n35043));
    SB_LUT4 mult_10_add_2137_4_lut (.I0(GND_net), .I1(n6542[1]), .I2(n292), 
            .I3(n34702), .O(n61[3])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_2137_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_11_add_2_9 (.CI(n34197), .I0(\PID_CONTROLLER.err_prev[7] ), 
            .I1(n64[7]), .CO(n34198));
    SB_LUT4 add_3067_6_lut (.I0(GND_net), .I1(n8274[3]), .I2(n522), .I3(n35481), 
            .O(n8253[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3067_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_11_add_2_8_lut (.I0(GND_net), .I1(\PID_CONTROLLER.err_prev[6] ), 
            .I2(n64[6]), .I3(n34196), .O(n57[6])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_11_add_2_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3056_13_lut (.I0(GND_net), .I1(n7988[10]), .I2(GND_net), 
            .I3(n35041), .O(n7956[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3056_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i392_2_lut (.I0(\Kp[6] ), .I1(\PID_CONTROLLER.err[0] ), 
            .I2(GND_net), .I3(GND_net), .O(n583_adj_3434));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i392_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i457_2_lut (.I0(\Kp[7] ), .I1(\PID_CONTROLLER.err[0] ), 
            .I2(GND_net), .I3(GND_net), .O(n680));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i457_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i81_2_lut (.I0(\Kd[1] ), .I1(n57[7]), .I2(GND_net), 
            .I3(GND_net), .O(n119_adj_3433));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i81_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i18_2_lut (.I0(\Kd[0] ), .I1(n57[8]), .I2(GND_net), 
            .I3(GND_net), .O(n26_adj_3432));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i18_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 state_23__I_0_inv_0_i9_1_lut (.I0(setpoint[8]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n58[8]));   // verilog/motorControl.v(39[14:30])
    defparam state_23__I_0_inv_0_i9_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_11_inv_0_i9_1_lut (.I0(\PID_CONTROLLER.err[8] ), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n64[8]));   // verilog/motorControl.v(43[31:45])
    defparam sub_11_inv_0_i9_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY sub_11_add_2_8 (.CI(n34196), .I0(\PID_CONTROLLER.err_prev[6] ), 
            .I1(n64[6]), .CO(n34197));
    SB_CARRY mult_10_add_2137_4 (.CI(n34702), .I0(n6542[1]), .I1(n292), 
            .CO(n34703));
    SB_LUT4 add_3248_18_lut (.I0(GND_net), .I1(n13109[15]), .I2(GND_net), 
            .I3(n34436), .O(n12575[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3248_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3315_16_lut (.I0(GND_net), .I1(n14434[13]), .I2(GND_net), 
            .I3(n34355), .O(n14035[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3315_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3315_16 (.CI(n34355), .I0(n14434[13]), .I1(GND_net), 
            .CO(n34356));
    SB_LUT4 add_3315_15_lut (.I0(GND_net), .I1(n14434[12]), .I2(GND_net), 
            .I3(n34354), .O(n14035[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3315_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3248_18 (.CI(n34436), .I0(n13109[15]), .I1(GND_net), 
            .CO(n34437));
    SB_LUT4 mult_10_i270_2_lut (.I0(\Kp[4] ), .I1(\PID_CONTROLLER.err[4] ), 
            .I2(GND_net), .I3(GND_net), .O(n401));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i270_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_add_2137_3_lut (.I0(GND_net), .I1(n6542[0]), .I2(n195), 
            .I3(n34701), .O(n61[2])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_2137_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3056_13 (.CI(n35041), .I0(n7988[10]), .I1(GND_net), .CO(n35042));
    SB_LUT4 add_3056_12_lut (.I0(GND_net), .I1(n7988[9]), .I2(GND_net), 
            .I3(n35040), .O(n7956[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3056_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_2137_3 (.CI(n34701), .I0(n6542[0]), .I1(n195), 
            .CO(n34702));
    SB_CARRY add_3064_21 (.CI(n35436), .I0(n8208[18]), .I1(GND_net), .CO(n35437));
    SB_LUT4 add_3248_17_lut (.I0(GND_net), .I1(n13109[14]), .I2(GND_net), 
            .I3(n34435), .O(n12575[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3248_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_11_add_2_7_lut (.I0(GND_net), .I1(\PID_CONTROLLER.err_prev[5] ), 
            .I2(n64[5]), .I3(n34195), .O(n57[5])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_11_add_2_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3061_26_lut (.I0(GND_net), .I1(n8133[23]), .I2(GND_net), 
            .I3(n35372), .O(n8106[24])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3061_26_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3061_25_lut (.I0(GND_net), .I1(n8133[22]), .I2(GND_net), 
            .I3(n35371), .O(n8106[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3061_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 state_23__I_0_inv_0_i10_1_lut (.I0(setpoint[9]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n58[9]));   // verilog/motorControl.v(39[14:30])
    defparam state_23__I_0_inv_0_i10_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_3248_17 (.CI(n34435), .I0(n13109[14]), .I1(GND_net), 
            .CO(n34436));
    SB_LUT4 mult_10_add_2137_2_lut (.I0(GND_net), .I1(n5), .I2(n98), .I3(GND_net), 
            .O(n61[1])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_2137_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3057_10 (.CI(n35250), .I0(n8019[7]), .I1(GND_net), .CO(n35251));
    SB_CARRY add_3061_25 (.CI(n35371), .I0(n8133[22]), .I1(GND_net), .CO(n35372));
    SB_LUT4 add_3057_9_lut (.I0(GND_net), .I1(n8019[6]), .I2(GND_net), 
            .I3(n35249), .O(n7988[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3057_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3056_12 (.CI(n35040), .I0(n7988[9]), .I1(GND_net), .CO(n35041));
    SB_CARRY add_3067_6 (.CI(n35481), .I0(n8274[3]), .I1(n522), .CO(n35482));
    SB_CARRY mult_10_add_2137_2 (.CI(GND_net), .I0(n5), .I1(n98), .CO(n34701));
    SB_LUT4 add_3067_5_lut (.I0(GND_net), .I1(n8274[2]), .I2(n425), .I3(n35480), 
            .O(n8253[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3067_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3061_24_lut (.I0(GND_net), .I1(n8133[21]), .I2(GND_net), 
            .I3(n35370), .O(n8106[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3061_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3064_20_lut (.I0(GND_net), .I1(n8208[17]), .I2(GND_net), 
            .I3(n35435), .O(n8184[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3064_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3067_5 (.CI(n35480), .I0(n8274[2]), .I1(n425), .CO(n35481));
    SB_CARRY add_3064_20 (.CI(n35435), .I0(n8208[17]), .I1(GND_net), .CO(n35436));
    SB_CARRY add_3061_24 (.CI(n35370), .I0(n8133[21]), .I1(GND_net), .CO(n35371));
    SB_LUT4 add_3064_19_lut (.I0(GND_net), .I1(n8208[16]), .I2(GND_net), 
            .I3(n35434), .O(n8184[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3064_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3067_4_lut (.I0(GND_net), .I1(n8274[1]), .I2(n328), .I3(n35479), 
            .O(n8253[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3067_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3069_13_lut (.I0(GND_net), .I1(n8313[10]), .I2(GND_net), 
            .I3(n35523), .O(n8294[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3069_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3248_16_lut (.I0(GND_net), .I1(n13109[13]), .I2(GND_net), 
            .I3(n34434), .O(n12575[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3248_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3067_4 (.CI(n35479), .I0(n8274[1]), .I1(n328), .CO(n35480));
    SB_LUT4 add_3067_3_lut (.I0(GND_net), .I1(n8274[0]), .I2(n231), .I3(n35478), 
            .O(n8253[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3067_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3069_13 (.CI(n35523), .I0(n8313[10]), .I1(GND_net), .CO(n35524));
    SB_LUT4 add_3073_12_lut (.I0(GND_net), .I1(n8379[9]), .I2(GND_net), 
            .I3(n35580), .O(n8364[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3073_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3057_9 (.CI(n35249), .I0(n8019[6]), .I1(GND_net), .CO(n35250));
    SB_LUT4 add_3061_23_lut (.I0(GND_net), .I1(n8133[20]), .I2(GND_net), 
            .I3(n35369), .O(n8106[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3061_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3073_12 (.CI(n35580), .I0(n8379[9]), .I1(GND_net), .CO(n35581));
    SB_LUT4 add_3069_12_lut (.I0(GND_net), .I1(n8313[9]), .I2(GND_net), 
            .I3(n35522), .O(n8294[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3069_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_11_inv_0_i10_1_lut (.I0(\PID_CONTROLLER.err[9] ), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n64[9]));   // verilog/motorControl.v(43[31:45])
    defparam sub_11_inv_0_i10_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_3057_8_lut (.I0(GND_net), .I1(n8019[5]), .I2(n686), .I3(n35248), 
            .O(n7988[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3057_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i29032_3_lut_4_lut (.I0(\PWMLimit[3] ), .I1(\PID_CONTROLLER.result [3]), 
            .I2(\PID_CONTROLLER.result [2]), .I3(\PWMLimit[2] ), .O(n44552));   // verilog/motorControl.v(45[12:27])
    defparam i29032_3_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_CARRY add_3067_3 (.CI(n35478), .I0(n8274[0]), .I1(n231), .CO(n35479));
    SB_LUT4 add_3067_2_lut (.I0(GND_net), .I1(n41), .I2(n134), .I3(GND_net), 
            .O(n8253[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3067_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3431_9_lut (.I0(GND_net), .I1(n16185[6]), .I2(GND_net), 
            .I3(n35672), .O(n16031[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3431_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3064_19 (.CI(n35434), .I0(n8208[16]), .I1(GND_net), .CO(n35435));
    SB_LUT4 add_3073_11_lut (.I0(GND_net), .I1(n8379[8]), .I2(GND_net), 
            .I3(n35579), .O(n8364[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3073_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3248_16 (.CI(n34434), .I0(n13109[13]), .I1(GND_net), 
            .CO(n34435));
    SB_CARRY add_3061_23 (.CI(n35369), .I0(n8133[20]), .I1(GND_net), .CO(n35370));
    SB_LUT4 mult_14_i49_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral [9]), 
            .I2(GND_net), .I3(GND_net), .O(n72));   // verilog/motorControl.v(43[48:59])
    defparam mult_14_i49_2_lut.LUT_INIT = 16'h4444;
    SB_CARRY add_3057_8 (.CI(n35248), .I0(n8019[5]), .I1(n686), .CO(n35249));
    SB_CARRY add_3315_15 (.CI(n34354), .I0(n14434[12]), .I1(GND_net), 
            .CO(n34355));
    SB_CARRY add_3073_11 (.CI(n35579), .I0(n8379[8]), .I1(GND_net), .CO(n35580));
    SB_LUT4 add_3056_11_lut (.I0(GND_net), .I1(n7988[8]), .I2(GND_net), 
            .I3(n35039), .O(n7956[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3056_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3069_12 (.CI(n35522), .I0(n8313[9]), .I1(GND_net), .CO(n35523));
    SB_LUT4 state_23__I_0_inv_0_i11_1_lut (.I0(setpoint[10]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n58[10]));   // verilog/motorControl.v(39[14:30])
    defparam state_23__I_0_inv_0_i11_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_3056_11 (.CI(n35039), .I0(n7988[8]), .I1(GND_net), .CO(n35040));
    SB_LUT4 add_3056_10_lut (.I0(GND_net), .I1(n7988[7]), .I2(GND_net), 
            .I3(n35038), .O(n7956[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3056_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3069_11_lut (.I0(GND_net), .I1(n8313[8]), .I2(GND_net), 
            .I3(n35521), .O(n8294[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3069_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_11_add_2_7 (.CI(n34195), .I0(\PID_CONTROLLER.err_prev[5] ), 
            .I1(n64[5]), .CO(n34196));
    SB_LUT4 mult_12_i146_2_lut (.I0(\Kd[2] ), .I1(n57[7]), .I2(GND_net), 
            .I3(GND_net), .O(n216_adj_3429));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i146_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_3057_7_lut (.I0(GND_net), .I1(n8019[4]), .I2(n589), .I3(n35247), 
            .O(n7988[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3057_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3248_15_lut (.I0(GND_net), .I1(n13109[12]), .I2(GND_net), 
            .I3(n34433), .O(n12575[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3248_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_11_add_2_6_lut (.I0(GND_net), .I1(\PID_CONTROLLER.err_prev[4] ), 
            .I2(n64[4]), .I3(n34194), .O(n57[4])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_11_add_2_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3056_10 (.CI(n35038), .I0(n7988[7]), .I1(GND_net), .CO(n35039));
    SB_LUT4 add_3061_22_lut (.I0(GND_net), .I1(n8133[19]), .I2(GND_net), 
            .I3(n35368), .O(n8106[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3061_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 state_23__I_0_inv_0_i12_1_lut (.I0(setpoint[11]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n58[11]));   // verilog/motorControl.v(39[14:30])
    defparam state_23__I_0_inv_0_i12_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_3057_7 (.CI(n35247), .I0(n8019[4]), .I1(n589), .CO(n35248));
    SB_LUT4 LessThan_20_i6_3_lut_3_lut (.I0(\PWMLimit[3] ), .I1(\PID_CONTROLLER.result [3]), 
            .I2(\PID_CONTROLLER.result [2]), .I3(GND_net), .O(n6));   // verilog/motorControl.v(45[12:27])
    defparam LessThan_20_i6_3_lut_3_lut.LUT_INIT = 16'hd4d4;
    SB_CARRY add_3069_11 (.CI(n35521), .I0(n8313[8]), .I1(GND_net), .CO(n35522));
    SB_CARRY add_3248_15 (.CI(n34433), .I0(n13109[12]), .I1(GND_net), 
            .CO(n34434));
    SB_LUT4 add_3248_14_lut (.I0(GND_net), .I1(n13109[11]), .I2(GND_net), 
            .I3(n34432), .O(n12575[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3248_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3248_14 (.CI(n34432), .I0(n13109[11]), .I1(GND_net), 
            .CO(n34433));
    SB_LUT4 add_3073_10_lut (.I0(GND_net), .I1(n8379[7]), .I2(GND_net), 
            .I3(n35578), .O(n8364[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3073_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3073_10 (.CI(n35578), .I0(n8379[7]), .I1(GND_net), .CO(n35579));
    SB_LUT4 add_3056_9_lut (.I0(GND_net), .I1(n7988[6]), .I2(GND_net), 
            .I3(n35037), .O(n7956[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3056_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3057_6_lut (.I0(GND_net), .I1(n8019[3]), .I2(n492), .I3(n35246), 
            .O(n7988[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3057_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3431_9 (.CI(n35672), .I0(n16185[6]), .I1(GND_net), .CO(n35673));
    SB_LUT4 add_3431_8_lut (.I0(GND_net), .I1(n16185[5]), .I2(n734), .I3(n35671), 
            .O(n16031[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3431_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3067_2 (.CI(GND_net), .I0(n41), .I1(n134), .CO(n35478));
    SB_LUT4 add_3064_18_lut (.I0(GND_net), .I1(n8208[15]), .I2(GND_net), 
            .I3(n35433), .O(n8184[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3064_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3248_13_lut (.I0(GND_net), .I1(n13109[10]), .I2(GND_net), 
            .I3(n34431), .O(n12575[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3248_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3248_13 (.CI(n34431), .I0(n13109[10]), .I1(GND_net), 
            .CO(n34432));
    SB_LUT4 add_3315_14_lut (.I0(GND_net), .I1(n14434[11]), .I2(GND_net), 
            .I3(n34353), .O(n14035[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3315_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3057_6 (.CI(n35246), .I0(n8019[3]), .I1(n492), .CO(n35247));
    SB_CARRY sub_11_add_2_6 (.CI(n34194), .I0(\PID_CONTROLLER.err_prev[4] ), 
            .I1(n64[4]), .CO(n34195));
    SB_CARRY add_3431_8 (.CI(n35671), .I0(n16185[5]), .I1(n734), .CO(n35672));
    SB_LUT4 add_3057_5_lut (.I0(GND_net), .I1(n8019[2]), .I2(n395), .I3(n35245), 
            .O(n7988[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3057_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3061_22 (.CI(n35368), .I0(n8133[19]), .I1(GND_net), .CO(n35369));
    SB_CARRY add_3064_18 (.CI(n35433), .I0(n8208[15]), .I1(GND_net), .CO(n35434));
    SB_CARRY add_3315_14 (.CI(n34353), .I0(n14434[11]), .I1(GND_net), 
            .CO(n34354));
    SB_CARRY add_3057_5 (.CI(n35245), .I0(n8019[2]), .I1(n395), .CO(n35246));
    SB_LUT4 add_3248_12_lut (.I0(GND_net), .I1(n13109[9]), .I2(GND_net), 
            .I3(n34430), .O(n12575[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3248_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3431_7_lut (.I0(GND_net), .I1(n16185[4]), .I2(n637), .I3(n35670), 
            .O(n16031[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3431_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3057_4_lut (.I0(GND_net), .I1(n8019[1]), .I2(n298), .I3(n35244), 
            .O(n7988[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3057_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3431_7 (.CI(n35670), .I0(n16185[4]), .I1(n637), .CO(n35671));
    SB_LUT4 add_3431_6_lut (.I0(GND_net), .I1(n16185[3]), .I2(n540), .I3(n35669), 
            .O(n16031[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3431_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_i98_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral [9]), 
            .I2(GND_net), .I3(GND_net), .O(n145));   // verilog/motorControl.v(43[48:59])
    defparam mult_14_i98_2_lut.LUT_INIT = 16'h4444;
    SB_CARRY add_3431_6 (.CI(n35669), .I0(n16185[3]), .I1(n540), .CO(n35670));
    SB_LUT4 add_3431_5_lut (.I0(GND_net), .I1(n16185[2]), .I2(n443), .I3(n35668), 
            .O(n16031[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3431_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_i147_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral [9]), 
            .I2(GND_net), .I3(GND_net), .O(n218));   // verilog/motorControl.v(43[48:59])
    defparam mult_14_i147_2_lut.LUT_INIT = 16'h4444;
    SB_CARRY add_3056_9 (.CI(n35037), .I0(n7988[6]), .I1(GND_net), .CO(n35038));
    SB_CARRY add_3248_12 (.CI(n34430), .I0(n13109[9]), .I1(GND_net), .CO(n34431));
    SB_LUT4 add_3248_11_lut (.I0(GND_net), .I1(n13109[8]), .I2(GND_net), 
            .I3(n34429), .O(n12575[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3248_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3431_5 (.CI(n35668), .I0(n16185[2]), .I1(n443), .CO(n35669));
    SB_LUT4 add_3431_4_lut (.I0(GND_net), .I1(n16185[1]), .I2(n346), .I3(n35667), 
            .O(n16031[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3431_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_11_add_2_5_lut (.I0(GND_net), .I1(\PID_CONTROLLER.err_prev[3] ), 
            .I2(n64[3]), .I3(n34193), .O(n57[3])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_11_add_2_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3431_4 (.CI(n35667), .I0(n16185[1]), .I1(n346), .CO(n35668));
    SB_LUT4 add_3056_8_lut (.I0(GND_net), .I1(n7988[5]), .I2(n683), .I3(n35036), 
            .O(n7956[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3056_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3069_10_lut (.I0(GND_net), .I1(n8313[7]), .I2(GND_net), 
            .I3(n35520), .O(n8294[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3069_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3056_8 (.CI(n35036), .I0(n7988[5]), .I1(n683), .CO(n35037));
    SB_LUT4 add_3315_13_lut (.I0(GND_net), .I1(n14434[10]), .I2(GND_net), 
            .I3(n34352), .O(n14035[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3315_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3431_3_lut (.I0(GND_net), .I1(n16185[0]), .I2(n249), .I3(n35666), 
            .O(n16031[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3431_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3073_9_lut (.I0(GND_net), .I1(n8379[6]), .I2(GND_net), 
            .I3(n35577), .O(n8364[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3073_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3431_3 (.CI(n35666), .I0(n16185[0]), .I1(n249), .CO(n35667));
    SB_CARRY add_3248_11 (.CI(n34429), .I0(n13109[8]), .I1(GND_net), .CO(n34430));
    SB_LUT4 add_3056_7_lut (.I0(GND_net), .I1(n7988[4]), .I2(n586), .I3(n35035), 
            .O(n7956[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3056_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3431_2_lut (.I0(GND_net), .I1(n59), .I2(n152_adj_3435), 
            .I3(GND_net), .O(n16031[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3431_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3061_21_lut (.I0(GND_net), .I1(n8133[18]), .I2(GND_net), 
            .I3(n35367), .O(n8106[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3061_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3061_21 (.CI(n35367), .I0(n8133[18]), .I1(GND_net), .CO(n35368));
    SB_CARRY add_3057_4 (.CI(n35244), .I0(n8019[1]), .I1(n298), .CO(n35245));
    SB_LUT4 add_3248_10_lut (.I0(GND_net), .I1(n13109[7]), .I2(GND_net), 
            .I3(n34428), .O(n12575[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3248_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3057_3_lut (.I0(GND_net), .I1(n8019[0]), .I2(n201), .I3(n35243), 
            .O(n7988[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3057_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3248_10 (.CI(n34428), .I0(n13109[7]), .I1(GND_net), .CO(n34429));
    SB_CARRY add_3056_7 (.CI(n35035), .I0(n7988[4]), .I1(n586), .CO(n35036));
    SB_LUT4 add_3061_20_lut (.I0(GND_net), .I1(n8133[17]), .I2(GND_net), 
            .I3(n35366), .O(n8106[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3061_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3056_6_lut (.I0(GND_net), .I1(n7988[3]), .I2(n489), .I3(n35034), 
            .O(n7956[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3056_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3057_3 (.CI(n35243), .I0(n8019[0]), .I1(n201), .CO(n35244));
    SB_CARRY add_3431_2 (.CI(GND_net), .I0(n59), .I1(n152_adj_3435), .CO(n35666));
    SB_CARRY add_3069_10 (.CI(n35520), .I0(n8313[7]), .I1(GND_net), .CO(n35521));
    SB_CARRY add_3061_20 (.CI(n35366), .I0(n8133[17]), .I1(GND_net), .CO(n35367));
    SB_CARRY add_3056_6 (.CI(n35034), .I0(n7988[3]), .I1(n489), .CO(n35035));
    SB_LUT4 add_2982_31_lut (.I0(GND_net), .I1(n7760[28]), .I2(GND_net), 
            .I3(n34693), .O(n6542[29])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2982_31_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2982_30_lut (.I0(GND_net), .I1(n7760[27]), .I2(GND_net), 
            .I3(n34692), .O(n6542[28])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2982_30_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3061_19_lut (.I0(GND_net), .I1(n8133[16]), .I2(GND_net), 
            .I3(n35365), .O(n8106[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3061_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2982_30 (.CI(n34692), .I0(n7760[27]), .I1(GND_net), .CO(n34693));
    SB_LUT4 add_3056_5_lut (.I0(GND_net), .I1(n7988[2]), .I2(n392), .I3(n35033), 
            .O(n7956[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3056_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i335_2_lut (.I0(\Kp[5] ), .I1(\PID_CONTROLLER.err[4] ), 
            .I2(GND_net), .I3(GND_net), .O(n498));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i335_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_3073_9 (.CI(n35577), .I0(n8379[6]), .I1(GND_net), .CO(n35578));
    SB_LUT4 add_3073_8_lut (.I0(GND_net), .I1(n8379[5]), .I2(n734_adj_3436), 
            .I3(n35576), .O(n8364[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3073_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3069_9_lut (.I0(GND_net), .I1(n8313[6]), .I2(GND_net), 
            .I3(n35519), .O(n8294[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3069_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3064_17_lut (.I0(GND_net), .I1(n8208[14]), .I2(GND_net), 
            .I3(n35432), .O(n8184[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3064_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3315_13 (.CI(n34352), .I0(n14434[10]), .I1(GND_net), 
            .CO(n34353));
    SB_CARRY add_3073_8 (.CI(n35576), .I0(n8379[5]), .I1(n734_adj_3436), 
            .CO(n35577));
    SB_CARRY add_3061_19 (.CI(n35365), .I0(n8133[16]), .I1(GND_net), .CO(n35366));
    SB_LUT4 add_3073_7_lut (.I0(GND_net), .I1(n8379[4]), .I2(n637_adj_3437), 
            .I3(n35575), .O(n8364[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3073_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3443_13_lut (.I0(GND_net), .I1(n16314[10]), .I2(GND_net), 
            .I3(n35665), .O(n16185[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3443_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3073_7 (.CI(n35575), .I0(n8379[4]), .I1(n637_adj_3437), 
            .CO(n35576));
    SB_LUT4 add_3248_9_lut (.I0(GND_net), .I1(n13109[6]), .I2(GND_net), 
            .I3(n34427), .O(n12575[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3248_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3061_18_lut (.I0(GND_net), .I1(n8133[15]), .I2(GND_net), 
            .I3(n35364), .O(n8106[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3061_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2982_29_lut (.I0(GND_net), .I1(n7760[26]), .I2(GND_net), 
            .I3(n34691), .O(n6542[27])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2982_29_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3069_9 (.CI(n35519), .I0(n8313[6]), .I1(GND_net), .CO(n35520));
    SB_LUT4 mult_14_i196_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral [9]), 
            .I2(GND_net), .I3(GND_net), .O(n291));   // verilog/motorControl.v(43[48:59])
    defparam mult_14_i196_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 mult_10_i400_2_lut (.I0(\Kp[6] ), .I1(\PID_CONTROLLER.err[4] ), 
            .I2(GND_net), .I3(GND_net), .O(n595));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i400_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_3066_21_lut (.I0(GND_net), .I1(n8253[18]), .I2(GND_net), 
            .I3(n35477), .O(n8231[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3066_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3057_2_lut (.I0(GND_net), .I1(n11_adj_3438), .I2(n104), 
            .I3(GND_net), .O(n7988[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3057_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3443_12_lut (.I0(GND_net), .I1(n16314[9]), .I2(GND_net), 
            .I3(n35664), .O(n16185[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3443_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3064_17 (.CI(n35432), .I0(n8208[14]), .I1(GND_net), .CO(n35433));
    SB_CARRY add_3061_18 (.CI(n35364), .I0(n8133[15]), .I1(GND_net), .CO(n35365));
    SB_LUT4 add_3069_8_lut (.I0(GND_net), .I1(n8313[5]), .I2(n722), .I3(n35518), 
            .O(n8294[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3069_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3061_17_lut (.I0(GND_net), .I1(n8133[14]), .I2(GND_net), 
            .I3(n35363), .O(n8106[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3061_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3064_16_lut (.I0(GND_net), .I1(n8208[13]), .I2(GND_net), 
            .I3(n35431), .O(n8184[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3064_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3248_9 (.CI(n34427), .I0(n13109[6]), .I1(GND_net), .CO(n34428));
    SB_CARRY add_2982_29 (.CI(n34691), .I0(n7760[26]), .I1(GND_net), .CO(n34692));
    SB_CARRY add_3061_17 (.CI(n35363), .I0(n8133[14]), .I1(GND_net), .CO(n35364));
    SB_CARRY add_3057_2 (.CI(GND_net), .I0(n11_adj_3438), .I1(n104), .CO(n35243));
    SB_LUT4 add_3248_8_lut (.I0(GND_net), .I1(n13109[5]), .I2(n704), .I3(n34426), 
            .O(n12575[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3248_8_lut.LUT_INIT = 16'hC33C;
    SB_DFF Kd_delay_counter_1015__i0 (.Q(Kd_delay_counter[0]), .C(clk32MHz), 
           .D(n69[0]));   // verilog/motorControl.v(55[27:47])
    SB_CARRY add_3248_8 (.CI(n34426), .I0(n13109[5]), .I1(n704), .CO(n34427));
    SB_LUT4 add_2982_28_lut (.I0(GND_net), .I1(n7760[25]), .I2(GND_net), 
            .I3(n34690), .O(n6542[26])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2982_28_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2982_28 (.CI(n34690), .I0(n7760[25]), .I1(GND_net), .CO(n34691));
    SB_LUT4 mult_12_add_2137_32_lut (.I0(n57[25]), .I1(n7956[29]), .I2(GND_net), 
            .I3(n35242), .O(n7061[0])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_12_add_2137_32_lut.LUT_INIT = 16'h6996;
    SB_CARRY add_3443_12 (.CI(n35664), .I0(n16314[9]), .I1(GND_net), .CO(n35665));
    SB_LUT4 add_3061_16_lut (.I0(GND_net), .I1(n8133[13]), .I2(GND_net), 
            .I3(n35362), .O(n8106[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3061_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3069_8 (.CI(n35518), .I0(n8313[5]), .I1(n722), .CO(n35519));
    SB_CARRY add_3061_16 (.CI(n35362), .I0(n8133[13]), .I1(GND_net), .CO(n35363));
    SB_CARRY add_3056_5 (.CI(n35033), .I0(n7988[2]), .I1(n392), .CO(n35034));
    SB_LUT4 add_3056_4_lut (.I0(GND_net), .I1(n7988[1]), .I2(n295), .I3(n35032), 
            .O(n7956[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3056_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3056_4 (.CI(n35032), .I0(n7988[1]), .I1(n295), .CO(n35033));
    SB_LUT4 add_3443_11_lut (.I0(GND_net), .I1(n16314[8]), .I2(GND_net), 
            .I3(n35663), .O(n16185[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3443_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3073_6_lut (.I0(GND_net), .I1(n8379[3]), .I2(n540_adj_3439), 
            .I3(n35574), .O(n8364[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3073_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3073_6 (.CI(n35574), .I0(n8379[3]), .I1(n540_adj_3439), 
            .CO(n35575));
    SB_LUT4 add_3069_7_lut (.I0(GND_net), .I1(n8313[4]), .I2(n625), .I3(n35517), 
            .O(n8294[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3069_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3443_11 (.CI(n35663), .I0(n16314[8]), .I1(GND_net), .CO(n35664));
    SB_LUT4 mult_12_add_2137_31_lut (.I0(GND_net), .I1(n7956[28]), .I2(GND_net), 
            .I3(n35241), .O(n191[30])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_12_add_2137_31_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3069_7 (.CI(n35517), .I0(n8313[4]), .I1(n625), .CO(n35518));
    SB_LUT4 add_3066_20_lut (.I0(GND_net), .I1(n8253[17]), .I2(GND_net), 
            .I3(n35476), .O(n8231[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3066_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3066_20 (.CI(n35476), .I0(n8253[17]), .I1(GND_net), .CO(n35477));
    SB_CARRY mult_12_add_2137_31 (.CI(n35241), .I0(n7956[28]), .I1(GND_net), 
            .CO(n35242));
    SB_LUT4 add_3066_19_lut (.I0(GND_net), .I1(n8253[16]), .I2(GND_net), 
            .I3(n35475), .O(n8231[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3066_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3056_3_lut (.I0(GND_net), .I1(n7988[0]), .I2(n198), .I3(n35031), 
            .O(n7956[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3056_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_12_add_2137_30_lut (.I0(GND_net), .I1(n7956[27]), .I2(GND_net), 
            .I3(n35240), .O(n191[29])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_12_add_2137_30_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_12_add_2137_30 (.CI(n35240), .I0(n7956[27]), .I1(GND_net), 
            .CO(n35241));
    SB_CARRY add_3064_16 (.CI(n35431), .I0(n8208[13]), .I1(GND_net), .CO(n35432));
    SB_LUT4 add_3443_10_lut (.I0(GND_net), .I1(n16314[7]), .I2(GND_net), 
            .I3(n35662), .O(n16185[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3443_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3248_7_lut (.I0(GND_net), .I1(n13109[4]), .I2(n607), .I3(n34425), 
            .O(n12575[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3248_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3248_7 (.CI(n34425), .I0(n13109[4]), .I1(n607), .CO(n34426));
    SB_CARRY add_3443_10 (.CI(n35662), .I0(n16314[7]), .I1(GND_net), .CO(n35663));
    SB_LUT4 add_2982_27_lut (.I0(GND_net), .I1(n7760[24]), .I2(GND_net), 
            .I3(n34689), .O(n6542[25])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2982_27_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_4_lut_4_lut (.I0(pwm[23]), .I1(hall1), .I2(hall2), .I3(GATES_5__N_3048[5]), 
            .O(n5_adj_3441));   // verilog/motorControl.v(86[38:44])
    defparam i1_4_lut_4_lut.LUT_INIT = 16'h55fd;
    SB_LUT4 add_3443_9_lut (.I0(GND_net), .I1(n16314[6]), .I2(GND_net), 
            .I3(n35661), .O(n16185[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3443_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i465_2_lut (.I0(\Kp[7] ), .I1(\PID_CONTROLLER.err[4] ), 
            .I2(GND_net), .I3(GND_net), .O(n692));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i465_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_14_i245_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral [9]), 
            .I2(GND_net), .I3(GND_net), .O(n364));   // verilog/motorControl.v(43[48:59])
    defparam mult_14_i245_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 add_3248_6_lut (.I0(GND_net), .I1(n13109[3]), .I2(n510_adj_3442), 
            .I3(n34424), .O(n12575[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3248_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3056_3 (.CI(n35031), .I0(n7988[0]), .I1(n198), .CO(n35032));
    SB_CARRY add_2982_27 (.CI(n34689), .I0(n7760[24]), .I1(GND_net), .CO(n34690));
    SB_CARRY add_3248_6 (.CI(n34424), .I0(n13109[3]), .I1(n510_adj_3442), 
            .CO(n34425));
    SB_LUT4 add_2982_26_lut (.I0(GND_net), .I1(n7760[23]), .I2(GND_net), 
            .I3(n34688), .O(n6542[24])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2982_26_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3069_6_lut (.I0(GND_net), .I1(n8313[3]), .I2(n528), .I3(n35516), 
            .O(n8294[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3069_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2982_26 (.CI(n34688), .I0(n7760[23]), .I1(GND_net), .CO(n34689));
    SB_CARRY add_3443_9 (.CI(n35661), .I0(n16314[6]), .I1(GND_net), .CO(n35662));
    SB_LUT4 add_3064_15_lut (.I0(GND_net), .I1(n8208[12]), .I2(GND_net), 
            .I3(n35430), .O(n8184[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3064_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3073_5_lut (.I0(GND_net), .I1(n8379[2]), .I2(n443_adj_3443), 
            .I3(n35573), .O(n8364[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3073_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3064_15 (.CI(n35430), .I0(n8208[12]), .I1(GND_net), .CO(n35431));
    SB_LUT4 add_3061_15_lut (.I0(GND_net), .I1(n8133[12]), .I2(GND_net), 
            .I3(n35361), .O(n8106[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3061_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3069_6 (.CI(n35516), .I0(n8313[3]), .I1(n528), .CO(n35517));
    SB_LUT4 add_2982_25_lut (.I0(GND_net), .I1(n7760[22]), .I2(GND_net), 
            .I3(n34687), .O(n6542[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2982_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3443_8_lut (.I0(GND_net), .I1(n16314[5]), .I2(n737), .I3(n35660), 
            .O(n16185[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3443_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3315_12_lut (.I0(GND_net), .I1(n14434[9]), .I2(GND_net), 
            .I3(n34351), .O(n14035[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3315_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3315_12 (.CI(n34351), .I0(n14434[9]), .I1(GND_net), .CO(n34352));
    SB_LUT4 mult_14_i294_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral [9]), 
            .I2(GND_net), .I3(GND_net), .O(n437));   // verilog/motorControl.v(43[48:59])
    defparam mult_14_i294_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 add_3248_5_lut (.I0(GND_net), .I1(n13109[2]), .I2(n413), .I3(n34423), 
            .O(n12575[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3248_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3073_5 (.CI(n35573), .I0(n8379[2]), .I1(n443_adj_3443), 
            .CO(n35574));
    SB_LUT4 mult_12_add_2137_29_lut (.I0(GND_net), .I1(n7956[26]), .I2(GND_net), 
            .I3(n35239), .O(n191[28])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_12_add_2137_29_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_12_add_2137_29 (.CI(n35239), .I0(n7956[26]), .I1(GND_net), 
            .CO(n35240));
    SB_LUT4 add_3056_2_lut (.I0(GND_net), .I1(n8), .I2(n101), .I3(GND_net), 
            .O(n7956[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3056_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3061_15 (.CI(n35361), .I0(n8133[12]), .I1(GND_net), .CO(n35362));
    SB_CARRY add_3443_8 (.CI(n35660), .I0(n16314[5]), .I1(n737), .CO(n35661));
    SB_CARRY add_3056_2 (.CI(GND_net), .I0(n8), .I1(n101), .CO(n35031));
    SB_CARRY add_3248_5 (.CI(n34423), .I0(n13109[2]), .I1(n413), .CO(n34424));
    SB_LUT4 add_3069_5_lut (.I0(GND_net), .I1(n8313[2]), .I2(n431), .I3(n35515), 
            .O(n8294[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3069_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3073_4_lut (.I0(GND_net), .I1(n8379[1]), .I2(n346_adj_3445), 
            .I3(n35572), .O(n8364[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3073_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_12_add_2137_28_lut (.I0(GND_net), .I1(n7956[25]), .I2(GND_net), 
            .I3(n35238), .O(n191[27])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_12_add_2137_28_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_11_add_2_5 (.CI(n34193), .I0(\PID_CONTROLLER.err_prev[3] ), 
            .I1(n64[3]), .CO(n34194));
    SB_CARRY add_2982_25 (.CI(n34687), .I0(n7760[22]), .I1(GND_net), .CO(n34688));
    SB_LUT4 add_3443_7_lut (.I0(GND_net), .I1(n16314[4]), .I2(n640), .I3(n35659), 
            .O(n16185[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3443_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3069_5 (.CI(n35515), .I0(n8313[2]), .I1(n431), .CO(n35516));
    SB_LUT4 add_3315_11_lut (.I0(GND_net), .I1(n14434[8]), .I2(GND_net), 
            .I3(n34350), .O(n14035[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3315_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3315_11 (.CI(n34350), .I0(n14434[8]), .I1(GND_net), .CO(n34351));
    SB_CARRY add_3443_7 (.CI(n35659), .I0(n16314[4]), .I1(n640), .CO(n35660));
    SB_LUT4 add_3443_6_lut (.I0(GND_net), .I1(n16314[3]), .I2(n543), .I3(n35658), 
            .O(n16185[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3443_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3073_4 (.CI(n35572), .I0(n8379[1]), .I1(n346_adj_3445), 
            .CO(n35573));
    SB_LUT4 add_3069_4_lut (.I0(GND_net), .I1(n8313[1]), .I2(n334), .I3(n35514), 
            .O(n8294[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3069_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_11_add_2_4_lut (.I0(GND_net), .I1(\PID_CONTROLLER.err_prev[2] ), 
            .I2(n64[2]), .I3(n34192), .O(n57[2])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_11_add_2_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3443_6 (.CI(n35658), .I0(n16314[3]), .I1(n543), .CO(n35659));
    SB_LUT4 add_3061_14_lut (.I0(GND_net), .I1(n8133[11]), .I2(GND_net), 
            .I3(n35360), .O(n8106[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3061_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3443_5_lut (.I0(GND_net), .I1(n16314[2]), .I2(n446_adj_3446), 
            .I3(n35657), .O(n16185[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3443_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3066_19 (.CI(n35475), .I0(n8253[16]), .I1(GND_net), .CO(n35476));
    SB_LUT4 mult_14_i343_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral [9]), 
            .I2(GND_net), .I3(GND_net), .O(n510));   // verilog/motorControl.v(43[48:59])
    defparam mult_14_i343_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 mult_14_i95_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral [9]), 
            .I2(GND_net), .I3(GND_net), .O(n107));   // verilog/motorControl.v(43[48:59])
    defparam mult_14_i95_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_3064_14_lut (.I0(GND_net), .I1(n8208[11]), .I2(GND_net), 
            .I3(n35429), .O(n8184[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3064_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3064_14 (.CI(n35429), .I0(n8208[11]), .I1(GND_net), .CO(n35430));
    SB_CARRY add_3061_14 (.CI(n35360), .I0(n8133[11]), .I1(GND_net), .CO(n35361));
    SB_LUT4 add_3061_13_lut (.I0(GND_net), .I1(n8133[10]), .I2(GND_net), 
            .I3(n35359), .O(n8106[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3061_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_i46_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral [9]), 
            .I2(GND_net), .I3(GND_net), .O(n35));   // verilog/motorControl.v(43[48:59])
    defparam mult_14_i46_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_14_i392_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral [9]), 
            .I2(GND_net), .I3(GND_net), .O(n583));   // verilog/motorControl.v(43[48:59])
    defparam mult_14_i392_2_lut.LUT_INIT = 16'h4444;
    SB_CARRY mult_12_add_2137_28 (.CI(n35238), .I0(n7956[25]), .I1(GND_net), 
            .CO(n35239));
    SB_LUT4 mult_12_add_2137_27_lut (.I0(GND_net), .I1(n7956[24]), .I2(GND_net), 
            .I3(n35237), .O(n191[26])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_12_add_2137_27_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3256_16_lut (.I0(GND_net), .I1(n13256[13]), .I2(GND_net), 
            .I3(n35030), .O(n12732[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3256_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_12_add_2137_27 (.CI(n35237), .I0(n7956[24]), .I1(GND_net), 
            .CO(n35238));
    SB_CARRY add_3443_5 (.CI(n35657), .I0(n16314[2]), .I1(n446_adj_3446), 
            .CO(n35658));
    SB_CARRY sub_11_add_2_4 (.CI(n34192), .I0(\PID_CONTROLLER.err_prev[2] ), 
            .I1(n64[2]), .CO(n34193));
    SB_LUT4 add_2982_24_lut (.I0(GND_net), .I1(n7760[21]), .I2(GND_net), 
            .I3(n34686), .O(n6542[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2982_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3248_4_lut (.I0(GND_net), .I1(n13109[1]), .I2(n316_adj_3447), 
            .I3(n34422), .O(n12575[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3248_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2982_24 (.CI(n34686), .I0(n7760[21]), .I1(GND_net), .CO(n34687));
    SB_CARRY add_3248_4 (.CI(n34422), .I0(n13109[1]), .I1(n316_adj_3447), 
            .CO(n34423));
    SB_LUT4 add_3248_3_lut (.I0(GND_net), .I1(n13109[0]), .I2(n219_adj_3448), 
            .I3(n34421), .O(n12575[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3248_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_12_add_2137_26_lut (.I0(GND_net), .I1(n7956[23]), .I2(GND_net), 
            .I3(n35236), .O(n191[25])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_12_add_2137_26_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3248_3 (.CI(n34421), .I0(n13109[0]), .I1(n219_adj_3448), 
            .CO(n34422));
    SB_LUT4 add_2982_23_lut (.I0(GND_net), .I1(n7760[20]), .I2(GND_net), 
            .I3(n34685), .O(n6542[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2982_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3256_15_lut (.I0(GND_net), .I1(n13256[12]), .I2(GND_net), 
            .I3(n35029), .O(n12732[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3256_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3248_2_lut (.I0(GND_net), .I1(n29_adj_3449), .I2(n122_adj_3450), 
            .I3(GND_net), .O(n12575[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3248_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2982_23 (.CI(n34685), .I0(n7760[20]), .I1(GND_net), .CO(n34686));
    SB_LUT4 add_2982_22_lut (.I0(GND_net), .I1(n7760[19]), .I2(GND_net), 
            .I3(n34684), .O(n6542[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2982_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3248_2 (.CI(GND_net), .I0(n29_adj_3449), .I1(n122_adj_3450), 
            .CO(n34421));
    SB_LUT4 add_3454_12_lut (.I0(GND_net), .I1(n16420[9]), .I2(GND_net), 
            .I3(n34420), .O(n16314[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3454_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3454_11_lut (.I0(GND_net), .I1(n16420[8]), .I2(GND_net), 
            .I3(n34419), .O(n16314[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3454_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_12_add_2137_26 (.CI(n35236), .I0(n7956[23]), .I1(GND_net), 
            .CO(n35237));
    SB_CARRY add_2982_22 (.CI(n34684), .I0(n7760[19]), .I1(GND_net), .CO(n34685));
    SB_CARRY add_3256_15 (.CI(n35029), .I0(n13256[12]), .I1(GND_net), 
            .CO(n35030));
    SB_CARRY add_3454_11 (.CI(n34419), .I0(n16420[8]), .I1(GND_net), .CO(n34420));
    SB_LUT4 add_2982_21_lut (.I0(GND_net), .I1(n7760[18]), .I2(GND_net), 
            .I3(n34683), .O(n6542[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2982_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3454_10_lut (.I0(GND_net), .I1(n16420[7]), .I2(GND_net), 
            .I3(n34418), .O(n16314[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3454_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_i144_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral [9]), 
            .I2(GND_net), .I3(GND_net), .O(n180));   // verilog/motorControl.v(43[48:59])
    defparam mult_14_i144_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_2982_21 (.CI(n34683), .I0(n7760[18]), .I1(GND_net), .CO(n34684));
    SB_LUT4 add_3066_18_lut (.I0(GND_net), .I1(n8253[15]), .I2(GND_net), 
            .I3(n35474), .O(n8231[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3066_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3454_10 (.CI(n34418), .I0(n16420[7]), .I1(GND_net), .CO(n34419));
    SB_LUT4 add_3064_13_lut (.I0(GND_net), .I1(n8208[10]), .I2(GND_net), 
            .I3(n35428), .O(n8184[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3064_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_12_i211_2_lut (.I0(\Kd[3] ), .I1(n57[7]), .I2(GND_net), 
            .I3(GND_net), .O(n313_adj_3426));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i211_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_3454_9_lut (.I0(GND_net), .I1(n16420[6]), .I2(GND_net), 
            .I3(n34417), .O(n16314[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3454_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3061_13 (.CI(n35359), .I0(n8133[10]), .I1(GND_net), .CO(n35360));
    SB_LUT4 add_3256_14_lut (.I0(GND_net), .I1(n13256[11]), .I2(GND_net), 
            .I3(n35028), .O(n12732[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3256_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2982_20_lut (.I0(GND_net), .I1(n7760[17]), .I2(GND_net), 
            .I3(n34682), .O(n6542[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2982_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3256_14 (.CI(n35028), .I0(n13256[11]), .I1(GND_net), 
            .CO(n35029));
    SB_CARRY add_2982_20 (.CI(n34682), .I0(n7760[17]), .I1(GND_net), .CO(n34683));
    SB_LUT4 add_2982_19_lut (.I0(GND_net), .I1(n7760[16]), .I2(GND_net), 
            .I3(n34681), .O(n6542[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2982_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3315_10_lut (.I0(GND_net), .I1(n14434[7]), .I2(GND_net), 
            .I3(n34349), .O(n14035[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3315_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_12_add_2137_25_lut (.I0(GND_net), .I1(n7956[22]), .I2(GND_net), 
            .I3(n35235), .O(n191[24])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_12_add_2137_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3454_9 (.CI(n34417), .I0(n16420[6]), .I1(GND_net), .CO(n34418));
    SB_LUT4 add_3256_13_lut (.I0(GND_net), .I1(n13256[10]), .I2(GND_net), 
            .I3(n35027), .O(n12732[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3256_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3454_8_lut (.I0(GND_net), .I1(n16420[5]), .I2(n740), .I3(n34416), 
            .O(n16314[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3454_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2982_19 (.CI(n34681), .I0(n7760[16]), .I1(GND_net), .CO(n34682));
    SB_LUT4 add_3061_12_lut (.I0(GND_net), .I1(n8133[9]), .I2(GND_net), 
            .I3(n35358), .O(n8106[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3061_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2982_18_lut (.I0(GND_net), .I1(n7760[15]), .I2(GND_net), 
            .I3(n34680), .O(n6542[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2982_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_12_add_2137_25 (.CI(n35235), .I0(n7956[22]), .I1(GND_net), 
            .CO(n35236));
    SB_CARRY add_3454_8 (.CI(n34416), .I0(n16420[5]), .I1(n740), .CO(n34417));
    SB_CARRY add_3256_13 (.CI(n35027), .I0(n13256[10]), .I1(GND_net), 
            .CO(n35028));
    SB_LUT4 mult_10_i81_2_lut (.I0(\Kp[1] ), .I1(\PID_CONTROLLER.err[7] ), 
            .I2(GND_net), .I3(GND_net), .O(n119));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i81_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_2982_18 (.CI(n34680), .I0(n7760[15]), .I1(GND_net), .CO(n34681));
    SB_LUT4 mult_10_i18_2_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err[8] ), 
            .I2(GND_net), .I3(GND_net), .O(n26_adj_3425));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i18_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_2982_17_lut (.I0(GND_net), .I1(n7760[14]), .I2(GND_net), 
            .I3(n34679), .O(n6542[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2982_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3256_12_lut (.I0(GND_net), .I1(n13256[9]), .I2(GND_net), 
            .I3(n35026), .O(n12732[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3256_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3454_7_lut (.I0(GND_net), .I1(n16420[4]), .I2(n643), .I3(n34415), 
            .O(n16314[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3454_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2982_17 (.CI(n34679), .I0(n7760[14]), .I1(GND_net), .CO(n34680));
    SB_CARRY add_3454_7 (.CI(n34415), .I0(n16420[4]), .I1(n643), .CO(n34416));
    SB_LUT4 add_2982_16_lut (.I0(GND_net), .I1(n7760[13]), .I2(GND_net), 
            .I3(n34678), .O(n6542[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2982_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3256_12 (.CI(n35026), .I0(n13256[9]), .I1(GND_net), .CO(n35027));
    SB_LUT4 add_3454_6_lut (.I0(GND_net), .I1(n16420[3]), .I2(n546), .I3(n34414), 
            .O(n16314[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3454_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2982_16 (.CI(n34678), .I0(n7760[13]), .I1(GND_net), .CO(n34679));
    SB_CARRY add_3454_6 (.CI(n34414), .I0(n16420[3]), .I1(n546), .CO(n34415));
    SB_LUT4 add_2982_15_lut (.I0(GND_net), .I1(n7760[12]), .I2(GND_net), 
            .I3(n34677), .O(n6542[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2982_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_12_add_2137_24_lut (.I0(GND_net), .I1(n7956[21]), .I2(GND_net), 
            .I3(n35234), .O(n191[23])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_12_add_2137_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_11_inv_0_i11_1_lut (.I0(\PID_CONTROLLER.err[10] ), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n64[10]));   // verilog/motorControl.v(43[31:45])
    defparam sub_11_inv_0_i11_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY mult_12_add_2137_24 (.CI(n35234), .I0(n7956[21]), .I1(GND_net), 
            .CO(n35235));
    SB_LUT4 add_3454_5_lut (.I0(GND_net), .I1(n16420[2]), .I2(n449), .I3(n34413), 
            .O(n16314[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3454_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_11_add_2_3_lut (.I0(GND_net), .I1(\PID_CONTROLLER.err_prev[1] ), 
            .I2(n64[1]), .I3(n34191), .O(n57[1])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_11_add_2_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3454_5 (.CI(n34413), .I0(n16420[2]), .I1(n449), .CO(n34414));
    SB_LUT4 mult_12_add_2137_23_lut (.I0(GND_net), .I1(n7956[20]), .I2(GND_net), 
            .I3(n35233), .O(n191[22])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_12_add_2137_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3256_11_lut (.I0(GND_net), .I1(n13256[8]), .I2(GND_net), 
            .I3(n35025), .O(n12732[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3256_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3256_11 (.CI(n35025), .I0(n13256[8]), .I1(GND_net), .CO(n35026));
    SB_CARRY add_2982_15 (.CI(n34677), .I0(n7760[12]), .I1(GND_net), .CO(n34678));
    SB_LUT4 add_2982_14_lut (.I0(GND_net), .I1(n7760[11]), .I2(GND_net), 
            .I3(n34676), .O(n6542[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2982_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2982_14 (.CI(n34676), .I0(n7760[11]), .I1(GND_net), .CO(n34677));
    SB_LUT4 add_2982_13_lut (.I0(GND_net), .I1(n7760[10]), .I2(GND_net), 
            .I3(n34675), .O(n6542[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2982_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3454_4_lut (.I0(GND_net), .I1(n16420[1]), .I2(n352), .I3(n34412), 
            .O(n16314[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3454_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3454_4 (.CI(n34412), .I0(n16420[1]), .I1(n352), .CO(n34413));
    SB_LUT4 add_3454_3_lut (.I0(GND_net), .I1(n16420[0]), .I2(n255), .I3(n34411), 
            .O(n16314[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3454_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3256_10_lut (.I0(GND_net), .I1(n13256[7]), .I2(GND_net), 
            .I3(n35024), .O(n12732[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3256_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_12_add_2137_23 (.CI(n35233), .I0(n7956[20]), .I1(GND_net), 
            .CO(n35234));
    SB_CARRY add_3315_10 (.CI(n34349), .I0(n14434[7]), .I1(GND_net), .CO(n34350));
    SB_LUT4 i29313_3_lut_3_lut (.I0(n70[10]), .I1(n421), .I2(\PID_CONTROLLER.result [17]), 
            .I3(GND_net), .O(n44153));   // verilog/motorControl.v(47[28:37])
    defparam i29313_3_lut_3_lut.LUT_INIT = 16'hb8b8;
    SB_CARRY add_2982_13 (.CI(n34675), .I0(n7760[10]), .I1(GND_net), .CO(n34676));
    SB_LUT4 add_2982_12_lut (.I0(GND_net), .I1(n7760[9]), .I2(GND_net), 
            .I3(n34674), .O(n6542[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2982_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3256_10 (.CI(n35024), .I0(n13256[7]), .I1(GND_net), .CO(n35025));
    SB_CARRY add_2982_12 (.CI(n34674), .I0(n7760[9]), .I1(GND_net), .CO(n34675));
    SB_CARRY add_3454_3 (.CI(n34411), .I0(n16420[0]), .I1(n255), .CO(n34412));
    SB_LUT4 add_3315_9_lut (.I0(GND_net), .I1(n14434[6]), .I2(GND_net), 
            .I3(n34348), .O(n14035[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3315_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3454_2_lut (.I0(GND_net), .I1(n65), .I2(n158), .I3(GND_net), 
            .O(n16314[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3454_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3315_9 (.CI(n34348), .I0(n14434[6]), .I1(GND_net), .CO(n34349));
    SB_CARRY add_3069_4 (.CI(n35514), .I0(n8313[1]), .I1(n334), .CO(n35515));
    SB_CARRY sub_11_add_2_3 (.CI(n34191), .I0(\PID_CONTROLLER.err_prev[1] ), 
            .I1(n64[1]), .CO(n34192));
    SB_CARRY add_3066_18 (.CI(n35474), .I0(n8253[15]), .I1(GND_net), .CO(n35475));
    SB_LUT4 mult_12_add_2137_22_lut (.I0(GND_net), .I1(n7956[19]), .I2(GND_net), 
            .I3(n35232), .O(n191[21])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_12_add_2137_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3256_9_lut (.I0(GND_net), .I1(n13256[6]), .I2(GND_net), 
            .I3(n35023), .O(n12732[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3256_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3064_13 (.CI(n35428), .I0(n8208[10]), .I1(GND_net), .CO(n35429));
    SB_CARRY add_3256_9 (.CI(n35023), .I0(n13256[6]), .I1(GND_net), .CO(n35024));
    SB_CARRY add_3061_12 (.CI(n35358), .I0(n8133[9]), .I1(GND_net), .CO(n35359));
    SB_LUT4 add_3256_8_lut (.I0(GND_net), .I1(n13256[5]), .I2(n545), .I3(n35022), 
            .O(n12732[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3256_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3061_11_lut (.I0(GND_net), .I1(n8133[8]), .I2(GND_net), 
            .I3(n35357), .O(n8106[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3061_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2982_11_lut (.I0(GND_net), .I1(n7760[8]), .I2(GND_net), 
            .I3(n34673), .O(n6542[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2982_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3066_17_lut (.I0(GND_net), .I1(n8253[14]), .I2(GND_net), 
            .I3(n35473), .O(n8231[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3066_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_12_add_2137_22 (.CI(n35232), .I0(n7956[19]), .I1(GND_net), 
            .CO(n35233));
    SB_LUT4 add_3443_4_lut (.I0(GND_net), .I1(n16314[1]), .I2(n349_adj_3453), 
            .I3(n35656), .O(n16185[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3443_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3315_8_lut (.I0(GND_net), .I1(n14434[5]), .I2(n713), .I3(n34347), 
            .O(n14035[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3315_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3064_12_lut (.I0(GND_net), .I1(n8208[9]), .I2(GND_net), 
            .I3(n35427), .O(n8184[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3064_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2982_11 (.CI(n34673), .I0(n7760[8]), .I1(GND_net), .CO(n34674));
    SB_LUT4 add_2982_10_lut (.I0(GND_net), .I1(n7760[7]), .I2(GND_net), 
            .I3(n34672), .O(n6542[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2982_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_11_add_2_2_lut (.I0(GND_net), .I1(\PID_CONTROLLER.err_prev[0] ), 
            .I2(n64[0]), .I3(VCC_net), .O(n57[0])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_11_add_2_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_12_add_2137_21_lut (.I0(GND_net), .I1(n7956[18]), .I2(GND_net), 
            .I3(n35231), .O(n191[20])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_12_add_2137_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3315_8 (.CI(n34347), .I0(n14434[5]), .I1(n713), .CO(n34348));
    SB_CARRY add_2982_10 (.CI(n34672), .I0(n7760[7]), .I1(GND_net), .CO(n34673));
    SB_CARRY sub_11_add_2_2 (.CI(VCC_net), .I0(\PID_CONTROLLER.err_prev[0] ), 
            .I1(n64[0]), .CO(n34191));
    SB_LUT4 add_2982_9_lut (.I0(GND_net), .I1(n7760[6]), .I2(GND_net), 
            .I3(n34671), .O(n6542[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2982_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3256_8 (.CI(n35022), .I0(n13256[5]), .I1(n545), .CO(n35023));
    SB_CARRY add_3061_11 (.CI(n35357), .I0(n8133[8]), .I1(GND_net), .CO(n35358));
    SB_CARRY add_2982_9 (.CI(n34671), .I0(n7760[6]), .I1(GND_net), .CO(n34672));
    SB_LUT4 add_3315_7_lut (.I0(GND_net), .I1(n14434[4]), .I2(n616), .I3(n34346), 
            .O(n14035[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3315_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_12_add_2137_21 (.CI(n35231), .I0(n7956[18]), .I1(GND_net), 
            .CO(n35232));
    SB_LUT4 add_2982_8_lut (.I0(GND_net), .I1(n7760[5]), .I2(n683_adj_3454), 
            .I3(n34670), .O(n6542[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2982_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2982_8 (.CI(n34670), .I0(n7760[5]), .I1(n683_adj_3454), 
            .CO(n34671));
    SB_CARRY add_3315_7 (.CI(n34346), .I0(n14434[4]), .I1(n616), .CO(n34347));
    SB_LUT4 add_2982_7_lut (.I0(GND_net), .I1(n7760[4]), .I2(n586_adj_3455), 
            .I3(n34669), .O(n6542[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2982_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_12_add_2137_20_lut (.I0(GND_net), .I1(n7956[17]), .I2(GND_net), 
            .I3(n35230), .O(n191[19])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_12_add_2137_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i23_4_lut_4_lut (.I0(hall3), .I1(hall1), .I2(n878), .I3(n17_adj_3456), 
            .O(GATES_5__N_2788[0]));   // verilog/motorControl.v(86[14] 109[8])
    defparam i23_4_lut_4_lut.LUT_INIT = 16'h2044;
    SB_CARRY add_2982_7 (.CI(n34669), .I0(n7760[4]), .I1(n586_adj_3455), 
            .CO(n34670));
    SB_LUT4 add_3061_10_lut (.I0(GND_net), .I1(n8133[7]), .I2(GND_net), 
            .I3(n35356), .O(n8106[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3061_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2982_6_lut (.I0(GND_net), .I1(n7760[3]), .I2(n489_adj_3457), 
            .I3(n34668), .O(n6542[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2982_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_12_add_2137_20 (.CI(n35230), .I0(n7956[17]), .I1(GND_net), 
            .CO(n35231));
    SB_CARRY add_3064_12 (.CI(n35427), .I0(n8208[9]), .I1(GND_net), .CO(n35428));
    SB_LUT4 add_3256_7_lut (.I0(GND_net), .I1(n13256[4]), .I2(n472), .I3(n35021), 
            .O(n12732[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3256_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3061_10 (.CI(n35356), .I0(n8133[7]), .I1(GND_net), .CO(n35357));
    SB_CARRY add_2982_6 (.CI(n34668), .I0(n7760[3]), .I1(n489_adj_3457), 
            .CO(n34669));
    SB_LUT4 mult_12_add_2137_19_lut (.I0(GND_net), .I1(n7956[16]), .I2(GND_net), 
            .I3(n35229), .O(n191[18])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_12_add_2137_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3315_6_lut (.I0(GND_net), .I1(n14434[3]), .I2(n519), .I3(n34345), 
            .O(n14035[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3315_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3256_7 (.CI(n35021), .I0(n13256[4]), .I1(n472), .CO(n35022));
    SB_LUT4 i29054_3_lut_3_lut (.I0(n70[10]), .I1(n421), .I2(\PID_CONTROLLER.result [18]), 
            .I3(GND_net), .O(n44151));   // verilog/motorControl.v(47[28:37])
    defparam i29054_3_lut_3_lut.LUT_INIT = 16'hb8b8;
    SB_CARRY add_3315_6 (.CI(n34345), .I0(n14434[3]), .I1(n519), .CO(n34346));
    SB_LUT4 add_2982_5_lut (.I0(GND_net), .I1(n7760[2]), .I2(n392_adj_3458), 
            .I3(n34667), .O(n6542[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2982_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3256_6_lut (.I0(GND_net), .I1(n13256[3]), .I2(n399), .I3(n35020), 
            .O(n12732[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3256_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_12_add_2137_19 (.CI(n35229), .I0(n7956[16]), .I1(GND_net), 
            .CO(n35230));
    SB_CARRY add_3443_4 (.CI(n35656), .I0(n16314[1]), .I1(n349_adj_3453), 
            .CO(n35657));
    SB_LUT4 add_3073_3_lut (.I0(GND_net), .I1(n8379[0]), .I2(n249_adj_3459), 
            .I3(n35571), .O(n8364[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3073_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3064_11_lut (.I0(GND_net), .I1(n8208[8]), .I2(GND_net), 
            .I3(n35426), .O(n8184[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3064_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3443_3_lut (.I0(GND_net), .I1(n16314[0]), .I2(n252_adj_3460), 
            .I3(n35655), .O(n16185[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3443_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i29015_3_lut_3_lut (.I0(n70[10]), .I1(n421), .I2(\PID_CONTROLLER.result [19]), 
            .I3(GND_net), .O(n44109));   // verilog/motorControl.v(47[28:37])
    defparam i29015_3_lut_3_lut.LUT_INIT = 16'hb8b8;
    SB_LUT4 add_3315_5_lut (.I0(GND_net), .I1(n14434[2]), .I2(n422), .I3(n34344), 
            .O(n14035[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3315_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2982_5 (.CI(n34667), .I0(n7760[2]), .I1(n392_adj_3458), 
            .CO(n34668));
    SB_CARRY add_3315_5 (.CI(n34344), .I0(n14434[2]), .I1(n422), .CO(n34345));
    SB_LUT4 add_3315_4_lut (.I0(GND_net), .I1(n14434[1]), .I2(n325), .I3(n34343), 
            .O(n14035[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3315_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3256_6 (.CI(n35020), .I0(n13256[3]), .I1(n399), .CO(n35021));
    SB_CARRY add_3315_4 (.CI(n34343), .I0(n14434[1]), .I1(n325), .CO(n34344));
    SB_LUT4 add_2982_4_lut (.I0(GND_net), .I1(n7760[1]), .I2(n295_adj_3461), 
            .I3(n34666), .O(n6542[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2982_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_12_add_2137_18_lut (.I0(GND_net), .I1(n7956[15]), .I2(GND_net), 
            .I3(n35228), .O(n191[17])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_12_add_2137_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3315_3_lut (.I0(GND_net), .I1(n14434[0]), .I2(n228_adj_3462), 
            .I3(n34342), .O(n14035[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3315_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3256_5_lut (.I0(GND_net), .I1(n13256[2]), .I2(n326), .I3(n35019), 
            .O(n12732[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3256_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i28834_3_lut_3_lut (.I0(n70[10]), .I1(n421), .I2(\PID_CONTROLLER.result [20]), 
            .I3(GND_net), .O(n44111));   // verilog/motorControl.v(47[28:37])
    defparam i28834_3_lut_3_lut.LUT_INIT = 16'hb8b8;
    SB_LUT4 add_3061_9_lut (.I0(GND_net), .I1(n8133[6]), .I2(GND_net), 
            .I3(n35355), .O(n8106[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3061_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3315_3 (.CI(n34342), .I0(n14434[0]), .I1(n228_adj_3462), 
            .CO(n34343));
    SB_CARRY mult_12_add_2137_18 (.CI(n35228), .I0(n7956[15]), .I1(GND_net), 
            .CO(n35229));
    SB_LUT4 add_3069_3_lut (.I0(GND_net), .I1(n8313[0]), .I2(n237), .I3(n35513), 
            .O(n8294[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3069_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3069_3 (.CI(n35513), .I0(n8313[0]), .I1(n237), .CO(n35514));
    SB_LUT4 add_3315_2_lut (.I0(GND_net), .I1(n38), .I2(n131_adj_3463), 
            .I3(GND_net), .O(n14035[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3315_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3073_3 (.CI(n35571), .I0(n8379[0]), .I1(n249_adj_3459), 
            .CO(n35572));
    SB_LUT4 mult_12_add_2137_17_lut (.I0(GND_net), .I1(n7956[14]), .I2(GND_net), 
            .I3(n35227), .O(n191[16])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_12_add_2137_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3256_5 (.CI(n35019), .I0(n13256[2]), .I1(n326), .CO(n35020));
    SB_LUT4 add_3256_4_lut (.I0(GND_net), .I1(n13256[1]), .I2(n253), .I3(n35018), 
            .O(n12732[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3256_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2982_4 (.CI(n34666), .I0(n7760[1]), .I1(n295_adj_3461), 
            .CO(n34667));
    SB_CARRY add_3256_4 (.CI(n35018), .I0(n13256[1]), .I1(n253), .CO(n35019));
    SB_CARRY add_3315_2 (.CI(GND_net), .I0(n38), .I1(n131_adj_3463), .CO(n34342));
    SB_LUT4 add_3073_2_lut (.I0(GND_net), .I1(n59_adj_3465), .I2(n152_adj_3466), 
            .I3(GND_net), .O(n8364[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3073_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3443_3 (.CI(n35655), .I0(n16314[0]), .I1(n252_adj_3460), 
            .CO(n35656));
    SB_LUT4 add_3335_20_lut (.I0(GND_net), .I1(n14793[17]), .I2(GND_net), 
            .I3(n34341), .O(n14434[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3335_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3335_19_lut (.I0(GND_net), .I1(n14793[16]), .I2(GND_net), 
            .I3(n34340), .O(n14434[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3335_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3073_2 (.CI(GND_net), .I0(n59_adj_3465), .I1(n152_adj_3466), 
            .CO(n35571));
    SB_CARRY add_3061_9 (.CI(n35355), .I0(n8133[6]), .I1(GND_net), .CO(n35356));
    SB_LUT4 add_3256_3_lut (.I0(GND_net), .I1(n13256[0]), .I2(n180), .I3(n35017), 
            .O(n12732[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3256_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3443_2_lut (.I0(GND_net), .I1(n62_adj_3467), .I2(n155_adj_3468), 
            .I3(GND_net), .O(n16185[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3443_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2982_3_lut (.I0(GND_net), .I1(n7760[0]), .I2(n198_adj_3469), 
            .I3(n34665), .O(n6542[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2982_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2982_3 (.CI(n34665), .I0(n7760[0]), .I1(n198_adj_3469), 
            .CO(n34666));
    SB_CARRY add_3335_19 (.CI(n34340), .I0(n14793[16]), .I1(GND_net), 
            .CO(n34341));
    SB_CARRY mult_12_add_2137_17 (.CI(n35227), .I0(n7956[14]), .I1(GND_net), 
            .CO(n35228));
    SB_LUT4 mult_12_add_2137_16_lut (.I0(GND_net), .I1(n7956[13]), .I2(GND_net), 
            .I3(n35226), .O(n191[15])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_12_add_2137_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3443_2 (.CI(GND_net), .I0(n62_adj_3467), .I1(n155_adj_3468), 
            .CO(n35655));
    SB_CARRY add_3454_2 (.CI(GND_net), .I0(n65), .I1(n158), .CO(n34411));
    SB_CARRY add_3064_11 (.CI(n35426), .I0(n8208[8]), .I1(GND_net), .CO(n35427));
    SB_LUT4 mult_10_i146_2_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err[7] ), 
            .I2(GND_net), .I3(GND_net), .O(n216));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i146_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_3335_18_lut (.I0(GND_net), .I1(n14793[15]), .I2(GND_net), 
            .I3(n34339), .O(n14434[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3335_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3272_23_lut (.I0(GND_net), .I1(n13594[20]), .I2(GND_net), 
            .I3(n34410), .O(n13109[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3272_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2982_2_lut (.I0(GND_net), .I1(n8_adj_3470), .I2(n101_adj_3471), 
            .I3(GND_net), .O(n6542[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2982_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3335_18 (.CI(n34339), .I0(n14793[15]), .I1(GND_net), 
            .CO(n34340));
    SB_CARRY add_3256_3 (.CI(n35017), .I0(n13256[0]), .I1(n180), .CO(n35018));
    SB_LUT4 i28836_3_lut_3_lut (.I0(n70[10]), .I1(n421), .I2(\PID_CONTROLLER.result [23]), 
            .I3(GND_net), .O(n44117));   // verilog/motorControl.v(47[28:37])
    defparam i28836_3_lut_3_lut.LUT_INIT = 16'hb8b8;
    SB_LUT4 add_3335_17_lut (.I0(GND_net), .I1(n14793[14]), .I2(GND_net), 
            .I3(n34338), .O(n14434[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3335_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3061_8_lut (.I0(GND_net), .I1(n8133[5]), .I2(n698_adj_3472), 
            .I3(n35354), .O(n8106[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3061_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_12_add_2137_16 (.CI(n35226), .I0(n7956[13]), .I1(GND_net), 
            .CO(n35227));
    SB_LUT4 add_3256_2_lut (.I0(GND_net), .I1(n35), .I2(n107), .I3(GND_net), 
            .O(n12732[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3256_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_12_add_2137_15_lut (.I0(GND_net), .I1(n7956[12]), .I2(GND_net), 
            .I3(n35225), .O(n191[14])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_12_add_2137_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2982_2 (.CI(GND_net), .I0(n8_adj_3470), .I1(n101_adj_3471), 
            .CO(n34665));
    SB_CARRY add_3335_17 (.CI(n34338), .I0(n14793[14]), .I1(GND_net), 
            .CO(n34339));
    SB_LUT4 add_3335_16_lut (.I0(GND_net), .I1(n14793[13]), .I2(GND_net), 
            .I3(n34337), .O(n14434[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3335_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3335_16 (.CI(n34337), .I0(n14793[13]), .I1(GND_net), 
            .CO(n34338));
    SB_CARRY add_3066_17 (.CI(n35473), .I0(n8253[14]), .I1(GND_net), .CO(n35474));
    SB_CARRY add_3256_2 (.CI(GND_net), .I0(n35), .I1(n107), .CO(n35017));
    SB_LUT4 add_3066_16_lut (.I0(GND_net), .I1(n8253[13]), .I2(GND_net), 
            .I3(n35472), .O(n8231[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3066_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3066_16 (.CI(n35472), .I0(n8253[13]), .I1(GND_net), .CO(n35473));
    SB_LUT4 add_3072_15_lut (.I0(GND_net), .I1(n8364[12]), .I2(GND_net), 
            .I3(n35570), .O(n8348[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3072_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3069_2_lut (.I0(GND_net), .I1(n47_adj_3473), .I2(n140_adj_3474), 
            .I3(GND_net), .O(n8294[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3069_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3066_15_lut (.I0(GND_net), .I1(n8253[12]), .I2(GND_net), 
            .I3(n35471), .O(n8231[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3066_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3066_15 (.CI(n35471), .I0(n8253[12]), .I1(GND_net), .CO(n35472));
    SB_LUT4 add_3049_30_lut (.I0(GND_net), .I1(n9125[27]), .I2(GND_net), 
            .I3(n34664), .O(n7760[28])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3049_30_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3335_15_lut (.I0(GND_net), .I1(n14793[12]), .I2(GND_net), 
            .I3(n34336), .O(n14434[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3335_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3049_29_lut (.I0(GND_net), .I1(n9125[26]), .I2(GND_net), 
            .I3(n34663), .O(n7760[27])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3049_29_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3335_15 (.CI(n34336), .I0(n14793[12]), .I1(GND_net), 
            .CO(n34337));
    SB_LUT4 add_3335_14_lut (.I0(GND_net), .I1(n14793[11]), .I2(GND_net), 
            .I3(n34335), .O(n14434[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3335_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3066_14_lut (.I0(GND_net), .I1(n8253[11]), .I2(GND_net), 
            .I3(n35470), .O(n8231[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3066_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3066_14 (.CI(n35470), .I0(n8253[11]), .I1(GND_net), .CO(n35471));
    SB_CARRY add_3049_29 (.CI(n34663), .I0(n9125[26]), .I1(GND_net), .CO(n34664));
    SB_CARRY add_3069_2 (.CI(GND_net), .I0(n47_adj_3473), .I1(n140_adj_3474), 
            .CO(n35513));
    SB_CARRY add_3335_14 (.CI(n34335), .I0(n14793[11]), .I1(GND_net), 
            .CO(n34336));
    SB_LUT4 add_3072_14_lut (.I0(GND_net), .I1(n8364[11]), .I2(GND_net), 
            .I3(n35569), .O(n8348[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3072_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3072_14 (.CI(n35569), .I0(n8364[11]), .I1(GND_net), .CO(n35570));
    SB_LUT4 add_3335_13_lut (.I0(GND_net), .I1(n14793[10]), .I2(GND_net), 
            .I3(n34334), .O(n14434[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3335_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3080_23_lut (.I0(GND_net), .I1(n8472[20]), .I2(GND_net), 
            .I3(n35654), .O(n8448[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3080_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3066_13_lut (.I0(GND_net), .I1(n8253[10]), .I2(GND_net), 
            .I3(n35469), .O(n8231[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3066_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3072_13_lut (.I0(GND_net), .I1(n8364[10]), .I2(GND_net), 
            .I3(n35568), .O(n8348[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3072_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3066_13 (.CI(n35469), .I0(n8253[10]), .I1(GND_net), .CO(n35470));
    SB_CARRY add_3072_13 (.CI(n35568), .I0(n8364[10]), .I1(GND_net), .CO(n35569));
    SB_LUT4 add_3068_19_lut (.I0(GND_net), .I1(n8294[16]), .I2(GND_net), 
            .I3(n35512), .O(n8274[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3068_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3068_18_lut (.I0(GND_net), .I1(n8294[15]), .I2(GND_net), 
            .I3(n35511), .O(n8274[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3068_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3072_12_lut (.I0(GND_net), .I1(n8364[9]), .I2(GND_net), 
            .I3(n35567), .O(n8348[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3072_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3068_18 (.CI(n35511), .I0(n8294[15]), .I1(GND_net), .CO(n35512));
    SB_LUT4 add_3080_22_lut (.I0(GND_net), .I1(n8472[19]), .I2(GND_net), 
            .I3(n35653), .O(n8448[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3080_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3066_12_lut (.I0(GND_net), .I1(n8253[9]), .I2(GND_net), 
            .I3(n35468), .O(n8231[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3066_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3068_17_lut (.I0(GND_net), .I1(n8294[14]), .I2(GND_net), 
            .I3(n35510), .O(n8274[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3068_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 Kd_delay_counter_1015_add_4_8_lut (.I0(GND_net), .I1(GND_net), 
            .I2(Kd_delay_counter[6]), .I3(n35016), .O(n69[6])) /* synthesis syn_instantiated=1 */ ;
    defparam Kd_delay_counter_1015_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3066_12 (.CI(n35468), .I0(n8253[9]), .I1(GND_net), .CO(n35469));
    SB_CARRY add_3072_12 (.CI(n35567), .I0(n8364[9]), .I1(GND_net), .CO(n35568));
    SB_CARRY add_3335_13 (.CI(n34334), .I0(n14793[10]), .I1(GND_net), 
            .CO(n34335));
    SB_LUT4 Kd_delay_counter_1015_add_4_7_lut (.I0(GND_net), .I1(GND_net), 
            .I2(Kd_delay_counter[5]), .I3(n35015), .O(n69[5])) /* synthesis syn_instantiated=1 */ ;
    defparam Kd_delay_counter_1015_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3080_22 (.CI(n35653), .I0(n8472[19]), .I1(GND_net), .CO(n35654));
    SB_LUT4 add_3080_21_lut (.I0(GND_net), .I1(n8472[18]), .I2(GND_net), 
            .I3(n35652), .O(n8448[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3080_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3066_11_lut (.I0(GND_net), .I1(n8253[8]), .I2(GND_net), 
            .I3(n35467), .O(n8231[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3066_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_12_add_2137_15 (.CI(n35225), .I0(n7956[12]), .I1(GND_net), 
            .CO(n35226));
    SB_CARRY add_3080_21 (.CI(n35652), .I0(n8472[18]), .I1(GND_net), .CO(n35653));
    SB_LUT4 i28842_3_lut_3_lut (.I0(n70[10]), .I1(n421), .I2(\PID_CONTROLLER.result [21]), 
            .I3(GND_net), .O(n44113));   // verilog/motorControl.v(47[28:37])
    defparam i28842_3_lut_3_lut.LUT_INIT = 16'hb8b8;
    SB_CARRY Kd_delay_counter_1015_add_4_7 (.CI(n35015), .I0(GND_net), .I1(Kd_delay_counter[5]), 
            .CO(n35016));
    SB_LUT4 add_3335_12_lut (.I0(GND_net), .I1(n14793[9]), .I2(GND_net), 
            .I3(n34333), .O(n14434[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3335_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3072_11_lut (.I0(GND_net), .I1(n8364[8]), .I2(GND_net), 
            .I3(n35566), .O(n8348[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3072_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3049_28_lut (.I0(GND_net), .I1(n9125[25]), .I2(GND_net), 
            .I3(n34662), .O(n7760[26])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3049_28_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3080_20_lut (.I0(GND_net), .I1(n8472[17]), .I2(GND_net), 
            .I3(n35651), .O(n8448[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3080_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3072_11 (.CI(n35566), .I0(n8364[8]), .I1(GND_net), .CO(n35567));
    SB_CARRY add_3080_20 (.CI(n35651), .I0(n8472[17]), .I1(GND_net), .CO(n35652));
    SB_LUT4 add_3072_10_lut (.I0(GND_net), .I1(n8364[7]), .I2(GND_net), 
            .I3(n35565), .O(n8348[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3072_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3080_19_lut (.I0(GND_net), .I1(n8472[16]), .I2(GND_net), 
            .I3(n35650), .O(n8448[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3080_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3072_10 (.CI(n35565), .I0(n8364[7]), .I1(GND_net), .CO(n35566));
    SB_CARRY add_3080_19 (.CI(n35650), .I0(n8472[16]), .I1(GND_net), .CO(n35651));
    SB_LUT4 add_3072_9_lut (.I0(GND_net), .I1(n8364[6]), .I2(GND_net), 
            .I3(n35564), .O(n8348[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3072_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3072_9 (.CI(n35564), .I0(n8364[6]), .I1(GND_net), .CO(n35565));
    SB_LUT4 add_3072_8_lut (.I0(GND_net), .I1(n8364[5]), .I2(n731), .I3(n35563), 
            .O(n8348[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3072_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3335_12 (.CI(n34333), .I0(n14793[9]), .I1(GND_net), .CO(n34334));
    SB_LUT4 add_3080_18_lut (.I0(GND_net), .I1(n8472[15]), .I2(GND_net), 
            .I3(n35649), .O(n8448[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3080_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3072_8 (.CI(n35563), .I0(n8364[5]), .I1(n731), .CO(n35564));
    SB_CARRY add_3068_17 (.CI(n35510), .I0(n8294[14]), .I1(GND_net), .CO(n35511));
    SB_LUT4 add_3335_11_lut (.I0(GND_net), .I1(n14793[8]), .I2(GND_net), 
            .I3(n34332), .O(n14434[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3335_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3335_11 (.CI(n34332), .I0(n14793[8]), .I1(GND_net), .CO(n34333));
    SB_CARRY add_3080_18 (.CI(n35649), .I0(n8472[15]), .I1(GND_net), .CO(n35650));
    SB_LUT4 i28831_3_lut_3_lut (.I0(n70[10]), .I1(n421), .I2(\PID_CONTROLLER.result [22]), 
            .I3(GND_net), .O(n44115));   // verilog/motorControl.v(47[28:37])
    defparam i28831_3_lut_3_lut.LUT_INIT = 16'hb8b8;
    SB_LUT4 Kd_delay_counter_1015_add_4_6_lut (.I0(GND_net), .I1(GND_net), 
            .I2(Kd_delay_counter[4]), .I3(n35014), .O(n69[4])) /* synthesis syn_instantiated=1 */ ;
    defparam Kd_delay_counter_1015_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3080_17_lut (.I0(GND_net), .I1(n8472[14]), .I2(GND_net), 
            .I3(n35648), .O(n8448[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3080_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3068_16_lut (.I0(GND_net), .I1(n8294[13]), .I2(GND_net), 
            .I3(n35509), .O(n8274[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3068_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3061_8 (.CI(n35354), .I0(n8133[5]), .I1(n698_adj_3472), 
            .CO(n35355));
    SB_CARRY add_3066_11 (.CI(n35467), .I0(n8253[8]), .I1(GND_net), .CO(n35468));
    SB_CARRY add_3080_17 (.CI(n35648), .I0(n8472[14]), .I1(GND_net), .CO(n35649));
    SB_LUT4 add_3080_16_lut (.I0(GND_net), .I1(n8472[13]), .I2(GND_net), 
            .I3(n35647), .O(n8448[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3080_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3080_16 (.CI(n35647), .I0(n8472[13]), .I1(GND_net), .CO(n35648));
    SB_LUT4 add_3080_15_lut (.I0(GND_net), .I1(n8472[12]), .I2(GND_net), 
            .I3(n35646), .O(n8448[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3080_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3064_10_lut (.I0(GND_net), .I1(n8208[7]), .I2(GND_net), 
            .I3(n35425), .O(n8184[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3064_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3080_15 (.CI(n35646), .I0(n8472[12]), .I1(GND_net), .CO(n35647));
    SB_LUT4 add_3080_14_lut (.I0(GND_net), .I1(n8472[11]), .I2(GND_net), 
            .I3(n35645), .O(n8448[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3080_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3080_14 (.CI(n35645), .I0(n8472[11]), .I1(GND_net), .CO(n35646));
    SB_CARRY add_3049_28 (.CI(n34662), .I0(n9125[25]), .I1(GND_net), .CO(n34663));
    SB_CARRY add_3068_16 (.CI(n35509), .I0(n8294[13]), .I1(GND_net), .CO(n35510));
    SB_CARRY add_3064_10 (.CI(n35425), .I0(n8208[7]), .I1(GND_net), .CO(n35426));
    SB_LUT4 add_3080_13_lut (.I0(GND_net), .I1(n8472[10]), .I2(GND_net), 
            .I3(n35644), .O(n8448[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3080_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3335_10_lut (.I0(GND_net), .I1(n14793[7]), .I2(GND_net), 
            .I3(n34331), .O(n14434[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3335_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3080_13 (.CI(n35644), .I0(n8472[10]), .I1(GND_net), .CO(n35645));
    SB_LUT4 add_3080_12_lut (.I0(GND_net), .I1(n8472[9]), .I2(GND_net), 
            .I3(n35643), .O(n8448[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3080_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_12_add_2137_14_lut (.I0(GND_net), .I1(n7956[11]), .I2(GND_net), 
            .I3(n35224), .O(n191[13])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_12_add_2137_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3080_12 (.CI(n35643), .I0(n8472[9]), .I1(GND_net), .CO(n35644));
    SB_LUT4 add_3049_27_lut (.I0(GND_net), .I1(n9125[24]), .I2(GND_net), 
            .I3(n34661), .O(n7760[25])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3049_27_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3049_27 (.CI(n34661), .I0(n9125[24]), .I1(GND_net), .CO(n34662));
    SB_LUT4 add_3080_11_lut (.I0(GND_net), .I1(n8472[8]), .I2(GND_net), 
            .I3(n35642), .O(n8448[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3080_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3335_10 (.CI(n34331), .I0(n14793[7]), .I1(GND_net), .CO(n34332));
    SB_CARRY Kd_delay_counter_1015_add_4_6 (.CI(n35014), .I0(GND_net), .I1(Kd_delay_counter[4]), 
            .CO(n35015));
    SB_CARRY add_3080_11 (.CI(n35642), .I0(n8472[8]), .I1(GND_net), .CO(n35643));
    SB_LUT4 add_3064_9_lut (.I0(GND_net), .I1(n8208[6]), .I2(GND_net), 
            .I3(n35424), .O(n8184[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3064_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3049_26_lut (.I0(GND_net), .I1(n9125[23]), .I2(GND_net), 
            .I3(n34660), .O(n7760[24])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3049_26_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3080_10_lut (.I0(GND_net), .I1(n8472[7]), .I2(GND_net), 
            .I3(n35641), .O(n8448[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3080_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3335_9_lut (.I0(GND_net), .I1(n14793[6]), .I2(GND_net), 
            .I3(n34330), .O(n14434[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3335_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3080_10 (.CI(n35641), .I0(n8472[7]), .I1(GND_net), .CO(n35642));
    SB_CARRY add_3335_9 (.CI(n34330), .I0(n14793[6]), .I1(GND_net), .CO(n34331));
    SB_LUT4 Kd_delay_counter_1015_add_4_5_lut (.I0(GND_net), .I1(GND_net), 
            .I2(Kd_delay_counter[3]), .I3(n35013), .O(n69[3])) /* synthesis syn_instantiated=1 */ ;
    defparam Kd_delay_counter_1015_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3061_7_lut (.I0(GND_net), .I1(n8133[4]), .I2(n601_adj_3476), 
            .I3(n35353), .O(n8106[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3061_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_12_add_2137_14 (.CI(n35224), .I0(n7956[11]), .I1(GND_net), 
            .CO(n35225));
    SB_LUT4 mult_12_add_2137_13_lut (.I0(GND_net), .I1(n7956[10]), .I2(GND_net), 
            .I3(n35223), .O(n191[12])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_12_add_2137_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Kd_delay_counter_1015_add_4_5 (.CI(n35013), .I0(GND_net), .I1(Kd_delay_counter[3]), 
            .CO(n35014));
    SB_LUT4 mult_12_i416_2_lut (.I0(\Kd[6] ), .I1(n57[12]), .I2(GND_net), 
            .I3(GND_net), .O(n619));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i416_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i211_2_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err[7] ), 
            .I2(GND_net), .I3(GND_net), .O(n313_adj_3423));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i211_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_3335_8_lut (.I0(GND_net), .I1(n14793[5]), .I2(n716_adj_3477), 
            .I3(n34329), .O(n14434[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3335_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i78_2_lut (.I0(hall1), .I1(hall2), .I2(GND_net), .I3(GND_net), 
            .O(GATES_5__N_3048[5]));   // verilog/motorControl.v(91[19:34])
    defparam i78_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i20070_2_lut_3_lut (.I0(\Kp[0] ), .I1(\Kp[1] ), .I2(\PID_CONTROLLER.err[31] ), 
            .I3(GND_net), .O(n16637[0]));   // verilog/motorControl.v(43[17:23])
    defparam i20070_2_lut_3_lut.LUT_INIT = 16'h6060;
    SB_CARRY add_3049_26 (.CI(n34660), .I0(n9125[23]), .I1(GND_net), .CO(n34661));
    SB_LUT4 add_3066_10_lut (.I0(GND_net), .I1(n8253[7]), .I2(GND_net), 
            .I3(n35466), .O(n8231[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3066_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3064_9 (.CI(n35424), .I0(n8208[6]), .I1(GND_net), .CO(n35425));
    SB_CARRY add_3061_7 (.CI(n35353), .I0(n8133[4]), .I1(n601_adj_3476), 
            .CO(n35354));
    SB_LUT4 i20270_2_lut_3_lut (.I0(\Kp[0] ), .I1(\Kp[1] ), .I2(\Kp[2] ), 
            .I3(GND_net), .O(n35990));   // verilog/motorControl.v(43[17:23])
    defparam i20270_2_lut_3_lut.LUT_INIT = 16'h9696;
    SB_CARRY mult_12_add_2137_13 (.CI(n35223), .I0(n7956[10]), .I1(GND_net), 
            .CO(n35224));
    SB_LUT4 Kd_delay_counter_1015_add_4_4_lut (.I0(GND_net), .I1(GND_net), 
            .I2(Kd_delay_counter[2]), .I3(n35012), .O(n69[2])) /* synthesis syn_instantiated=1 */ ;
    defparam Kd_delay_counter_1015_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Kd_delay_counter_1015_add_4_4 (.CI(n35012), .I0(GND_net), .I1(Kd_delay_counter[2]), 
            .CO(n35013));
    SB_CARRY add_3335_8 (.CI(n34329), .I0(n14793[5]), .I1(n716_adj_3477), 
            .CO(n34330));
    SB_LUT4 add_3049_25_lut (.I0(GND_net), .I1(n9125[22]), .I2(GND_net), 
            .I3(n34659), .O(n7760[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3049_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3080_9_lut (.I0(GND_net), .I1(n8472[6]), .I2(GND_net), 
            .I3(n35640), .O(n8448[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3080_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3080_9 (.CI(n35640), .I0(n8472[6]), .I1(GND_net), .CO(n35641));
    SB_CARRY add_3049_25 (.CI(n34659), .I0(n9125[22]), .I1(GND_net), .CO(n34660));
    SB_LUT4 add_3064_8_lut (.I0(GND_net), .I1(n8208[5]), .I2(n707), .I3(n35423), 
            .O(n8184[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3064_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3068_15_lut (.I0(GND_net), .I1(n8294[12]), .I2(GND_net), 
            .I3(n35508), .O(n8274[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3068_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3072_7_lut (.I0(GND_net), .I1(n8364[4]), .I2(n634), .I3(n35562), 
            .O(n8348[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3072_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3072_7 (.CI(n35562), .I0(n8364[4]), .I1(n634), .CO(n35563));
    SB_LUT4 add_3080_8_lut (.I0(GND_net), .I1(n8472[5]), .I2(n545), .I3(n35639), 
            .O(n8448[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3080_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3072_6_lut (.I0(GND_net), .I1(n8364[3]), .I2(n537), .I3(n35561), 
            .O(n8348[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3072_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3080_8 (.CI(n35639), .I0(n8472[5]), .I1(n545), .CO(n35640));
    SB_CARRY add_3072_6 (.CI(n35561), .I0(n8364[3]), .I1(n537), .CO(n35562));
    SB_LUT4 add_3072_5_lut (.I0(GND_net), .I1(n8364[2]), .I2(n440), .I3(n35560), 
            .O(n8348[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3072_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3080_7_lut (.I0(GND_net), .I1(n8472[4]), .I2(n472), .I3(n35638), 
            .O(n8448[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3080_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3080_7 (.CI(n35638), .I0(n8472[4]), .I1(n472), .CO(n35639));
    SB_LUT4 add_3080_6_lut (.I0(GND_net), .I1(n8472[3]), .I2(n399), .I3(n35637), 
            .O(n8448[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3080_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3072_5 (.CI(n35560), .I0(n8364[2]), .I1(n440), .CO(n35561));
    SB_LUT4 add_3072_4_lut (.I0(GND_net), .I1(n8364[1]), .I2(n343), .I3(n35559), 
            .O(n8348[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3072_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3072_4 (.CI(n35559), .I0(n8364[1]), .I1(n343), .CO(n35560));
    SB_CARRY add_3080_6 (.CI(n35637), .I0(n8472[3]), .I1(n399), .CO(n35638));
    SB_LUT4 add_3072_3_lut (.I0(GND_net), .I1(n8364[0]), .I2(n246), .I3(n35558), 
            .O(n8348[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3072_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3068_15 (.CI(n35508), .I0(n8294[12]), .I1(GND_net), .CO(n35509));
    SB_CARRY add_3072_3 (.CI(n35558), .I0(n8364[0]), .I1(n246), .CO(n35559));
    SB_LUT4 add_3080_5_lut (.I0(GND_net), .I1(n8472[2]), .I2(n326), .I3(n35636), 
            .O(n8448[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3080_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3080_5 (.CI(n35636), .I0(n8472[2]), .I1(n326), .CO(n35637));
    SB_LUT4 add_3080_4_lut (.I0(GND_net), .I1(n8472[1]), .I2(n253), .I3(n35635), 
            .O(n8448[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3080_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3049_24_lut (.I0(GND_net), .I1(n9125[21]), .I2(GND_net), 
            .I3(n34658), .O(n7760[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3049_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_12_add_2137_12_lut (.I0(GND_net), .I1(n7956[9]), .I2(GND_net), 
            .I3(n35222), .O(n191[11])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_12_add_2137_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3049_24 (.CI(n34658), .I0(n9125[21]), .I1(GND_net), .CO(n34659));
    SB_LUT4 add_3049_23_lut (.I0(GND_net), .I1(n9125[20]), .I2(GND_net), 
            .I3(n34657), .O(n7760[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3049_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3061_6_lut (.I0(GND_net), .I1(n8133[3]), .I2(n504_adj_3479), 
            .I3(n35352), .O(n8106[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3061_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_12_add_2137_12 (.CI(n35222), .I0(n7956[9]), .I1(GND_net), 
            .CO(n35223));
    SB_CARRY add_3049_23 (.CI(n34657), .I0(n9125[20]), .I1(GND_net), .CO(n34658));
    SB_LUT4 add_3049_22_lut (.I0(GND_net), .I1(n9125[19]), .I2(GND_net), 
            .I3(n34656), .O(n7760[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3049_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3335_7_lut (.I0(GND_net), .I1(n14793[4]), .I2(n619_adj_3480), 
            .I3(n34328), .O(n14434[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3335_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_12_add_2137_11_lut (.I0(GND_net), .I1(n7956[8]), .I2(GND_net), 
            .I3(n35221), .O(n191[10])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_12_add_2137_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3049_22 (.CI(n34656), .I0(n9125[19]), .I1(GND_net), .CO(n34657));
    SB_CARRY add_3080_4 (.CI(n35635), .I0(n8472[1]), .I1(n253), .CO(n35636));
    SB_LUT4 add_3049_21_lut (.I0(GND_net), .I1(n9125[18]), .I2(GND_net), 
            .I3(n34655), .O(n7760[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3049_21_lut.LUT_INIT = 16'hC33C;
    SB_DFF pwm_count_1016__i0 (.Q(pwm_count[0]), .C(clk32MHz), .D(n67[0]));   // verilog/motorControl.v(110[18:29])
    SB_CARRY add_3061_6 (.CI(n35352), .I0(n8133[3]), .I1(n504_adj_3479), 
            .CO(n35353));
    SB_CARRY add_3335_7 (.CI(n34328), .I0(n14793[4]), .I1(n619_adj_3480), 
            .CO(n34329));
    SB_LUT4 add_3272_22_lut (.I0(GND_net), .I1(n13594[19]), .I2(GND_net), 
            .I3(n34409), .O(n13109[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3272_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3064_8 (.CI(n35423), .I0(n8208[5]), .I1(n707), .CO(n35424));
    SB_LUT4 add_3080_3_lut (.I0(GND_net), .I1(n8472[0]), .I2(n180), .I3(n35634), 
            .O(n8448[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3080_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3061_5_lut (.I0(GND_net), .I1(n8133[2]), .I2(n407_adj_3482), 
            .I3(n35351), .O(n8106[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3061_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3080_3 (.CI(n35634), .I0(n8472[0]), .I1(n180), .CO(n35635));
    SB_LUT4 add_3080_2_lut (.I0(GND_net), .I1(n35), .I2(n107), .I3(GND_net), 
            .O(n8448[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3080_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3072_2_lut (.I0(GND_net), .I1(n56), .I2(n149_adj_3483), 
            .I3(GND_net), .O(n8348[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3072_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_12_add_2137_11 (.CI(n35221), .I0(n7956[8]), .I1(GND_net), 
            .CO(n35222));
    SB_CARRY add_3080_2 (.CI(GND_net), .I0(n35), .I1(n107), .CO(n35634));
    SB_CARRY add_3072_2 (.CI(GND_net), .I0(n56), .I1(n149_adj_3483), .CO(n35558));
    SB_LUT4 Kd_delay_counter_1015_add_4_3_lut (.I0(GND_net), .I1(GND_net), 
            .I2(Kd_delay_counter[1]), .I3(n35011), .O(n69[1])) /* synthesis syn_instantiated=1 */ ;
    defparam Kd_delay_counter_1015_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3272_22 (.CI(n34409), .I0(n13594[19]), .I1(GND_net), 
            .CO(n34410));
    SB_CARRY add_3049_21 (.CI(n34655), .I0(n9125[18]), .I1(GND_net), .CO(n34656));
    SB_LUT4 add_3071_16_lut (.I0(GND_net), .I1(n8348[13]), .I2(GND_net), 
            .I3(n35557), .O(n8331[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3071_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3335_6_lut (.I0(GND_net), .I1(n14793[3]), .I2(n522_adj_3484), 
            .I3(n34327), .O(n14434[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3335_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3272_21_lut (.I0(GND_net), .I1(n13594[18]), .I2(GND_net), 
            .I3(n34408), .O(n13109[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3272_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3079_8_lut (.I0(GND_net), .I1(n9319[5]), .I2(n752), .I3(n35633), 
            .O(n8439[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3079_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3335_6 (.CI(n34327), .I0(n14793[3]), .I1(n522_adj_3484), 
            .CO(n34328));
    SB_LUT4 add_3049_20_lut (.I0(GND_net), .I1(n9125[17]), .I2(GND_net), 
            .I3(n34654), .O(n7760[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3049_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Kd_delay_counter_1015_add_4_3 (.CI(n35011), .I0(GND_net), .I1(Kd_delay_counter[1]), 
            .CO(n35012));
    SB_CARRY add_3049_20 (.CI(n34654), .I0(n9125[17]), .I1(GND_net), .CO(n34655));
    SB_LUT4 add_3049_19_lut (.I0(GND_net), .I1(n9125[16]), .I2(GND_net), 
            .I3(n34653), .O(n7760[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3049_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3335_5_lut (.I0(GND_net), .I1(n14793[2]), .I2(n425_adj_3485), 
            .I3(n34326), .O(n14434[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3335_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3335_5 (.CI(n34326), .I0(n14793[2]), .I1(n425_adj_3485), 
            .CO(n34327));
    SB_LUT4 add_3071_15_lut (.I0(GND_net), .I1(n8348[12]), .I2(GND_net), 
            .I3(n35556), .O(n8331[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3071_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 Kd_delay_counter_1015_add_4_2_lut (.I0(GND_net), .I1(GND_net), 
            .I2(Kd_delay_counter[0]), .I3(VCC_net), .O(n69[0])) /* synthesis syn_instantiated=1 */ ;
    defparam Kd_delay_counter_1015_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3335_4_lut (.I0(GND_net), .I1(n14793[1]), .I2(n328_adj_3486), 
            .I3(n34325), .O(n14434[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3335_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3049_19 (.CI(n34653), .I0(n9125[16]), .I1(GND_net), .CO(n34654));
    SB_LUT4 add_3064_7_lut (.I0(GND_net), .I1(n8208[4]), .I2(n610), .I3(n35422), 
            .O(n8184[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3064_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3064_7 (.CI(n35422), .I0(n8208[4]), .I1(n610), .CO(n35423));
    SB_CARRY add_3335_4 (.CI(n34325), .I0(n14793[1]), .I1(n328_adj_3486), 
            .CO(n34326));
    SB_CARRY add_3272_21 (.CI(n34408), .I0(n13594[18]), .I1(GND_net), 
            .CO(n34409));
    SB_LUT4 add_3272_20_lut (.I0(GND_net), .I1(n13594[17]), .I2(GND_net), 
            .I3(n34407), .O(n13109[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3272_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3335_3_lut (.I0(GND_net), .I1(n14793[0]), .I2(n231_adj_3487), 
            .I3(n34324), .O(n14434[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3335_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3079_7_lut (.I0(GND_net), .I1(n9319[4]), .I2(n655), .I3(n35632), 
            .O(n8439[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3079_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3071_15 (.CI(n35556), .I0(n8348[12]), .I1(GND_net), .CO(n35557));
    SB_LUT4 mult_12_add_2137_10_lut (.I0(GND_net), .I1(n7956[7]), .I2(GND_net), 
            .I3(n35220), .O(n191[9])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_12_add_2137_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3335_3 (.CI(n34324), .I0(n14793[0]), .I1(n231_adj_3487), 
            .CO(n34325));
    SB_LUT4 add_3335_2_lut (.I0(GND_net), .I1(n41_adj_3488), .I2(n134_adj_3489), 
            .I3(GND_net), .O(n14434[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3335_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3068_14_lut (.I0(GND_net), .I1(n8294[11]), .I2(GND_net), 
            .I3(n35507), .O(n8274[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3068_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3335_2 (.CI(GND_net), .I0(n41_adj_3488), .I1(n134_adj_3489), 
            .CO(n34324));
    SB_CARRY mult_12_add_2137_10 (.CI(n35220), .I0(n7956[7]), .I1(GND_net), 
            .CO(n35221));
    SB_CARRY Kd_delay_counter_1015_add_4_2 (.CI(VCC_net), .I0(GND_net), 
            .I1(Kd_delay_counter[0]), .CO(n35011));
    SB_CARRY add_3079_7 (.CI(n35632), .I0(n9319[4]), .I1(n655), .CO(n35633));
    SB_LUT4 add_3071_14_lut (.I0(GND_net), .I1(n8348[11]), .I2(GND_net), 
            .I3(n35555), .O(n8331[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3071_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3049_18_lut (.I0(GND_net), .I1(n9125[15]), .I2(GND_net), 
            .I3(n34652), .O(n7760[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3049_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i73_4_lut (.I0(pwm[23]), .I1(n25), .I2(n30), .I3(n26), .O(n878));   // verilog/motorControl.v(86[19:44])
    defparam i73_4_lut.LUT_INIT = 16'haaa8;
    SB_CARRY add_3049_18 (.CI(n34652), .I0(n9125[15]), .I1(GND_net), .CO(n34653));
    SB_LUT4 add_3473_10_lut (.I0(GND_net), .I1(n16571[7]), .I2(GND_net), 
            .I3(n34323), .O(n16505[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3473_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3473_9_lut (.I0(GND_net), .I1(n16571[6]), .I2(GND_net), 
            .I3(n34322), .O(n16505[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3473_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3066_10 (.CI(n35466), .I0(n8253[7]), .I1(GND_net), .CO(n35467));
    SB_CARRY add_3473_9 (.CI(n34322), .I0(n16571[6]), .I1(GND_net), .CO(n34323));
    SB_LUT4 add_3473_8_lut (.I0(GND_net), .I1(n16571[5]), .I2(n746), .I3(n34321), 
            .O(n16505[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3473_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3066_9_lut (.I0(GND_net), .I1(n8253[6]), .I2(GND_net), 
            .I3(n35465), .O(n8231[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3066_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3064_6_lut (.I0(GND_net), .I1(n8208[3]), .I2(n513), .I3(n35421), 
            .O(n8184[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3064_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_2_lut (.I0(hall3), .I1(n878), .I2(GND_net), .I3(GND_net), 
            .O(n40121));   // verilog/motorControl.v(86[14] 109[8])
    defparam i1_2_lut.LUT_INIT = 16'h4444;
    SB_CARRY add_3061_5 (.CI(n35351), .I0(n8133[2]), .I1(n407_adj_3482), 
            .CO(n35352));
    SB_LUT4 add_3049_17_lut (.I0(GND_net), .I1(n9125[14]), .I2(GND_net), 
            .I3(n34651), .O(n7760[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3049_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3473_8 (.CI(n34321), .I0(n16571[5]), .I1(n746), .CO(n34322));
    SB_LUT4 mult_12_add_2137_9_lut (.I0(GND_net), .I1(n7956[6]), .I2(GND_net), 
            .I3(n35219), .O(n191[8])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_12_add_2137_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3049_17 (.CI(n34651), .I0(n9125[14]), .I1(GND_net), .CO(n34652));
    SB_LUT4 add_3049_16_lut (.I0(GND_net), .I1(n9125[13]), .I2(GND_net), 
            .I3(n34650), .O(n7760[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3049_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3473_7_lut (.I0(GND_net), .I1(n16571[4]), .I2(n649), .I3(n34320), 
            .O(n16505[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3473_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_70_add_3_25_lut (.I0(GND_net), .I1(GND_net), .I2(GATES_5__N_3055), 
            .I3(n34166), .O(n853)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_70_add_3_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3473_7 (.CI(n34320), .I0(n16571[4]), .I1(n649), .CO(n34321));
    SB_LUT4 unary_minus_70_add_3_24_lut (.I0(n852[18]), .I1(GND_net), .I2(n73[22]), 
            .I3(n34165), .O(n21)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_70_add_3_24_lut.LUT_INIT = 16'hebbe;
    SB_CARRY add_3064_6 (.CI(n35421), .I0(n8208[3]), .I1(n513), .CO(n35422));
    SB_CARRY mult_12_add_2137_9 (.CI(n35219), .I0(n7956[6]), .I1(GND_net), 
            .CO(n35220));
    SB_LUT4 add_3473_6_lut (.I0(GND_net), .I1(n16571[3]), .I2(n552), .I3(n34319), 
            .O(n16505[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3473_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3061_4_lut (.I0(GND_net), .I1(n8133[1]), .I2(n310_adj_3494), 
            .I3(n35350), .O(n8106[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3061_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_12_add_2137_8_lut (.I0(GND_net), .I1(n7956[5]), .I2(n680_adj_3495), 
            .I3(n35218), .O(n191[7])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_12_add_2137_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3473_6 (.CI(n34319), .I0(n16571[3]), .I1(n552), .CO(n34320));
    SB_CARRY mult_12_add_2137_8 (.CI(n35218), .I0(n7956[5]), .I1(n680_adj_3495), 
            .CO(n35219));
    SB_LUT4 add_3473_5_lut (.I0(GND_net), .I1(n16571[2]), .I2(n455_c), 
            .I3(n34318), .O(n16505[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3473_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3049_16 (.CI(n34650), .I0(n9125[13]), .I1(GND_net), .CO(n34651));
    SB_CARRY add_3473_5 (.CI(n34318), .I0(n16571[2]), .I1(n455_c), .CO(n34319));
    SB_LUT4 add_3473_4_lut (.I0(GND_net), .I1(n16571[1]), .I2(n358), .I3(n34317), 
            .O(n16505[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3473_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3049_15_lut (.I0(GND_net), .I1(n9125[12]), .I2(GND_net), 
            .I3(n34649), .O(n7760[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3049_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3473_4 (.CI(n34317), .I0(n16571[1]), .I1(n358), .CO(n34318));
    SB_LUT4 add_3473_3_lut (.I0(GND_net), .I1(n16571[0]), .I2(n261), .I3(n34316), 
            .O(n16505[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3473_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_70_add_3_24 (.CI(n34165), .I0(GND_net), .I1(n73[22]), 
            .CO(n34166));
    SB_CARRY add_3061_4 (.CI(n35350), .I0(n8133[1]), .I1(n310_adj_3494), 
            .CO(n35351));
    SB_LUT4 mult_12_add_2137_7_lut (.I0(GND_net), .I1(n7956[4]), .I2(n583_adj_3496), 
            .I3(n35217), .O(n191[6])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_12_add_2137_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3068_14 (.CI(n35507), .I0(n8294[11]), .I1(GND_net), .CO(n35508));
    SB_CARRY add_3049_15 (.CI(n34649), .I0(n9125[12]), .I1(GND_net), .CO(n34650));
    SB_LUT4 add_3049_14_lut (.I0(GND_net), .I1(n9125[11]), .I2(GND_net), 
            .I3(n34648), .O(n7760[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3049_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3473_3 (.CI(n34316), .I0(n16571[0]), .I1(n261), .CO(n34317));
    SB_LUT4 add_3473_2_lut (.I0(GND_net), .I1(n71), .I2(n164), .I3(GND_net), 
            .O(n16505[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3473_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3049_14 (.CI(n34648), .I0(n9125[11]), .I1(GND_net), .CO(n34649));
    SB_CARRY add_3473_2 (.CI(GND_net), .I0(n71), .I1(n164), .CO(n34316));
    SB_LUT4 unary_minus_70_add_3_23_lut (.I0(GND_net), .I1(GND_net), .I2(n73[21]), 
            .I3(n34164), .O(n855)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_70_add_3_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3071_14 (.CI(n35555), .I0(n8348[11]), .I1(GND_net), .CO(n35556));
    SB_CARRY mult_12_add_2137_7 (.CI(n35217), .I0(n7956[4]), .I1(n583_adj_3496), 
            .CO(n35218));
    SB_LUT4 add_3049_13_lut (.I0(GND_net), .I1(n9125[10]), .I2(GND_net), 
            .I3(n34647), .O(n7760[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3049_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_70_add_3_23 (.CI(n34164), .I0(GND_net), .I1(n73[21]), 
            .CO(n34165));
    SB_CARRY add_3049_13 (.CI(n34647), .I0(n9125[10]), .I1(GND_net), .CO(n34648));
    SB_LUT4 mult_12_add_2137_6_lut (.I0(GND_net), .I1(n7956[3]), .I2(n486_adj_3497), 
            .I3(n35216), .O(n191[5])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_12_add_2137_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3049_12_lut (.I0(GND_net), .I1(n9125[9]), .I2(GND_net), 
            .I3(n34646), .O(n7760[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3049_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_70_add_3_22_lut (.I0(GND_net), .I1(GND_net), .I2(n73[20]), 
            .I3(n34163), .O(n856)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_70_add_3_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3079_6_lut (.I0(GND_net), .I1(n9319[3]), .I2(n558), .I3(n35631), 
            .O(n8439[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3079_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3079_6 (.CI(n35631), .I0(n9319[3]), .I1(n558), .CO(n35632));
    SB_LUT4 add_3079_5_lut (.I0(GND_net), .I1(n9319[2]), .I2(n461_c), 
            .I3(n35630), .O(n8439[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3079_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_70_add_3_22 (.CI(n34163), .I0(GND_net), .I1(n73[20]), 
            .CO(n34164));
    SB_LUT4 unary_minus_70_add_3_21_lut (.I0(GND_net), .I1(GND_net), .I2(n73[19]), 
            .I3(n34162), .O(n857)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_70_add_3_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_70_add_3_21 (.CI(n34162), .I0(GND_net), .I1(n73[19]), 
            .CO(n34163));
    SB_LUT4 unary_minus_70_add_3_20_lut (.I0(GND_net), .I1(GND_net), .I2(n73[18]), 
            .I3(n34161), .O(n852[18])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_70_add_3_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_70_add_3_20 (.CI(n34161), .I0(GND_net), .I1(n73[18]), 
            .CO(n34162));
    SB_CARRY add_3049_12 (.CI(n34646), .I0(n9125[9]), .I1(GND_net), .CO(n34647));
    SB_LUT4 unary_minus_70_add_3_19_lut (.I0(GND_net), .I1(GND_net), .I2(n73[17]), 
            .I3(n34160), .O(n859)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_70_add_3_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_70_add_3_19 (.CI(n34160), .I0(GND_net), .I1(n73[17]), 
            .CO(n34161));
    SB_LUT4 add_3049_11_lut (.I0(GND_net), .I1(n9125[8]), .I2(GND_net), 
            .I3(n34645), .O(n7760[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3049_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3061_3_lut (.I0(GND_net), .I1(n8133[0]), .I2(n213_adj_3502), 
            .I3(n35349), .O(n8106[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3061_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_70_add_3_18_lut (.I0(GND_net), .I1(GND_net), .I2(n73[16]), 
            .I3(n34159), .O(n860)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_70_add_3_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_20061_33_lut (.I0(GND_net), .I1(n63[31]), .I2(n7061[0]), 
            .I3(n34310), .O(\PID_CONTROLLER.result_31__N_3003 [31])) /* synthesis syn_instantiated=1 */ ;
    defparam add_20061_33_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_12_add_2137_6 (.CI(n35216), .I0(n7956[3]), .I1(n486_adj_3497), 
            .CO(n35217));
    SB_CARRY unary_minus_70_add_3_18 (.CI(n34159), .I0(GND_net), .I1(n73[16]), 
            .CO(n34160));
    SB_CARRY add_3049_11 (.CI(n34645), .I0(n9125[8]), .I1(GND_net), .CO(n34646));
    SB_LUT4 add_20061_32_lut (.I0(GND_net), .I1(n63[30]), .I2(n191[30]), 
            .I3(n34309), .O(\PID_CONTROLLER.result_31__N_3003 [30])) /* synthesis syn_instantiated=1 */ ;
    defparam add_20061_32_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3049_10_lut (.I0(GND_net), .I1(n9125[7]), .I2(GND_net), 
            .I3(n34644), .O(n7760[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3049_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3049_10 (.CI(n34644), .I0(n9125[7]), .I1(GND_net), .CO(n34645));
    SB_CARRY add_20061_32 (.CI(n34309), .I0(n63[30]), .I1(n191[30]), .CO(n34310));
    SB_LUT4 add_20061_31_lut (.I0(GND_net), .I1(n63[29]), .I2(n191[29]), 
            .I3(n34308), .O(\PID_CONTROLLER.result_31__N_3003 [29])) /* synthesis syn_instantiated=1 */ ;
    defparam add_20061_31_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_20061_31 (.CI(n34308), .I0(n63[29]), .I1(n191[29]), .CO(n34309));
    SB_LUT4 add_20061_30_lut (.I0(GND_net), .I1(n63[28]), .I2(n191[28]), 
            .I3(n34307), .O(\PID_CONTROLLER.result_31__N_3003 [28])) /* synthesis syn_instantiated=1 */ ;
    defparam add_20061_30_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_70_add_3_17_lut (.I0(GND_net), .I1(GND_net), .I2(n73[15]), 
            .I3(n34158), .O(n861)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_70_add_3_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3066_9 (.CI(n35465), .I0(n8253[6]), .I1(GND_net), .CO(n35466));
    SB_LUT4 add_3064_5_lut (.I0(GND_net), .I1(n8208[2]), .I2(n416), .I3(n35420), 
            .O(n8184[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3064_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3079_5 (.CI(n35630), .I0(n9319[2]), .I1(n461_c), .CO(n35631));
    SB_CARRY add_3061_3 (.CI(n35349), .I0(n8133[0]), .I1(n213_adj_3502), 
            .CO(n35350));
    SB_LUT4 mult_12_add_2137_5_lut (.I0(GND_net), .I1(n7956[2]), .I2(n389_adj_3504), 
            .I3(n35215), .O(n191[4])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_12_add_2137_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3049_9_lut (.I0(GND_net), .I1(n9125[6]), .I2(GND_net), 
            .I3(n34643), .O(n7760[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3049_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3049_9 (.CI(n34643), .I0(n9125[6]), .I1(GND_net), .CO(n34644));
    SB_CARRY add_20061_30 (.CI(n34307), .I0(n63[28]), .I1(n191[28]), .CO(n34308));
    SB_CARRY unary_minus_70_add_3_17 (.CI(n34158), .I0(GND_net), .I1(n73[15]), 
            .CO(n34159));
    SB_LUT4 add_20061_29_lut (.I0(GND_net), .I1(n63[27]), .I2(n191[27]), 
            .I3(n34306), .O(\PID_CONTROLLER.result_31__N_3003 [27])) /* synthesis syn_instantiated=1 */ ;
    defparam add_20061_29_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_70_add_3_16_lut (.I0(GND_net), .I1(GND_net), .I2(n73[14]), 
            .I3(n34157), .O(n862)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_70_add_3_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3049_8_lut (.I0(GND_net), .I1(n9125[5]), .I2(n686_adj_3506), 
            .I3(n34642), .O(n7760[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3049_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_70_add_3_16 (.CI(n34157), .I0(GND_net), .I1(n73[14]), 
            .CO(n34158));
    SB_CARRY add_20061_29 (.CI(n34306), .I0(n63[27]), .I1(n191[27]), .CO(n34307));
    SB_LUT4 add_3079_4_lut (.I0(GND_net), .I1(n9319[1]), .I2(n364_adj_3507), 
            .I3(n35629), .O(n8439[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3079_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3079_4 (.CI(n35629), .I0(n9319[1]), .I1(n364_adj_3507), 
            .CO(n35630));
    SB_LUT4 add_3079_3_lut (.I0(GND_net), .I1(n9319[0]), .I2(n267), .I3(n35628), 
            .O(n8439[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3079_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_70_add_3_15_lut (.I0(GND_net), .I1(GND_net), .I2(n73[13]), 
            .I3(n34156), .O(n863)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_70_add_3_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_12_add_2137_5 (.CI(n35215), .I0(n7956[2]), .I1(n389_adj_3504), 
            .CO(n35216));
    SB_LUT4 add_20061_28_lut (.I0(GND_net), .I1(n63[26]), .I2(n191[26]), 
            .I3(n34305), .O(\PID_CONTROLLER.result_31__N_3003 [26])) /* synthesis syn_instantiated=1 */ ;
    defparam add_20061_28_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_70_add_3_15 (.CI(n34156), .I0(GND_net), .I1(n73[13]), 
            .CO(n34157));
    SB_CARRY add_20061_28 (.CI(n34305), .I0(n63[26]), .I1(n191[26]), .CO(n34306));
    SB_CARRY add_3049_8 (.CI(n34642), .I0(n9125[5]), .I1(n686_adj_3506), 
            .CO(n34643));
    SB_LUT4 unary_minus_70_add_3_14_lut (.I0(GND_net), .I1(GND_net), .I2(n73[12]), 
            .I3(n34155), .O(n864)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_70_add_3_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3061_2_lut (.I0(GND_net), .I1(n23_adj_3510), .I2(n116_adj_3511), 
            .I3(GND_net), .O(n8106[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3061_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_20061_27_lut (.I0(GND_net), .I1(n63[25]), .I2(n191[25]), 
            .I3(n34304), .O(\PID_CONTROLLER.result_31__N_3003 [25])) /* synthesis syn_instantiated=1 */ ;
    defparam add_20061_27_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_20061_27 (.CI(n34304), .I0(n63[25]), .I1(n191[25]), .CO(n34305));
    SB_LUT4 mult_12_add_2137_4_lut (.I0(GND_net), .I1(n7956[1]), .I2(n292_adj_3512), 
            .I3(n35214), .O(n191[3])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_12_add_2137_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_70_add_3_14 (.CI(n34155), .I0(GND_net), .I1(n73[12]), 
            .CO(n34156));
    SB_LUT4 add_3049_7_lut (.I0(GND_net), .I1(n9125[4]), .I2(n589_adj_3513), 
            .I3(n34641), .O(n7760[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3049_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_20061_26_lut (.I0(GND_net), .I1(n63[24]), .I2(n191[24]), 
            .I3(n34303), .O(\PID_CONTROLLER.result_31__N_3003 [24])) /* synthesis syn_instantiated=1 */ ;
    defparam add_20061_26_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3061_2 (.CI(GND_net), .I0(n23_adj_3510), .I1(n116_adj_3511), 
            .CO(n35349));
    SB_CARRY mult_12_add_2137_4 (.CI(n35214), .I0(n7956[1]), .I1(n292_adj_3512), 
            .CO(n35215));
    SB_LUT4 unary_minus_70_add_3_13_lut (.I0(GND_net), .I1(GND_net), .I2(n73[11]), 
            .I3(n34154), .O(n865)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_70_add_3_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_20061_26 (.CI(n34303), .I0(n63[24]), .I1(n191[24]), .CO(n34304));
    SB_CARRY unary_minus_70_add_3_13 (.CI(n34154), .I0(GND_net), .I1(n73[11]), 
            .CO(n34155));
    SB_CARRY add_3049_7 (.CI(n34641), .I0(n9125[4]), .I1(n589_adj_3513), 
            .CO(n34642));
    SB_LUT4 add_3049_6_lut (.I0(GND_net), .I1(n9125[3]), .I2(n492_adj_3515), 
            .I3(n34640), .O(n7760[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3049_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_20061_25_lut (.I0(GND_net), .I1(n63[23]), .I2(n191[23]), 
            .I3(n34302), .O(\PID_CONTROLLER.result_31__N_3003 [23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_20061_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_20061_25 (.CI(n34302), .I0(n63[23]), .I1(n191[23]), .CO(n34303));
    SB_LUT4 add_20061_24_lut (.I0(GND_net), .I1(n63[22]), .I2(n191[22]), 
            .I3(n34301), .O(\PID_CONTROLLER.result_31__N_3003 [22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_20061_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_70_add_3_12_lut (.I0(GND_net), .I1(GND_net), .I2(n73[10]), 
            .I3(n34153), .O(n866)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_70_add_3_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_70_add_3_12 (.CI(n34153), .I0(GND_net), .I1(n73[10]), 
            .CO(n34154));
    SB_LUT4 unary_minus_70_add_3_11_lut (.I0(GND_net), .I1(GND_net), .I2(n73[9]), 
            .I3(n34152), .O(n867)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_70_add_3_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_20061_24 (.CI(n34301), .I0(n63[22]), .I1(n191[22]), .CO(n34302));
    SB_LUT4 add_20061_23_lut (.I0(GND_net), .I1(n63[21]), .I2(n191[21]), 
            .I3(n34300), .O(\PID_CONTROLLER.result_31__N_3003 [21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_20061_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_70_add_3_11 (.CI(n34152), .I0(GND_net), .I1(n73[9]), 
            .CO(n34153));
    SB_LUT4 unary_minus_70_add_3_10_lut (.I0(GND_net), .I1(GND_net), .I2(n73[8]), 
            .I3(n34151), .O(n868)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_70_add_3_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_70_add_3_10 (.CI(n34151), .I0(GND_net), .I1(n73[8]), 
            .CO(n34152));
    SB_CARRY add_3049_6 (.CI(n34640), .I0(n9125[3]), .I1(n492_adj_3515), 
            .CO(n34641));
    SB_CARRY add_20061_23 (.CI(n34300), .I0(n63[21]), .I1(n191[21]), .CO(n34301));
    SB_LUT4 i1_2_lut_adj_1402 (.I0(hall3), .I1(hall1), .I2(GND_net), .I3(GND_net), 
            .O(n40176));   // verilog/motorControl.v(86[14] 109[8])
    defparam i1_2_lut_adj_1402.LUT_INIT = 16'h2222;
    SB_LUT4 unary_minus_70_add_3_9_lut (.I0(GND_net), .I1(GND_net), .I2(n73[7]), 
            .I3(n34150), .O(n869)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_70_add_3_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3049_5_lut (.I0(GND_net), .I1(n9125[2]), .I2(n395_adj_3520), 
            .I3(n34639), .O(n7760[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3049_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3079_3 (.CI(n35628), .I0(n9319[0]), .I1(n267), .CO(n35629));
    SB_LUT4 add_3079_2_lut (.I0(GND_net), .I1(n86), .I2(n170_adj_3521), 
            .I3(GND_net), .O(n8439[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3079_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_20061_22_lut (.I0(GND_net), .I1(n63[20]), .I2(n191[20]), 
            .I3(n34299), .O(\PID_CONTROLLER.result_31__N_3003 [20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_20061_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3079_2 (.CI(GND_net), .I0(n86), .I1(n170_adj_3521), .CO(n35628));
    SB_LUT4 add_3078_9_lut (.I0(GND_net), .I1(n8439[6]), .I2(GND_net), 
            .I3(n35627), .O(n8429[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3078_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3078_8_lut (.I0(GND_net), .I1(n8439[5]), .I2(n749), .I3(n35626), 
            .O(n8429[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3078_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3078_8 (.CI(n35626), .I0(n8439[5]), .I1(n749), .CO(n35627));
    SB_CARRY unary_minus_70_add_3_9 (.CI(n34150), .I0(GND_net), .I1(n73[7]), 
            .CO(n34151));
    SB_CARRY add_20061_22 (.CI(n34299), .I0(n63[20]), .I1(n191[20]), .CO(n34300));
    SB_LUT4 unary_minus_70_add_3_8_lut (.I0(GND_net), .I1(GND_net), .I2(n73[6]), 
            .I3(n34149), .O(n870)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_70_add_3_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_70_add_3_8 (.CI(n34149), .I0(GND_net), .I1(n73[6]), 
            .CO(n34150));
    SB_CARRY add_3049_5 (.CI(n34639), .I0(n9125[2]), .I1(n395_adj_3520), 
            .CO(n34640));
    SB_LUT4 add_20061_21_lut (.I0(GND_net), .I1(n63[19]), .I2(n191[19]), 
            .I3(n34298), .O(\PID_CONTROLLER.result_31__N_3003 [19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_20061_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_70_add_3_7_lut (.I0(GND_net), .I1(GND_net), .I2(n73[5]), 
            .I3(n34148), .O(n871)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_70_add_3_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_70_add_3_7 (.CI(n34148), .I0(GND_net), .I1(n73[5]), 
            .CO(n34149));
    SB_CARRY add_20061_21 (.CI(n34298), .I0(n63[19]), .I1(n191[19]), .CO(n34299));
    SB_LUT4 unary_minus_70_add_3_6_lut (.I0(GND_net), .I1(GND_net), .I2(n73[4]), 
            .I3(n34147), .O(n872)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_70_add_3_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_70_add_3_6 (.CI(n34147), .I0(GND_net), .I1(n73[4]), 
            .CO(n34148));
    SB_LUT4 mult_12_add_2137_3_lut (.I0(GND_net), .I1(n7956[0]), .I2(n195_adj_3525), 
            .I3(n35213), .O(n191[2])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_12_add_2137_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3049_4_lut (.I0(GND_net), .I1(n9125[1]), .I2(n298_adj_3526), 
            .I3(n34638), .O(n7760[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3049_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_20061_20_lut (.I0(GND_net), .I1(n63[18]), .I2(n191[18]), 
            .I3(n34297), .O(\PID_CONTROLLER.result_31__N_3003 [18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_20061_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_70_add_3_5_lut (.I0(GND_net), .I1(GND_net), .I2(n73[3]), 
            .I3(n34146), .O(n873)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_70_add_3_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_70_add_3_5 (.CI(n34146), .I0(GND_net), .I1(n73[3]), 
            .CO(n34147));
    SB_CARRY add_20061_20 (.CI(n34297), .I0(n63[18]), .I1(n191[18]), .CO(n34298));
    SB_LUT4 unary_minus_70_add_3_4_lut (.I0(GND_net), .I1(GND_net), .I2(n73[2]), 
            .I3(n34145), .O(n874)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_70_add_3_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_70_add_3_4 (.CI(n34145), .I0(GND_net), .I1(n73[2]), 
            .CO(n34146));
    SB_CARRY add_3049_4 (.CI(n34638), .I0(n9125[1]), .I1(n298_adj_3526), 
            .CO(n34639));
    SB_LUT4 add_3071_13_lut (.I0(GND_net), .I1(n8348[10]), .I2(GND_net), 
            .I3(n35554), .O(n8331[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3071_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3078_7_lut (.I0(GND_net), .I1(n8439[4]), .I2(n652), .I3(n35625), 
            .O(n8429[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3078_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3071_13 (.CI(n35554), .I0(n8348[10]), .I1(GND_net), .CO(n35555));
    SB_LUT4 add_3068_13_lut (.I0(GND_net), .I1(n8294[10]), .I2(GND_net), 
            .I3(n35506), .O(n8274[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3068_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3066_8_lut (.I0(GND_net), .I1(n8253[5]), .I2(n713_adj_3529), 
            .I3(n35464), .O(n8231[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3066_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3064_5 (.CI(n35420), .I0(n8208[2]), .I1(n416), .CO(n35421));
    SB_LUT4 add_3060_27_lut (.I0(GND_net), .I1(n8106[24]), .I2(GND_net), 
            .I3(n35348), .O(n8078[25])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3060_27_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_12_add_2137_3 (.CI(n35213), .I0(n7956[0]), .I1(n195_adj_3525), 
            .CO(n35214));
    SB_LUT4 mult_12_add_2137_2_lut (.I0(GND_net), .I1(n5_adj_3531), .I2(n98_adj_3532), 
            .I3(GND_net), .O(n191[1])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_12_add_2137_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3078_7 (.CI(n35625), .I0(n8439[4]), .I1(n652), .CO(n35626));
    SB_LUT4 add_20061_19_lut (.I0(GND_net), .I1(n63[17]), .I2(n191[17]), 
            .I3(n34296), .O(\PID_CONTROLLER.result_31__N_3003 [17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_20061_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3049_3_lut (.I0(GND_net), .I1(n9125[0]), .I2(n201_adj_3533), 
            .I3(n34637), .O(n7760[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3049_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_70_add_3_3_lut (.I0(GND_net), .I1(GND_net), .I2(n73[1]), 
            .I3(n34144), .O(n875)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_70_add_3_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_12_add_2137_2 (.CI(GND_net), .I0(n5_adj_3531), .I1(n98_adj_3532), 
            .CO(n35213));
    SB_CARRY add_3049_3 (.CI(n34637), .I0(n9125[0]), .I1(n201_adj_3533), 
            .CO(n34638));
    SB_CARRY unary_minus_70_add_3_3 (.CI(n34144), .I0(GND_net), .I1(n73[1]), 
            .CO(n34145));
    SB_CARRY add_20061_19 (.CI(n34296), .I0(n63[17]), .I1(n191[17]), .CO(n34297));
    SB_LUT4 add_20061_18_lut (.I0(GND_net), .I1(n63[16]), .I2(n191[16]), 
            .I3(n34295), .O(\PID_CONTROLLER.result_31__N_3003 [16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_20061_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_70_add_3_2_lut (.I0(n25474), .I1(GND_net), .I2(n73[0]), 
            .I3(VCC_net), .O(n44074)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_70_add_3_2_lut.LUT_INIT = 16'h8228;
    SB_CARRY unary_minus_70_add_3_2 (.CI(VCC_net), .I0(GND_net), .I1(n73[0]), 
            .CO(n34144));
    SB_CARRY add_20061_18 (.CI(n34295), .I0(n63[16]), .I1(n191[16]), .CO(n34296));
    SB_LUT4 unary_minus_21_add_3_12_lut (.I0(GND_net), .I1(GND_net), .I2(n6_adj_3536), 
            .I3(n34143), .O(n70[10])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_21_add_3_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3049_2_lut (.I0(GND_net), .I1(n11_adj_3537), .I2(n104_adj_3538), 
            .I3(GND_net), .O(n7760[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3049_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_20061_17_lut (.I0(GND_net), .I1(n63[15]), .I2(n191[15]), 
            .I3(n34294), .O(\PID_CONTROLLER.result_31__N_3003 [15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_20061_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_20061_17 (.CI(n34294), .I0(n63[15]), .I1(n191[15]), .CO(n34295));
    SB_LUT4 add_20061_16_lut (.I0(GND_net), .I1(n63[14]), .I2(n191[14]), 
            .I3(n34293), .O(\PID_CONTROLLER.result_31__N_3003 [14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_20061_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_21_add_3_11_lut (.I0(GND_net), .I1(GND_net), .I2(n6_adj_3536), 
            .I3(n34142), .O(n70[9])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_21_add_3_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_21_add_3_11 (.CI(n34142), .I0(GND_net), .I1(n6_adj_3536), 
            .CO(n34143));
    SB_LUT4 unary_minus_21_add_3_10_lut (.I0(GND_net), .I1(GND_net), .I2(n75[8]), 
            .I3(n34141), .O(n70[8])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_21_add_3_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_21_add_3_10 (.CI(n34141), .I0(GND_net), .I1(n75[8]), 
            .CO(n34142));
    SB_LUT4 add_3078_6_lut (.I0(GND_net), .I1(n8439[3]), .I2(n555), .I3(n35624), 
            .O(n8429[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3078_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3078_6 (.CI(n35624), .I0(n8439[3]), .I1(n555), .CO(n35625));
    SB_LUT4 add_3078_5_lut (.I0(GND_net), .I1(n8439[2]), .I2(n458_c), 
            .I3(n35623), .O(n8429[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3078_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3068_13 (.CI(n35506), .I0(n8294[10]), .I1(GND_net), .CO(n35507));
    SB_LUT4 add_3060_26_lut (.I0(GND_net), .I1(n8106[23]), .I2(GND_net), 
            .I3(n35347), .O(n8078[24])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3060_26_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3121_21_lut (.I0(GND_net), .I1(n10118[18]), .I2(GND_net), 
            .I3(n35212), .O(n9327[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3121_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3024_10_lut (.I0(GND_net), .I1(n1804[22]), .I2(n1711), 
            .I3(n35987), .O(n7065[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3024_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3024_9_lut (.I0(GND_net), .I1(n1803[22]), .I2(n1707), 
            .I3(n35986), .O(n7065[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3024_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3024_9 (.CI(n35986), .I0(n1803[22]), .I1(n1707), .CO(n35987));
    SB_LUT4 add_3024_8_lut (.I0(GND_net), .I1(n1802[22]), .I2(n1703), 
            .I3(n35985), .O(n7065[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3024_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3024_8 (.CI(n35985), .I0(n1802[22]), .I1(n1703), .CO(n35986));
    SB_LUT4 add_3024_7_lut (.I0(GND_net), .I1(n1801[22]), .I2(n1699), 
            .I3(n35984), .O(n7065[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3024_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3024_7 (.CI(n35984), .I0(n1801[22]), .I1(n1699), .CO(n35985));
    SB_LUT4 add_3024_6_lut (.I0(GND_net), .I1(n1800[22]), .I2(n1695), 
            .I3(n35983), .O(n7065[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3024_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3024_6 (.CI(n35983), .I0(n1800[22]), .I1(n1695), .CO(n35984));
    SB_CARRY add_3049_2 (.CI(GND_net), .I0(n11_adj_3537), .I1(n104_adj_3538), 
            .CO(n34637));
    SB_CARRY add_20061_16 (.CI(n34293), .I0(n63[14]), .I1(n191[14]), .CO(n34294));
    SB_LUT4 add_3024_5_lut (.I0(GND_net), .I1(n1799[22]), .I2(n1691), 
            .I3(n35982), .O(n7065[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3024_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3024_5 (.CI(n35982), .I0(n1799[22]), .I1(n1691), .CO(n35983));
    SB_LUT4 add_3024_4_lut (.I0(GND_net), .I1(n1798[22]), .I2(n1687), 
            .I3(n35981), .O(n7065[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3024_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3071_12_lut (.I0(GND_net), .I1(n8348[9]), .I2(GND_net), 
            .I3(n35553), .O(n8331[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3071_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3071_12 (.CI(n35553), .I0(n8348[9]), .I1(GND_net), .CO(n35554));
    SB_CARRY add_3078_5 (.CI(n35623), .I0(n8439[2]), .I1(n458_c), .CO(n35624));
    SB_LUT4 add_3071_11_lut (.I0(GND_net), .I1(n8348[8]), .I2(GND_net), 
            .I3(n35552), .O(n8331[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3071_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3024_4 (.CI(n35981), .I0(n1798[22]), .I1(n1687), .CO(n35982));
    SB_LUT4 add_3024_3_lut (.I0(GND_net), .I1(n1797[22]), .I2(n1683), 
            .I3(n35980), .O(n7065[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3024_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3024_3 (.CI(n35980), .I0(n1797[22]), .I1(n1683), .CO(n35981));
    SB_LUT4 add_3024_2_lut (.I0(GND_net), .I1(n1796[22]), .I2(\PID_CONTROLLER.integral [9]), 
            .I3(GND_net), .O(n7065[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3024_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3024_2 (.CI(GND_net), .I0(n1796[22]), .I1(\PID_CONTROLLER.integral [9]), 
            .CO(n35980));
    SB_LUT4 add_3081_22_lut (.I0(GND_net), .I1(n9327[19]), .I2(GND_net), 
            .I3(n35979), .O(n8472[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3081_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_20061_15_lut (.I0(GND_net), .I1(n63[13]), .I2(n191[13]), 
            .I3(n34292), .O(\PID_CONTROLLER.result_31__N_3003 [13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_20061_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_21_add_3_9_lut (.I0(GND_net), .I1(GND_net), .I2(n75[7]), 
            .I3(n34140), .O(n70[7])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_21_add_3_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3081_21_lut (.I0(GND_net), .I1(n9327[18]), .I2(GND_net), 
            .I3(n35978), .O(n8472[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3081_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_21_add_3_9 (.CI(n34140), .I0(GND_net), .I1(n75[7]), 
            .CO(n34141));
    SB_LUT4 add_3121_20_lut (.I0(GND_net), .I1(n10118[17]), .I2(GND_net), 
            .I3(n35211), .O(n9327[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3121_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3081_21 (.CI(n35978), .I0(n9327[18]), .I1(GND_net), .CO(n35979));
    SB_LUT4 add_3081_20_lut (.I0(GND_net), .I1(n9327[17]), .I2(GND_net), 
            .I3(n35977), .O(n8472[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3081_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3081_20 (.CI(n35977), .I0(n9327[17]), .I1(GND_net), .CO(n35978));
    SB_LUT4 add_3081_19_lut (.I0(GND_net), .I1(n9327[16]), .I2(GND_net), 
            .I3(n35976), .O(n8472[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3081_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3081_19 (.CI(n35976), .I0(n9327[16]), .I1(GND_net), .CO(n35977));
    SB_LUT4 add_3081_18_lut (.I0(GND_net), .I1(n9327[15]), .I2(GND_net), 
            .I3(n35975), .O(n8472[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3081_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3081_18 (.CI(n35975), .I0(n9327[15]), .I1(GND_net), .CO(n35976));
    SB_LUT4 add_3081_17_lut (.I0(GND_net), .I1(n9327[14]), .I2(GND_net), 
            .I3(n35974), .O(n8472[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3081_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3071_11 (.CI(n35552), .I0(n8348[8]), .I1(GND_net), .CO(n35553));
    SB_LUT4 add_3068_12_lut (.I0(GND_net), .I1(n8294[9]), .I2(GND_net), 
            .I3(n35505), .O(n8274[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3068_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3068_12 (.CI(n35505), .I0(n8294[9]), .I1(GND_net), .CO(n35506));
    SB_LUT4 add_3071_10_lut (.I0(GND_net), .I1(n8348[7]), .I2(GND_net), 
            .I3(n35551), .O(n8331[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3071_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3078_4_lut (.I0(GND_net), .I1(n8439[1]), .I2(n361), .I3(n35622), 
            .O(n8429[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3078_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3068_11_lut (.I0(GND_net), .I1(n8294[8]), .I2(GND_net), 
            .I3(n35504), .O(n8274[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3068_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3068_11 (.CI(n35504), .I0(n8294[8]), .I1(GND_net), .CO(n35505));
    SB_CARRY add_3071_10 (.CI(n35551), .I0(n8348[7]), .I1(GND_net), .CO(n35552));
    SB_CARRY add_3078_4 (.CI(n35622), .I0(n8439[1]), .I1(n361), .CO(n35623));
    SB_LUT4 add_3078_3_lut (.I0(GND_net), .I1(n8439[0]), .I2(n264), .I3(n35621), 
            .O(n8429[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3078_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3078_3 (.CI(n35621), .I0(n8439[0]), .I1(n264), .CO(n35622));
    SB_LUT4 add_3068_10_lut (.I0(GND_net), .I1(n8294[7]), .I2(GND_net), 
            .I3(n35503), .O(n8274[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3068_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3060_26 (.CI(n35347), .I0(n8106[23]), .I1(GND_net), .CO(n35348));
    SB_CARRY add_3066_8 (.CI(n35464), .I0(n8253[5]), .I1(n713_adj_3529), 
            .CO(n35465));
    SB_CARRY add_3121_20 (.CI(n35211), .I0(n10118[17]), .I1(GND_net), 
            .CO(n35212));
    SB_LUT4 add_3071_9_lut (.I0(GND_net), .I1(n8348[6]), .I2(GND_net), 
            .I3(n35550), .O(n8331[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3071_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3078_2_lut (.I0(GND_net), .I1(n74), .I2(n167_adj_3542), 
            .I3(GND_net), .O(n8429[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3078_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3078_2 (.CI(GND_net), .I0(n74), .I1(n167_adj_3542), .CO(n35621));
    SB_LUT4 add_3121_19_lut (.I0(GND_net), .I1(n10118[16]), .I2(GND_net), 
            .I3(n35210), .O(n9327[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3121_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3077_10_lut (.I0(GND_net), .I1(n8429[7]), .I2(GND_net), 
            .I3(n35620), .O(n8418[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3077_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3077_9_lut (.I0(GND_net), .I1(n8429[6]), .I2(GND_net), 
            .I3(n35619), .O(n8418[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3077_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3077_9 (.CI(n35619), .I0(n8429[6]), .I1(GND_net), .CO(n35620));
    SB_LUT4 add_3077_8_lut (.I0(GND_net), .I1(n8429[5]), .I2(n746_adj_3543), 
            .I3(n35618), .O(n8418[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3077_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3064_4_lut (.I0(GND_net), .I1(n8208[1]), .I2(n319), .I3(n35419), 
            .O(n8184[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3064_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3060_25_lut (.I0(GND_net), .I1(n8106[22]), .I2(GND_net), 
            .I3(n35346), .O(n8078[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3060_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3068_10 (.CI(n35503), .I0(n8294[7]), .I1(GND_net), .CO(n35504));
    SB_CARRY add_3121_19 (.CI(n35210), .I0(n10118[16]), .I1(GND_net), 
            .CO(n35211));
    SB_CARRY add_3077_8 (.CI(n35618), .I0(n8429[5]), .I1(n746_adj_3543), 
            .CO(n35619));
    SB_LUT4 add_3077_7_lut (.I0(GND_net), .I1(n8429[4]), .I2(n649_adj_3544), 
            .I3(n35617), .O(n8418[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3077_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3081_17 (.CI(n35974), .I0(n9327[14]), .I1(GND_net), .CO(n35975));
    SB_LUT4 add_3121_18_lut (.I0(GND_net), .I1(n10118[15]), .I2(GND_net), 
            .I3(n35209), .O(n9327[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3121_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3081_16_lut (.I0(GND_net), .I1(n9327[13]), .I2(GND_net), 
            .I3(n35973), .O(n8472[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3081_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3081_16 (.CI(n35973), .I0(n9327[13]), .I1(GND_net), .CO(n35974));
    SB_LUT4 add_3081_15_lut (.I0(GND_net), .I1(n9327[12]), .I2(GND_net), 
            .I3(n35972), .O(n8472[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3081_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3081_15 (.CI(n35972), .I0(n9327[12]), .I1(GND_net), .CO(n35973));
    SB_CARRY add_3060_25 (.CI(n35346), .I0(n8106[22]), .I1(GND_net), .CO(n35347));
    SB_CARRY add_3121_18 (.CI(n35209), .I0(n10118[15]), .I1(GND_net), 
            .CO(n35210));
    SB_LUT4 add_3081_14_lut (.I0(GND_net), .I1(n9327[11]), .I2(GND_net), 
            .I3(n35971), .O(n8472[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3081_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3081_14 (.CI(n35971), .I0(n9327[11]), .I1(GND_net), .CO(n35972));
    SB_LUT4 add_3081_13_lut (.I0(GND_net), .I1(n9327[10]), .I2(GND_net), 
            .I3(n35970), .O(n8472[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3081_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3081_13 (.CI(n35970), .I0(n9327[10]), .I1(GND_net), .CO(n35971));
    SB_LUT4 add_3081_12_lut (.I0(GND_net), .I1(n9327[9]), .I2(GND_net), 
            .I3(n35969), .O(n8472[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3081_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3121_17_lut (.I0(GND_net), .I1(n10118[14]), .I2(GND_net), 
            .I3(n35208), .O(n9327[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3121_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3081_12 (.CI(n35969), .I0(n9327[9]), .I1(GND_net), .CO(n35970));
    SB_CARRY add_20061_15 (.CI(n34292), .I0(n63[13]), .I1(n191[13]), .CO(n34293));
    SB_LUT4 unary_minus_21_add_3_8_lut (.I0(GND_net), .I1(GND_net), .I2(n75[6]), 
            .I3(n34139), .O(n414)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_21_add_3_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_21_add_3_8 (.CI(n34139), .I0(GND_net), .I1(n75[6]), 
            .CO(n34140));
    SB_LUT4 add_3081_11_lut (.I0(GND_net), .I1(n9327[8]), .I2(GND_net), 
            .I3(n35968), .O(n8472[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3081_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3081_11 (.CI(n35968), .I0(n9327[8]), .I1(GND_net), .CO(n35969));
    SB_LUT4 unary_minus_21_add_3_7_lut (.I0(GND_net), .I1(GND_net), .I2(n75[5]), 
            .I3(n34138), .O(n415)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_21_add_3_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3081_10_lut (.I0(GND_net), .I1(n9327[7]), .I2(GND_net), 
            .I3(n35967), .O(n8472[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3081_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3081_10 (.CI(n35967), .I0(n9327[7]), .I1(GND_net), .CO(n35968));
    SB_LUT4 add_3081_9_lut (.I0(GND_net), .I1(n9327[6]), .I2(GND_net), 
            .I3(n35966), .O(n8472[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3081_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3081_9 (.CI(n35966), .I0(n9327[6]), .I1(GND_net), .CO(n35967));
    SB_LUT4 add_3081_8_lut (.I0(GND_net), .I1(n9327[5]), .I2(n545), .I3(n35965), 
            .O(n8472[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3081_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3066_7_lut (.I0(GND_net), .I1(n8253[4]), .I2(n616_adj_3547), 
            .I3(n35463), .O(n8231[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3066_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3077_7 (.CI(n35617), .I0(n8429[4]), .I1(n649_adj_3544), 
            .CO(n35618));
    SB_CARRY add_3071_9 (.CI(n35550), .I0(n8348[6]), .I1(GND_net), .CO(n35551));
    SB_CARRY add_3081_8 (.CI(n35965), .I0(n9327[5]), .I1(n545), .CO(n35966));
    SB_LUT4 add_3081_7_lut (.I0(GND_net), .I1(n9327[4]), .I2(n472), .I3(n35964), 
            .O(n8472[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3081_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3081_7 (.CI(n35964), .I0(n9327[4]), .I1(n472), .CO(n35965));
    SB_LUT4 add_3081_6_lut (.I0(GND_net), .I1(n9327[3]), .I2(n399), .I3(n35963), 
            .O(n8472[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3081_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3081_6 (.CI(n35963), .I0(n9327[3]), .I1(n399), .CO(n35964));
    SB_LUT4 add_3081_5_lut (.I0(GND_net), .I1(n9327[2]), .I2(n326), .I3(n35962), 
            .O(n8472[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3081_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3077_6_lut (.I0(GND_net), .I1(n8429[3]), .I2(n552_adj_3548), 
            .I3(n35616), .O(n8418[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3077_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3081_5 (.CI(n35962), .I0(n9327[2]), .I1(n326), .CO(n35963));
    SB_LUT4 add_3068_9_lut (.I0(GND_net), .I1(n8294[6]), .I2(GND_net), 
            .I3(n35502), .O(n8274[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3068_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3081_4_lut (.I0(GND_net), .I1(n9327[1]), .I2(n253), .I3(n35961), 
            .O(n8472[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3081_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3081_4 (.CI(n35961), .I0(n9327[1]), .I1(n253), .CO(n35962));
    SB_CARRY add_3066_7 (.CI(n35463), .I0(n8253[4]), .I1(n616_adj_3547), 
            .CO(n35464));
    SB_LUT4 add_3081_3_lut (.I0(GND_net), .I1(n9327[0]), .I2(n180), .I3(n35960), 
            .O(n8472[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3081_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3064_4 (.CI(n35419), .I0(n8208[1]), .I1(n319), .CO(n35420));
    SB_CARRY add_3081_3 (.CI(n35960), .I0(n9327[0]), .I1(n180), .CO(n35961));
    SB_LUT4 add_3081_2_lut (.I0(GND_net), .I1(n35), .I2(n107), .I3(GND_net), 
            .O(n8472[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3081_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3060_24_lut (.I0(GND_net), .I1(n8106[21]), .I2(GND_net), 
            .I3(n35345), .O(n8078[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3060_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3077_6 (.CI(n35616), .I0(n8429[3]), .I1(n552_adj_3548), 
            .CO(n35617));
    SB_CARRY add_3121_17 (.CI(n35208), .I0(n10118[14]), .I1(GND_net), 
            .CO(n35209));
    SB_CARRY add_3081_2 (.CI(GND_net), .I0(n35), .I1(n107), .CO(n35960));
    SB_LUT4 add_3071_8_lut (.I0(GND_net), .I1(n8348[5]), .I2(n728), .I3(n35549), 
            .O(n8331[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3071_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3077_5_lut (.I0(GND_net), .I1(n8429[2]), .I2(n455_adj_3549), 
            .I3(n35615), .O(n8418[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3077_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1219_24_lut (.I0(GND_net), .I1(n8448[21]), .I2(GND_net), 
            .I3(n35959), .O(n1804[22])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1219_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3077_5 (.CI(n35615), .I0(n8429[2]), .I1(n455_adj_3549), 
            .CO(n35616));
    SB_LUT4 add_3121_16_lut (.I0(GND_net), .I1(n10118[13]), .I2(GND_net), 
            .I3(n35207), .O(n9327[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3121_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3068_9 (.CI(n35502), .I0(n8294[6]), .I1(GND_net), .CO(n35503));
    SB_LUT4 add_3077_4_lut (.I0(GND_net), .I1(n8429[1]), .I2(n358_adj_3550), 
            .I3(n35614), .O(n8418[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3077_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1219_23_lut (.I0(GND_net), .I1(n8448[20]), .I2(GND_net), 
            .I3(n35958), .O(n1804[21])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1219_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3068_8_lut (.I0(GND_net), .I1(n8294[5]), .I2(n719), .I3(n35501), 
            .O(n8274[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3068_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3077_4 (.CI(n35614), .I0(n8429[1]), .I1(n358_adj_3550), 
            .CO(n35615));
    SB_CARRY add_3060_24 (.CI(n35345), .I0(n8106[21]), .I1(GND_net), .CO(n35346));
    SB_CARRY mult_14_add_1219_23 (.CI(n35958), .I0(n8448[20]), .I1(GND_net), 
            .CO(n35959));
    SB_CARRY add_3071_8 (.CI(n35549), .I0(n8348[5]), .I1(n728), .CO(n35550));
    SB_CARRY add_3121_16 (.CI(n35207), .I0(n10118[13]), .I1(GND_net), 
            .CO(n35208));
    SB_LUT4 add_3279_15_lut (.I0(GND_net), .I1(n13734[12]), .I2(GND_net), 
            .I3(n34636), .O(n13256[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3279_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3279_14_lut (.I0(GND_net), .I1(n13734[11]), .I2(GND_net), 
            .I3(n34635), .O(n13256[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3279_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3066_6_lut (.I0(GND_net), .I1(n8253[3]), .I2(n519_adj_3551), 
            .I3(n35462), .O(n8231[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3066_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_20061_14_lut (.I0(GND_net), .I1(n63[12]), .I2(n191[12]), 
            .I3(n34291), .O(\PID_CONTROLLER.result_31__N_3003 [12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_20061_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3272_20 (.CI(n34407), .I0(n13594[17]), .I1(GND_net), 
            .CO(n34408));
    SB_CARRY add_20061_14 (.CI(n34291), .I0(n63[12]), .I1(n191[12]), .CO(n34292));
    SB_CARRY unary_minus_21_add_3_7 (.CI(n34138), .I0(GND_net), .I1(n75[5]), 
            .CO(n34139));
    SB_LUT4 unary_minus_21_add_3_6_lut (.I0(GND_net), .I1(GND_net), .I2(n75[4]), 
            .I3(n34137), .O(n70[4])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_21_add_3_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i5_4_lut (.I0(n45714), .I1(pwm[21]), .I2(pwm[8]), .I3(pwm_count[8]), 
            .O(n20_adj_3554));
    defparam i5_4_lut.LUT_INIT = 16'hecfe;
    SB_CARRY add_3279_14 (.CI(n34635), .I0(n13734[11]), .I1(GND_net), 
            .CO(n34636));
    SB_CARRY unary_minus_21_add_3_6 (.CI(n34137), .I0(GND_net), .I1(n75[4]), 
            .CO(n34138));
    SB_LUT4 unary_minus_21_add_3_5_lut (.I0(GND_net), .I1(GND_net), .I2(n75[3]), 
            .I3(n34136), .O(n70[3])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_21_add_3_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_20061_13_lut (.I0(GND_net), .I1(n63[11]), .I2(n191[11]), 
            .I3(n34290), .O(\PID_CONTROLLER.result_31__N_3003 [11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_20061_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1219_22_lut (.I0(GND_net), .I1(n8448[19]), .I2(GND_net), 
            .I3(n35957), .O(n1804[20])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1219_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_21_add_3_5 (.CI(n34136), .I0(GND_net), .I1(n75[3]), 
            .CO(n34137));
    SB_LUT4 add_3077_3_lut (.I0(GND_net), .I1(n8429[0]), .I2(n261_adj_3556), 
            .I3(n35613), .O(n8418[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3077_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1219_22 (.CI(n35957), .I0(n8448[19]), .I1(GND_net), 
            .CO(n35958));
    SB_LUT4 mult_14_add_1219_21_lut (.I0(GND_net), .I1(n8448[18]), .I2(GND_net), 
            .I3(n35956), .O(n1804[19])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1219_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_21_add_3_4_lut (.I0(GND_net), .I1(GND_net), .I2(n75[2]), 
            .I3(n34135), .O(n70[2])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_21_add_3_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3071_7_lut (.I0(GND_net), .I1(n8348[4]), .I2(n631), .I3(n35548), 
            .O(n8331[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3071_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1219_21 (.CI(n35956), .I0(n8448[18]), .I1(GND_net), 
            .CO(n35957));
    SB_LUT4 add_3064_3_lut (.I0(GND_net), .I1(n8208[0]), .I2(n222_adj_3558), 
            .I3(n35418), .O(n8184[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3064_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_20061_13 (.CI(n34290), .I0(n63[11]), .I1(n191[11]), .CO(n34291));
    SB_LUT4 mult_14_add_1219_20_lut (.I0(GND_net), .I1(n8448[17]), .I2(GND_net), 
            .I3(n35955), .O(n1804[18])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1219_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_20061_12_lut (.I0(GND_net), .I1(n63[10]), .I2(n191[10]), 
            .I3(n34289), .O(\PID_CONTROLLER.result_31__N_3003 [10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_20061_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1219_20 (.CI(n35955), .I0(n8448[17]), .I1(GND_net), 
            .CO(n35956));
    SB_LUT4 add_3279_13_lut (.I0(GND_net), .I1(n13734[10]), .I2(GND_net), 
            .I3(n34634), .O(n13256[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3279_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1219_19_lut (.I0(GND_net), .I1(n8448[16]), .I2(GND_net), 
            .I3(n35954), .O(n1804[17])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1219_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1219_19 (.CI(n35954), .I0(n8448[16]), .I1(GND_net), 
            .CO(n35955));
    SB_CARRY add_3071_7 (.CI(n35548), .I0(n8348[4]), .I1(n631), .CO(n35549));
    SB_LUT4 mult_14_add_1219_18_lut (.I0(GND_net), .I1(n8448[15]), .I2(GND_net), 
            .I3(n35953), .O(n1804[16])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1219_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1219_18 (.CI(n35953), .I0(n8448[15]), .I1(GND_net), 
            .CO(n35954));
    SB_LUT4 mult_14_add_1219_17_lut (.I0(GND_net), .I1(n8448[14]), .I2(GND_net), 
            .I3(n35952), .O(n1804[15])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1219_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3068_8 (.CI(n35501), .I0(n8294[5]), .I1(n719), .CO(n35502));
    SB_CARRY mult_14_add_1219_17 (.CI(n35952), .I0(n8448[14]), .I1(GND_net), 
            .CO(n35953));
    SB_LUT4 mult_14_add_1219_16_lut (.I0(GND_net), .I1(n8448[13]), .I2(GND_net), 
            .I3(n35951), .O(n1804[14])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1219_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1219_16 (.CI(n35951), .I0(n8448[13]), .I1(GND_net), 
            .CO(n35952));
    SB_LUT4 mult_14_add_1219_15_lut (.I0(GND_net), .I1(n8448[12]), .I2(GND_net), 
            .I3(n35950), .O(n1804[13])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1219_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1219_15 (.CI(n35950), .I0(n8448[12]), .I1(GND_net), 
            .CO(n35951));
    SB_CARRY add_3066_6 (.CI(n35462), .I0(n8253[3]), .I1(n519_adj_3551), 
            .CO(n35463));
    SB_LUT4 mult_14_add_1219_14_lut (.I0(GND_net), .I1(n8448[11]), .I2(GND_net), 
            .I3(n35949), .O(n1804[12])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1219_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1219_14 (.CI(n35949), .I0(n8448[11]), .I1(GND_net), 
            .CO(n35950));
    SB_LUT4 mult_14_add_1219_13_lut (.I0(GND_net), .I1(n8448[10]), .I2(GND_net), 
            .I3(n35948), .O(n1804[11])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1219_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3064_3 (.CI(n35418), .I0(n8208[0]), .I1(n222_adj_3558), 
            .CO(n35419));
    SB_CARRY mult_14_add_1219_13 (.CI(n35948), .I0(n8448[10]), .I1(GND_net), 
            .CO(n35949));
    SB_LUT4 mult_14_add_1219_12_lut (.I0(GND_net), .I1(n8448[9]), .I2(GND_net), 
            .I3(n35947), .O(n1804[10])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1219_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3060_23_lut (.I0(GND_net), .I1(n8106[20]), .I2(GND_net), 
            .I3(n35344), .O(n8078[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3060_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1219_12 (.CI(n35947), .I0(n8448[9]), .I1(GND_net), 
            .CO(n35948));
    SB_LUT4 mult_14_add_1219_11_lut (.I0(GND_net), .I1(n8448[8]), .I2(GND_net), 
            .I3(n35946), .O(n1804[9])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1219_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i11_4_lut (.I0(pwm[11]), .I1(pwm[17]), .I2(pwm[19]), .I3(pwm[12]), 
            .O(n26_adj_3559));
    defparam i11_4_lut.LUT_INIT = 16'hfffe;
    SB_CARRY add_3060_23 (.CI(n35344), .I0(n8106[20]), .I1(GND_net), .CO(n35345));
    SB_CARRY unary_minus_21_add_3_4 (.CI(n34135), .I0(GND_net), .I1(n75[2]), 
            .CO(n34136));
    SB_CARRY add_20061_12 (.CI(n34289), .I0(n63[10]), .I1(n191[10]), .CO(n34290));
    SB_LUT4 unary_minus_21_add_3_3_lut (.I0(GND_net), .I1(GND_net), .I2(n75[1]), 
            .I3(n34134), .O(n70[1])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_21_add_3_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1219_11 (.CI(n35946), .I0(n8448[8]), .I1(GND_net), 
            .CO(n35947));
    SB_LUT4 add_3064_2_lut (.I0(GND_net), .I1(n32_adj_3562), .I2(n125), 
            .I3(GND_net), .O(n8184[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3064_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1219_10_lut (.I0(GND_net), .I1(n8448[7]), .I2(GND_net), 
            .I3(n35945), .O(n1804[8])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1219_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3060_22_lut (.I0(GND_net), .I1(n8106[19]), .I2(GND_net), 
            .I3(n35343), .O(n8078[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3060_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1219_10 (.CI(n35945), .I0(n8448[7]), .I1(GND_net), 
            .CO(n35946));
    SB_LUT4 add_3121_15_lut (.I0(GND_net), .I1(n10118[12]), .I2(GND_net), 
            .I3(n35206), .O(n9327[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3121_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1219_9_lut (.I0(GND_net), .I1(n8448[6]), .I2(GND_net), 
            .I3(n35944), .O(n1804[7])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1219_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1219_9 (.CI(n35944), .I0(n8448[6]), .I1(GND_net), 
            .CO(n35945));
    SB_CARRY add_3060_22 (.CI(n35343), .I0(n8106[19]), .I1(GND_net), .CO(n35344));
    SB_LUT4 mult_14_add_1219_8_lut (.I0(GND_net), .I1(n8448[5]), .I2(n536), 
            .I3(n35943), .O(n1804[6])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1219_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1219_8 (.CI(n35943), .I0(n8448[5]), .I1(n536), 
            .CO(n35944));
    SB_LUT4 mult_14_add_1219_7_lut (.I0(GND_net), .I1(n8448[4]), .I2(n463_c), 
            .I3(n35942), .O(n1804[5])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1219_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1219_7 (.CI(n35942), .I0(n8448[4]), .I1(n463_c), 
            .CO(n35943));
    SB_LUT4 mult_14_add_1219_6_lut (.I0(GND_net), .I1(n8448[3]), .I2(n390), 
            .I3(n35941), .O(n1804[4])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1219_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3060_21_lut (.I0(GND_net), .I1(n8106[18]), .I2(GND_net), 
            .I3(n35342), .O(n8078[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3060_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3077_3 (.CI(n35613), .I0(n8429[0]), .I1(n261_adj_3556), 
            .CO(n35614));
    SB_CARRY add_3121_15 (.CI(n35206), .I0(n10118[12]), .I1(GND_net), 
            .CO(n35207));
    SB_LUT4 add_3071_6_lut (.I0(GND_net), .I1(n8348[3]), .I2(n534), .I3(n35547), 
            .O(n8331[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3071_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3066_5_lut (.I0(GND_net), .I1(n8253[2]), .I2(n422_adj_3566), 
            .I3(n35461), .O(n8231[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3066_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3077_2_lut (.I0(GND_net), .I1(n71_adj_3567), .I2(n164_adj_3568), 
            .I3(GND_net), .O(n8418[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3077_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3071_6 (.CI(n35547), .I0(n8348[3]), .I1(n534), .CO(n35548));
    SB_CARRY add_3064_2 (.CI(GND_net), .I0(n32_adj_3562), .I1(n125), .CO(n35418));
    SB_CARRY mult_14_add_1219_6 (.CI(n35941), .I0(n8448[3]), .I1(n390), 
            .CO(n35942));
    SB_LUT4 mult_14_add_1219_5_lut (.I0(GND_net), .I1(n8448[2]), .I2(n317), 
            .I3(n35940), .O(n1804[3])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1219_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3060_21 (.CI(n35342), .I0(n8106[18]), .I1(GND_net), .CO(n35343));
    SB_CARRY mult_14_add_1219_5 (.CI(n35940), .I0(n8448[2]), .I1(n317), 
            .CO(n35941));
    SB_CARRY add_3279_13 (.CI(n34634), .I0(n13734[10]), .I1(GND_net), 
            .CO(n34635));
    SB_LUT4 add_20061_11_lut (.I0(GND_net), .I1(n63[9]), .I2(n191[9]), 
            .I3(n34288), .O(\PID_CONTROLLER.result_31__N_3003 [9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_20061_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_21_add_3_3 (.CI(n34134), .I0(GND_net), .I1(n75[1]), 
            .CO(n34135));
    SB_LUT4 unary_minus_21_add_3_2_lut (.I0(GND_net), .I1(GND_net), .I2(n75[0]), 
            .I3(VCC_net), .O(n70[0])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_21_add_3_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1219_4_lut (.I0(GND_net), .I1(n8448[1]), .I2(n244_adj_3571), 
            .I3(n35939), .O(n1804[2])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1219_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_20061_11 (.CI(n34288), .I0(n63[9]), .I1(n191[9]), .CO(n34289));
    SB_CARRY unary_minus_21_add_3_2 (.CI(VCC_net), .I0(GND_net), .I1(n75[0]), 
            .CO(n34134));
    SB_LUT4 unary_minus_5_add_3_25_lut (.I0(GND_net), .I1(GND_net), .I2(n79[23]), 
            .I3(n34133), .O(n76[23])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3121_14_lut (.I0(GND_net), .I1(n10118[11]), .I2(GND_net), 
            .I3(n35205), .O(n9327[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3121_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3279_12_lut (.I0(GND_net), .I1(n13734[9]), .I2(GND_net), 
            .I3(n34633), .O(n13256[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3279_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_20061_10_lut (.I0(GND_net), .I1(n63[8]), .I2(n191[8]), 
            .I3(n34287), .O(\PID_CONTROLLER.result_31__N_3003 [8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_20061_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_5_add_3_24_lut (.I0(\PID_CONTROLLER.integral [9]), 
            .I1(GND_net), .I2(n79[22]), .I3(n34132), .O(n45_adj_3573)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_24_lut.LUT_INIT = 16'h6996;
    SB_CARRY unary_minus_5_add_3_24 (.CI(n34132), .I0(GND_net), .I1(n79[22]), 
            .CO(n34133));
    SB_CARRY add_20061_10 (.CI(n34287), .I0(n63[8]), .I1(n191[8]), .CO(n34288));
    SB_LUT4 unary_minus_5_add_3_23_lut (.I0(\PID_CONTROLLER.integral [9]), 
            .I1(GND_net), .I2(n79[21]), .I3(n34131), .O(n43_adj_3575)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_23_lut.LUT_INIT = 16'h6996;
    SB_CARRY add_3121_14 (.CI(n35205), .I0(n10118[11]), .I1(GND_net), 
            .CO(n35206));
    SB_CARRY unary_minus_5_add_3_23 (.CI(n34131), .I0(GND_net), .I1(n79[21]), 
            .CO(n34132));
    SB_LUT4 add_3060_20_lut (.I0(GND_net), .I1(n8106[17]), .I2(GND_net), 
            .I3(n35341), .O(n8078[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3060_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3063_24_lut (.I0(GND_net), .I1(n8184[21]), .I2(GND_net), 
            .I3(n35417), .O(n8159[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3063_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3060_20 (.CI(n35341), .I0(n8106[17]), .I1(GND_net), .CO(n35342));
    SB_CARRY mult_14_add_1219_4 (.CI(n35939), .I0(n8448[1]), .I1(n244_adj_3571), 
            .CO(n35940));
    SB_LUT4 add_3121_13_lut (.I0(GND_net), .I1(n10118[10]), .I2(GND_net), 
            .I3(n35204), .O(n9327[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3121_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3077_2 (.CI(GND_net), .I0(n71_adj_3567), .I1(n164_adj_3568), 
            .CO(n35613));
    SB_CARRY add_3121_13 (.CI(n35204), .I0(n10118[10]), .I1(GND_net), 
            .CO(n35205));
    SB_LUT4 add_3121_12_lut (.I0(GND_net), .I1(n10118[9]), .I2(GND_net), 
            .I3(n35203), .O(n9327[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3121_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3076_11_lut (.I0(GND_net), .I1(n8418[8]), .I2(GND_net), 
            .I3(n35612), .O(n8406[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3076_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3076_10_lut (.I0(GND_net), .I1(n8418[7]), .I2(GND_net), 
            .I3(n35611), .O(n8406[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3076_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3076_10 (.CI(n35611), .I0(n8418[7]), .I1(GND_net), .CO(n35612));
    SB_LUT4 add_3076_9_lut (.I0(GND_net), .I1(n8418[6]), .I2(GND_net), 
            .I3(n35610), .O(n8406[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3076_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i9_4_lut (.I0(pwm[16]), .I1(pwm[10]), .I2(pwm[14]), .I3(pwm[9]), 
            .O(n24_adj_3577));
    defparam i9_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 mult_14_add_1219_3_lut (.I0(GND_net), .I1(n8448[0]), .I2(n171_adj_3579), 
            .I3(n35938), .O(n1804[1])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1219_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1219_3 (.CI(n35938), .I0(n8448[0]), .I1(n171_adj_3579), 
            .CO(n35939));
    SB_LUT4 mult_14_add_1219_2_lut (.I0(GND_net), .I1(n35), .I2(n98_adj_3580), 
            .I3(GND_net), .O(n1804[0])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1219_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1219_2 (.CI(GND_net), .I0(n35), .I1(n98_adj_3580), 
            .CO(n35938));
    SB_LUT4 mult_14_add_1218_24_lut (.I0(GND_net), .I1(n1804[21]), .I2(GND_net), 
            .I3(n35936), .O(n1803[22])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1218_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1218_24 (.CI(n35936), .I0(n1804[21]), .I1(GND_net), 
            .CO(n1711));
    SB_LUT4 mult_14_add_1218_23_lut (.I0(GND_net), .I1(n1804[20]), .I2(GND_net), 
            .I3(n35935), .O(n1803[21])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1218_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1218_23 (.CI(n35935), .I0(n1804[20]), .I1(GND_net), 
            .CO(n35936));
    SB_LUT4 mult_14_add_1218_22_lut (.I0(GND_net), .I1(n1804[19]), .I2(GND_net), 
            .I3(n35934), .O(n1803[20])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1218_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1218_22 (.CI(n35934), .I0(n1804[19]), .I1(GND_net), 
            .CO(n35935));
    SB_LUT4 mult_14_add_1218_21_lut (.I0(GND_net), .I1(n1804[18]), .I2(GND_net), 
            .I3(n35933), .O(n1803[19])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1218_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1218_21 (.CI(n35933), .I0(n1804[18]), .I1(GND_net), 
            .CO(n35934));
    SB_LUT4 mult_14_add_1218_20_lut (.I0(GND_net), .I1(n1804[17]), .I2(GND_net), 
            .I3(n35932), .O(n1803[18])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1218_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1218_20 (.CI(n35932), .I0(n1804[17]), .I1(GND_net), 
            .CO(n35933));
    SB_LUT4 mult_14_add_1218_19_lut (.I0(GND_net), .I1(n1804[16]), .I2(GND_net), 
            .I3(n35931), .O(n1803[17])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1218_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1218_19 (.CI(n35931), .I0(n1804[16]), .I1(GND_net), 
            .CO(n35932));
    SB_CARRY add_3076_9 (.CI(n35610), .I0(n8418[6]), .I1(GND_net), .CO(n35611));
    SB_LUT4 add_3071_5_lut (.I0(GND_net), .I1(n8348[2]), .I2(n437_adj_3581), 
            .I3(n35546), .O(n8331[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3071_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3076_8_lut (.I0(GND_net), .I1(n8418[5]), .I2(n743_adj_3582), 
            .I3(n35609), .O(n8406[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3076_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3076_8 (.CI(n35609), .I0(n8418[5]), .I1(n743_adj_3582), 
            .CO(n35610));
    SB_CARRY add_3071_5 (.CI(n35546), .I0(n8348[2]), .I1(n437_adj_3581), 
            .CO(n35547));
    SB_LUT4 add_3076_7_lut (.I0(GND_net), .I1(n8418[4]), .I2(n646_adj_3583), 
            .I3(n35608), .O(n8406[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3076_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3076_7 (.CI(n35608), .I0(n8418[4]), .I1(n646_adj_3583), 
            .CO(n35609));
    SB_LUT4 add_3076_6_lut (.I0(GND_net), .I1(n8418[3]), .I2(n549_adj_3584), 
            .I3(n35607), .O(n8406[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3076_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3076_6 (.CI(n35607), .I0(n8418[3]), .I1(n549_adj_3584), 
            .CO(n35608));
    SB_LUT4 add_3076_5_lut (.I0(GND_net), .I1(n8418[2]), .I2(n452_adj_3585), 
            .I3(n35606), .O(n8406[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3076_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3076_5 (.CI(n35606), .I0(n8418[2]), .I1(n452_adj_3585), 
            .CO(n35607));
    SB_LUT4 add_3076_4_lut (.I0(GND_net), .I1(n8418[1]), .I2(n355_adj_3586), 
            .I3(n35605), .O(n8406[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3076_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3076_4 (.CI(n35605), .I0(n8418[1]), .I1(n355_adj_3586), 
            .CO(n35606));
    SB_LUT4 add_3076_3_lut (.I0(GND_net), .I1(n8418[0]), .I2(n258_adj_3587), 
            .I3(n35604), .O(n8406[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3076_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3076_3 (.CI(n35604), .I0(n8418[0]), .I1(n258_adj_3587), 
            .CO(n35605));
    SB_LUT4 add_3076_2_lut (.I0(GND_net), .I1(n68_adj_3588), .I2(n161_adj_3589), 
            .I3(GND_net), .O(n8406[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3076_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3068_7_lut (.I0(GND_net), .I1(n8294[4]), .I2(n622), .I3(n35500), 
            .O(n8274[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3068_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1218_18_lut (.I0(GND_net), .I1(n1804[15]), .I2(GND_net), 
            .I3(n35930), .O(n1803[16])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1218_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1218_18 (.CI(n35930), .I0(n1804[15]), .I1(GND_net), 
            .CO(n35931));
    SB_LUT4 mult_14_add_1218_17_lut (.I0(GND_net), .I1(n1804[14]), .I2(GND_net), 
            .I3(n35929), .O(n1803[15])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1218_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1218_17 (.CI(n35929), .I0(n1804[14]), .I1(GND_net), 
            .CO(n35930));
    SB_LUT4 mult_14_add_1218_16_lut (.I0(GND_net), .I1(n1804[13]), .I2(GND_net), 
            .I3(n35928), .O(n1803[14])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1218_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1218_16 (.CI(n35928), .I0(n1804[13]), .I1(GND_net), 
            .CO(n35929));
    SB_LUT4 mult_14_add_1218_15_lut (.I0(GND_net), .I1(n1804[12]), .I2(GND_net), 
            .I3(n35927), .O(n1803[13])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1218_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1218_15 (.CI(n35927), .I0(n1804[12]), .I1(GND_net), 
            .CO(n35928));
    SB_LUT4 mult_14_add_1218_14_lut (.I0(GND_net), .I1(n1804[11]), .I2(GND_net), 
            .I3(n35926), .O(n1803[12])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1218_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1218_14 (.CI(n35926), .I0(n1804[11]), .I1(GND_net), 
            .CO(n35927));
    SB_LUT4 mult_14_add_1218_13_lut (.I0(GND_net), .I1(n1804[10]), .I2(GND_net), 
            .I3(n35925), .O(n1803[11])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1218_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1218_13 (.CI(n35925), .I0(n1804[10]), .I1(GND_net), 
            .CO(n35926));
    SB_LUT4 mult_14_add_1218_12_lut (.I0(GND_net), .I1(n1804[9]), .I2(GND_net), 
            .I3(n35924), .O(n1803[10])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1218_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1218_12 (.CI(n35924), .I0(n1804[9]), .I1(GND_net), 
            .CO(n35925));
    SB_LUT4 mult_14_add_1218_11_lut (.I0(GND_net), .I1(n1804[8]), .I2(GND_net), 
            .I3(n35923), .O(n1803[9])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1218_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1218_11 (.CI(n35923), .I0(n1804[8]), .I1(GND_net), 
            .CO(n35924));
    SB_LUT4 add_3071_4_lut (.I0(GND_net), .I1(n8348[1]), .I2(n340), .I3(n35545), 
            .O(n8331[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3071_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3071_4 (.CI(n35545), .I0(n8348[1]), .I1(n340), .CO(n35546));
    SB_LUT4 add_3071_3_lut (.I0(GND_net), .I1(n8348[0]), .I2(n243_adj_3590), 
            .I3(n35544), .O(n8331[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3071_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i13_4_lut (.I0(pwm[13]), .I1(n26_adj_3559), .I2(n20_adj_3554), 
            .I3(pwm[22]), .O(n28_adj_3591));
    defparam i13_4_lut.LUT_INIT = 16'hfffe;
    SB_CARRY add_3279_12 (.CI(n34633), .I0(n13734[9]), .I1(GND_net), .CO(n34634));
    SB_LUT4 add_20061_9_lut (.I0(GND_net), .I1(n63[7]), .I2(n191[7]), 
            .I3(n34286), .O(\PID_CONTROLLER.result_31__N_3003 [7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_20061_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_5_add_3_22_lut (.I0(\PID_CONTROLLER.integral [9]), 
            .I1(GND_net), .I2(n79[20]), .I3(n34130), .O(n41_adj_3592)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_22_lut.LUT_INIT = 16'h6996;
    SB_CARRY unary_minus_5_add_3_22 (.CI(n34130), .I0(GND_net), .I1(n79[20]), 
            .CO(n34131));
    SB_CARRY add_20061_9 (.CI(n34286), .I0(n63[7]), .I1(n191[7]), .CO(n34287));
    SB_DFFE \PID_CONTROLLER.integral_1017__i0  (.Q(\PID_CONTROLLER.integral [0]), 
            .C(clk32MHz), .E(n55_adj_3594), .D(n66[0]));   // verilog/motorControl.v(41[21:33])
    SB_LUT4 mult_14_add_1218_10_lut (.I0(GND_net), .I1(n1804[7]), .I2(GND_net), 
            .I3(n35922), .O(n1803[8])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1218_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_i242_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral [9]), 
            .I2(GND_net), .I3(GND_net), .O(n326));   // verilog/motorControl.v(43[48:59])
    defparam mult_14_i242_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i8_3_lut (.I0(pwm[15]), .I1(pwm[18]), .I2(pwm[20]), .I3(GND_net), 
            .O(n23_adj_3596));
    defparam i8_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 unary_minus_5_add_3_21_lut (.I0(\PID_CONTROLLER.integral [9]), 
            .I1(GND_net), .I2(n79[19]), .I3(n34129), .O(n39_adj_3597)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_21_lut.LUT_INIT = 16'h6996;
    SB_LUT4 mult_12_i75_2_lut (.I0(\Kd[1] ), .I1(n57[4]), .I2(GND_net), 
            .I3(GND_net), .O(n110));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i75_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i12_2_lut (.I0(\Kd[0] ), .I1(n57[5]), .I2(GND_net), 
            .I3(GND_net), .O(n17));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i12_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i83_2_lut (.I0(\Kd[1] ), .I1(n57[8]), .I2(GND_net), 
            .I3(GND_net), .O(n122));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i83_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_3071_3 (.CI(n35544), .I0(n8348[0]), .I1(n243_adj_3590), 
            .CO(n35545));
    SB_LUT4 add_3060_19_lut (.I0(GND_net), .I1(n8106[16]), .I2(GND_net), 
            .I3(n35340), .O(n8078[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3060_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3121_12 (.CI(n35203), .I0(n10118[9]), .I1(GND_net), .CO(n35204));
    SB_LUT4 add_3121_11_lut (.I0(GND_net), .I1(n10118[8]), .I2(GND_net), 
            .I3(n35202), .O(n9327[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3121_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3071_2_lut (.I0(GND_net), .I1(n53_adj_3599), .I2(n146_adj_3600), 
            .I3(GND_net), .O(n8331[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3071_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3068_7 (.CI(n35500), .I0(n8294[4]), .I1(n622), .CO(n35501));
    SB_CARRY add_3066_5 (.CI(n35461), .I0(n8253[2]), .I1(n422_adj_3566), 
            .CO(n35462));
    SB_LUT4 add_3063_23_lut (.I0(GND_net), .I1(n8184[20]), .I2(GND_net), 
            .I3(n35416), .O(n8159[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3063_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3060_19 (.CI(n35340), .I0(n8106[16]), .I1(GND_net), .CO(n35341));
    SB_CARRY add_3121_11 (.CI(n35202), .I0(n10118[8]), .I1(GND_net), .CO(n35203));
    SB_LUT4 add_3068_6_lut (.I0(GND_net), .I1(n8294[3]), .I2(n525), .I3(n35499), 
            .O(n8274[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3068_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3121_10_lut (.I0(GND_net), .I1(n10118[7]), .I2(GND_net), 
            .I3(n35201), .O(n9327[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3121_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_4_lut (.I0(pwm[23]), .I1(n23_adj_3596), .I2(n28_adj_3591), 
            .I3(n24_adj_3577), .O(n17_adj_3456));   // verilog/motorControl.v(65[9:32])
    defparam i1_4_lut.LUT_INIT = 16'haaab;
    SB_CARRY unary_minus_5_add_3_21 (.CI(n34129), .I0(GND_net), .I1(n79[19]), 
            .CO(n34130));
    SB_LUT4 i25457_2_lut (.I0(hall2), .I1(hall3), .I2(GND_net), .I3(GND_net), 
            .O(n40975));
    defparam i25457_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 add_3279_11_lut (.I0(GND_net), .I1(n13734[8]), .I2(GND_net), 
            .I3(n34632), .O(n13256[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3279_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3060_18_lut (.I0(GND_net), .I1(n8106[15]), .I2(GND_net), 
            .I3(n35339), .O(n8078[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3060_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i29338_3_lut (.I0(n40121), .I1(hall1), .I2(hall2), .I3(GND_net), 
            .O(n44158));   // verilog/motorControl.v(86[14] 109[8])
    defparam i29338_3_lut.LUT_INIT = 16'h8080;
    SB_CARRY add_3121_10 (.CI(n35201), .I0(n10118[7]), .I1(GND_net), .CO(n35202));
    SB_LUT4 unary_minus_5_add_3_20_lut (.I0(\PID_CONTROLLER.integral [9]), 
            .I1(GND_net), .I2(n79[18]), .I3(n34128), .O(n37_adj_3601)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_20_lut.LUT_INIT = 16'h6996;
    SB_CARRY add_3063_23 (.CI(n35416), .I0(n8184[20]), .I1(GND_net), .CO(n35417));
    SB_LUT4 add_20061_8_lut (.I0(GND_net), .I1(n63[6]), .I2(n191[6]), 
            .I3(n34285), .O(\PID_CONTROLLER.result_31__N_3003 [6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_20061_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3060_18 (.CI(n35339), .I0(n8106[15]), .I1(GND_net), .CO(n35340));
    SB_LUT4 i34_4_lut (.I0(n44158), .I1(n40975), .I2(n17_adj_3456), .I3(n40176), 
            .O(n18_adj_3603));   // verilog/motorControl.v(86[14] 109[8])
    defparam i34_4_lut.LUT_INIT = 16'ha3a0;
    SB_LUT4 add_3121_9_lut (.I0(GND_net), .I1(n10118[6]), .I2(GND_net), 
            .I3(n35200), .O(n9327[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3121_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3121_9 (.CI(n35200), .I0(n10118[6]), .I1(GND_net), .CO(n35201));
    SB_CARRY add_3279_11 (.CI(n34632), .I0(n13734[8]), .I1(GND_net), .CO(n34633));
    SB_CARRY add_20061_8 (.CI(n34285), .I0(n63[6]), .I1(n191[6]), .CO(n34286));
    SB_LUT4 add_20061_7_lut (.I0(GND_net), .I1(n63[5]), .I2(n191[5]), 
            .I3(n34284), .O(\PID_CONTROLLER.result_31__N_3003 [5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_20061_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_5_add_3_20 (.CI(n34128), .I0(GND_net), .I1(n79[18]), 
            .CO(n34129));
    SB_LUT4 add_3063_22_lut (.I0(GND_net), .I1(n8184[19]), .I2(GND_net), 
            .I3(n35415), .O(n8159[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3063_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_20061_7 (.CI(n34284), .I0(n63[5]), .I1(n191[5]), .CO(n34285));
    SB_LUT4 add_3060_17_lut (.I0(GND_net), .I1(n8106[14]), .I2(GND_net), 
            .I3(n35338), .O(n8078[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3060_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_5_add_3_19_lut (.I0(\PID_CONTROLLER.integral [9]), 
            .I1(GND_net), .I2(n79[17]), .I3(n34127), .O(n35_adj_3604)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_19_lut.LUT_INIT = 16'h6996;
    SB_CARRY mult_14_add_1218_10 (.CI(n35922), .I0(n1804[7]), .I1(GND_net), 
            .CO(n35923));
    SB_LUT4 add_3121_8_lut (.I0(GND_net), .I1(n10118[5]), .I2(n545), .I3(n35199), 
            .O(n9327[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3121_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3279_10_lut (.I0(GND_net), .I1(n13734[7]), .I2(GND_net), 
            .I3(n34631), .O(n13256[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3279_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1218_9_lut (.I0(GND_net), .I1(n1804[6]), .I2(GND_net), 
            .I3(n35921), .O(n1803[7])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1218_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3279_10 (.CI(n34631), .I0(n13734[7]), .I1(GND_net), .CO(n34632));
    SB_LUT4 add_20061_6_lut (.I0(GND_net), .I1(n63[4]), .I2(n191[4]), 
            .I3(n34283), .O(\PID_CONTROLLER.result_31__N_3003 [4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_20061_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1218_9 (.CI(n35921), .I0(n1804[6]), .I1(GND_net), 
            .CO(n35922));
    SB_LUT4 i33_4_lut (.I0(n18_adj_3603), .I1(n17_adj_3456), .I2(GATES_5__N_3048[5]), 
            .I3(n40121), .O(GATES_5__N_2788[1]));   // verilog/motorControl.v(86[14] 109[8])
    defparam i33_4_lut.LUT_INIT = 16'hca0a;
    SB_CARRY unary_minus_5_add_3_19 (.CI(n34127), .I0(GND_net), .I1(n79[17]), 
            .CO(n34128));
    SB_LUT4 mult_14_add_1218_8_lut (.I0(GND_net), .I1(n1804[5]), .I2(n533), 
            .I3(n35920), .O(n1803[6])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1218_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3121_8 (.CI(n35199), .I0(n10118[5]), .I1(n545), .CO(n35200));
    SB_CARRY add_20061_6 (.CI(n34283), .I0(n63[4]), .I1(n191[4]), .CO(n34284));
    SB_LUT4 add_20061_5_lut (.I0(GND_net), .I1(n63[3]), .I2(n191[3]), 
            .I3(n34282), .O(\PID_CONTROLLER.result_31__N_3003 [3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_20061_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1218_8 (.CI(n35920), .I0(n1804[5]), .I1(n533), 
            .CO(n35921));
    SB_LUT4 unary_minus_5_add_3_18_lut (.I0(\PID_CONTROLLER.integral [9]), 
            .I1(GND_net), .I2(n79[16]), .I3(n34126), .O(n33_adj_3608)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_18_lut.LUT_INIT = 16'h6996;
    SB_LUT4 add_3121_7_lut (.I0(GND_net), .I1(n10118[4]), .I2(n472), .I3(n35198), 
            .O(n9327[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3121_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3060_17 (.CI(n35338), .I0(n8106[14]), .I1(GND_net), .CO(n35339));
    SB_CARRY add_3121_7 (.CI(n35198), .I0(n10118[4]), .I1(n472), .CO(n35199));
    SB_LUT4 add_3121_6_lut (.I0(GND_net), .I1(n10118[3]), .I2(n399), .I3(n35197), 
            .O(n9327[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3121_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3279_9_lut (.I0(GND_net), .I1(n13734[6]), .I2(GND_net), 
            .I3(n34630), .O(n13256[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3279_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_5_add_3_18 (.CI(n34126), .I0(GND_net), .I1(n79[16]), 
            .CO(n34127));
    SB_LUT4 mult_14_add_1218_7_lut (.I0(GND_net), .I1(n1804[4]), .I2(n460_c), 
            .I3(n35919), .O(n1803[5])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1218_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_20061_5 (.CI(n34282), .I0(n63[3]), .I1(n191[3]), .CO(n34283));
    SB_CARRY mult_14_add_1218_7 (.CI(n35919), .I0(n1804[4]), .I1(n460_c), 
            .CO(n35920));
    SB_CARRY add_3121_6 (.CI(n35197), .I0(n10118[3]), .I1(n399), .CO(n35198));
    SB_LUT4 unary_minus_5_add_3_17_lut (.I0(\PID_CONTROLLER.integral [9]), 
            .I1(GND_net), .I2(n79[15]), .I3(n34125), .O(n31_adj_3611)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_17_lut.LUT_INIT = 16'h6996;
    SB_LUT4 add_20061_4_lut (.I0(GND_net), .I1(n63[2]), .I2(n191[2]), 
            .I3(n34281), .O(\PID_CONTROLLER.result_31__N_3003 [2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_20061_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1218_6_lut (.I0(GND_net), .I1(n1804[3]), .I2(n387_c), 
            .I3(n35918), .O(n1803[4])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1218_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3121_5_lut (.I0(GND_net), .I1(n10118[2]), .I2(n326), .I3(n35196), 
            .O(n9327[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3121_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3068_6 (.CI(n35499), .I0(n8294[3]), .I1(n525), .CO(n35500));
    SB_CARRY mult_14_add_1218_6 (.CI(n35918), .I0(n1804[3]), .I1(n387_c), 
            .CO(n35919));
    SB_LUT4 add_3068_5_lut (.I0(GND_net), .I1(n8294[2]), .I2(n428), .I3(n35498), 
            .O(n8274[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3068_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3066_4_lut (.I0(GND_net), .I1(n8253[1]), .I2(n325_adj_3613), 
            .I3(n35460), .O(n8231[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3066_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i276_2_lut (.I0(\Kp[4] ), .I1(\PID_CONTROLLER.err[7] ), 
            .I2(GND_net), .I3(GND_net), .O(n410_adj_3422));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i276_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_14_add_1218_5_lut (.I0(GND_net), .I1(n1804[2]), .I2(n314_adj_3615), 
            .I3(n35917), .O(n1803[3])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1218_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1218_5 (.CI(n35917), .I0(n1804[2]), .I1(n314_adj_3615), 
            .CO(n35918));
    SB_CARRY add_3063_22 (.CI(n35415), .I0(n8184[19]), .I1(GND_net), .CO(n35416));
    SB_CARRY add_3121_5 (.CI(n35196), .I0(n10118[2]), .I1(n326), .CO(n35197));
    SB_LUT4 add_3060_16_lut (.I0(GND_net), .I1(n8106[13]), .I2(GND_net), 
            .I3(n35337), .O(n8078[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3060_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1218_4_lut (.I0(GND_net), .I1(n1804[1]), .I2(n241_adj_3617), 
            .I3(n35916), .O(n1803[2])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1218_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3121_4_lut (.I0(GND_net), .I1(n10118[1]), .I2(n253), .I3(n35195), 
            .O(n9327[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3121_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3121_4 (.CI(n35195), .I0(n10118[1]), .I1(n253), .CO(n35196));
    SB_CARRY mult_14_add_1218_4 (.CI(n35916), .I0(n1804[1]), .I1(n241_adj_3617), 
            .CO(n35917));
    SB_LUT4 add_3121_3_lut (.I0(GND_net), .I1(n10118[0]), .I2(n180), .I3(n35194), 
            .O(n9327[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3121_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1218_3_lut (.I0(GND_net), .I1(n1804[0]), .I2(n168_adj_3619), 
            .I3(n35915), .O(n1803[1])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1218_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_20061_4 (.CI(n34281), .I0(n63[2]), .I1(n191[2]), .CO(n34282));
    SB_CARRY add_3121_3 (.CI(n35194), .I0(n10118[0]), .I1(n180), .CO(n35195));
    SB_CARRY mult_14_add_1218_3 (.CI(n35915), .I0(n1804[0]), .I1(n168_adj_3619), 
            .CO(n35916));
    SB_LUT4 mult_14_add_1218_2_lut (.I0(GND_net), .I1(n26_adj_3620), .I2(n95), 
            .I3(GND_net), .O(n1803[0])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1218_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3076_2 (.CI(GND_net), .I0(n68_adj_3588), .I1(n161_adj_3589), 
            .CO(n35604));
    SB_LUT4 add_3075_12_lut (.I0(GND_net), .I1(n8406[9]), .I2(GND_net), 
            .I3(n35603), .O(n8393[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3075_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_5_add_3_17 (.CI(n34125), .I0(GND_net), .I1(n79[15]), 
            .CO(n34126));
    SB_CARRY mult_14_add_1218_2 (.CI(GND_net), .I0(n26_adj_3620), .I1(n95), 
            .CO(n35915));
    SB_LUT4 add_3075_11_lut (.I0(GND_net), .I1(n8406[8]), .I2(GND_net), 
            .I3(n35602), .O(n8393[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3075_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1217_24_lut (.I0(GND_net), .I1(n1803[21]), .I2(GND_net), 
            .I3(n35913), .O(n1802[22])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1217_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3279_9 (.CI(n34630), .I0(n13734[6]), .I1(GND_net), .CO(n34631));
    SB_CARRY add_3075_11 (.CI(n35602), .I0(n8406[8]), .I1(GND_net), .CO(n35603));
    SB_CARRY mult_14_add_1217_24 (.CI(n35913), .I0(n1803[21]), .I1(GND_net), 
            .CO(n1707));
    SB_LUT4 add_3075_10_lut (.I0(GND_net), .I1(n8406[7]), .I2(GND_net), 
            .I3(n35601), .O(n8393[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3075_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3075_10 (.CI(n35601), .I0(n8406[7]), .I1(GND_net), .CO(n35602));
    SB_LUT4 add_3279_8_lut (.I0(GND_net), .I1(n13734[5]), .I2(n545), .I3(n34629), 
            .O(n13256[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3279_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i109_2_lut (.I0(\Kp[1] ), .I1(\PID_CONTROLLER.err[21] ), 
            .I2(GND_net), .I3(GND_net), .O(n161));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i109_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_3279_8 (.CI(n34629), .I0(n13734[5]), .I1(n545), .CO(n34630));
    SB_LUT4 add_20061_3_lut (.I0(GND_net), .I1(n63[1]), .I2(n191[1]), 
            .I3(n34280), .O(\PID_CONTROLLER.result_31__N_3003 [1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_20061_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3075_9_lut (.I0(GND_net), .I1(n8406[6]), .I2(GND_net), 
            .I3(n35600), .O(n8393[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3075_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i46_2_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err[22] ), 
            .I2(GND_net), .I3(GND_net), .O(n68));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i46_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_3071_2 (.CI(GND_net), .I0(n53_adj_3599), .I1(n146_adj_3600), 
            .CO(n35544));
    SB_CARRY add_20061_3 (.CI(n34280), .I0(n63[1]), .I1(n191[1]), .CO(n34281));
    SB_LUT4 mult_14_add_1217_23_lut (.I0(GND_net), .I1(n1803[20]), .I2(GND_net), 
            .I3(n35912), .O(n1802[21])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1217_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_5_add_3_16_lut (.I0(\PID_CONTROLLER.integral [9]), 
            .I1(GND_net), .I2(n79[14]), .I3(n34124), .O(n29_adj_3621)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_16_lut.LUT_INIT = 16'h6996;
    SB_CARRY add_3075_9 (.CI(n35600), .I0(n8406[6]), .I1(GND_net), .CO(n35601));
    SB_LUT4 add_3070_17_lut (.I0(GND_net), .I1(n8331[14]), .I2(GND_net), 
            .I3(n35543), .O(n8313[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3070_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_20061_2_lut (.I0(GND_net), .I1(n63[0]), .I2(n191[0]), 
            .I3(GND_net), .O(\PID_CONTROLLER.result_31__N_3003 [0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_20061_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3068_5 (.CI(n35498), .I0(n8294[2]), .I1(n428), .CO(n35499));
    SB_LUT4 add_3070_16_lut (.I0(GND_net), .I1(n8331[13]), .I2(GND_net), 
            .I3(n35542), .O(n8313[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3070_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_20061_2 (.CI(GND_net), .I0(n63[0]), .I1(n191[0]), .CO(n34280));
    SB_CARRY add_3066_4 (.CI(n35460), .I0(n8253[1]), .I1(n325_adj_3613), 
            .CO(n35461));
    SB_LUT4 add_3063_21_lut (.I0(GND_net), .I1(n8184[18]), .I2(GND_net), 
            .I3(n35414), .O(n8159[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3063_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3060_16 (.CI(n35337), .I0(n8106[13]), .I1(GND_net), .CO(n35338));
    SB_LUT4 add_3279_7_lut (.I0(GND_net), .I1(n13734[4]), .I2(n472), .I3(n34628), 
            .O(n13256[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3279_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_5_add_3_16 (.CI(n34124), .I0(GND_net), .I1(n79[14]), 
            .CO(n34125));
    SB_LUT4 add_3121_2_lut (.I0(GND_net), .I1(n35), .I2(n107), .I3(GND_net), 
            .O(n9327[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3121_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_5_add_3_15_lut (.I0(\PID_CONTROLLER.integral [9]), 
            .I1(GND_net), .I2(n79[13]), .I3(n34123), .O(n27_adj_3623)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_15_lut.LUT_INIT = 16'h6996;
    SB_CARRY add_3279_7 (.CI(n34628), .I0(n13734[4]), .I1(n472), .CO(n34629));
    SB_LUT4 add_3354_19_lut (.I0(GND_net), .I1(n15114[16]), .I2(GND_net), 
            .I3(n34279), .O(n14793[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3354_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3121_2 (.CI(GND_net), .I0(n35), .I1(n107), .CO(n35194));
    SB_LUT4 mult_10_i341_2_lut (.I0(\Kp[5] ), .I1(\PID_CONTROLLER.err[7] ), 
            .I2(GND_net), .I3(GND_net), .O(n507_adj_3421));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i341_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_3354_18_lut (.I0(GND_net), .I1(n15114[15]), .I2(GND_net), 
            .I3(n34278), .O(n14793[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3354_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3354_18 (.CI(n34278), .I0(n15114[15]), .I1(GND_net), 
            .CO(n34279));
    SB_CARRY unary_minus_5_add_3_15 (.CI(n34123), .I0(GND_net), .I1(n79[13]), 
            .CO(n34124));
    SB_LUT4 add_3060_15_lut (.I0(GND_net), .I1(n8106[12]), .I2(GND_net), 
            .I3(n35336), .O(n8078[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3060_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3120_7_lut (.I0(GND_net), .I1(n41372), .I2(n658), .I3(n35193), 
            .O(n9319[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3120_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3354_17_lut (.I0(GND_net), .I1(n15114[14]), .I2(GND_net), 
            .I3(n34277), .O(n14793[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3354_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3068_4_lut (.I0(GND_net), .I1(n8294[1]), .I2(n331), .I3(n35497), 
            .O(n8274[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3068_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1217_23 (.CI(n35912), .I0(n1803[20]), .I1(GND_net), 
            .CO(n35913));
    SB_CARRY add_3060_15 (.CI(n35336), .I0(n8106[12]), .I1(GND_net), .CO(n35337));
    SB_LUT4 add_3060_14_lut (.I0(GND_net), .I1(n8106[11]), .I2(GND_net), 
            .I3(n35335), .O(n8078[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3060_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3120_6_lut (.I0(GND_net), .I1(n10111[3]), .I2(n564), .I3(n35192), 
            .O(n9319[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3120_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3120_6 (.CI(n35192), .I0(n10111[3]), .I1(n564), .CO(n35193));
    SB_LUT4 add_3075_8_lut (.I0(GND_net), .I1(n8406[5]), .I2(n740_adj_3625), 
            .I3(n35599), .O(n8393[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3075_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1217_22_lut (.I0(GND_net), .I1(n1803[19]), .I2(GND_net), 
            .I3(n35911), .O(n1802[20])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1217_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3075_8 (.CI(n35599), .I0(n8406[5]), .I1(n740_adj_3625), 
            .CO(n35600));
    SB_LUT4 add_3066_3_lut (.I0(GND_net), .I1(n8253[0]), .I2(n228_adj_3626), 
            .I3(n35459), .O(n8231[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3066_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3066_3 (.CI(n35459), .I0(n8253[0]), .I1(n228_adj_3626), 
            .CO(n35460));
    SB_CARRY add_3070_16 (.CI(n35542), .I0(n8331[13]), .I1(GND_net), .CO(n35543));
    SB_LUT4 add_3075_7_lut (.I0(GND_net), .I1(n8406[4]), .I2(n643_adj_3627), 
            .I3(n35598), .O(n8393[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3075_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3063_21 (.CI(n35414), .I0(n8184[18]), .I1(GND_net), .CO(n35415));
    SB_CARRY add_3060_14 (.CI(n35335), .I0(n8106[11]), .I1(GND_net), .CO(n35336));
    SB_LUT4 add_3120_5_lut (.I0(GND_net), .I1(n10111[2]), .I2(n464_adj_3628), 
            .I3(n35191), .O(n9319[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3120_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_5_add_3_14_lut (.I0(\PID_CONTROLLER.integral [9]), 
            .I1(GND_net), .I2(n79[12]), .I3(n34122), .O(n25_adj_3629)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_14_lut.LUT_INIT = 16'h6996;
    SB_CARRY add_3354_17 (.CI(n34277), .I0(n15114[14]), .I1(GND_net), 
            .CO(n34278));
    SB_CARRY unary_minus_5_add_3_14 (.CI(n34122), .I0(GND_net), .I1(n79[12]), 
            .CO(n34123));
    SB_LUT4 unary_minus_5_add_3_13_lut (.I0(\PID_CONTROLLER.integral [9]), 
            .I1(GND_net), .I2(n79[11]), .I3(n34121), .O(n23_adj_3631)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_13_lut.LUT_INIT = 16'h6996;
    SB_LUT4 add_3354_16_lut (.I0(GND_net), .I1(n15114[13]), .I2(GND_net), 
            .I3(n34276), .O(n14793[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3354_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3120_5 (.CI(n35191), .I0(n10111[2]), .I1(n464_adj_3628), 
            .CO(n35192));
    SB_LUT4 add_3279_6_lut (.I0(GND_net), .I1(n13734[3]), .I2(n399), .I3(n34627), 
            .O(n13256[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3279_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3075_7 (.CI(n35598), .I0(n8406[4]), .I1(n643_adj_3627), 
            .CO(n35599));
    SB_CARRY add_3354_16 (.CI(n34276), .I0(n15114[13]), .I1(GND_net), 
            .CO(n34277));
    SB_LUT4 add_3070_15_lut (.I0(GND_net), .I1(n8331[12]), .I2(GND_net), 
            .I3(n35541), .O(n8313[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3070_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_5_add_3_13 (.CI(n34121), .I0(GND_net), .I1(n79[11]), 
            .CO(n34122));
    SB_LUT4 unary_minus_5_add_3_12_lut (.I0(\PID_CONTROLLER.integral [9]), 
            .I1(GND_net), .I2(n79[10]), .I3(n34120), .O(n21_adj_3633)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_12_lut.LUT_INIT = 16'h6996;
    SB_LUT4 add_3060_13_lut (.I0(GND_net), .I1(n8106[10]), .I2(GND_net), 
            .I3(n35334), .O(n8078[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3060_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_5_add_3_12 (.CI(n34120), .I0(GND_net), .I1(n79[10]), 
            .CO(n34121));
    SB_LUT4 add_3120_4_lut (.I0(GND_net), .I1(n10111[1]), .I2(n370), .I3(n35190), 
            .O(n9319[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3120_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3075_6_lut (.I0(GND_net), .I1(n8406[3]), .I2(n546_adj_3635), 
            .I3(n35597), .O(n8393[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3075_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3120_4 (.CI(n35190), .I0(n10111[1]), .I1(n370), .CO(n35191));
    SB_CARRY add_3279_6 (.CI(n34627), .I0(n13734[3]), .I1(n399), .CO(n34628));
    SB_LUT4 add_3354_15_lut (.I0(GND_net), .I1(n15114[12]), .I2(GND_net), 
            .I3(n34275), .O(n14793[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3354_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_5_add_3_11_lut (.I0(\PID_CONTROLLER.integral [9]), 
            .I1(GND_net), .I2(n79[9]), .I3(n34119), .O(n19_adj_3636)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_11_lut.LUT_INIT = 16'h6996;
    SB_LUT4 add_3120_3_lut (.I0(GND_net), .I1(n10111[0]), .I2(n276), .I3(n35189), 
            .O(n9319[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3120_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_5_add_3_11 (.CI(n34119), .I0(GND_net), .I1(n79[9]), 
            .CO(n34120));
    SB_CARRY add_3354_15 (.CI(n34275), .I0(n15114[12]), .I1(GND_net), 
            .CO(n34276));
    SB_LUT4 add_3063_20_lut (.I0(GND_net), .I1(n8184[17]), .I2(GND_net), 
            .I3(n35413), .O(n8159[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3063_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_5_add_3_10_lut (.I0(\PID_CONTROLLER.integral [8]), 
            .I1(GND_net), .I2(n79[8]), .I3(n34118), .O(n17_adj_3638)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_10_lut.LUT_INIT = 16'h6996;
    SB_CARRY unary_minus_5_add_3_10 (.CI(n34118), .I0(GND_net), .I1(n79[8]), 
            .CO(n34119));
    SB_CARRY add_3060_13 (.CI(n35334), .I0(n8106[10]), .I1(GND_net), .CO(n35335));
    SB_LUT4 add_3060_12_lut (.I0(GND_net), .I1(n8106[9]), .I2(GND_net), 
            .I3(n35333), .O(n8078[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3060_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3120_3 (.CI(n35189), .I0(n10111[0]), .I1(n276), .CO(n35190));
    SB_LUT4 add_3120_2_lut (.I0(GND_net), .I1(n86), .I2(n182_adj_3640), 
            .I3(GND_net), .O(n9319[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3120_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3120_2 (.CI(GND_net), .I0(n86), .I1(n182_adj_3640), .CO(n35189));
    SB_CARRY add_3068_4 (.CI(n35497), .I0(n8294[1]), .I1(n331), .CO(n35498));
    SB_LUT4 add_3066_2_lut (.I0(GND_net), .I1(n38_adj_3641), .I2(n131_adj_3642), 
            .I3(GND_net), .O(n8231[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3066_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3063_20 (.CI(n35413), .I0(n8184[17]), .I1(GND_net), .CO(n35414));
    SB_LUT4 add_3150_20_lut (.I0(GND_net), .I1(n10852[17]), .I2(GND_net), 
            .I3(n35188), .O(n10118[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3150_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3060_12 (.CI(n35333), .I0(n8106[9]), .I1(GND_net), .CO(n35334));
    SB_LUT4 add_3150_19_lut (.I0(GND_net), .I1(n10852[16]), .I2(GND_net), 
            .I3(n35187), .O(n10118[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3150_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3150_19 (.CI(n35187), .I0(n10852[16]), .I1(GND_net), 
            .CO(n35188));
    SB_LUT4 mult_12_i276_2_lut (.I0(\Kd[4] ), .I1(n57[7]), .I2(GND_net), 
            .I3(GND_net), .O(n410));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i276_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_3060_11_lut (.I0(GND_net), .I1(n8106[8]), .I2(GND_net), 
            .I3(n35332), .O(n8078[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3060_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3150_18_lut (.I0(GND_net), .I1(n10852[15]), .I2(GND_net), 
            .I3(n35186), .O(n10118[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3150_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3060_11 (.CI(n35332), .I0(n8106[8]), .I1(GND_net), .CO(n35333));
    SB_CARRY add_3150_18 (.CI(n35186), .I0(n10852[15]), .I1(GND_net), 
            .CO(n35187));
    SB_CARRY add_3075_6 (.CI(n35597), .I0(n8406[3]), .I1(n546_adj_3635), 
            .CO(n35598));
    SB_CARRY mult_14_add_1217_22 (.CI(n35911), .I0(n1803[19]), .I1(GND_net), 
            .CO(n35912));
    SB_LUT4 sub_11_inv_0_i12_1_lut (.I0(\PID_CONTROLLER.err[11] ), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n64[11]));   // verilog/motorControl.v(43[31:45])
    defparam sub_11_inv_0_i12_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_14_add_1217_21_lut (.I0(GND_net), .I1(n1803[18]), .I2(GND_net), 
            .I3(n35910), .O(n1802[19])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1217_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3068_3_lut (.I0(GND_net), .I1(n8294[0]), .I2(n234_adj_3643), 
            .I3(n35496), .O(n8274[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3068_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1217_21 (.CI(n35910), .I0(n1803[18]), .I1(GND_net), 
            .CO(n35911));
    SB_LUT4 mult_14_add_1217_20_lut (.I0(GND_net), .I1(n1803[17]), .I2(GND_net), 
            .I3(n35909), .O(n1802[18])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1217_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1217_20 (.CI(n35909), .I0(n1803[17]), .I1(GND_net), 
            .CO(n35910));
    SB_CARRY add_3068_3 (.CI(n35496), .I0(n8294[0]), .I1(n234_adj_3643), 
            .CO(n35497));
    SB_LUT4 mult_14_add_1217_19_lut (.I0(GND_net), .I1(n1803[16]), .I2(GND_net), 
            .I3(n35908), .O(n1802[17])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1217_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1217_19 (.CI(n35908), .I0(n1803[16]), .I1(GND_net), 
            .CO(n35909));
    SB_LUT4 mult_14_add_1217_18_lut (.I0(GND_net), .I1(n1803[15]), .I2(GND_net), 
            .I3(n35907), .O(n1802[16])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1217_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3279_5_lut (.I0(GND_net), .I1(n13734[2]), .I2(n326), .I3(n34626), 
            .O(n13256[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3279_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3354_14_lut (.I0(GND_net), .I1(n15114[11]), .I2(GND_net), 
            .I3(n34274), .O(n14793[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3354_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_5_add_3_9_lut (.I0(\PID_CONTROLLER.integral [7]), 
            .I1(GND_net), .I2(n79[7]), .I3(n34117), .O(n15_adj_3644)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_9_lut.LUT_INIT = 16'h6996;
    SB_CARRY add_3354_14 (.CI(n34274), .I0(n15114[11]), .I1(GND_net), 
            .CO(n34275));
    SB_CARRY unary_minus_5_add_3_9 (.CI(n34117), .I0(GND_net), .I1(n79[7]), 
            .CO(n34118));
    SB_LUT4 add_3150_17_lut (.I0(GND_net), .I1(n10852[14]), .I2(GND_net), 
            .I3(n35185), .O(n10118[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3150_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3070_15 (.CI(n35541), .I0(n8331[12]), .I1(GND_net), .CO(n35542));
    SB_CARRY mult_14_add_1217_18 (.CI(n35907), .I0(n1803[15]), .I1(GND_net), 
            .CO(n35908));
    SB_LUT4 unary_minus_5_add_3_8_lut (.I0(\PID_CONTROLLER.integral [6]), 
            .I1(GND_net), .I2(n79[6]), .I3(n34116), .O(n13_adj_3646)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_8_lut.LUT_INIT = 16'h6996;
    SB_LUT4 mult_14_add_1217_17_lut (.I0(GND_net), .I1(n1803[14]), .I2(GND_net), 
            .I3(n35906), .O(n1802[15])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1217_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3279_5 (.CI(n34626), .I0(n13734[2]), .I1(n326), .CO(n34627));
    SB_LUT4 add_3354_13_lut (.I0(GND_net), .I1(n15114[10]), .I2(GND_net), 
            .I3(n34273), .O(n14793[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3354_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_5_add_3_8 (.CI(n34116), .I0(GND_net), .I1(n79[6]), 
            .CO(n34117));
    SB_CARRY add_3354_13 (.CI(n34273), .I0(n15114[10]), .I1(GND_net), 
            .CO(n34274));
    SB_LUT4 unary_minus_5_add_3_7_lut (.I0(\PID_CONTROLLER.integral [5]), 
            .I1(GND_net), .I2(n79[5]), .I3(n34115), .O(n11_adj_3648)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_7_lut.LUT_INIT = 16'h6996;
    SB_CARRY mult_14_add_1217_17 (.CI(n35906), .I0(n1803[14]), .I1(GND_net), 
            .CO(n35907));
    SB_LUT4 mult_14_add_1217_16_lut (.I0(GND_net), .I1(n1803[13]), .I2(GND_net), 
            .I3(n35905), .O(n1802[14])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1217_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3150_17 (.CI(n35185), .I0(n10852[14]), .I1(GND_net), 
            .CO(n35186));
    SB_LUT4 add_3279_4_lut (.I0(GND_net), .I1(n13734[1]), .I2(n253), .I3(n34625), 
            .O(n13256[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3279_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3354_12_lut (.I0(GND_net), .I1(n15114[9]), .I2(GND_net), 
            .I3(n34272), .O(n14793[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3354_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_5_add_3_7 (.CI(n34115), .I0(GND_net), .I1(n79[5]), 
            .CO(n34116));
    SB_LUT4 unary_minus_5_add_3_6_lut (.I0(\PID_CONTROLLER.integral [4]), 
            .I1(GND_net), .I2(n79[4]), .I3(n34114), .O(n9_adj_3650)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_6_lut.LUT_INIT = 16'h6996;
    SB_CARRY add_3354_12 (.CI(n34272), .I0(n15114[9]), .I1(GND_net), .CO(n34273));
    SB_CARRY unary_minus_5_add_3_6 (.CI(n34114), .I0(GND_net), .I1(n79[4]), 
            .CO(n34115));
    SB_LUT4 unary_minus_5_add_3_5_lut (.I0(\PID_CONTROLLER.integral [3]), 
            .I1(GND_net), .I2(n79[3]), .I3(n34113), .O(n7_adj_3652)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_5_lut.LUT_INIT = 16'h6996;
    SB_CARRY mult_14_add_1217_16 (.CI(n35905), .I0(n1803[13]), .I1(GND_net), 
            .CO(n35906));
    SB_CARRY add_3279_4 (.CI(n34625), .I0(n13734[1]), .I1(n253), .CO(n34626));
    SB_LUT4 add_3354_11_lut (.I0(GND_net), .I1(n15114[8]), .I2(GND_net), 
            .I3(n34271), .O(n14793[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3354_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_5_add_3_5 (.CI(n34113), .I0(GND_net), .I1(n79[3]), 
            .CO(n34114));
    SB_LUT4 unary_minus_5_add_3_4_lut (.I0(\PID_CONTROLLER.integral [2]), 
            .I1(GND_net), .I2(n79[2]), .I3(n34112), .O(n5_adj_3654)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 add_3068_2_lut (.I0(GND_net), .I1(n44_adj_3656), .I2(n137_adj_3657), 
            .I3(GND_net), .O(n8274[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3068_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3354_11 (.CI(n34271), .I0(n15114[8]), .I1(GND_net), .CO(n34272));
    SB_CARRY add_3066_2 (.CI(GND_net), .I0(n38_adj_3641), .I1(n131_adj_3642), 
            .CO(n35459));
    SB_LUT4 mult_14_add_1217_15_lut (.I0(GND_net), .I1(n1803[12]), .I2(GND_net), 
            .I3(n35904), .O(n1802[13])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1217_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1217_15 (.CI(n35904), .I0(n1803[12]), .I1(GND_net), 
            .CO(n35905));
    SB_LUT4 add_3063_19_lut (.I0(GND_net), .I1(n8184[16]), .I2(GND_net), 
            .I3(n35412), .O(n8159[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3063_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3060_10_lut (.I0(GND_net), .I1(n8106[7]), .I2(GND_net), 
            .I3(n35331), .O(n8078[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3060_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3150_16_lut (.I0(GND_net), .I1(n10852[13]), .I2(GND_net), 
            .I3(n35184), .O(n10118[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3150_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1217_14_lut (.I0(GND_net), .I1(n1803[11]), .I2(GND_net), 
            .I3(n35903), .O(n1802[12])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1217_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3354_10_lut (.I0(GND_net), .I1(n15114[7]), .I2(GND_net), 
            .I3(n34270), .O(n14793[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3354_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1217_14 (.CI(n35903), .I0(n1803[11]), .I1(GND_net), 
            .CO(n35904));
    SB_CARRY unary_minus_5_add_3_4 (.CI(n34112), .I0(GND_net), .I1(n79[2]), 
            .CO(n34113));
    SB_LUT4 unary_minus_5_add_3_3_lut (.I0(\PID_CONTROLLER.integral [1]), 
            .I1(GND_net), .I2(n79[1]), .I3(n34111), .O(n3_adj_3658)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_3_lut.LUT_INIT = 16'h6996;
    SB_LUT4 mult_14_add_1217_13_lut (.I0(GND_net), .I1(n1803[10]), .I2(GND_net), 
            .I3(n35902), .O(n1802[11])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1217_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3354_10 (.CI(n34270), .I0(n15114[7]), .I1(GND_net), .CO(n34271));
    SB_CARRY mult_14_add_1217_13 (.CI(n35902), .I0(n1803[10]), .I1(GND_net), 
            .CO(n35903));
    SB_LUT4 mult_14_add_1217_12_lut (.I0(GND_net), .I1(n1803[9]), .I2(GND_net), 
            .I3(n35901), .O(n1802[10])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1217_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3068_2 (.CI(GND_net), .I0(n44_adj_3656), .I1(n137_adj_3657), 
            .CO(n35496));
    SB_LUT4 add_3065_22_lut (.I0(GND_net), .I1(n8231[19]), .I2(GND_net), 
            .I3(n35458), .O(n8208[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3065_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3063_19 (.CI(n35412), .I0(n8184[16]), .I1(GND_net), .CO(n35413));
    SB_CARRY add_3060_10 (.CI(n35331), .I0(n8106[7]), .I1(GND_net), .CO(n35332));
    SB_CARRY add_3150_16 (.CI(n35184), .I0(n10852[13]), .I1(GND_net), 
            .CO(n35185));
    SB_CARRY mult_14_add_1217_12 (.CI(n35901), .I0(n1803[9]), .I1(GND_net), 
            .CO(n35902));
    SB_LUT4 add_3279_3_lut (.I0(GND_net), .I1(n13734[0]), .I2(n180), .I3(n34624), 
            .O(n13256[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3279_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1217_11_lut (.I0(GND_net), .I1(n1803[8]), .I2(GND_net), 
            .I3(n35900), .O(n1802[9])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1217_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3354_9_lut (.I0(GND_net), .I1(n15114[6]), .I2(GND_net), 
            .I3(n34269), .O(n14793[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3354_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3354_9 (.CI(n34269), .I0(n15114[6]), .I1(GND_net), .CO(n34270));
    SB_CARRY add_3279_3 (.CI(n34624), .I0(n13734[0]), .I1(n180), .CO(n34625));
    SB_CARRY mult_14_add_1217_11 (.CI(n35900), .I0(n1803[8]), .I1(GND_net), 
            .CO(n35901));
    SB_LUT4 add_3354_8_lut (.I0(GND_net), .I1(n15114[5]), .I2(n719_adj_3660), 
            .I3(n34268), .O(n14793[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3354_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3354_8 (.CI(n34268), .I0(n15114[5]), .I1(n719_adj_3660), 
            .CO(n34269));
    SB_CARRY unary_minus_5_add_3_3 (.CI(n34111), .I0(GND_net), .I1(n79[1]), 
            .CO(n34112));
    SB_LUT4 add_3150_15_lut (.I0(GND_net), .I1(n10852[12]), .I2(GND_net), 
            .I3(n35183), .O(n10118[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3150_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3279_2_lut (.I0(GND_net), .I1(n35), .I2(n107), .I3(GND_net), 
            .O(n13256[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3279_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3354_7_lut (.I0(GND_net), .I1(n15114[4]), .I2(n622_adj_3661), 
            .I3(n34267), .O(n14793[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3354_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1217_10_lut (.I0(GND_net), .I1(n1803[7]), .I2(GND_net), 
            .I3(n35899), .O(n1802[8])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1217_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_5_add_3_2_lut (.I0(GND_net), .I1(GND_net), .I2(n79[0]), 
            .I3(VCC_net), .O(n76[0])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1217_10 (.CI(n35899), .I0(n1803[7]), .I1(GND_net), 
            .CO(n35900));
    SB_CARRY add_3354_7 (.CI(n34267), .I0(n15114[4]), .I1(n622_adj_3661), 
            .CO(n34268));
    SB_CARRY unary_minus_5_add_3_2 (.CI(VCC_net), .I0(GND_net), .I1(n79[0]), 
            .CO(n34111));
    SB_CARRY add_3279_2 (.CI(GND_net), .I0(n35), .I1(n107), .CO(n34624));
    SB_LUT4 add_3354_6_lut (.I0(GND_net), .I1(n15114[3]), .I2(n525_adj_3664), 
            .I3(n34266), .O(n14793[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3354_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1217_9_lut (.I0(GND_net), .I1(n1803[6]), .I2(GND_net), 
            .I3(n35898), .O(n1802[7])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1217_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3103_29_lut (.I0(GND_net), .I1(n9929[26]), .I2(GND_net), 
            .I3(n34623), .O(n9125[27])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3103_29_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_17_add_3_12_lut (.I0(GND_net), .I1(GND_net), .I2(n82[31]), 
            .I3(n34110), .O(pwm_23__N_2960[10])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_17_add_3_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_17_add_3_11_lut (.I0(GND_net), .I1(GND_net), .I2(n82[31]), 
            .I3(n34109), .O(pwm_23__N_2960[9])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_17_add_3_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3354_6 (.CI(n34266), .I0(n15114[3]), .I1(n525_adj_3664), 
            .CO(n34267));
    SB_CARRY unary_minus_17_add_3_11 (.CI(n34109), .I0(GND_net), .I1(n82[31]), 
            .CO(n34110));
    SB_LUT4 unary_minus_17_add_3_10_lut (.I0(GND_net), .I1(GND_net), .I2(n82[8]), 
            .I3(n34108), .O(pwm_23__N_2960[8])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_17_add_3_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3060_9_lut (.I0(GND_net), .I1(n8106[6]), .I2(GND_net), 
            .I3(n35330), .O(n8078[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3060_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3150_15 (.CI(n35183), .I0(n10852[12]), .I1(GND_net), 
            .CO(n35184));
    SB_LUT4 add_3103_28_lut (.I0(GND_net), .I1(n9929[25]), .I2(GND_net), 
            .I3(n34622), .O(n9125[26])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3103_28_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3354_5_lut (.I0(GND_net), .I1(n15114[2]), .I2(n428_adj_3668), 
            .I3(n34265), .O(n14793[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3354_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3354_5 (.CI(n34265), .I0(n15114[2]), .I1(n428_adj_3668), 
            .CO(n34266));
    SB_LUT4 add_3354_4_lut (.I0(GND_net), .I1(n15114[1]), .I2(n331_adj_3669), 
            .I3(n34264), .O(n14793[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3354_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3067_20_lut (.I0(GND_net), .I1(n8274[17]), .I2(GND_net), 
            .I3(n35495), .O(n8253[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3067_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3065_21_lut (.I0(GND_net), .I1(n8231[18]), .I2(GND_net), 
            .I3(n35457), .O(n8208[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3065_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3063_18_lut (.I0(GND_net), .I1(n8184[15]), .I2(GND_net), 
            .I3(n35411), .O(n8159[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3063_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3354_4 (.CI(n34264), .I0(n15114[1]), .I1(n331_adj_3669), 
            .CO(n34265));
    SB_CARRY mult_14_add_1217_9 (.CI(n35898), .I0(n1803[6]), .I1(GND_net), 
            .CO(n35899));
    SB_LUT4 add_3150_14_lut (.I0(GND_net), .I1(n10852[11]), .I2(GND_net), 
            .I3(n35182), .O(n10118[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3150_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3103_28 (.CI(n34622), .I0(n9929[25]), .I1(GND_net), .CO(n34623));
    SB_LUT4 add_3354_3_lut (.I0(GND_net), .I1(n15114[0]), .I2(n234_adj_3670), 
            .I3(n34263), .O(n14793[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3354_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3060_9 (.CI(n35330), .I0(n8106[6]), .I1(GND_net), .CO(n35331));
    SB_CARRY add_3354_3 (.CI(n34263), .I0(n15114[0]), .I1(n234_adj_3670), 
            .CO(n34264));
    SB_LUT4 add_3103_27_lut (.I0(GND_net), .I1(n9929[24]), .I2(GND_net), 
            .I3(n34621), .O(n9125[25])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3103_27_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3354_2_lut (.I0(GND_net), .I1(n44_adj_3671), .I2(n137_adj_3672), 
            .I3(GND_net), .O(n14793[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3354_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3150_14 (.CI(n35182), .I0(n10852[11]), .I1(GND_net), 
            .CO(n35183));
    SB_CARRY add_3103_27 (.CI(n34621), .I0(n9929[24]), .I1(GND_net), .CO(n34622));
    SB_CARRY unary_minus_17_add_3_10 (.CI(n34108), .I0(GND_net), .I1(n82[8]), 
            .CO(n34109));
    SB_LUT4 unary_minus_17_add_3_9_lut (.I0(GND_net), .I1(GND_net), .I2(n82[7]), 
            .I3(n34107), .O(pwm_23__N_2960[7])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_17_add_3_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1217_8_lut (.I0(GND_net), .I1(n1803[5]), .I2(n530), 
            .I3(n35897), .O(n1802[6])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1217_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3103_26_lut (.I0(GND_net), .I1(n9929[23]), .I2(GND_net), 
            .I3(n34620), .O(n9125[24])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3103_26_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3354_2 (.CI(GND_net), .I0(n44_adj_3671), .I1(n137_adj_3672), 
            .CO(n34263));
    SB_CARRY unary_minus_17_add_3_9 (.CI(n34107), .I0(GND_net), .I1(n82[7]), 
            .CO(n34108));
    SB_LUT4 add_3150_13_lut (.I0(GND_net), .I1(n10852[10]), .I2(GND_net), 
            .I3(n35181), .O(n10118[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3150_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3103_26 (.CI(n34620), .I0(n9929[23]), .I1(GND_net), .CO(n34621));
    SB_LUT4 unary_minus_17_add_3_8_lut (.I0(GND_net), .I1(GND_net), .I2(n82[6]), 
            .I3(n34106), .O(\pwm_23__N_2960[6] )) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_17_add_3_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_17_add_3_8 (.CI(n34106), .I0(GND_net), .I1(n82[6]), 
            .CO(n34107));
    SB_LUT4 unary_minus_17_add_3_7_lut (.I0(GND_net), .I1(GND_net), .I2(n82[5]), 
            .I3(n34105), .O(\pwm_23__N_2960[5] )) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_17_add_3_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3103_25_lut (.I0(GND_net), .I1(n9929[22]), .I2(GND_net), 
            .I3(n34619), .O(n9125[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3103_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1217_8 (.CI(n35897), .I0(n1803[5]), .I1(n530), 
            .CO(n35898));
    SB_CARRY add_3103_25 (.CI(n34619), .I0(n9929[22]), .I1(GND_net), .CO(n34620));
    SB_CARRY unary_minus_17_add_3_7 (.CI(n34105), .I0(GND_net), .I1(n82[5]), 
            .CO(n34106));
    SB_LUT4 unary_minus_17_add_3_6_lut (.I0(GND_net), .I1(GND_net), .I2(n82[4]), 
            .I3(n34104), .O(pwm_23__N_2960[4])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_17_add_3_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_17_add_3_6 (.CI(n34104), .I0(GND_net), .I1(n82[4]), 
            .CO(n34105));
    SB_CARRY add_3063_18 (.CI(n35411), .I0(n8184[15]), .I1(GND_net), .CO(n35412));
    SB_LUT4 add_3060_8_lut (.I0(GND_net), .I1(n8106[5]), .I2(n695_adj_3677), 
            .I3(n35329), .O(n8078[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3060_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3150_13 (.CI(n35181), .I0(n10852[10]), .I1(GND_net), 
            .CO(n35182));
    SB_LUT4 add_3103_24_lut (.I0(GND_net), .I1(n9929[21]), .I2(GND_net), 
            .I3(n34618), .O(n9125[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3103_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1217_7_lut (.I0(GND_net), .I1(n1803[4]), .I2(n457_c), 
            .I3(n35896), .O(n1802[5])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1217_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_11_inv_0_i13_1_lut (.I0(\PID_CONTROLLER.err[12] ), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n64[12]));   // verilog/motorControl.v(43[31:45])
    defparam sub_11_inv_0_i13_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_3150_12_lut (.I0(GND_net), .I1(n10852[9]), .I2(GND_net), 
            .I3(n35180), .O(n10118[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3150_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1217_7 (.CI(n35896), .I0(n1803[4]), .I1(n457_c), 
            .CO(n35897));
    SB_LUT4 mult_10_i406_2_lut (.I0(\Kp[6] ), .I1(\PID_CONTROLLER.err[7] ), 
            .I2(GND_net), .I3(GND_net), .O(n604_adj_3417));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i406_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i20_2_lut (.I0(\Kd[0] ), .I1(n57[9]), .I2(GND_net), 
            .I3(GND_net), .O(n29));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i20_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i174_2_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err[21] ), 
            .I2(GND_net), .I3(GND_net), .O(n258));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i174_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_3070_14_lut (.I0(GND_net), .I1(n8331[11]), .I2(GND_net), 
            .I3(n35540), .O(n8313[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3070_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3070_14 (.CI(n35540), .I0(n8331[11]), .I1(GND_net), .CO(n35541));
    SB_CARRY add_3150_12 (.CI(n35180), .I0(n10852[9]), .I1(GND_net), .CO(n35181));
    SB_CARRY add_3065_21 (.CI(n35457), .I0(n8231[18]), .I1(GND_net), .CO(n35458));
    SB_LUT4 add_3063_17_lut (.I0(GND_net), .I1(n8184[14]), .I2(GND_net), 
            .I3(n35410), .O(n8159[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3063_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i239_2_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err[21] ), 
            .I2(GND_net), .I3(GND_net), .O(n355));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i239_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_14_add_1217_6_lut (.I0(GND_net), .I1(n1803[3]), .I2(n384), 
            .I3(n35895), .O(n1802[4])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1217_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3103_24 (.CI(n34618), .I0(n9929[21]), .I1(GND_net), .CO(n34619));
    SB_LUT4 unary_minus_17_add_3_5_lut (.I0(GND_net), .I1(GND_net), .I2(n82[3]), 
            .I3(n34103), .O(pwm_23__N_2960[3])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_17_add_3_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3150_11_lut (.I0(GND_net), .I1(n10852[8]), .I2(GND_net), 
            .I3(n35179), .O(n10118[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3150_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3103_23_lut (.I0(GND_net), .I1(n9929[20]), .I2(GND_net), 
            .I3(n34617), .O(n9125[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3103_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1217_6 (.CI(n35895), .I0(n1803[3]), .I1(n384), 
            .CO(n35896));
    SB_LUT4 sub_11_inv_0_i14_1_lut (.I0(\PID_CONTROLLER.err[13] ), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n64[13]));   // verilog/motorControl.v(43[31:45])
    defparam sub_11_inv_0_i14_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_3103_23 (.CI(n34617), .I0(n9929[20]), .I1(GND_net), .CO(n34618));
    SB_LUT4 mult_14_add_1217_5_lut (.I0(GND_net), .I1(n1803[2]), .I2(n311_adj_3681), 
            .I3(n35894), .O(n1802[3])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1217_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_17_add_3_5 (.CI(n34103), .I0(GND_net), .I1(n82[3]), 
            .CO(n34104));
    SB_CARRY add_3060_8 (.CI(n35329), .I0(n8106[5]), .I1(n695_adj_3677), 
            .CO(n35330));
    SB_CARRY add_3150_11 (.CI(n35179), .I0(n10852[8]), .I1(GND_net), .CO(n35180));
    SB_LUT4 add_3150_10_lut (.I0(GND_net), .I1(n10852[7]), .I2(GND_net), 
            .I3(n35178), .O(n10118[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3150_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3060_7_lut (.I0(GND_net), .I1(n8106[4]), .I2(n598_adj_3682), 
            .I3(n35328), .O(n8078[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3060_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3060_7 (.CI(n35328), .I0(n8106[4]), .I1(n598_adj_3682), 
            .CO(n35329));
    SB_CARRY add_3150_10 (.CI(n35178), .I0(n10852[7]), .I1(GND_net), .CO(n35179));
    SB_LUT4 add_3150_9_lut (.I0(GND_net), .I1(n10852[6]), .I2(GND_net), 
            .I3(n35177), .O(n10118[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3150_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3150_9 (.CI(n35177), .I0(n10852[6]), .I1(GND_net), .CO(n35178));
    SB_CARRY mult_14_add_1217_5 (.CI(n35894), .I0(n1803[2]), .I1(n311_adj_3681), 
            .CO(n35895));
    SB_LUT4 add_3065_20_lut (.I0(GND_net), .I1(n8231[17]), .I2(GND_net), 
            .I3(n35456), .O(n8208[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3065_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3060_6_lut (.I0(GND_net), .I1(n8106[3]), .I2(n501_adj_3683), 
            .I3(n35327), .O(n8078[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3060_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3063_17 (.CI(n35410), .I0(n8184[14]), .I1(GND_net), .CO(n35411));
    SB_CARRY add_3060_6 (.CI(n35327), .I0(n8106[3]), .I1(n501_adj_3683), 
            .CO(n35328));
    SB_LUT4 mult_14_add_1217_4_lut (.I0(GND_net), .I1(n1803[1]), .I2(n238_adj_3685), 
            .I3(n35893), .O(n1802[2])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1217_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3067_19_lut (.I0(GND_net), .I1(n8274[16]), .I2(GND_net), 
            .I3(n35494), .O(n8253[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3067_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1217_4 (.CI(n35893), .I0(n1803[1]), .I1(n238_adj_3685), 
            .CO(n35894));
    SB_LUT4 mult_14_add_1217_3_lut (.I0(GND_net), .I1(n1803[0]), .I2(n165_adj_3687), 
            .I3(n35892), .O(n1802[1])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1217_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3070_13_lut (.I0(GND_net), .I1(n8331[10]), .I2(GND_net), 
            .I3(n35539), .O(n8313[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3070_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3150_8_lut (.I0(GND_net), .I1(n10852[5]), .I2(n545), .I3(n35176), 
            .O(n10118[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3150_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1217_3 (.CI(n35892), .I0(n1803[0]), .I1(n165_adj_3687), 
            .CO(n35893));
    SB_LUT4 mult_14_add_1217_2_lut (.I0(GND_net), .I1(n23_adj_3688), .I2(n92), 
            .I3(GND_net), .O(n1802[0])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1217_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1217_2 (.CI(GND_net), .I0(n23_adj_3688), .I1(n92), 
            .CO(n35892));
    SB_LUT4 add_3075_5_lut (.I0(GND_net), .I1(n8406[2]), .I2(n449_adj_3689), 
            .I3(n35596), .O(n8393[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3075_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3103_22_lut (.I0(GND_net), .I1(n9929[19]), .I2(GND_net), 
            .I3(n34616), .O(n9125[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3103_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1216_24_lut (.I0(GND_net), .I1(n1802[21]), .I2(GND_net), 
            .I3(n35890), .O(n1801[22])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1216_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1216_24 (.CI(n35890), .I0(n1802[21]), .I1(GND_net), 
            .CO(n1703));
    SB_LUT4 mult_14_add_1216_23_lut (.I0(GND_net), .I1(n1802[20]), .I2(GND_net), 
            .I3(n35889), .O(n1801[21])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1216_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1216_23 (.CI(n35889), .I0(n1802[20]), .I1(GND_net), 
            .CO(n35890));
    SB_CARRY add_3150_8 (.CI(n35176), .I0(n10852[5]), .I1(n545), .CO(n35177));
    SB_CARRY add_3103_22 (.CI(n34616), .I0(n9929[19]), .I1(GND_net), .CO(n34617));
    SB_CARRY add_3067_19 (.CI(n35494), .I0(n8274[16]), .I1(GND_net), .CO(n35495));
    SB_CARRY add_3075_5 (.CI(n35596), .I0(n8406[2]), .I1(n449_adj_3689), 
            .CO(n35597));
    SB_LUT4 mult_14_add_1216_22_lut (.I0(GND_net), .I1(n1802[19]), .I2(GND_net), 
            .I3(n35888), .O(n1801[20])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1216_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3075_4_lut (.I0(GND_net), .I1(n8406[1]), .I2(n352_adj_3690), 
            .I3(n35595), .O(n8393[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3075_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1216_22 (.CI(n35888), .I0(n1802[19]), .I1(GND_net), 
            .CO(n35889));
    SB_LUT4 mult_14_add_1216_21_lut (.I0(GND_net), .I1(n1802[18]), .I2(GND_net), 
            .I3(n35887), .O(n1801[19])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1216_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1216_21 (.CI(n35887), .I0(n1802[18]), .I1(GND_net), 
            .CO(n35888));
    SB_LUT4 mult_14_add_1216_20_lut (.I0(GND_net), .I1(n1802[17]), .I2(GND_net), 
            .I3(n35886), .O(n1801[18])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1216_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_17_add_3_4_lut (.I0(GND_net), .I1(GND_net), .I2(n82[2]), 
            .I3(n34102), .O(pwm_23__N_2960[2])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_17_add_3_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3150_7_lut (.I0(GND_net), .I1(n10852[4]), .I2(n472), .I3(n35175), 
            .O(n10118[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3150_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1216_20 (.CI(n35886), .I0(n1802[17]), .I1(GND_net), 
            .CO(n35887));
    SB_LUT4 add_3103_21_lut (.I0(GND_net), .I1(n9929[18]), .I2(GND_net), 
            .I3(n34615), .O(n9125[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3103_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1216_19_lut (.I0(GND_net), .I1(n1802[16]), .I2(GND_net), 
            .I3(n35885), .O(n1801[17])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1216_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1216_19 (.CI(n35885), .I0(n1802[16]), .I1(GND_net), 
            .CO(n35886));
    SB_CARRY add_3070_13 (.CI(n35539), .I0(n8331[10]), .I1(GND_net), .CO(n35540));
    SB_CARRY add_3075_4 (.CI(n35595), .I0(n8406[1]), .I1(n352_adj_3690), 
            .CO(n35596));
    SB_CARRY add_3103_21 (.CI(n34615), .I0(n9929[18]), .I1(GND_net), .CO(n34616));
    SB_CARRY unary_minus_17_add_3_4 (.CI(n34102), .I0(GND_net), .I1(n82[2]), 
            .CO(n34103));
    SB_CARRY add_3150_7 (.CI(n35175), .I0(n10852[4]), .I1(n472), .CO(n35176));
    SB_LUT4 add_3103_20_lut (.I0(GND_net), .I1(n9929[17]), .I2(GND_net), 
            .I3(n34614), .O(n9125[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3103_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3103_20 (.CI(n34614), .I0(n9929[17]), .I1(GND_net), .CO(n34615));
    SB_LUT4 add_3103_19_lut (.I0(GND_net), .I1(n9929[16]), .I2(GND_net), 
            .I3(n34613), .O(n9125[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3103_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3070_12_lut (.I0(GND_net), .I1(n8331[9]), .I2(GND_net), 
            .I3(n35538), .O(n8313[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3070_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3067_18_lut (.I0(GND_net), .I1(n8274[15]), .I2(GND_net), 
            .I3(n35493), .O(n8253[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3067_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3065_20 (.CI(n35456), .I0(n8231[17]), .I1(GND_net), .CO(n35457));
    SB_CARRY add_3070_12 (.CI(n35538), .I0(n8331[9]), .I1(GND_net), .CO(n35539));
    SB_LUT4 add_3063_16_lut (.I0(GND_net), .I1(n8184[13]), .I2(GND_net), 
            .I3(n35409), .O(n8159[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3063_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3060_5_lut (.I0(GND_net), .I1(n8106[2]), .I2(n404_adj_3692), 
            .I3(n35326), .O(n8078[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3060_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3150_6_lut (.I0(GND_net), .I1(n10852[3]), .I2(n399), .I3(n35174), 
            .O(n10118[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3150_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3150_6 (.CI(n35174), .I0(n10852[3]), .I1(n399), .CO(n35175));
    SB_CARRY add_3060_5 (.CI(n35326), .I0(n8106[2]), .I1(n404_adj_3692), 
            .CO(n35327));
    SB_LUT4 add_3150_5_lut (.I0(GND_net), .I1(n10852[2]), .I2(n326), .I3(n35173), 
            .O(n10118[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3150_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3150_5 (.CI(n35173), .I0(n10852[2]), .I1(n326), .CO(n35174));
    SB_LUT4 add_3150_4_lut (.I0(GND_net), .I1(n10852[1]), .I2(n253), .I3(n35172), 
            .O(n10118[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3150_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3065_19_lut (.I0(GND_net), .I1(n8231[16]), .I2(GND_net), 
            .I3(n35455), .O(n8208[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3065_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3063_16 (.CI(n35409), .I0(n8184[13]), .I1(GND_net), .CO(n35410));
    SB_LUT4 add_3060_4_lut (.I0(GND_net), .I1(n8106[1]), .I2(n307_adj_3693), 
            .I3(n35325), .O(n8078[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3060_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3150_4 (.CI(n35172), .I0(n10852[1]), .I1(n253), .CO(n35173));
    SB_LUT4 add_3150_3_lut (.I0(GND_net), .I1(n10852[0]), .I2(n180), .I3(n35171), 
            .O(n10118[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3150_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1216_18_lut (.I0(GND_net), .I1(n1802[15]), .I2(GND_net), 
            .I3(n35884), .O(n1801[16])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1216_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3060_4 (.CI(n35325), .I0(n8106[1]), .I1(n307_adj_3693), 
            .CO(n35326));
    SB_CARRY add_3150_3 (.CI(n35171), .I0(n10852[0]), .I1(n180), .CO(n35172));
    SB_CARRY mult_14_add_1216_18 (.CI(n35884), .I0(n1802[15]), .I1(GND_net), 
            .CO(n35885));
    SB_LUT4 add_3150_2_lut (.I0(GND_net), .I1(n35), .I2(n107), .I3(GND_net), 
            .O(n10118[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3150_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3067_18 (.CI(n35493), .I0(n8274[15]), .I1(GND_net), .CO(n35494));
    SB_LUT4 mult_14_add_1216_17_lut (.I0(GND_net), .I1(n1802[14]), .I2(GND_net), 
            .I3(n35883), .O(n1801[15])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1216_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3065_19 (.CI(n35455), .I0(n8231[16]), .I1(GND_net), .CO(n35456));
    SB_LUT4 add_3063_15_lut (.I0(GND_net), .I1(n8184[12]), .I2(GND_net), 
            .I3(n35408), .O(n8159[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3063_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3060_3_lut (.I0(GND_net), .I1(n8106[0]), .I2(n210_adj_3694), 
            .I3(n35324), .O(n8078[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3060_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3150_2 (.CI(GND_net), .I0(n35), .I1(n107), .CO(n35171));
    SB_CARRY mult_14_add_1216_17 (.CI(n35883), .I0(n1802[14]), .I1(GND_net), 
            .CO(n35884));
    SB_LUT4 add_3070_11_lut (.I0(GND_net), .I1(n8331[8]), .I2(GND_net), 
            .I3(n35537), .O(n8313[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3070_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1216_16_lut (.I0(GND_net), .I1(n1802[13]), .I2(GND_net), 
            .I3(n35882), .O(n1801[14])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1216_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1216_16 (.CI(n35882), .I0(n1802[13]), .I1(GND_net), 
            .CO(n35883));
    SB_LUT4 add_3075_3_lut (.I0(GND_net), .I1(n8406[0]), .I2(n255_adj_3695), 
            .I3(n35594), .O(n8393[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3075_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3070_11 (.CI(n35537), .I0(n8331[8]), .I1(GND_net), .CO(n35538));
    SB_LUT4 mult_14_add_1216_15_lut (.I0(GND_net), .I1(n1802[12]), .I2(GND_net), 
            .I3(n35881), .O(n1801[13])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1216_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3070_10_lut (.I0(GND_net), .I1(n8331[7]), .I2(GND_net), 
            .I3(n35536), .O(n8313[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3070_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1216_15 (.CI(n35881), .I0(n1802[12]), .I1(GND_net), 
            .CO(n35882));
    SB_LUT4 unary_minus_17_add_3_3_lut (.I0(GND_net), .I1(GND_net), .I2(n82[1]), 
            .I3(n34101), .O(pwm_23__N_2960[1])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_17_add_3_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1216_14_lut (.I0(GND_net), .I1(n1802[11]), .I2(GND_net), 
            .I3(n35880), .O(n1801[12])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1216_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1216_14 (.CI(n35880), .I0(n1802[11]), .I1(GND_net), 
            .CO(n35881));
    SB_CARRY unary_minus_17_add_3_3 (.CI(n34101), .I0(GND_net), .I1(n82[1]), 
            .CO(n34102));
    SB_CARRY add_3070_10 (.CI(n35536), .I0(n8331[7]), .I1(GND_net), .CO(n35537));
    SB_LUT4 mult_14_add_1216_13_lut (.I0(GND_net), .I1(n1802[10]), .I2(GND_net), 
            .I3(n35879), .O(n1801[11])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1216_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3178_19_lut (.I0(GND_net), .I1(n11531[16]), .I2(GND_net), 
            .I3(n35170), .O(n10852[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3178_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1216_13 (.CI(n35879), .I0(n1802[10]), .I1(GND_net), 
            .CO(n35880));
    SB_CARRY add_3060_3 (.CI(n35324), .I0(n8106[0]), .I1(n210_adj_3694), 
            .CO(n35325));
    SB_LUT4 add_3178_18_lut (.I0(GND_net), .I1(n11531[15]), .I2(GND_net), 
            .I3(n35169), .O(n10852[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3178_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3178_18 (.CI(n35169), .I0(n11531[15]), .I1(GND_net), 
            .CO(n35170));
    SB_LUT4 add_3065_18_lut (.I0(GND_net), .I1(n8231[15]), .I2(GND_net), 
            .I3(n35454), .O(n8208[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3065_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3063_15 (.CI(n35408), .I0(n8184[12]), .I1(GND_net), .CO(n35409));
    SB_LUT4 add_3060_2_lut (.I0(GND_net), .I1(n20_adj_3697), .I2(n113_adj_3698), 
            .I3(GND_net), .O(n8078[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3060_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3178_17_lut (.I0(GND_net), .I1(n11531[14]), .I2(GND_net), 
            .I3(n35168), .O(n10852[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3178_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3178_17 (.CI(n35168), .I0(n11531[14]), .I1(GND_net), 
            .CO(n35169));
    SB_CARRY add_3060_2 (.CI(GND_net), .I0(n20_adj_3697), .I1(n113_adj_3698), 
            .CO(n35324));
    SB_LUT4 add_3178_16_lut (.I0(GND_net), .I1(n11531[13]), .I2(GND_net), 
            .I3(n35167), .O(n10852[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3178_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3178_16 (.CI(n35167), .I0(n11531[13]), .I1(GND_net), 
            .CO(n35168));
    SB_LUT4 sub_11_inv_0_i15_1_lut (.I0(\PID_CONTROLLER.err[14] ), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n64[14]));   // verilog/motorControl.v(43[31:45])
    defparam sub_11_inv_0_i15_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_3075_3 (.CI(n35594), .I0(n8406[0]), .I1(n255_adj_3695), 
            .CO(n35595));
    SB_LUT4 add_3070_9_lut (.I0(GND_net), .I1(n8331[6]), .I2(GND_net), 
            .I3(n35535), .O(n8313[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3070_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3063_14_lut (.I0(GND_net), .I1(n8184[11]), .I2(GND_net), 
            .I3(n35407), .O(n8159[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3063_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3059_28_lut (.I0(GND_net), .I1(n8078[25]), .I2(GND_net), 
            .I3(n35323), .O(n8049[26])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3059_28_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3067_17_lut (.I0(GND_net), .I1(n8274[14]), .I2(GND_net), 
            .I3(n35492), .O(n8253[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3067_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3065_18 (.CI(n35454), .I0(n8231[15]), .I1(GND_net), .CO(n35455));
    SB_LUT4 add_3178_15_lut (.I0(GND_net), .I1(n11531[12]), .I2(GND_net), 
            .I3(n35166), .O(n10852[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3178_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3063_14 (.CI(n35407), .I0(n8184[11]), .I1(GND_net), .CO(n35408));
    SB_LUT4 add_3059_27_lut (.I0(GND_net), .I1(n8078[24]), .I2(GND_net), 
            .I3(n35322), .O(n8049[25])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3059_27_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3178_15 (.CI(n35166), .I0(n11531[12]), .I1(GND_net), 
            .CO(n35167));
    SB_LUT4 add_3178_14_lut (.I0(GND_net), .I1(n11531[11]), .I2(GND_net), 
            .I3(n35165), .O(n10852[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3178_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3178_14 (.CI(n35165), .I0(n11531[11]), .I1(GND_net), 
            .CO(n35166));
    SB_CARRY add_3059_27 (.CI(n35322), .I0(n8078[24]), .I1(GND_net), .CO(n35323));
    SB_LUT4 add_3059_26_lut (.I0(GND_net), .I1(n8078[23]), .I2(GND_net), 
            .I3(n35321), .O(n8049[24])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3059_26_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3178_13_lut (.I0(GND_net), .I1(n11531[10]), .I2(GND_net), 
            .I3(n35164), .O(n10852[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3178_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3178_13 (.CI(n35164), .I0(n11531[10]), .I1(GND_net), 
            .CO(n35165));
    SB_LUT4 add_3075_2_lut (.I0(GND_net), .I1(n65_adj_3699), .I2(n158_adj_3700), 
            .I3(GND_net), .O(n8393[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3075_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3178_12_lut (.I0(GND_net), .I1(n11531[9]), .I2(GND_net), 
            .I3(n35163), .O(n10852[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3178_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_17_add_3_2_lut (.I0(n28200), .I1(GND_net), .I2(n82[0]), 
            .I3(VCC_net), .O(n44044)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_17_add_3_2_lut.LUT_INIT = 16'h8228;
    SB_LUT4 add_3063_13_lut (.I0(GND_net), .I1(n8184[10]), .I2(GND_net), 
            .I3(n35406), .O(n8159[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3063_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1216_12_lut (.I0(GND_net), .I1(n1802[9]), .I2(GND_net), 
            .I3(n35878), .O(n1801[10])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1216_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_17_add_3_2 (.CI(VCC_net), .I0(GND_net), .I1(n82[0]), 
            .CO(n34101));
    SB_CARRY mult_14_add_1216_12 (.CI(n35878), .I0(n1802[9]), .I1(GND_net), 
            .CO(n35879));
    SB_LUT4 mult_14_add_1216_11_lut (.I0(GND_net), .I1(n1802[8]), .I2(GND_net), 
            .I3(n35877), .O(n1801[9])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1216_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3070_9 (.CI(n35535), .I0(n8331[6]), .I1(GND_net), .CO(n35536));
    SB_CARRY mult_14_add_1216_11 (.CI(n35877), .I0(n1802[8]), .I1(GND_net), 
            .CO(n35878));
    SB_LUT4 mult_14_add_1216_10_lut (.I0(GND_net), .I1(n1802[7]), .I2(GND_net), 
            .I3(n35876), .O(n1801[8])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1216_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3065_17_lut (.I0(GND_net), .I1(n8231[14]), .I2(GND_net), 
            .I3(n35453), .O(n8208[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3065_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3075_2 (.CI(GND_net), .I0(n65_adj_3699), .I1(n158_adj_3700), 
            .CO(n35594));
    SB_CARRY mult_14_add_1216_10 (.CI(n35876), .I0(n1802[7]), .I1(GND_net), 
            .CO(n35877));
    SB_LUT4 mult_14_add_1216_9_lut (.I0(GND_net), .I1(n1802[6]), .I2(GND_net), 
            .I3(n35875), .O(n1801[7])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1216_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3067_17 (.CI(n35492), .I0(n8274[14]), .I1(GND_net), .CO(n35493));
    SB_LUT4 add_3074_13_lut (.I0(GND_net), .I1(n8393[10]), .I2(GND_net), 
            .I3(n35593), .O(n8379[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3074_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1216_9 (.CI(n35875), .I0(n1802[6]), .I1(GND_net), 
            .CO(n35876));
    SB_LUT4 add_3074_12_lut (.I0(GND_net), .I1(n8393[9]), .I2(GND_net), 
            .I3(n35592), .O(n8379[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3074_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1216_8_lut (.I0(GND_net), .I1(n1802[5]), .I2(n527), 
            .I3(n35874), .O(n1801[6])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1216_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3059_26 (.CI(n35321), .I0(n8078[23]), .I1(GND_net), .CO(n35322));
    SB_CARRY mult_14_add_1216_8 (.CI(n35874), .I0(n1802[5]), .I1(n527), 
            .CO(n35875));
    SB_LUT4 add_3067_16_lut (.I0(GND_net), .I1(n8274[13]), .I2(GND_net), 
            .I3(n35491), .O(n8253[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3067_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1216_7_lut (.I0(GND_net), .I1(n1802[4]), .I2(n454), 
            .I3(n35873), .O(n1801[5])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1216_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1216_7 (.CI(n35873), .I0(n1802[4]), .I1(n454), 
            .CO(n35874));
    SB_LUT4 mult_14_add_1216_6_lut (.I0(GND_net), .I1(n1802[3]), .I2(n381), 
            .I3(n35872), .O(n1801[4])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1216_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1216_6 (.CI(n35872), .I0(n1802[3]), .I1(n381), 
            .CO(n35873));
    SB_CARRY add_3063_13 (.CI(n35406), .I0(n8184[10]), .I1(GND_net), .CO(n35407));
    SB_LUT4 mult_14_add_1216_5_lut (.I0(GND_net), .I1(n1802[2]), .I2(n308_adj_3706), 
            .I3(n35871), .O(n1801[3])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1216_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1216_5 (.CI(n35871), .I0(n1802[2]), .I1(n308_adj_3706), 
            .CO(n35872));
    SB_LUT4 mult_14_add_1216_4_lut (.I0(GND_net), .I1(n1802[1]), .I2(n235_adj_3708), 
            .I3(n35870), .O(n1801[2])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1216_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3070_8_lut (.I0(GND_net), .I1(n8331[5]), .I2(n725), .I3(n35534), 
            .O(n8313[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3070_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1216_4 (.CI(n35870), .I0(n1802[1]), .I1(n235_adj_3708), 
            .CO(n35871));
    SB_LUT4 mult_14_add_1216_3_lut (.I0(GND_net), .I1(n1802[0]), .I2(n162), 
            .I3(n35869), .O(n1801[1])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1216_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3103_19 (.CI(n34613), .I0(n9929[16]), .I1(GND_net), .CO(n34614));
    SB_CARRY add_3074_12 (.CI(n35592), .I0(n8393[9]), .I1(GND_net), .CO(n35593));
    SB_CARRY mult_14_add_1216_3 (.CI(n35869), .I0(n1802[0]), .I1(n162), 
            .CO(n35870));
    SB_LUT4 mult_14_add_1216_2_lut (.I0(GND_net), .I1(n20_adj_3709), .I2(n89), 
            .I3(GND_net), .O(n1801[0])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1216_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1216_2 (.CI(GND_net), .I0(n20_adj_3709), .I1(n89), 
            .CO(n35869));
    SB_LUT4 mult_14_add_1215_24_lut (.I0(GND_net), .I1(n1801[21]), .I2(GND_net), 
            .I3(n35867), .O(n1800[22])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1215_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3070_8 (.CI(n35534), .I0(n8331[5]), .I1(n725), .CO(n35535));
    SB_CARRY mult_14_add_1215_24 (.CI(n35867), .I0(n1801[21]), .I1(GND_net), 
            .CO(n1699));
    SB_LUT4 add_3074_11_lut (.I0(GND_net), .I1(n8393[8]), .I2(GND_net), 
            .I3(n35591), .O(n8379[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3074_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1215_23_lut (.I0(GND_net), .I1(n1801[20]), .I2(GND_net), 
            .I3(n35866), .O(n1800[21])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1215_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3103_18_lut (.I0(GND_net), .I1(n9929[15]), .I2(GND_net), 
            .I3(n34612), .O(n9125[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3103_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3074_11 (.CI(n35591), .I0(n8393[8]), .I1(GND_net), .CO(n35592));
    SB_CARRY mult_14_add_1215_23 (.CI(n35866), .I0(n1801[20]), .I1(GND_net), 
            .CO(n35867));
    SB_LUT4 mult_14_add_1215_22_lut (.I0(GND_net), .I1(n1801[19]), .I2(GND_net), 
            .I3(n35865), .O(n1800[20])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1215_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3059_25_lut (.I0(GND_net), .I1(n8078[22]), .I2(GND_net), 
            .I3(n35320), .O(n8049[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3059_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1215_22 (.CI(n35865), .I0(n1801[19]), .I1(GND_net), 
            .CO(n35866));
    SB_LUT4 mult_14_add_1215_21_lut (.I0(GND_net), .I1(n1801[18]), .I2(GND_net), 
            .I3(n35864), .O(n1800[19])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1215_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3074_10_lut (.I0(GND_net), .I1(n8393[7]), .I2(GND_net), 
            .I3(n35590), .O(n8379[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3074_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1215_21 (.CI(n35864), .I0(n1801[18]), .I1(GND_net), 
            .CO(n35865));
    SB_CARRY add_3067_16 (.CI(n35491), .I0(n8274[13]), .I1(GND_net), .CO(n35492));
    SB_LUT4 mult_14_add_1215_20_lut (.I0(GND_net), .I1(n1801[17]), .I2(GND_net), 
            .I3(n35863), .O(n1800[18])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1215_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3178_12 (.CI(n35163), .I0(n11531[9]), .I1(GND_net), .CO(n35164));
    SB_LUT4 add_3067_15_lut (.I0(GND_net), .I1(n8274[12]), .I2(GND_net), 
            .I3(n35490), .O(n8253[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3067_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1215_20 (.CI(n35863), .I0(n1801[17]), .I1(GND_net), 
            .CO(n35864));
    SB_LUT4 mult_14_add_1215_19_lut (.I0(GND_net), .I1(n1801[16]), .I2(GND_net), 
            .I3(n35862), .O(n1800[17])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1215_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1215_19 (.CI(n35862), .I0(n1801[16]), .I1(GND_net), 
            .CO(n35863));
    SB_LUT4 mult_14_add_1215_18_lut (.I0(GND_net), .I1(n1801[15]), .I2(GND_net), 
            .I3(n35861), .O(n1800[16])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1215_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3178_11_lut (.I0(GND_net), .I1(n11531[8]), .I2(GND_net), 
            .I3(n35162), .O(n10852[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3178_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1215_18 (.CI(n35861), .I0(n1801[15]), .I1(GND_net), 
            .CO(n35862));
    SB_LUT4 mult_14_add_1215_17_lut (.I0(GND_net), .I1(n1801[14]), .I2(GND_net), 
            .I3(n35860), .O(n1800[15])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1215_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1215_17 (.CI(n35860), .I0(n1801[14]), .I1(GND_net), 
            .CO(n35861));
    SB_LUT4 mult_14_add_1215_16_lut (.I0(GND_net), .I1(n1801[13]), .I2(GND_net), 
            .I3(n35859), .O(n1800[14])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1215_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1215_16 (.CI(n35859), .I0(n1801[13]), .I1(GND_net), 
            .CO(n35860));
    SB_LUT4 mult_14_add_1215_15_lut (.I0(GND_net), .I1(n1801[12]), .I2(GND_net), 
            .I3(n35858), .O(n1800[13])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1215_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1215_15 (.CI(n35858), .I0(n1801[12]), .I1(GND_net), 
            .CO(n35859));
    SB_LUT4 mult_14_add_1215_14_lut (.I0(GND_net), .I1(n1801[11]), .I2(GND_net), 
            .I3(n35857), .O(n1800[12])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1215_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3178_11 (.CI(n35162), .I0(n11531[8]), .I1(GND_net), .CO(n35163));
    SB_CARRY add_3065_17 (.CI(n35453), .I0(n8231[14]), .I1(GND_net), .CO(n35454));
    SB_LUT4 add_3063_12_lut (.I0(GND_net), .I1(n8184[9]), .I2(GND_net), 
            .I3(n35405), .O(n8159[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3063_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3059_25 (.CI(n35320), .I0(n8078[22]), .I1(GND_net), .CO(n35321));
    SB_LUT4 add_3178_10_lut (.I0(GND_net), .I1(n11531[7]), .I2(GND_net), 
            .I3(n35161), .O(n10852[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3178_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3103_18 (.CI(n34612), .I0(n9929[15]), .I1(GND_net), .CO(n34613));
    SB_CARRY add_3178_10 (.CI(n35161), .I0(n11531[7]), .I1(GND_net), .CO(n35162));
    SB_CARRY mult_14_add_1215_14 (.CI(n35857), .I0(n1801[11]), .I1(GND_net), 
            .CO(n35858));
    SB_LUT4 add_3103_17_lut (.I0(GND_net), .I1(n9929[14]), .I2(GND_net), 
            .I3(n34611), .O(n9125[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3103_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1215_13_lut (.I0(GND_net), .I1(n1801[10]), .I2(GND_net), 
            .I3(n35856), .O(n1800[11])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1215_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1215_13 (.CI(n35856), .I0(n1801[10]), .I1(GND_net), 
            .CO(n35857));
    SB_CARRY add_3103_17 (.CI(n34611), .I0(n9929[14]), .I1(GND_net), .CO(n34612));
    SB_LUT4 add_3059_24_lut (.I0(GND_net), .I1(n8078[21]), .I2(GND_net), 
            .I3(n35319), .O(n8049[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3059_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1215_12_lut (.I0(GND_net), .I1(n1801[9]), .I2(GND_net), 
            .I3(n35855), .O(n1800[10])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1215_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3178_9_lut (.I0(GND_net), .I1(n11531[6]), .I2(GND_net), 
            .I3(n35160), .O(n10852[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3178_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1215_12 (.CI(n35855), .I0(n1801[9]), .I1(GND_net), 
            .CO(n35856));
    SB_LUT4 mult_14_add_1215_11_lut (.I0(GND_net), .I1(n1801[8]), .I2(GND_net), 
            .I3(n35854), .O(n1800[9])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1215_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3103_16_lut (.I0(GND_net), .I1(n9929[13]), .I2(GND_net), 
            .I3(n34610), .O(n9125[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3103_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3103_16 (.CI(n34610), .I0(n9929[13]), .I1(GND_net), .CO(n34611));
    SB_CARRY add_3178_9 (.CI(n35160), .I0(n11531[6]), .I1(GND_net), .CO(n35161));
    SB_LUT4 add_3103_15_lut (.I0(GND_net), .I1(n9929[12]), .I2(GND_net), 
            .I3(n34609), .O(n9125[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3103_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3103_15 (.CI(n34609), .I0(n9929[12]), .I1(GND_net), .CO(n34610));
    SB_CARRY add_3063_12 (.CI(n35405), .I0(n8184[9]), .I1(GND_net), .CO(n35406));
    SB_CARRY add_3059_24 (.CI(n35319), .I0(n8078[21]), .I1(GND_net), .CO(n35320));
    SB_LUT4 add_3103_14_lut (.I0(GND_net), .I1(n9929[11]), .I2(GND_net), 
            .I3(n34608), .O(n9125[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3103_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3178_8_lut (.I0(GND_net), .I1(n11531[5]), .I2(n545), .I3(n35159), 
            .O(n10852[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3178_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3103_14 (.CI(n34608), .I0(n9929[11]), .I1(GND_net), .CO(n34609));
    SB_LUT4 add_3103_13_lut (.I0(GND_net), .I1(n9929[10]), .I2(GND_net), 
            .I3(n34607), .O(n9125[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3103_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3059_23_lut (.I0(GND_net), .I1(n8078[20]), .I2(GND_net), 
            .I3(n35318), .O(n8049[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3059_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3178_8 (.CI(n35159), .I0(n11531[5]), .I1(n545), .CO(n35160));
    SB_CARRY add_3103_13 (.CI(n34607), .I0(n9929[10]), .I1(GND_net), .CO(n34608));
    SB_LUT4 add_3103_12_lut (.I0(GND_net), .I1(n9929[9]), .I2(GND_net), 
            .I3(n34606), .O(n9125[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3103_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3178_7_lut (.I0(GND_net), .I1(n11531[4]), .I2(n472), .I3(n35158), 
            .O(n10852[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3178_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3103_12 (.CI(n34606), .I0(n9929[9]), .I1(GND_net), .CO(n34607));
    SB_LUT4 add_3103_11_lut (.I0(GND_net), .I1(n9929[8]), .I2(GND_net), 
            .I3(n34605), .O(n9125[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3103_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3065_16_lut (.I0(GND_net), .I1(n8231[13]), .I2(GND_net), 
            .I3(n35452), .O(n8208[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3065_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3063_11_lut (.I0(GND_net), .I1(n8184[8]), .I2(GND_net), 
            .I3(n35404), .O(n8159[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3063_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3059_23 (.CI(n35318), .I0(n8078[20]), .I1(GND_net), .CO(n35319));
    SB_CARRY add_3178_7 (.CI(n35158), .I0(n11531[4]), .I1(n472), .CO(n35159));
    SB_LUT4 add_3178_6_lut (.I0(GND_net), .I1(n11531[3]), .I2(n399), .I3(n35157), 
            .O(n10852[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3178_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3059_22_lut (.I0(GND_net), .I1(n8078[19]), .I2(GND_net), 
            .I3(n35317), .O(n8049[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3059_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3178_6 (.CI(n35157), .I0(n11531[3]), .I1(n399), .CO(n35158));
    SB_CARRY mult_14_add_1215_11 (.CI(n35854), .I0(n1801[8]), .I1(GND_net), 
            .CO(n35855));
    SB_LUT4 add_3178_5_lut (.I0(GND_net), .I1(n11531[2]), .I2(n326), .I3(n35156), 
            .O(n10852[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3178_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3103_11 (.CI(n34605), .I0(n9929[8]), .I1(GND_net), .CO(n34606));
    SB_LUT4 add_3103_10_lut (.I0(GND_net), .I1(n9929[7]), .I2(GND_net), 
            .I3(n34604), .O(n9125[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3103_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3178_5 (.CI(n35156), .I0(n11531[2]), .I1(n326), .CO(n35157));
    SB_LUT4 add_3178_4_lut (.I0(GND_net), .I1(n11531[1]), .I2(n253), .I3(n35155), 
            .O(n10852[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3178_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1215_10_lut (.I0(GND_net), .I1(n1801[7]), .I2(GND_net), 
            .I3(n35853), .O(n1800[8])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1215_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3103_10 (.CI(n34604), .I0(n9929[7]), .I1(GND_net), .CO(n34605));
    SB_CARRY add_3063_11 (.CI(n35404), .I0(n8184[8]), .I1(GND_net), .CO(n35405));
    SB_CARRY add_3059_22 (.CI(n35317), .I0(n8078[19]), .I1(GND_net), .CO(n35318));
    SB_CARRY add_3178_4 (.CI(n35155), .I0(n11531[1]), .I1(n253), .CO(n35156));
    SB_LUT4 add_3103_9_lut (.I0(GND_net), .I1(n9929[6]), .I2(GND_net), 
            .I3(n34603), .O(n9125[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3103_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3103_9 (.CI(n34603), .I0(n9929[6]), .I1(GND_net), .CO(n34604));
    SB_LUT4 add_3059_21_lut (.I0(GND_net), .I1(n8078[18]), .I2(GND_net), 
            .I3(n35316), .O(n8049[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3059_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3103_8_lut (.I0(GND_net), .I1(n9929[5]), .I2(n689_adj_3710), 
            .I3(n34602), .O(n9125[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3103_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3178_3_lut (.I0(GND_net), .I1(n11531[0]), .I2(n180), .I3(n35154), 
            .O(n10852[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3178_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3178_3 (.CI(n35154), .I0(n11531[0]), .I1(n180), .CO(n35155));
    SB_CARRY add_3103_8 (.CI(n34602), .I0(n9929[5]), .I1(n689_adj_3710), 
            .CO(n34603));
    SB_LUT4 add_3103_7_lut (.I0(GND_net), .I1(n9929[4]), .I2(n592_adj_3711), 
            .I3(n34601), .O(n9125[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3103_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3103_7 (.CI(n34601), .I0(n9929[4]), .I1(n592_adj_3711), 
            .CO(n34602));
    SB_CARRY add_3059_21 (.CI(n35316), .I0(n8078[18]), .I1(GND_net), .CO(n35317));
    SB_LUT4 add_3178_2_lut (.I0(GND_net), .I1(n35), .I2(n107), .I3(GND_net), 
            .O(n10852[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3178_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3103_6_lut (.I0(GND_net), .I1(n9929[3]), .I2(n495_adj_3712), 
            .I3(n34600), .O(n9125[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3103_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3103_6 (.CI(n34600), .I0(n9929[3]), .I1(n495_adj_3712), 
            .CO(n34601));
    SB_CARRY add_3178_2 (.CI(GND_net), .I0(n35), .I1(n107), .CO(n35154));
    SB_LUT4 add_3103_5_lut (.I0(GND_net), .I1(n9929[2]), .I2(n398_adj_3713), 
            .I3(n34599), .O(n9125[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3103_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3059_20_lut (.I0(GND_net), .I1(n8078[17]), .I2(GND_net), 
            .I3(n35315), .O(n8049[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3059_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3103_5 (.CI(n34599), .I0(n9929[2]), .I1(n398_adj_3713), 
            .CO(n34600));
    SB_CARRY add_3065_16 (.CI(n35452), .I0(n8231[13]), .I1(GND_net), .CO(n35453));
    SB_CARRY add_3067_15 (.CI(n35490), .I0(n8274[12]), .I1(GND_net), .CO(n35491));
    SB_CARRY mult_14_add_1215_10 (.CI(n35853), .I0(n1801[7]), .I1(GND_net), 
            .CO(n35854));
    SB_LUT4 add_3065_15_lut (.I0(GND_net), .I1(n8231[12]), .I2(GND_net), 
            .I3(n35451), .O(n8208[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3065_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1215_9_lut (.I0(GND_net), .I1(n1801[6]), .I2(GND_net), 
            .I3(n35852), .O(n1800[7])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1215_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3063_10_lut (.I0(GND_net), .I1(n8184[7]), .I2(GND_net), 
            .I3(n35403), .O(n8159[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3063_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1215_9 (.CI(n35852), .I0(n1801[6]), .I1(GND_net), 
            .CO(n35853));
    SB_CARRY add_3059_20 (.CI(n35315), .I0(n8078[17]), .I1(GND_net), .CO(n35316));
    SB_LUT4 mult_14_add_1215_8_lut (.I0(GND_net), .I1(n1801[5]), .I2(n524), 
            .I3(n35851), .O(n1800[6])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1215_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3205_18_lut (.I0(GND_net), .I1(n12157[15]), .I2(GND_net), 
            .I3(n35153), .O(n11531[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3205_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1215_8 (.CI(n35851), .I0(n1801[5]), .I1(n524), 
            .CO(n35852));
    SB_LUT4 add_3205_17_lut (.I0(GND_net), .I1(n12157[14]), .I2(GND_net), 
            .I3(n35152), .O(n11531[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3205_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3059_19_lut (.I0(GND_net), .I1(n8078[16]), .I2(GND_net), 
            .I3(n35314), .O(n8049[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3059_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3205_17 (.CI(n35152), .I0(n12157[14]), .I1(GND_net), 
            .CO(n35153));
    SB_LUT4 add_3205_16_lut (.I0(GND_net), .I1(n12157[13]), .I2(GND_net), 
            .I3(n35151), .O(n11531[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3205_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3063_10 (.CI(n35403), .I0(n8184[7]), .I1(GND_net), .CO(n35404));
    SB_LUT4 add_3063_9_lut (.I0(GND_net), .I1(n8184[6]), .I2(GND_net), 
            .I3(n35402), .O(n8159[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3063_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1215_7_lut (.I0(GND_net), .I1(n1801[4]), .I2(n451), 
            .I3(n35850), .O(n1800[5])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1215_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3059_19 (.CI(n35314), .I0(n8078[16]), .I1(GND_net), .CO(n35315));
    SB_CARRY mult_14_add_1215_7 (.CI(n35850), .I0(n1801[4]), .I1(n451), 
            .CO(n35851));
    SB_CARRY add_3205_16 (.CI(n35151), .I0(n12157[13]), .I1(GND_net), 
            .CO(n35152));
    SB_LUT4 mult_14_add_1215_6_lut (.I0(GND_net), .I1(n1801[3]), .I2(n378), 
            .I3(n35849), .O(n1800[4])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1215_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3205_15_lut (.I0(GND_net), .I1(n12157[12]), .I2(GND_net), 
            .I3(n35150), .O(n11531[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3205_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1215_6 (.CI(n35849), .I0(n1801[3]), .I1(n378), 
            .CO(n35850));
    SB_LUT4 add_3059_18_lut (.I0(GND_net), .I1(n8078[15]), .I2(GND_net), 
            .I3(n35313), .O(n8049[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3059_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1215_5_lut (.I0(GND_net), .I1(n1801[2]), .I2(n305), 
            .I3(n35848), .O(n1800[3])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1215_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3205_15 (.CI(n35150), .I0(n12157[12]), .I1(GND_net), 
            .CO(n35151));
    SB_LUT4 add_3205_14_lut (.I0(GND_net), .I1(n12157[11]), .I2(GND_net), 
            .I3(n35149), .O(n11531[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3205_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3065_15 (.CI(n35451), .I0(n8231[12]), .I1(GND_net), .CO(n35452));
    SB_CARRY add_3063_9 (.CI(n35402), .I0(n8184[6]), .I1(GND_net), .CO(n35403));
    SB_CARRY add_3059_18 (.CI(n35313), .I0(n8078[15]), .I1(GND_net), .CO(n35314));
    SB_LUT4 add_3059_17_lut (.I0(GND_net), .I1(n8078[14]), .I2(GND_net), 
            .I3(n35312), .O(n8049[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3059_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3205_14 (.CI(n35149), .I0(n12157[11]), .I1(GND_net), 
            .CO(n35150));
    SB_CARRY mult_14_add_1215_5 (.CI(n35848), .I0(n1801[2]), .I1(n305), 
            .CO(n35849));
    SB_LUT4 mult_14_add_1215_4_lut (.I0(GND_net), .I1(n1801[1]), .I2(n232_adj_3718), 
            .I3(n35847), .O(n1800[2])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1215_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1215_4 (.CI(n35847), .I0(n1801[1]), .I1(n232_adj_3718), 
            .CO(n35848));
    SB_LUT4 add_3205_13_lut (.I0(GND_net), .I1(n12157[10]), .I2(GND_net), 
            .I3(n35148), .O(n11531[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3205_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1215_3_lut (.I0(GND_net), .I1(n1801[0]), .I2(n159), 
            .I3(n35846), .O(n1800[1])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1215_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1215_3 (.CI(n35846), .I0(n1801[0]), .I1(n159), 
            .CO(n35847));
    SB_CARRY add_3059_17 (.CI(n35312), .I0(n8078[14]), .I1(GND_net), .CO(n35313));
    SB_LUT4 mult_14_add_1215_2_lut (.I0(GND_net), .I1(n17_adj_3719), .I2(n86_adj_3720), 
            .I3(GND_net), .O(n1800[0])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1215_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3205_13 (.CI(n35148), .I0(n12157[10]), .I1(GND_net), 
            .CO(n35149));
    SB_LUT4 add_3059_16_lut (.I0(GND_net), .I1(n8078[13]), .I2(GND_net), 
            .I3(n35311), .O(n8049[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3059_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3205_12_lut (.I0(GND_net), .I1(n12157[9]), .I2(GND_net), 
            .I3(n35147), .O(n11531[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3205_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1215_2 (.CI(GND_net), .I0(n17_adj_3719), .I1(n86_adj_3720), 
            .CO(n35846));
    SB_LUT4 mult_14_add_1214_24_lut (.I0(GND_net), .I1(n1800[21]), .I2(GND_net), 
            .I3(n35844), .O(n1799[22])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1214_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_12_i140_2_lut (.I0(\Kd[2] ), .I1(n57[4]), .I2(GND_net), 
            .I3(GND_net), .O(n207));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i140_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY mult_14_add_1214_24 (.CI(n35844), .I0(n1800[21]), .I1(GND_net), 
            .CO(n1695));
    SB_LUT4 add_3063_8_lut (.I0(GND_net), .I1(n8184[5]), .I2(n704_adj_3721), 
            .I3(n35401), .O(n8159[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3063_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3103_4_lut (.I0(GND_net), .I1(n9929[1]), .I2(n301_adj_3722), 
            .I3(n34598), .O(n9125[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3103_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1214_23_lut (.I0(GND_net), .I1(n1800[20]), .I2(GND_net), 
            .I3(n35843), .O(n1799[21])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1214_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3103_4 (.CI(n34598), .I0(n9929[1]), .I1(n301_adj_3722), 
            .CO(n34599));
    SB_CARRY add_3059_16 (.CI(n35311), .I0(n8078[13]), .I1(GND_net), .CO(n35312));
    SB_CARRY add_3205_12 (.CI(n35147), .I0(n12157[9]), .I1(GND_net), .CO(n35148));
    SB_LUT4 add_3070_7_lut (.I0(GND_net), .I1(n8331[4]), .I2(n628), .I3(n35533), 
            .O(n8313[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3070_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3205_11_lut (.I0(GND_net), .I1(n12157[8]), .I2(GND_net), 
            .I3(n35146), .O(n11531[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3205_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3103_3_lut (.I0(GND_net), .I1(n9929[0]), .I2(n204_adj_3723), 
            .I3(n34597), .O(n9125[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3103_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1214_23 (.CI(n35843), .I0(n1800[20]), .I1(GND_net), 
            .CO(n35844));
    SB_LUT4 mult_14_add_1214_22_lut (.I0(GND_net), .I1(n1800[19]), .I2(GND_net), 
            .I3(n35842), .O(n1799[20])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1214_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1214_22 (.CI(n35842), .I0(n1800[19]), .I1(GND_net), 
            .CO(n35843));
    SB_LUT4 mult_14_add_1214_21_lut (.I0(GND_net), .I1(n1800[18]), .I2(GND_net), 
            .I3(n35841), .O(n1799[19])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1214_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_12_i105_2_lut (.I0(\Kd[1] ), .I1(n57[19]), .I2(GND_net), 
            .I3(GND_net), .O(n155_adj_3414));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i105_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i42_2_lut (.I0(\Kd[0] ), .I1(n57[20]), .I2(GND_net), 
            .I3(GND_net), .O(n62));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i42_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY mult_14_add_1214_21 (.CI(n35841), .I0(n1800[18]), .I1(GND_net), 
            .CO(n35842));
    SB_CARRY add_3205_11 (.CI(n35146), .I0(n12157[8]), .I1(GND_net), .CO(n35147));
    SB_LUT4 add_3205_10_lut (.I0(GND_net), .I1(n12157[7]), .I2(GND_net), 
            .I3(n35145), .O(n11531[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3205_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3059_15_lut (.I0(GND_net), .I1(n8078[12]), .I2(GND_net), 
            .I3(n35310), .O(n8049[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3059_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3205_10 (.CI(n35145), .I0(n12157[7]), .I1(GND_net), .CO(n35146));
    SB_LUT4 add_13_add_1_20061_add_1_33_lut (.I0(GND_net), .I1(n7065[8]), 
            .I2(n5786[0]), .I3(n34886), .O(n63[31])) /* synthesis syn_instantiated=1 */ ;
    defparam add_13_add_1_20061_add_1_33_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_13_add_1_20061_add_1_32_lut (.I0(GND_net), .I1(n7065[7]), 
            .I2(n61[30]), .I3(n34885), .O(n63[30])) /* synthesis syn_instantiated=1 */ ;
    defparam add_13_add_1_20061_add_1_32_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_13_add_1_20061_add_1_32 (.CI(n34885), .I0(n7065[7]), .I1(n61[30]), 
            .CO(n34886));
    SB_LUT4 add_3205_9_lut (.I0(GND_net), .I1(n12157[6]), .I2(GND_net), 
            .I3(n35144), .O(n11531[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3205_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3103_3 (.CI(n34597), .I0(n9929[0]), .I1(n204_adj_3723), 
            .CO(n34598));
    SB_LUT4 add_13_add_1_20061_add_1_31_lut (.I0(GND_net), .I1(n7065[6]), 
            .I2(n61[29]), .I3(n34884), .O(n63[29])) /* synthesis syn_instantiated=1 */ ;
    defparam add_13_add_1_20061_add_1_31_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_13_add_1_20061_add_1_31 (.CI(n34884), .I0(n7065[6]), .I1(n61[29]), 
            .CO(n34885));
    SB_LUT4 add_3103_2_lut (.I0(GND_net), .I1(n14_adj_3724), .I2(n107_adj_3725), 
            .I3(GND_net), .O(n9125[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3103_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1214_20_lut (.I0(GND_net), .I1(n1800[17]), .I2(GND_net), 
            .I3(n35840), .O(n1799[18])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1214_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3067_14_lut (.I0(GND_net), .I1(n8274[11]), .I2(GND_net), 
            .I3(n35489), .O(n8253[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3067_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_13_add_1_20061_add_1_30_lut (.I0(GND_net), .I1(n7065[5]), 
            .I2(n61[28]), .I3(n34883), .O(n63[28])) /* synthesis syn_instantiated=1 */ ;
    defparam add_13_add_1_20061_add_1_30_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3065_14_lut (.I0(GND_net), .I1(n8231[11]), .I2(GND_net), 
            .I3(n35450), .O(n8208[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3065_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3063_8 (.CI(n35401), .I0(n8184[5]), .I1(n704_adj_3721), 
            .CO(n35402));
    SB_CARRY add_3059_15 (.CI(n35310), .I0(n8078[12]), .I1(GND_net), .CO(n35311));
    SB_CARRY add_3205_9 (.CI(n35144), .I0(n12157[6]), .I1(GND_net), .CO(n35145));
    SB_CARRY add_3070_7 (.CI(n35533), .I0(n8331[4]), .I1(n628), .CO(n35534));
    SB_LUT4 add_3205_8_lut (.I0(GND_net), .I1(n12157[5]), .I2(n545), .I3(n35143), 
            .O(n11531[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3205_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3067_14 (.CI(n35489), .I0(n8274[11]), .I1(GND_net), .CO(n35490));
    SB_CARRY mult_14_add_1214_20 (.CI(n35840), .I0(n1800[17]), .I1(GND_net), 
            .CO(n35841));
    SB_LUT4 mult_14_add_1214_19_lut (.I0(GND_net), .I1(n1800[16]), .I2(GND_net), 
            .I3(n35839), .O(n1799[17])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1214_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1214_19 (.CI(n35839), .I0(n1800[16]), .I1(GND_net), 
            .CO(n35840));
    SB_LUT4 mult_14_add_1214_18_lut (.I0(GND_net), .I1(n1800[15]), .I2(GND_net), 
            .I3(n35838), .O(n1799[16])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1214_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1214_18 (.CI(n35838), .I0(n1800[15]), .I1(GND_net), 
            .CO(n35839));
    SB_LUT4 mult_14_add_1214_17_lut (.I0(GND_net), .I1(n1800[14]), .I2(GND_net), 
            .I3(n35837), .O(n1799[15])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1214_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1214_17 (.CI(n35837), .I0(n1800[14]), .I1(GND_net), 
            .CO(n35838));
    SB_LUT4 mult_14_add_1214_16_lut (.I0(GND_net), .I1(n1800[13]), .I2(GND_net), 
            .I3(n35836), .O(n1799[14])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1214_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1214_16 (.CI(n35836), .I0(n1800[13]), .I1(GND_net), 
            .CO(n35837));
    SB_LUT4 mult_14_add_1214_15_lut (.I0(GND_net), .I1(n1800[12]), .I2(GND_net), 
            .I3(n35835), .O(n1799[13])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1214_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1214_15 (.CI(n35835), .I0(n1800[12]), .I1(GND_net), 
            .CO(n35836));
    SB_LUT4 mult_14_add_1214_14_lut (.I0(GND_net), .I1(n1800[11]), .I2(GND_net), 
            .I3(n35834), .O(n1799[12])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1214_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3059_14_lut (.I0(GND_net), .I1(n8078[11]), .I2(GND_net), 
            .I3(n35309), .O(n8049[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3059_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1214_14 (.CI(n35834), .I0(n1800[11]), .I1(GND_net), 
            .CO(n35835));
    SB_LUT4 mult_14_add_1214_13_lut (.I0(GND_net), .I1(n1800[10]), .I2(GND_net), 
            .I3(n35833), .O(n1799[11])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1214_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3205_8 (.CI(n35143), .I0(n12157[5]), .I1(n545), .CO(n35144));
    SB_CARRY mult_14_add_1214_13 (.CI(n35833), .I0(n1800[10]), .I1(GND_net), 
            .CO(n35834));
    SB_LUT4 mult_14_add_1214_12_lut (.I0(GND_net), .I1(n1800[9]), .I2(GND_net), 
            .I3(n35832), .O(n1799[10])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1214_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3205_7_lut (.I0(GND_net), .I1(n12157[4]), .I2(n472), .I3(n35142), 
            .O(n11531[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3205_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1214_12 (.CI(n35832), .I0(n1800[9]), .I1(GND_net), 
            .CO(n35833));
    SB_LUT4 mult_14_add_1214_11_lut (.I0(GND_net), .I1(n1800[8]), .I2(GND_net), 
            .I3(n35831), .O(n1799[9])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1214_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1214_11 (.CI(n35831), .I0(n1800[8]), .I1(GND_net), 
            .CO(n35832));
    SB_DFF \PID_CONTROLLER.err_prev__i2  (.Q(\PID_CONTROLLER.err_prev[1] ), 
           .C(clk32MHz), .D(n23746));   // verilog/motorControl.v(38[14] 59[8])
    SB_LUT4 mult_14_add_1214_10_lut (.I0(GND_net), .I1(n1800[7]), .I2(GND_net), 
            .I3(n35830), .O(n1799[8])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1214_10_lut.LUT_INIT = 16'hC33C;
    SB_DFF \PID_CONTROLLER.err_prev__i3  (.Q(\PID_CONTROLLER.err_prev[2] ), 
           .C(clk32MHz), .D(n23745));   // verilog/motorControl.v(38[14] 59[8])
    SB_DFF \PID_CONTROLLER.err_prev__i4  (.Q(\PID_CONTROLLER.err_prev[3] ), 
           .C(clk32MHz), .D(n23744));   // verilog/motorControl.v(38[14] 59[8])
    SB_LUT4 add_3070_6_lut (.I0(GND_net), .I1(n8331[3]), .I2(n531_adj_3726), 
            .I3(n35532), .O(n8313[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3070_6_lut.LUT_INIT = 16'hC33C;
    SB_DFF \PID_CONTROLLER.err_prev__i5  (.Q(\PID_CONTROLLER.err_prev[4] ), 
           .C(clk32MHz), .D(n23743));   // verilog/motorControl.v(38[14] 59[8])
    SB_CARRY mult_14_add_1214_10 (.CI(n35830), .I0(n1800[7]), .I1(GND_net), 
            .CO(n35831));
    SB_CARRY add_3205_7 (.CI(n35142), .I0(n12157[4]), .I1(n472), .CO(n35143));
    SB_LUT4 mult_14_add_1214_9_lut (.I0(GND_net), .I1(n1800[6]), .I2(GND_net), 
            .I3(n35829), .O(n1799[7])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1214_9_lut.LUT_INIT = 16'hC33C;
    SB_DFF \PID_CONTROLLER.err_prev__i6  (.Q(\PID_CONTROLLER.err_prev[5] ), 
           .C(clk32MHz), .D(n23742));   // verilog/motorControl.v(38[14] 59[8])
    SB_CARRY mult_14_add_1214_9 (.CI(n35829), .I0(n1800[6]), .I1(GND_net), 
            .CO(n35830));
    SB_DFF \PID_CONTROLLER.err_prev__i7  (.Q(\PID_CONTROLLER.err_prev[6] ), 
           .C(clk32MHz), .D(n23741));   // verilog/motorControl.v(38[14] 59[8])
    SB_DFF \PID_CONTROLLER.err_prev__i8  (.Q(\PID_CONTROLLER.err_prev[7] ), 
           .C(clk32MHz), .D(n23740));   // verilog/motorControl.v(38[14] 59[8])
    SB_DFF \PID_CONTROLLER.err_prev__i9  (.Q(\PID_CONTROLLER.err_prev[8] ), 
           .C(clk32MHz), .D(n23739));   // verilog/motorControl.v(38[14] 59[8])
    SB_LUT4 add_3063_7_lut (.I0(GND_net), .I1(n8184[4]), .I2(n607_adj_3728), 
            .I3(n35400), .O(n8159[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3063_7_lut.LUT_INIT = 16'hC33C;
    SB_DFF \PID_CONTROLLER.err_prev__i10  (.Q(\PID_CONTROLLER.err_prev[9] ), 
           .C(clk32MHz), .D(n23738));   // verilog/motorControl.v(38[14] 59[8])
    SB_DFF \PID_CONTROLLER.err_prev__i11  (.Q(\PID_CONTROLLER.err_prev[10] ), 
           .C(clk32MHz), .D(n23737));   // verilog/motorControl.v(38[14] 59[8])
    SB_LUT4 mult_14_add_1214_8_lut (.I0(GND_net), .I1(n1800[5]), .I2(n521), 
            .I3(n35828), .O(n1799[6])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1214_8_lut.LUT_INIT = 16'hC33C;
    SB_DFF \PID_CONTROLLER.err_prev__i12  (.Q(\PID_CONTROLLER.err_prev[11] ), 
           .C(clk32MHz), .D(n23736));   // verilog/motorControl.v(38[14] 59[8])
    SB_DFF \PID_CONTROLLER.err_prev__i13  (.Q(\PID_CONTROLLER.err_prev[12] ), 
           .C(clk32MHz), .D(n23735));   // verilog/motorControl.v(38[14] 59[8])
    SB_DFF \PID_CONTROLLER.err_prev__i14  (.Q(\PID_CONTROLLER.err_prev[13] ), 
           .C(clk32MHz), .D(n23734));   // verilog/motorControl.v(38[14] 59[8])
    SB_DFF \PID_CONTROLLER.err_prev__i15  (.Q(\PID_CONTROLLER.err_prev[14] ), 
           .C(clk32MHz), .D(n23733));   // verilog/motorControl.v(38[14] 59[8])
    SB_DFF \PID_CONTROLLER.err_prev__i16  (.Q(\PID_CONTROLLER.err_prev[15] ), 
           .C(clk32MHz), .D(n23732));   // verilog/motorControl.v(38[14] 59[8])
    SB_DFF \PID_CONTROLLER.err_prev__i17  (.Q(\PID_CONTROLLER.err_prev[16] ), 
           .C(clk32MHz), .D(n23731));   // verilog/motorControl.v(38[14] 59[8])
    SB_DFF \PID_CONTROLLER.err_prev__i18  (.Q(\PID_CONTROLLER.err_prev[17] ), 
           .C(clk32MHz), .D(n23730));   // verilog/motorControl.v(38[14] 59[8])
    SB_CARRY add_13_add_1_20061_add_1_30 (.CI(n34883), .I0(n7065[5]), .I1(n61[28]), 
            .CO(n34884));
    SB_DFF \PID_CONTROLLER.err_prev__i19  (.Q(\PID_CONTROLLER.err_prev[18] ), 
           .C(clk32MHz), .D(n23729));   // verilog/motorControl.v(38[14] 59[8])
    SB_CARRY add_3103_2 (.CI(GND_net), .I0(n14_adj_3724), .I1(n107_adj_3725), 
            .CO(n34597));
    SB_DFF \PID_CONTROLLER.err_prev__i20  (.Q(\PID_CONTROLLER.err_prev[19] ), 
           .C(clk32MHz), .D(n23728));   // verilog/motorControl.v(38[14] 59[8])
    SB_DFF \PID_CONTROLLER.err_prev__i21  (.Q(\PID_CONTROLLER.err_prev[20] ), 
           .C(clk32MHz), .D(n23727));   // verilog/motorControl.v(38[14] 59[8])
    SB_DFF \PID_CONTROLLER.err_prev__i22  (.Q(\PID_CONTROLLER.err_prev[21] ), 
           .C(clk32MHz), .D(n23726));   // verilog/motorControl.v(38[14] 59[8])
    SB_DFF \PID_CONTROLLER.err_prev__i23  (.Q(\PID_CONTROLLER.err_prev[22] ), 
           .C(clk32MHz), .D(n23725));   // verilog/motorControl.v(38[14] 59[8])
    SB_DFF \PID_CONTROLLER.err_prev__i24  (.Q(\PID_CONTROLLER.err_prev[23] ), 
           .C(clk32MHz), .D(n23724));   // verilog/motorControl.v(38[14] 59[8])
    SB_DFF \PID_CONTROLLER.err_prev__i25  (.Q(\PID_CONTROLLER.err_prev[31] ), 
           .C(clk32MHz), .D(n23723));   // verilog/motorControl.v(38[14] 59[8])
    SB_LUT4 add_3205_6_lut (.I0(GND_net), .I1(n12157[3]), .I2(n399), .I3(n35141), 
            .O(n11531[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3205_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_13_add_1_20061_add_1_29_lut (.I0(GND_net), .I1(n7065[4]), 
            .I2(n61[27]), .I3(n34882), .O(n63[27])) /* synthesis syn_instantiated=1 */ ;
    defparam add_13_add_1_20061_add_1_29_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3301_14_lut (.I0(GND_net), .I1(n14168[11]), .I2(GND_net), 
            .I3(n34596), .O(n13734[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3301_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3059_14 (.CI(n35309), .I0(n8078[11]), .I1(GND_net), .CO(n35310));
    SB_CARRY add_3205_6 (.CI(n35141), .I0(n12157[3]), .I1(n399), .CO(n35142));
    SB_LUT4 add_3205_5_lut (.I0(GND_net), .I1(n12157[2]), .I2(n326), .I3(n35140), 
            .O(n11531[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3205_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1214_8 (.CI(n35828), .I0(n1800[5]), .I1(n521), 
            .CO(n35829));
    SB_CARRY add_3063_7 (.CI(n35400), .I0(n8184[4]), .I1(n607_adj_3728), 
            .CO(n35401));
    SB_LUT4 add_3059_13_lut (.I0(GND_net), .I1(n8078[10]), .I2(GND_net), 
            .I3(n35308), .O(n8049[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3059_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3205_5 (.CI(n35140), .I0(n12157[2]), .I1(n326), .CO(n35141));
    SB_CARRY add_3059_13 (.CI(n35308), .I0(n8078[10]), .I1(GND_net), .CO(n35309));
    SB_CARRY add_13_add_1_20061_add_1_29 (.CI(n34882), .I0(n7065[4]), .I1(n61[27]), 
            .CO(n34883));
    SB_LUT4 add_13_add_1_20061_add_1_28_lut (.I0(GND_net), .I1(n7065[3]), 
            .I2(n61[26]), .I3(n34881), .O(n63[26])) /* synthesis syn_instantiated=1 */ ;
    defparam add_13_add_1_20061_add_1_28_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1214_7_lut (.I0(GND_net), .I1(n1800[4]), .I2(n448), 
            .I3(n35827), .O(n1799[5])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1214_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3205_4_lut (.I0(GND_net), .I1(n12157[1]), .I2(n253), .I3(n35139), 
            .O(n11531[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3205_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_13_add_1_20061_add_1_28 (.CI(n34881), .I0(n7065[3]), .I1(n61[26]), 
            .CO(n34882));
    SB_LUT4 add_13_add_1_20061_add_1_27_lut (.I0(GND_net), .I1(n7065[2]), 
            .I2(n61[25]), .I3(n34880), .O(n63[25])) /* synthesis syn_instantiated=1 */ ;
    defparam add_13_add_1_20061_add_1_27_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_13_add_1_20061_add_1_27 (.CI(n34880), .I0(n7065[2]), .I1(n61[25]), 
            .CO(n34881));
    SB_CARRY add_3205_4 (.CI(n35139), .I0(n12157[1]), .I1(n253), .CO(n35140));
    SB_LUT4 add_3059_12_lut (.I0(GND_net), .I1(n8078[9]), .I2(GND_net), 
            .I3(n35307), .O(n8049[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3059_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_13_add_1_20061_add_1_26_lut (.I0(GND_net), .I1(n7065[1]), 
            .I2(n61[24]), .I3(n34879), .O(n63[24])) /* synthesis syn_instantiated=1 */ ;
    defparam add_13_add_1_20061_add_1_26_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3065_14 (.CI(n35450), .I0(n8231[11]), .I1(GND_net), .CO(n35451));
    SB_DFF \PID_CONTROLLER.result_i1  (.Q(\PID_CONTROLLER.result [1]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.result_31__N_3003 [1]));   // verilog/motorControl.v(38[14] 59[8])
    SB_LUT4 add_3301_13_lut (.I0(GND_net), .I1(n14168[10]), .I2(GND_net), 
            .I3(n34595), .O(n13734[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3301_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3063_6_lut (.I0(GND_net), .I1(n8184[3]), .I2(n510_adj_3731), 
            .I3(n35399), .O(n8159[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3063_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1214_7 (.CI(n35827), .I0(n1800[4]), .I1(n448), 
            .CO(n35828));
    SB_CARRY add_3301_13 (.CI(n34595), .I0(n14168[10]), .I1(GND_net), 
            .CO(n34596));
    SB_CARRY add_3074_10 (.CI(n35590), .I0(n8393[7]), .I1(GND_net), .CO(n35591));
    SB_CARRY add_3059_12 (.CI(n35307), .I0(n8078[9]), .I1(GND_net), .CO(n35308));
    SB_LUT4 mult_14_add_1214_6_lut (.I0(GND_net), .I1(n1800[3]), .I2(n375), 
            .I3(n35826), .O(n1799[4])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1214_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1214_6 (.CI(n35826), .I0(n1800[3]), .I1(n375), 
            .CO(n35827));
    SB_LUT4 mult_14_add_1214_5_lut (.I0(GND_net), .I1(n1800[2]), .I2(n302), 
            .I3(n35825), .O(n1799[3])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1214_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1214_5 (.CI(n35825), .I0(n1800[2]), .I1(n302), 
            .CO(n35826));
    SB_LUT4 add_3301_12_lut (.I0(GND_net), .I1(n14168[9]), .I2(GND_net), 
            .I3(n34594), .O(n13734[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3301_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3205_3_lut (.I0(GND_net), .I1(n12157[0]), .I2(n180), .I3(n35138), 
            .O(n11531[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3205_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3074_9_lut (.I0(GND_net), .I1(n8393[6]), .I2(GND_net), 
            .I3(n35589), .O(n8379[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3074_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_13_add_1_20061_add_1_26 (.CI(n34879), .I0(n7065[1]), .I1(n61[24]), 
            .CO(n34880));
    SB_CARRY add_3301_12 (.CI(n34594), .I0(n14168[9]), .I1(GND_net), .CO(n34595));
    SB_LUT4 mult_14_add_1214_4_lut (.I0(GND_net), .I1(n1800[1]), .I2(n229_adj_3733), 
            .I3(n35824), .O(n1799[2])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1214_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1214_4 (.CI(n35824), .I0(n1800[1]), .I1(n229_adj_3733), 
            .CO(n35825));
    SB_LUT4 mult_14_add_1214_3_lut (.I0(GND_net), .I1(n1800[0]), .I2(n156_adj_3735), 
            .I3(n35823), .O(n1799[1])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1214_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3074_9 (.CI(n35589), .I0(n8393[6]), .I1(GND_net), .CO(n35590));
    SB_CARRY add_3070_6 (.CI(n35532), .I0(n8331[3]), .I1(n531_adj_3726), 
            .CO(n35533));
    SB_LUT4 state_23__I_0_add_2_26_lut (.I0(GND_net), .I1(\motor_state[23] ), 
            .I2(n58[23]), .I3(n34239), .O(\PID_CONTROLLER.err_31__N_2825 [24])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_26_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3205_3 (.CI(n35138), .I0(n12157[0]), .I1(n180), .CO(n35139));
    SB_LUT4 state_23__I_0_add_2_25_lut (.I0(GND_net), .I1(\motor_state[23] ), 
            .I2(n58[23]), .I3(n34238), .O(\PID_CONTROLLER.err_31__N_2825 [23])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_13_add_1_20061_add_1_25_lut (.I0(GND_net), .I1(n7065[0]), 
            .I2(n61[23]), .I3(n34878), .O(n63[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_13_add_1_20061_add_1_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_13_add_1_20061_add_1_25 (.CI(n34878), .I0(n7065[0]), .I1(n61[23]), 
            .CO(n34879));
    SB_LUT4 add_13_add_1_20061_add_1_24_lut (.I0(GND_net), .I1(n282[22]), 
            .I2(n61[22]), .I3(n34877), .O(n63[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_13_add_1_20061_add_1_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3205_2_lut (.I0(GND_net), .I1(n35), .I2(n107), .I3(GND_net), 
            .O(n11531[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3205_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3301_11_lut (.I0(GND_net), .I1(n14168[8]), .I2(GND_net), 
            .I3(n34593), .O(n13734[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3301_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_13_add_1_20061_add_1_24 (.CI(n34877), .I0(n282[22]), .I1(n61[22]), 
            .CO(n34878));
    SB_LUT4 add_13_add_1_20061_add_1_23_lut (.I0(GND_net), .I1(n282[21]), 
            .I2(n61[21]), .I3(n34876), .O(n63[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_13_add_1_20061_add_1_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1214_3 (.CI(n35823), .I0(n1800[0]), .I1(n156_adj_3735), 
            .CO(n35824));
    SB_LUT4 mult_14_add_1214_2_lut (.I0(GND_net), .I1(n14_adj_3738), .I2(n83), 
            .I3(GND_net), .O(n1799[0])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1214_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1214_2 (.CI(GND_net), .I0(n14_adj_3738), .I1(n83), 
            .CO(n35823));
    SB_LUT4 mult_14_add_1213_24_lut (.I0(GND_net), .I1(n1799[21]), .I2(GND_net), 
            .I3(n35821), .O(n1798[22])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1213_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1213_24 (.CI(n35821), .I0(n1799[21]), .I1(GND_net), 
            .CO(n1691));
    SB_LUT4 mult_14_add_1213_23_lut (.I0(GND_net), .I1(n1799[20]), .I2(GND_net), 
            .I3(n35820), .O(n1798[21])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1213_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1213_23 (.CI(n35820), .I0(n1799[20]), .I1(GND_net), 
            .CO(n35821));
    SB_LUT4 mult_14_add_1213_22_lut (.I0(GND_net), .I1(n1799[19]), .I2(GND_net), 
            .I3(n35819), .O(n1798[20])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1213_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1213_22 (.CI(n35819), .I0(n1799[19]), .I1(GND_net), 
            .CO(n35820));
    SB_LUT4 mult_14_add_1213_21_lut (.I0(GND_net), .I1(n1799[18]), .I2(GND_net), 
            .I3(n35818), .O(n1798[19])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1213_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_12_i148_2_lut (.I0(\Kd[2] ), .I1(n57[8]), .I2(GND_net), 
            .I3(GND_net), .O(n219));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i148_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY state_23__I_0_add_2_25 (.CI(n34238), .I0(\motor_state[23] ), 
            .I1(n58[23]), .CO(n34239));
    SB_CARRY mult_14_add_1213_21 (.CI(n35818), .I0(n1799[18]), .I1(GND_net), 
            .CO(n35819));
    SB_DFF \PID_CONTROLLER.result_i2  (.Q(\PID_CONTROLLER.result [2]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.result_31__N_3003 [2]));   // verilog/motorControl.v(38[14] 59[8])
    SB_DFF \PID_CONTROLLER.result_i3  (.Q(\PID_CONTROLLER.result [3]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.result_31__N_3003 [3]));   // verilog/motorControl.v(38[14] 59[8])
    SB_DFF \PID_CONTROLLER.result_i4  (.Q(\PID_CONTROLLER.result [4]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.result_31__N_3003 [4]));   // verilog/motorControl.v(38[14] 59[8])
    SB_DFF \PID_CONTROLLER.result_i5  (.Q(\PID_CONTROLLER.result[5] ), .C(clk32MHz), 
           .D(\PID_CONTROLLER.result_31__N_3003 [5]));   // verilog/motorControl.v(38[14] 59[8])
    SB_DFF \PID_CONTROLLER.result_i6  (.Q(\PID_CONTROLLER.result[6] ), .C(clk32MHz), 
           .D(\PID_CONTROLLER.result_31__N_3003 [6]));   // verilog/motorControl.v(38[14] 59[8])
    SB_DFF \PID_CONTROLLER.result_i7  (.Q(\PID_CONTROLLER.result [7]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.result_31__N_3003 [7]));   // verilog/motorControl.v(38[14] 59[8])
    SB_DFF \PID_CONTROLLER.result_i8  (.Q(\PID_CONTROLLER.result [8]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.result_31__N_3003 [8]));   // verilog/motorControl.v(38[14] 59[8])
    SB_DFF \PID_CONTROLLER.result_i9  (.Q(\PID_CONTROLLER.result [9]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.result_31__N_3003 [9]));   // verilog/motorControl.v(38[14] 59[8])
    SB_DFF \PID_CONTROLLER.result_i10  (.Q(\PID_CONTROLLER.result [10]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.result_31__N_3003 [10]));   // verilog/motorControl.v(38[14] 59[8])
    SB_DFF \PID_CONTROLLER.result_i11  (.Q(\PID_CONTROLLER.result [11]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.result_31__N_3003 [11]));   // verilog/motorControl.v(38[14] 59[8])
    SB_DFF \PID_CONTROLLER.result_i12  (.Q(\PID_CONTROLLER.result [12]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.result_31__N_3003 [12]));   // verilog/motorControl.v(38[14] 59[8])
    SB_DFF \PID_CONTROLLER.result_i13  (.Q(\PID_CONTROLLER.result [13]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.result_31__N_3003 [13]));   // verilog/motorControl.v(38[14] 59[8])
    SB_DFF \PID_CONTROLLER.result_i14  (.Q(\PID_CONTROLLER.result [14]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.result_31__N_3003 [14]));   // verilog/motorControl.v(38[14] 59[8])
    SB_DFF \PID_CONTROLLER.result_i15  (.Q(\PID_CONTROLLER.result [15]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.result_31__N_3003 [15]));   // verilog/motorControl.v(38[14] 59[8])
    SB_DFF \PID_CONTROLLER.result_i16  (.Q(\PID_CONTROLLER.result [16]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.result_31__N_3003 [16]));   // verilog/motorControl.v(38[14] 59[8])
    SB_DFF \PID_CONTROLLER.result_i17  (.Q(\PID_CONTROLLER.result [17]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.result_31__N_3003 [17]));   // verilog/motorControl.v(38[14] 59[8])
    SB_DFF \PID_CONTROLLER.result_i18  (.Q(\PID_CONTROLLER.result [18]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.result_31__N_3003 [18]));   // verilog/motorControl.v(38[14] 59[8])
    SB_DFF \PID_CONTROLLER.result_i19  (.Q(\PID_CONTROLLER.result [19]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.result_31__N_3003 [19]));   // verilog/motorControl.v(38[14] 59[8])
    SB_DFF \PID_CONTROLLER.result_i20  (.Q(\PID_CONTROLLER.result [20]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.result_31__N_3003 [20]));   // verilog/motorControl.v(38[14] 59[8])
    SB_DFF \PID_CONTROLLER.result_i21  (.Q(\PID_CONTROLLER.result [21]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.result_31__N_3003 [21]));   // verilog/motorControl.v(38[14] 59[8])
    SB_DFF \PID_CONTROLLER.result_i22  (.Q(\PID_CONTROLLER.result [22]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.result_31__N_3003 [22]));   // verilog/motorControl.v(38[14] 59[8])
    SB_DFF \PID_CONTROLLER.result_i23  (.Q(\PID_CONTROLLER.result [23]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.result_31__N_3003 [23]));   // verilog/motorControl.v(38[14] 59[8])
    SB_DFF \PID_CONTROLLER.result_i24  (.Q(\PID_CONTROLLER.result [24]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.result_31__N_3003 [24]));   // verilog/motorControl.v(38[14] 59[8])
    SB_DFF \PID_CONTROLLER.result_i25  (.Q(\PID_CONTROLLER.result [25]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.result_31__N_3003 [25]));   // verilog/motorControl.v(38[14] 59[8])
    SB_DFF \PID_CONTROLLER.result_i26  (.Q(\PID_CONTROLLER.result [26]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.result_31__N_3003 [26]));   // verilog/motorControl.v(38[14] 59[8])
    SB_DFF \PID_CONTROLLER.result_i27  (.Q(\PID_CONTROLLER.result [27]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.result_31__N_3003 [27]));   // verilog/motorControl.v(38[14] 59[8])
    SB_DFF \PID_CONTROLLER.result_i28  (.Q(\PID_CONTROLLER.result [28]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.result_31__N_3003 [28]));   // verilog/motorControl.v(38[14] 59[8])
    SB_DFF \PID_CONTROLLER.result_i29  (.Q(\PID_CONTROLLER.result [29]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.result_31__N_3003 [29]));   // verilog/motorControl.v(38[14] 59[8])
    SB_DFF \PID_CONTROLLER.result_i30  (.Q(\PID_CONTROLLER.result [30]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.result_31__N_3003 [30]));   // verilog/motorControl.v(38[14] 59[8])
    SB_DFF \PID_CONTROLLER.result_i31  (.Q(\PID_CONTROLLER.result [31]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.result_31__N_3003 [31]));   // verilog/motorControl.v(38[14] 59[8])
    SB_DFF \PID_CONTROLLER.err_i2  (.Q(\PID_CONTROLLER.err[1] ), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_31__N_2825 [1]));   // verilog/motorControl.v(38[14] 59[8])
    SB_DFF GATES_i3 (.Q(PIN_8_c_2), .C(clk32MHz), .D(GATES_5__N_2788[2]));   // verilog/motorControl.v(64[10] 111[6])
    SB_DFF GATES_i4 (.Q(PIN_9_c_3), .C(clk32MHz), .D(GATES_5__N_2788[3]));   // verilog/motorControl.v(64[10] 111[6])
    SB_DFF GATES_i5 (.Q(PIN_10_c_4), .C(clk32MHz), .D(GATES_5__N_2788[4]));   // verilog/motorControl.v(64[10] 111[6])
    SB_DFF GATES_i6 (.Q(PIN_11_c_5), .C(clk32MHz), .D(GATES_5__N_2788[5]));   // verilog/motorControl.v(64[10] 111[6])
    SB_DFF \PID_CONTROLLER.err_i3  (.Q(\PID_CONTROLLER.err[2] ), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_31__N_2825 [2]));   // verilog/motorControl.v(38[14] 59[8])
    SB_CARRY add_13_add_1_20061_add_1_23 (.CI(n34876), .I0(n282[21]), .I1(n61[21]), 
            .CO(n34877));
    SB_LUT4 state_23__I_0_add_2_24_lut (.I0(GND_net), .I1(\motor_state[22] ), 
            .I2(n58[22]), .I3(n34237), .O(\PID_CONTROLLER.err_31__N_2825 [22])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3065_13_lut (.I0(GND_net), .I1(n8231[10]), .I2(GND_net), 
            .I3(n35449), .O(n8208[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3065_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3063_6 (.CI(n35399), .I0(n8184[3]), .I1(n510_adj_3731), 
            .CO(n35400));
    SB_CARRY add_3065_13 (.CI(n35449), .I0(n8231[10]), .I1(GND_net), .CO(n35450));
    SB_LUT4 add_3059_11_lut (.I0(GND_net), .I1(n8078[8]), .I2(GND_net), 
            .I3(n35306), .O(n8049[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3059_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3205_2 (.CI(GND_net), .I0(n35), .I1(n107), .CO(n35138));
    SB_CARRY add_3059_11 (.CI(n35306), .I0(n8078[8]), .I1(GND_net), .CO(n35307));
    SB_LUT4 add_3231_17_lut (.I0(GND_net), .I1(n12732[14]), .I2(GND_net), 
            .I3(n35137), .O(n12157[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3231_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1213_20_lut (.I0(GND_net), .I1(n1799[17]), .I2(GND_net), 
            .I3(n35817), .O(n1798[18])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1213_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3059_10_lut (.I0(GND_net), .I1(n8078[7]), .I2(GND_net), 
            .I3(n35305), .O(n8049[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3059_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3231_16_lut (.I0(GND_net), .I1(n12732[13]), .I2(GND_net), 
            .I3(n35136), .O(n12157[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3231_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3231_16 (.CI(n35136), .I0(n12732[13]), .I1(GND_net), 
            .CO(n35137));
    SB_LUT4 add_3063_5_lut (.I0(GND_net), .I1(n8184[2]), .I2(n413_adj_3740), 
            .I3(n35398), .O(n8159[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3063_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1213_20 (.CI(n35817), .I0(n1799[17]), .I1(GND_net), 
            .CO(n35818));
    SB_CARRY add_3059_10 (.CI(n35305), .I0(n8078[7]), .I1(GND_net), .CO(n35306));
    SB_CARRY add_3063_5 (.CI(n35398), .I0(n8184[2]), .I1(n413_adj_3740), 
            .CO(n35399));
    SB_LUT4 add_3231_15_lut (.I0(GND_net), .I1(n12732[12]), .I2(GND_net), 
            .I3(n35135), .O(n12157[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3231_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3231_15 (.CI(n35135), .I0(n12732[12]), .I1(GND_net), 
            .CO(n35136));
    SB_LUT4 add_13_add_1_20061_add_1_22_lut (.I0(GND_net), .I1(n282[20]), 
            .I2(n61[20]), .I3(n34875), .O(n63[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_13_add_1_20061_add_1_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_13_add_1_20061_add_1_22 (.CI(n34875), .I0(n282[20]), .I1(n61[20]), 
            .CO(n34876));
    SB_LUT4 add_3231_14_lut (.I0(GND_net), .I1(n12732[11]), .I2(GND_net), 
            .I3(n35134), .O(n12157[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3231_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_13_add_1_20061_add_1_21_lut (.I0(GND_net), .I1(n282[19]), 
            .I2(n61[19]), .I3(n34874), .O(n63[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_13_add_1_20061_add_1_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_13_add_1_20061_add_1_21 (.CI(n34874), .I0(n282[19]), .I1(n61[19]), 
            .CO(n34875));
    SB_LUT4 mult_14_add_1213_19_lut (.I0(GND_net), .I1(n1799[16]), .I2(GND_net), 
            .I3(n35816), .O(n1798[17])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1213_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3059_9_lut (.I0(GND_net), .I1(n8078[6]), .I2(GND_net), 
            .I3(n35304), .O(n8049[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3059_9_lut.LUT_INIT = 16'hC33C;
    SB_DFF \PID_CONTROLLER.err_i4  (.Q(\PID_CONTROLLER.err[3] ), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_31__N_2825 [3]));   // verilog/motorControl.v(38[14] 59[8])
    SB_DFF \PID_CONTROLLER.err_i5  (.Q(\PID_CONTROLLER.err[4] ), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_31__N_2825 [4]));   // verilog/motorControl.v(38[14] 59[8])
    SB_DFF \PID_CONTROLLER.err_i6  (.Q(\PID_CONTROLLER.err[5] ), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_31__N_2825 [5]));   // verilog/motorControl.v(38[14] 59[8])
    SB_DFF \PID_CONTROLLER.err_i7  (.Q(\PID_CONTROLLER.err[6] ), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_31__N_2825 [6]));   // verilog/motorControl.v(38[14] 59[8])
    SB_DFF \PID_CONTROLLER.err_i8  (.Q(\PID_CONTROLLER.err[7] ), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_31__N_2825 [7]));   // verilog/motorControl.v(38[14] 59[8])
    SB_DFF \PID_CONTROLLER.err_i9  (.Q(\PID_CONTROLLER.err[8] ), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_31__N_2825 [8]));   // verilog/motorControl.v(38[14] 59[8])
    SB_DFF \PID_CONTROLLER.err_i10  (.Q(\PID_CONTROLLER.err[9] ), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_31__N_2825 [9]));   // verilog/motorControl.v(38[14] 59[8])
    SB_DFF \PID_CONTROLLER.err_i11  (.Q(\PID_CONTROLLER.err[10] ), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_31__N_2825 [10]));   // verilog/motorControl.v(38[14] 59[8])
    SB_DFF \PID_CONTROLLER.err_i12  (.Q(\PID_CONTROLLER.err[11] ), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_31__N_2825 [11]));   // verilog/motorControl.v(38[14] 59[8])
    SB_DFF \PID_CONTROLLER.err_i13  (.Q(\PID_CONTROLLER.err[12] ), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_31__N_2825 [12]));   // verilog/motorControl.v(38[14] 59[8])
    SB_DFF \PID_CONTROLLER.err_i14  (.Q(\PID_CONTROLLER.err[13] ), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_31__N_2825 [13]));   // verilog/motorControl.v(38[14] 59[8])
    SB_DFF \PID_CONTROLLER.err_i15  (.Q(\PID_CONTROLLER.err[14] ), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_31__N_2825 [14]));   // verilog/motorControl.v(38[14] 59[8])
    SB_DFF \PID_CONTROLLER.err_i16  (.Q(\PID_CONTROLLER.err[15] ), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_31__N_2825 [15]));   // verilog/motorControl.v(38[14] 59[8])
    SB_DFF \PID_CONTROLLER.err_i17  (.Q(\PID_CONTROLLER.err[16] ), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_31__N_2825 [16]));   // verilog/motorControl.v(38[14] 59[8])
    SB_DFF \PID_CONTROLLER.err_i18  (.Q(\PID_CONTROLLER.err[17] ), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_31__N_2825 [17]));   // verilog/motorControl.v(38[14] 59[8])
    SB_DFF \PID_CONTROLLER.err_i19  (.Q(\PID_CONTROLLER.err[18] ), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_31__N_2825 [18]));   // verilog/motorControl.v(38[14] 59[8])
    SB_DFF \PID_CONTROLLER.err_i20  (.Q(\PID_CONTROLLER.err[19] ), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_31__N_2825 [19]));   // verilog/motorControl.v(38[14] 59[8])
    SB_DFF \PID_CONTROLLER.err_i21  (.Q(\PID_CONTROLLER.err[20] ), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_31__N_2825 [20]));   // verilog/motorControl.v(38[14] 59[8])
    SB_DFF \PID_CONTROLLER.err_i22  (.Q(\PID_CONTROLLER.err[21] ), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_31__N_2825 [21]));   // verilog/motorControl.v(38[14] 59[8])
    SB_DFF \PID_CONTROLLER.err_i23  (.Q(\PID_CONTROLLER.err[22] ), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_31__N_2825 [22]));   // verilog/motorControl.v(38[14] 59[8])
    SB_DFF \PID_CONTROLLER.err_i24  (.Q(\PID_CONTROLLER.err[23] ), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_31__N_2825 [23]));   // verilog/motorControl.v(38[14] 59[8])
    SB_DFF \PID_CONTROLLER.err_i25  (.Q(\PID_CONTROLLER.err[31] ), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_31__N_2825 [24]));   // verilog/motorControl.v(38[14] 59[8])
    SB_CARRY mult_14_add_1213_19 (.CI(n35816), .I0(n1799[16]), .I1(GND_net), 
            .CO(n35817));
    SB_LUT4 mult_14_add_1213_18_lut (.I0(GND_net), .I1(n1799[15]), .I2(GND_net), 
            .I3(n35815), .O(n1798[16])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1213_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3231_14 (.CI(n35134), .I0(n12732[11]), .I1(GND_net), 
            .CO(n35135));
    SB_LUT4 add_13_add_1_20061_add_1_20_lut (.I0(GND_net), .I1(n282[18]), 
            .I2(n61[18]), .I3(n34873), .O(n63[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_13_add_1_20061_add_1_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_13_add_1_20061_add_1_20 (.CI(n34873), .I0(n282[18]), .I1(n61[18]), 
            .CO(n34874));
    SB_LUT4 add_3231_13_lut (.I0(GND_net), .I1(n12732[10]), .I2(GND_net), 
            .I3(n35133), .O(n12157[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3231_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_13_add_1_20061_add_1_19_lut (.I0(GND_net), .I1(n282[17]), 
            .I2(n61[17]), .I3(n34872), .O(n63[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_13_add_1_20061_add_1_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_13_add_1_20061_add_1_19 (.CI(n34872), .I0(n282[17]), .I1(n61[17]), 
            .CO(n34873));
    SB_LUT4 add_3070_5_lut (.I0(GND_net), .I1(n8331[2]), .I2(n434), .I3(n35531), 
            .O(n8313[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3070_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_13_add_1_20061_add_1_18_lut (.I0(GND_net), .I1(n282[16]), 
            .I2(n61[16]), .I3(n34871), .O(n63[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_13_add_1_20061_add_1_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3067_13_lut (.I0(GND_net), .I1(n8274[10]), .I2(GND_net), 
            .I3(n35488), .O(n8253[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3067_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3065_12_lut (.I0(GND_net), .I1(n8231[9]), .I2(GND_net), 
            .I3(n35448), .O(n8208[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3065_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3059_9 (.CI(n35304), .I0(n8078[6]), .I1(GND_net), .CO(n35305));
    SB_LUT4 add_3063_4_lut (.I0(GND_net), .I1(n8184[1]), .I2(n316_adj_3742), 
            .I3(n35397), .O(n8159[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3063_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3059_8_lut (.I0(GND_net), .I1(n8078[5]), .I2(n692_adj_3743), 
            .I3(n35303), .O(n8049[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3059_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3301_11 (.CI(n34593), .I0(n14168[8]), .I1(GND_net), .CO(n34594));
    SB_CARRY add_3231_13 (.CI(n35133), .I0(n12732[10]), .I1(GND_net), 
            .CO(n35134));
    SB_LUT4 add_3231_12_lut (.I0(GND_net), .I1(n12732[9]), .I2(GND_net), 
            .I3(n35132), .O(n12157[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3231_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1213_18 (.CI(n35815), .I0(n1799[15]), .I1(GND_net), 
            .CO(n35816));
    SB_LUT4 add_3301_10_lut (.I0(GND_net), .I1(n14168[7]), .I2(GND_net), 
            .I3(n34592), .O(n13734[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3301_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_13_add_1_20061_add_1_18 (.CI(n34871), .I0(n282[16]), .I1(n61[16]), 
            .CO(n34872));
    SB_LUT4 mult_14_add_1213_17_lut (.I0(GND_net), .I1(n1799[14]), .I2(GND_net), 
            .I3(n35814), .O(n1798[15])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1213_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY state_23__I_0_add_2_24 (.CI(n34237), .I0(\motor_state[22] ), 
            .I1(n58[22]), .CO(n34238));
    SB_CARRY add_3301_10 (.CI(n34592), .I0(n14168[7]), .I1(GND_net), .CO(n34593));
    SB_LUT4 state_23__I_0_add_2_23_lut (.I0(GND_net), .I1(\motor_state[21] ), 
            .I2(n58[21]), .I3(n34236), .O(\PID_CONTROLLER.err_31__N_2825 [21])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1213_17 (.CI(n35814), .I0(n1799[14]), .I1(GND_net), 
            .CO(n35815));
    SB_LUT4 mult_14_add_1213_16_lut (.I0(GND_net), .I1(n1799[13]), .I2(GND_net), 
            .I3(n35813), .O(n1798[14])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1213_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1213_16 (.CI(n35813), .I0(n1799[13]), .I1(GND_net), 
            .CO(n35814));
    SB_LUT4 mult_14_add_1213_15_lut (.I0(GND_net), .I1(n1799[12]), .I2(GND_net), 
            .I3(n35812), .O(n1798[13])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1213_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1213_15 (.CI(n35812), .I0(n1799[12]), .I1(GND_net), 
            .CO(n35813));
    SB_LUT4 mult_14_add_1213_14_lut (.I0(GND_net), .I1(n1799[11]), .I2(GND_net), 
            .I3(n35811), .O(n1798[12])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1213_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY state_23__I_0_add_2_23 (.CI(n34236), .I0(\motor_state[21] ), 
            .I1(n58[21]), .CO(n34237));
    SB_LUT4 add_13_add_1_20061_add_1_17_lut (.I0(GND_net), .I1(n282[15]), 
            .I2(n61[15]), .I3(n34870), .O(n63[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_13_add_1_20061_add_1_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 state_23__I_0_add_2_22_lut (.I0(GND_net), .I1(\motor_state[20] ), 
            .I2(n58[20]), .I3(n34235), .O(\PID_CONTROLLER.err_31__N_2825 [20])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3301_9_lut (.I0(GND_net), .I1(n14168[6]), .I2(GND_net), 
            .I3(n34591), .O(n13734[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3301_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_12_i170_2_lut (.I0(\Kd[2] ), .I1(n57[19]), .I2(GND_net), 
            .I3(GND_net), .O(n252));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i170_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY mult_14_add_1213_14 (.CI(n35811), .I0(n1799[11]), .I1(GND_net), 
            .CO(n35812));
    SB_CARRY state_23__I_0_add_2_22 (.CI(n34235), .I0(\motor_state[20] ), 
            .I1(n58[20]), .CO(n34236));
    SB_LUT4 add_3272_19_lut (.I0(GND_net), .I1(n13594[16]), .I2(GND_net), 
            .I3(n34406), .O(n13109[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3272_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1213_13_lut (.I0(GND_net), .I1(n1799[10]), .I2(GND_net), 
            .I3(n35810), .O(n1798[11])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1213_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1213_13 (.CI(n35810), .I0(n1799[10]), .I1(GND_net), 
            .CO(n35811));
    SB_LUT4 state_23__I_0_add_2_21_lut (.I0(GND_net), .I1(\motor_state[19] ), 
            .I2(n58[19]), .I3(n34234), .O(\PID_CONTROLLER.err_31__N_2825 [19])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1213_12_lut (.I0(GND_net), .I1(n1799[9]), .I2(GND_net), 
            .I3(n35809), .O(n1798[10])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1213_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3272_19 (.CI(n34406), .I0(n13594[16]), .I1(GND_net), 
            .CO(n34407));
    SB_CARRY mult_14_add_1213_12 (.CI(n35809), .I0(n1799[9]), .I1(GND_net), 
            .CO(n35810));
    SB_CARRY add_3301_9 (.CI(n34591), .I0(n14168[6]), .I1(GND_net), .CO(n34592));
    SB_LUT4 add_3272_18_lut (.I0(GND_net), .I1(n13594[15]), .I2(GND_net), 
            .I3(n34405), .O(n13109[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3272_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3272_18 (.CI(n34405), .I0(n13594[15]), .I1(GND_net), 
            .CO(n34406));
    SB_CARRY add_3231_12 (.CI(n35132), .I0(n12732[9]), .I1(GND_net), .CO(n35133));
    SB_LUT4 add_3301_8_lut (.I0(GND_net), .I1(n14168[5]), .I2(n545), .I3(n34590), 
            .O(n13734[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3301_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3272_17_lut (.I0(GND_net), .I1(n13594[14]), .I2(GND_net), 
            .I3(n34404), .O(n13109[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3272_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3272_17 (.CI(n34404), .I0(n13594[14]), .I1(GND_net), 
            .CO(n34405));
    SB_CARRY add_3301_8 (.CI(n34590), .I0(n14168[5]), .I1(n545), .CO(n34591));
    SB_LUT4 add_3272_16_lut (.I0(GND_net), .I1(n13594[13]), .I2(GND_net), 
            .I3(n34403), .O(n13109[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3272_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3059_8 (.CI(n35303), .I0(n8078[5]), .I1(n692_adj_3743), 
            .CO(n35304));
    SB_LUT4 add_3231_11_lut (.I0(GND_net), .I1(n12732[8]), .I2(GND_net), 
            .I3(n35131), .O(n12157[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3231_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3301_7_lut (.I0(GND_net), .I1(n14168[4]), .I2(n472), .I3(n34589), 
            .O(n13734[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3301_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3272_16 (.CI(n34403), .I0(n13594[13]), .I1(GND_net), 
            .CO(n34404));
    SB_LUT4 add_3272_15_lut (.I0(GND_net), .I1(n13594[12]), .I2(GND_net), 
            .I3(n34402), .O(n13109[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3272_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3301_7 (.CI(n34589), .I0(n14168[4]), .I1(n472), .CO(n34590));
    SB_CARRY add_3272_15 (.CI(n34402), .I0(n13594[12]), .I1(GND_net), 
            .CO(n34403));
    SB_CARRY add_3070_5 (.CI(n35531), .I0(n8331[2]), .I1(n434), .CO(n35532));
    SB_LUT4 add_3272_14_lut (.I0(GND_net), .I1(n13594[11]), .I2(GND_net), 
            .I3(n34401), .O(n13109[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3272_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3070_4_lut (.I0(GND_net), .I1(n8331[1]), .I2(n337), .I3(n35530), 
            .O(n8313[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3070_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3070_4 (.CI(n35530), .I0(n8331[1]), .I1(n337), .CO(n35531));
    SB_LUT4 add_3070_3_lut (.I0(GND_net), .I1(n8331[0]), .I2(n240_adj_3748), 
            .I3(n35529), .O(n8313[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3070_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3070_3 (.CI(n35529), .I0(n8331[0]), .I1(n240_adj_3748), 
            .CO(n35530));
    SB_LUT4 add_3070_2_lut (.I0(GND_net), .I1(n50_adj_3749), .I2(n143_adj_3750), 
            .I3(GND_net), .O(n8313[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3070_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3070_2 (.CI(GND_net), .I0(n50_adj_3749), .I1(n143_adj_3750), 
            .CO(n35529));
    SB_CARRY add_3231_11 (.CI(n35131), .I0(n12732[8]), .I1(GND_net), .CO(n35132));
    SB_LUT4 mult_14_add_1213_11_lut (.I0(GND_net), .I1(n1799[8]), .I2(GND_net), 
            .I3(n35808), .O(n1798[9])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1213_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1213_11 (.CI(n35808), .I0(n1799[8]), .I1(GND_net), 
            .CO(n35809));
    SB_LUT4 mult_14_add_1213_10_lut (.I0(GND_net), .I1(n1799[7]), .I2(GND_net), 
            .I3(n35807), .O(n1798[8])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1213_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1213_10 (.CI(n35807), .I0(n1799[7]), .I1(GND_net), 
            .CO(n35808));
    SB_LUT4 mult_14_add_1213_9_lut (.I0(GND_net), .I1(n1799[6]), .I2(GND_net), 
            .I3(n35806), .O(n1798[7])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1213_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1213_9 (.CI(n35806), .I0(n1799[6]), .I1(GND_net), 
            .CO(n35807));
    SB_LUT4 mult_14_add_1213_8_lut (.I0(GND_net), .I1(n1799[5]), .I2(n518), 
            .I3(n35805), .O(n1798[6])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1213_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1213_8 (.CI(n35805), .I0(n1799[5]), .I1(n518), 
            .CO(n35806));
    SB_LUT4 mult_14_add_1213_7_lut (.I0(GND_net), .I1(n1799[4]), .I2(n445), 
            .I3(n35804), .O(n1798[5])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1213_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1213_7 (.CI(n35804), .I0(n1799[4]), .I1(n445), 
            .CO(n35805));
    SB_LUT4 mult_14_add_1213_6_lut (.I0(GND_net), .I1(n1799[3]), .I2(n372), 
            .I3(n35803), .O(n1798[4])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1213_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1213_6 (.CI(n35803), .I0(n1799[3]), .I1(n372), 
            .CO(n35804));
    SB_LUT4 mult_14_add_1213_5_lut (.I0(GND_net), .I1(n1799[2]), .I2(n299_adj_3755), 
            .I3(n35802), .O(n1798[3])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1213_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1213_5 (.CI(n35802), .I0(n1799[2]), .I1(n299_adj_3755), 
            .CO(n35803));
    SB_LUT4 mult_14_add_1213_4_lut (.I0(GND_net), .I1(n1799[1]), .I2(n226_adj_3757), 
            .I3(n35801), .O(n1798[2])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1213_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1213_4 (.CI(n35801), .I0(n1799[1]), .I1(n226_adj_3757), 
            .CO(n35802));
    SB_LUT4 mult_14_add_1213_3_lut (.I0(GND_net), .I1(n1799[0]), .I2(n153_adj_3759), 
            .I3(n35800), .O(n1798[1])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1213_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1213_3 (.CI(n35800), .I0(n1799[0]), .I1(n153_adj_3759), 
            .CO(n35801));
    SB_LUT4 mult_14_add_1213_2_lut (.I0(GND_net), .I1(n11_adj_3760), .I2(n80), 
            .I3(GND_net), .O(n1798[0])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1213_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1213_2 (.CI(GND_net), .I0(n11_adj_3760), .I1(n80), 
            .CO(n35800));
    SB_LUT4 mult_14_add_1212_24_lut (.I0(GND_net), .I1(n1798[21]), .I2(GND_net), 
            .I3(n35798), .O(n1797[22])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1212_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1212_24 (.CI(n35798), .I0(n1798[21]), .I1(GND_net), 
            .CO(n1687));
    SB_LUT4 mult_14_add_1212_23_lut (.I0(GND_net), .I1(n1798[20]), .I2(GND_net), 
            .I3(n35797), .O(n1797[21])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1212_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1212_23 (.CI(n35797), .I0(n1798[20]), .I1(GND_net), 
            .CO(n35798));
    SB_LUT4 add_3301_6_lut (.I0(GND_net), .I1(n14168[3]), .I2(n399), .I3(n34588), 
            .O(n13734[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3301_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3272_14 (.CI(n34401), .I0(n13594[11]), .I1(GND_net), 
            .CO(n34402));
    SB_LUT4 add_3272_13_lut (.I0(GND_net), .I1(n13594[10]), .I2(GND_net), 
            .I3(n34400), .O(n13109[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3272_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3301_6 (.CI(n34588), .I0(n14168[3]), .I1(n399), .CO(n34589));
    SB_CARRY state_23__I_0_add_2_21 (.CI(n34234), .I0(\motor_state[19] ), 
            .I1(n58[19]), .CO(n34235));
    SB_LUT4 mult_14_add_1212_22_lut (.I0(GND_net), .I1(n1798[19]), .I2(GND_net), 
            .I3(n35796), .O(n1797[20])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1212_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1212_22 (.CI(n35796), .I0(n1798[19]), .I1(GND_net), 
            .CO(n35797));
    SB_CARRY add_3272_13 (.CI(n34400), .I0(n13594[10]), .I1(GND_net), 
            .CO(n34401));
    SB_LUT4 mult_14_add_1212_21_lut (.I0(GND_net), .I1(n1798[18]), .I2(GND_net), 
            .I3(n35795), .O(n1797[19])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1212_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3067_13 (.CI(n35488), .I0(n8274[10]), .I1(GND_net), .CO(n35489));
    SB_CARRY mult_14_add_1212_21 (.CI(n35795), .I0(n1798[18]), .I1(GND_net), 
            .CO(n35796));
    SB_LUT4 mult_14_add_1212_20_lut (.I0(GND_net), .I1(n1798[17]), .I2(GND_net), 
            .I3(n35794), .O(n1797[18])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1212_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1212_20 (.CI(n35794), .I0(n1798[17]), .I1(GND_net), 
            .CO(n35795));
    SB_LUT4 mult_14_add_1212_19_lut (.I0(GND_net), .I1(n1798[16]), .I2(GND_net), 
            .I3(n35793), .O(n1797[17])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1212_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1212_19 (.CI(n35793), .I0(n1798[16]), .I1(GND_net), 
            .CO(n35794));
    SB_LUT4 mult_14_add_1212_18_lut (.I0(GND_net), .I1(n1798[15]), .I2(GND_net), 
            .I3(n35792), .O(n1797[16])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1212_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1212_18 (.CI(n35792), .I0(n1798[15]), .I1(GND_net), 
            .CO(n35793));
    SB_LUT4 mult_14_add_1212_17_lut (.I0(GND_net), .I1(n1798[14]), .I2(GND_net), 
            .I3(n35791), .O(n1797[15])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1212_17_lut.LUT_INIT = 16'hC33C;
    SB_DFF Kd_delay_counter_1015__i1 (.Q(Kd_delay_counter[1]), .C(clk32MHz), 
           .D(n69[1]));   // verilog/motorControl.v(55[27:47])
    SB_CARRY mult_14_add_1212_17 (.CI(n35791), .I0(n1798[14]), .I1(GND_net), 
            .CO(n35792));
    SB_LUT4 mult_14_add_1212_16_lut (.I0(GND_net), .I1(n1798[13]), .I2(GND_net), 
            .I3(n35790), .O(n1797[14])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1212_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1212_16 (.CI(n35790), .I0(n1798[13]), .I1(GND_net), 
            .CO(n35791));
    SB_LUT4 mult_14_add_1212_15_lut (.I0(GND_net), .I1(n1798[12]), .I2(GND_net), 
            .I3(n35789), .O(n1797[13])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1212_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1212_15 (.CI(n35789), .I0(n1798[12]), .I1(GND_net), 
            .CO(n35790));
    SB_LUT4 mult_14_add_1212_14_lut (.I0(GND_net), .I1(n1798[11]), .I2(GND_net), 
            .I3(n35788), .O(n1797[12])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1212_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1212_14 (.CI(n35788), .I0(n1798[11]), .I1(GND_net), 
            .CO(n35789));
    SB_LUT4 mult_14_add_1212_13_lut (.I0(GND_net), .I1(n1798[10]), .I2(GND_net), 
            .I3(n35787), .O(n1797[11])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1212_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1212_13 (.CI(n35787), .I0(n1798[10]), .I1(GND_net), 
            .CO(n35788));
    SB_LUT4 mult_14_add_1212_12_lut (.I0(GND_net), .I1(n1798[9]), .I2(GND_net), 
            .I3(n35786), .O(n1797[10])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1212_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1212_12 (.CI(n35786), .I0(n1798[9]), .I1(GND_net), 
            .CO(n35787));
    SB_LUT4 mult_14_add_1212_11_lut (.I0(GND_net), .I1(n1798[8]), .I2(GND_net), 
            .I3(n35785), .O(n1797[9])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1212_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1212_11 (.CI(n35785), .I0(n1798[8]), .I1(GND_net), 
            .CO(n35786));
    SB_LUT4 mult_14_add_1212_10_lut (.I0(GND_net), .I1(n1798[7]), .I2(GND_net), 
            .I3(n35784), .O(n1797[8])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1212_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1212_10 (.CI(n35784), .I0(n1798[7]), .I1(GND_net), 
            .CO(n35785));
    SB_LUT4 mult_14_add_1212_9_lut (.I0(GND_net), .I1(n1798[6]), .I2(GND_net), 
            .I3(n35783), .O(n1797[7])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1212_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1212_9 (.CI(n35783), .I0(n1798[6]), .I1(GND_net), 
            .CO(n35784));
    SB_LUT4 mult_14_add_1212_8_lut (.I0(GND_net), .I1(n1798[5]), .I2(n515), 
            .I3(n35782), .O(n1797[6])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1212_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1212_8 (.CI(n35782), .I0(n1798[5]), .I1(n515), 
            .CO(n35783));
    SB_LUT4 mult_14_add_1212_7_lut (.I0(GND_net), .I1(n1798[4]), .I2(n442), 
            .I3(n35781), .O(n1797[5])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1212_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1212_7 (.CI(n35781), .I0(n1798[4]), .I1(n442), 
            .CO(n35782));
    SB_LUT4 mult_14_add_1212_6_lut (.I0(GND_net), .I1(n1798[3]), .I2(n369), 
            .I3(n35780), .O(n1797[4])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1212_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1212_6 (.CI(n35780), .I0(n1798[3]), .I1(n369), 
            .CO(n35781));
    SB_LUT4 mult_14_add_1212_5_lut (.I0(GND_net), .I1(n1798[2]), .I2(n296_adj_3766), 
            .I3(n35779), .O(n1797[3])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1212_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1212_5 (.CI(n35779), .I0(n1798[2]), .I1(n296_adj_3766), 
            .CO(n35780));
    SB_LUT4 mult_14_add_1212_4_lut (.I0(GND_net), .I1(n1798[1]), .I2(n223_adj_3768), 
            .I3(n35778), .O(n1797[2])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1212_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1212_4 (.CI(n35778), .I0(n1798[1]), .I1(n223_adj_3768), 
            .CO(n35779));
    SB_LUT4 mult_14_add_1212_3_lut (.I0(GND_net), .I1(n1798[0]), .I2(n150_adj_3770), 
            .I3(n35777), .O(n1797[1])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1212_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1212_3 (.CI(n35777), .I0(n1798[0]), .I1(n150_adj_3770), 
            .CO(n35778));
    SB_LUT4 mult_14_add_1212_2_lut (.I0(GND_net), .I1(n8_adj_3771), .I2(n77), 
            .I3(GND_net), .O(n1797[0])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1212_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1212_2 (.CI(GND_net), .I0(n8_adj_3771), .I1(n77), 
            .CO(n35777));
    SB_LUT4 mult_14_add_1211_24_lut (.I0(GND_net), .I1(n1797[21]), .I2(GND_net), 
            .I3(n35775), .O(n1796[22])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1211_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1211_24 (.CI(n35775), .I0(n1797[21]), .I1(GND_net), 
            .CO(n1683));
    SB_LUT4 mult_14_add_1211_23_lut (.I0(GND_net), .I1(n1797[20]), .I2(GND_net), 
            .I3(n35774), .O(n282[22])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1211_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1211_23 (.CI(n35774), .I0(n1797[20]), .I1(GND_net), 
            .CO(n35775));
    SB_LUT4 mult_14_add_1211_22_lut (.I0(GND_net), .I1(n1797[19]), .I2(GND_net), 
            .I3(n35773), .O(n282[21])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1211_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1211_22 (.CI(n35773), .I0(n1797[19]), .I1(GND_net), 
            .CO(n35774));
    SB_LUT4 mult_14_add_1211_21_lut (.I0(GND_net), .I1(n1797[18]), .I2(GND_net), 
            .I3(n35772), .O(n282[20])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1211_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1211_21 (.CI(n35772), .I0(n1797[18]), .I1(GND_net), 
            .CO(n35773));
    SB_LUT4 mult_14_add_1211_20_lut (.I0(GND_net), .I1(n1797[17]), .I2(GND_net), 
            .I3(n35771), .O(n282[19])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1211_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1211_20 (.CI(n35771), .I0(n1797[17]), .I1(GND_net), 
            .CO(n35772));
    SB_LUT4 mult_14_add_1211_19_lut (.I0(GND_net), .I1(n1797[16]), .I2(GND_net), 
            .I3(n35770), .O(n282[18])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1211_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1211_19 (.CI(n35770), .I0(n1797[16]), .I1(GND_net), 
            .CO(n35771));
    SB_LUT4 mult_14_add_1211_18_lut (.I0(GND_net), .I1(n1797[15]), .I2(GND_net), 
            .I3(n35769), .O(n282[17])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1211_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1211_18 (.CI(n35769), .I0(n1797[15]), .I1(GND_net), 
            .CO(n35770));
    SB_LUT4 mult_14_add_1211_17_lut (.I0(GND_net), .I1(n1797[14]), .I2(GND_net), 
            .I3(n35768), .O(n282[16])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1211_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1211_17 (.CI(n35768), .I0(n1797[14]), .I1(GND_net), 
            .CO(n35769));
    SB_LUT4 mult_14_add_1211_16_lut (.I0(GND_net), .I1(n1797[13]), .I2(GND_net), 
            .I3(n35767), .O(n282[15])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1211_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1211_16 (.CI(n35767), .I0(n1797[13]), .I1(GND_net), 
            .CO(n35768));
    SB_LUT4 mult_14_add_1211_15_lut (.I0(GND_net), .I1(n1797[12]), .I2(GND_net), 
            .I3(n35766), .O(n282[14])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1211_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1211_15 (.CI(n35766), .I0(n1797[12]), .I1(GND_net), 
            .CO(n35767));
    SB_LUT4 mult_14_add_1211_14_lut (.I0(GND_net), .I1(n1797[11]), .I2(GND_net), 
            .I3(n35765), .O(n282[13])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1211_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1211_14 (.CI(n35765), .I0(n1797[11]), .I1(GND_net), 
            .CO(n35766));
    SB_LUT4 mult_14_add_1211_13_lut (.I0(GND_net), .I1(n1797[10]), .I2(GND_net), 
            .I3(n35764), .O(n282[12])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1211_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1211_13 (.CI(n35764), .I0(n1797[10]), .I1(GND_net), 
            .CO(n35765));
    SB_LUT4 mult_14_add_1211_12_lut (.I0(GND_net), .I1(n1797[9]), .I2(GND_net), 
            .I3(n35763), .O(n282[11])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1211_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1211_12 (.CI(n35763), .I0(n1797[9]), .I1(GND_net), 
            .CO(n35764));
    SB_LUT4 mult_14_add_1211_11_lut (.I0(GND_net), .I1(n1797[8]), .I2(GND_net), 
            .I3(n35762), .O(n282[10])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1211_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1211_11 (.CI(n35762), .I0(n1797[8]), .I1(GND_net), 
            .CO(n35763));
    SB_LUT4 mult_14_add_1211_10_lut (.I0(GND_net), .I1(n1797[7]), .I2(GND_net), 
            .I3(n35761), .O(n282[9])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1211_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1211_10 (.CI(n35761), .I0(n1797[7]), .I1(GND_net), 
            .CO(n35762));
    SB_LUT4 mult_14_add_1211_9_lut (.I0(GND_net), .I1(n1797[6]), .I2(GND_net), 
            .I3(n35760), .O(n282[8])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1211_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1211_9 (.CI(n35760), .I0(n1797[6]), .I1(GND_net), 
            .CO(n35761));
    SB_LUT4 mult_14_add_1211_8_lut (.I0(GND_net), .I1(n1797[5]), .I2(n512), 
            .I3(n35759), .O(n282[7])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1211_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1211_8 (.CI(n35759), .I0(n1797[5]), .I1(n512), 
            .CO(n35760));
    SB_LUT4 mult_14_add_1211_7_lut (.I0(GND_net), .I1(n1797[4]), .I2(n439), 
            .I3(n35758), .O(n282[6])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1211_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1211_7 (.CI(n35758), .I0(n1797[4]), .I1(n439), 
            .CO(n35759));
    SB_LUT4 mult_14_add_1211_6_lut (.I0(GND_net), .I1(n1797[3]), .I2(n366), 
            .I3(n35757), .O(n282[5])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1211_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1211_6 (.CI(n35757), .I0(n1797[3]), .I1(n366), 
            .CO(n35758));
    SB_LUT4 mult_14_add_1211_5_lut (.I0(GND_net), .I1(n1797[2]), .I2(n293), 
            .I3(n35756), .O(n282[4])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1211_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1211_5 (.CI(n35756), .I0(n1797[2]), .I1(n293), 
            .CO(n35757));
    SB_LUT4 mult_14_add_1211_4_lut (.I0(GND_net), .I1(n1797[1]), .I2(n220_adj_3777), 
            .I3(n35755), .O(n282[3])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1211_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1211_4 (.CI(n35755), .I0(n1797[1]), .I1(n220_adj_3777), 
            .CO(n35756));
    SB_LUT4 mult_14_add_1211_3_lut (.I0(GND_net), .I1(n1797[0]), .I2(n147_adj_3778), 
            .I3(n35754), .O(n282[2])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1211_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1211_3 (.CI(n35754), .I0(n1797[0]), .I1(n147_adj_3778), 
            .CO(n35755));
    SB_LUT4 mult_14_add_1211_2_lut (.I0(GND_net), .I1(n5_adj_3779), .I2(n74_adj_3780), 
            .I3(GND_net), .O(n282[1])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1211_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1211_2 (.CI(GND_net), .I0(n5_adj_3779), .I1(n74_adj_3780), 
            .CO(n35754));
    SB_LUT4 add_3372_18_lut (.I0(GND_net), .I1(n15399[15]), .I2(GND_net), 
            .I3(n35753), .O(n15114[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3372_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3372_17_lut (.I0(GND_net), .I1(n15399[14]), .I2(GND_net), 
            .I3(n35752), .O(n15114[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3372_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3372_17 (.CI(n35752), .I0(n15399[14]), .I1(GND_net), 
            .CO(n35753));
    SB_LUT4 add_3372_16_lut (.I0(GND_net), .I1(n15399[13]), .I2(GND_net), 
            .I3(n35751), .O(n15114[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3372_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3372_16 (.CI(n35751), .I0(n15399[13]), .I1(GND_net), 
            .CO(n35752));
    SB_LUT4 add_3372_15_lut (.I0(GND_net), .I1(n15399[12]), .I2(GND_net), 
            .I3(n35750), .O(n15114[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3372_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3372_15 (.CI(n35750), .I0(n15399[12]), .I1(GND_net), 
            .CO(n35751));
    SB_LUT4 add_3372_14_lut (.I0(GND_net), .I1(n15399[11]), .I2(GND_net), 
            .I3(n35749), .O(n15114[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3372_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3372_14 (.CI(n35749), .I0(n15399[11]), .I1(GND_net), 
            .CO(n35750));
    SB_LUT4 add_3372_13_lut (.I0(GND_net), .I1(n15399[10]), .I2(GND_net), 
            .I3(n35748), .O(n15114[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3372_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3372_13 (.CI(n35748), .I0(n15399[10]), .I1(GND_net), 
            .CO(n35749));
    SB_LUT4 add_3372_12_lut (.I0(GND_net), .I1(n15399[9]), .I2(GND_net), 
            .I3(n35747), .O(n15114[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3372_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3372_12 (.CI(n35747), .I0(n15399[9]), .I1(GND_net), .CO(n35748));
    SB_LUT4 add_3372_11_lut (.I0(GND_net), .I1(n15399[8]), .I2(GND_net), 
            .I3(n35746), .O(n15114[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3372_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3372_11 (.CI(n35746), .I0(n15399[8]), .I1(GND_net), .CO(n35747));
    SB_LUT4 add_3372_10_lut (.I0(GND_net), .I1(n15399[7]), .I2(GND_net), 
            .I3(n35745), .O(n15114[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3372_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3372_10 (.CI(n35745), .I0(n15399[7]), .I1(GND_net), .CO(n35746));
    SB_LUT4 add_3372_9_lut (.I0(GND_net), .I1(n15399[6]), .I2(GND_net), 
            .I3(n35744), .O(n15114[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3372_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3372_9 (.CI(n35744), .I0(n15399[6]), .I1(GND_net), .CO(n35745));
    SB_LUT4 add_3372_8_lut (.I0(GND_net), .I1(n15399[5]), .I2(n722_adj_3781), 
            .I3(n35743), .O(n15114[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3372_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3372_8 (.CI(n35743), .I0(n15399[5]), .I1(n722_adj_3781), 
            .CO(n35744));
    SB_LUT4 add_3372_7_lut (.I0(GND_net), .I1(n15399[4]), .I2(n625_adj_3782), 
            .I3(n35742), .O(n15114[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3372_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3372_7 (.CI(n35742), .I0(n15399[4]), .I1(n625_adj_3782), 
            .CO(n35743));
    SB_LUT4 add_3372_6_lut (.I0(GND_net), .I1(n15399[3]), .I2(n528_adj_3783), 
            .I3(n35741), .O(n15114[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3372_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3372_6 (.CI(n35741), .I0(n15399[3]), .I1(n528_adj_3783), 
            .CO(n35742));
    SB_LUT4 add_3372_5_lut (.I0(GND_net), .I1(n15399[2]), .I2(n431_adj_3784), 
            .I3(n35740), .O(n15114[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3372_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3372_5 (.CI(n35740), .I0(n15399[2]), .I1(n431_adj_3784), 
            .CO(n35741));
    SB_LUT4 add_3372_4_lut (.I0(GND_net), .I1(n15399[1]), .I2(n334_adj_3785), 
            .I3(n35739), .O(n15114[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3372_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3372_4 (.CI(n35739), .I0(n15399[1]), .I1(n334_adj_3785), 
            .CO(n35740));
    SB_LUT4 add_3372_3_lut (.I0(GND_net), .I1(n15399[0]), .I2(n237_adj_3786), 
            .I3(n35738), .O(n15114[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3372_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3372_3 (.CI(n35738), .I0(n15399[0]), .I1(n237_adj_3786), 
            .CO(n35739));
    SB_LUT4 add_3372_2_lut (.I0(GND_net), .I1(n47_adj_3787), .I2(n140_adj_3788), 
            .I3(GND_net), .O(n15114[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3372_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3372_2 (.CI(GND_net), .I0(n47_adj_3787), .I1(n140_adj_3788), 
            .CO(n35738));
    SB_LUT4 add_3481_9_lut (.I0(GND_net), .I1(n16620[6]), .I2(GND_net), 
            .I3(n35737), .O(n16571[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3481_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3481_8_lut (.I0(GND_net), .I1(n16620[5]), .I2(n749_adj_3789), 
            .I3(n35736), .O(n16571[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3481_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3481_8 (.CI(n35736), .I0(n16620[5]), .I1(n749_adj_3789), 
            .CO(n35737));
    SB_LUT4 add_3481_7_lut (.I0(GND_net), .I1(n16620[4]), .I2(n652_adj_3790), 
            .I3(n35735), .O(n16571[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3481_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3059_7_lut (.I0(GND_net), .I1(n8078[4]), .I2(n595_adj_3791), 
            .I3(n35302), .O(n8049[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3059_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3272_12_lut (.I0(GND_net), .I1(n13594[9]), .I2(GND_net), 
            .I3(n34399), .O(n13109[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3272_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3481_7 (.CI(n35735), .I0(n16620[4]), .I1(n652_adj_3790), 
            .CO(n35736));
    SB_LUT4 add_3231_10_lut (.I0(GND_net), .I1(n12732[7]), .I2(GND_net), 
            .I3(n35130), .O(n12157[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3231_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3272_12 (.CI(n34399), .I0(n13594[9]), .I1(GND_net), .CO(n34400));
    SB_LUT4 add_3301_5_lut (.I0(GND_net), .I1(n14168[2]), .I2(n326), .I3(n34587), 
            .O(n13734[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3301_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3059_7 (.CI(n35302), .I0(n8078[4]), .I1(n595_adj_3791), 
            .CO(n35303));
    SB_LUT4 add_3272_11_lut (.I0(GND_net), .I1(n13594[8]), .I2(GND_net), 
            .I3(n34398), .O(n13109[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3272_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3481_6_lut (.I0(GND_net), .I1(n16620[3]), .I2(n555_adj_3792), 
            .I3(n35734), .O(n16571[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3481_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3481_6 (.CI(n35734), .I0(n16620[3]), .I1(n555_adj_3792), 
            .CO(n35735));
    SB_LUT4 add_3481_5_lut (.I0(GND_net), .I1(n16620[2]), .I2(n458_adj_3793), 
            .I3(n35733), .O(n16571[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3481_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3481_5 (.CI(n35733), .I0(n16620[2]), .I1(n458_adj_3793), 
            .CO(n35734));
    SB_LUT4 add_3481_4_lut (.I0(GND_net), .I1(n16620[1]), .I2(n361_adj_3794), 
            .I3(n35732), .O(n16571[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3481_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3481_4 (.CI(n35732), .I0(n16620[1]), .I1(n361_adj_3794), 
            .CO(n35733));
    SB_LUT4 add_3481_3_lut (.I0(GND_net), .I1(n16620[0]), .I2(n264_adj_3795), 
            .I3(n35731), .O(n16571[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3481_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3481_3 (.CI(n35731), .I0(n16620[0]), .I1(n264_adj_3795), 
            .CO(n35732));
    SB_LUT4 add_3481_2_lut (.I0(GND_net), .I1(n86_adj_3796), .I2(n167_adj_3797), 
            .I3(GND_net), .O(n16571[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3481_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3481_2 (.CI(GND_net), .I0(n86_adj_3796), .I1(n167_adj_3797), 
            .CO(n35731));
    SB_LUT4 add_3389_17_lut (.I0(GND_net), .I1(n15640[14]), .I2(GND_net), 
            .I3(n35730), .O(n15399[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3389_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3389_16_lut (.I0(GND_net), .I1(n15640[13]), .I2(GND_net), 
            .I3(n35729), .O(n15399[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3389_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3389_16 (.CI(n35729), .I0(n15640[13]), .I1(GND_net), 
            .CO(n35730));
    SB_LUT4 add_3389_15_lut (.I0(GND_net), .I1(n15640[12]), .I2(GND_net), 
            .I3(n35728), .O(n15399[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3389_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3389_15 (.CI(n35728), .I0(n15640[12]), .I1(GND_net), 
            .CO(n35729));
    SB_LUT4 add_3389_14_lut (.I0(GND_net), .I1(n15640[11]), .I2(GND_net), 
            .I3(n35727), .O(n15399[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3389_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3389_14 (.CI(n35727), .I0(n15640[11]), .I1(GND_net), 
            .CO(n35728));
    SB_LUT4 add_3389_13_lut (.I0(GND_net), .I1(n15640[10]), .I2(GND_net), 
            .I3(n35726), .O(n15399[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3389_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3389_13 (.CI(n35726), .I0(n15640[10]), .I1(GND_net), 
            .CO(n35727));
    SB_LUT4 add_3389_12_lut (.I0(GND_net), .I1(n15640[9]), .I2(GND_net), 
            .I3(n35725), .O(n15399[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3389_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3389_12 (.CI(n35725), .I0(n15640[9]), .I1(GND_net), .CO(n35726));
    SB_LUT4 add_3389_11_lut (.I0(GND_net), .I1(n15640[8]), .I2(GND_net), 
            .I3(n35724), .O(n15399[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3389_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3389_11 (.CI(n35724), .I0(n15640[8]), .I1(GND_net), .CO(n35725));
    SB_LUT4 add_3389_10_lut (.I0(GND_net), .I1(n15640[7]), .I2(GND_net), 
            .I3(n35723), .O(n15399[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3389_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3389_10 (.CI(n35723), .I0(n15640[7]), .I1(GND_net), .CO(n35724));
    SB_LUT4 add_3389_9_lut (.I0(GND_net), .I1(n15640[6]), .I2(GND_net), 
            .I3(n35722), .O(n15399[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3389_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3389_9 (.CI(n35722), .I0(n15640[6]), .I1(GND_net), .CO(n35723));
    SB_LUT4 add_3389_8_lut (.I0(GND_net), .I1(n15640[5]), .I2(n725_adj_3798), 
            .I3(n35721), .O(n15399[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3389_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3389_8 (.CI(n35721), .I0(n15640[5]), .I1(n725_adj_3798), 
            .CO(n35722));
    SB_LUT4 add_3389_7_lut (.I0(GND_net), .I1(n15640[4]), .I2(n628_adj_3799), 
            .I3(n35720), .O(n15399[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3389_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3389_7 (.CI(n35720), .I0(n15640[4]), .I1(n628_adj_3799), 
            .CO(n35721));
    SB_LUT4 add_3389_6_lut (.I0(GND_net), .I1(n15640[3]), .I2(n531_adj_3800), 
            .I3(n35719), .O(n15399[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3389_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3389_6 (.CI(n35719), .I0(n15640[3]), .I1(n531_adj_3800), 
            .CO(n35720));
    SB_LUT4 add_3389_5_lut (.I0(GND_net), .I1(n15640[2]), .I2(n434_adj_3801), 
            .I3(n35718), .O(n15399[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3389_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3389_5 (.CI(n35718), .I0(n15640[2]), .I1(n434_adj_3801), 
            .CO(n35719));
    SB_LUT4 add_3389_4_lut (.I0(GND_net), .I1(n15640[1]), .I2(n337_adj_3802), 
            .I3(n35717), .O(n15399[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3389_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3389_4 (.CI(n35717), .I0(n15640[1]), .I1(n337_adj_3802), 
            .CO(n35718));
    SB_LUT4 add_3389_3_lut (.I0(GND_net), .I1(n15640[0]), .I2(n240_adj_3803), 
            .I3(n35716), .O(n15399[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3389_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3389_3 (.CI(n35716), .I0(n15640[0]), .I1(n240_adj_3803), 
            .CO(n35717));
    SB_LUT4 add_3389_2_lut (.I0(GND_net), .I1(n50_adj_3804), .I2(n143_adj_3805), 
            .I3(GND_net), .O(n15399[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3389_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3389_2 (.CI(GND_net), .I0(n50_adj_3804), .I1(n143_adj_3805), 
            .CO(n35716));
    SB_LUT4 add_3489_7_lut (.I0(GND_net), .I1(n41719), .I2(n658_adj_3806), 
            .I3(n35715), .O(n16629[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3489_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3489_6_lut (.I0(GND_net), .I1(n16637[3]), .I2(n558_adj_3807), 
            .I3(n35714), .O(n16629[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3489_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3489_6 (.CI(n35714), .I0(n16637[3]), .I1(n558_adj_3807), 
            .CO(n35715));
    SB_LUT4 add_3489_5_lut (.I0(GND_net), .I1(n16637[2]), .I2(n464_adj_3808), 
            .I3(n35713), .O(n16629[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3489_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3489_5 (.CI(n35713), .I0(n16637[2]), .I1(n464_adj_3808), 
            .CO(n35714));
    SB_LUT4 add_3489_4_lut (.I0(GND_net), .I1(n16644[1]), .I2(n370_adj_3809), 
            .I3(n35712), .O(n16629[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3489_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3489_4 (.CI(n35712), .I0(n16644[1]), .I1(n370_adj_3809), 
            .CO(n35713));
    SB_LUT4 add_3489_3_lut (.I0(GND_net), .I1(n16637[0]), .I2(n276_adj_3810), 
            .I3(n35711), .O(n16629[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3489_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3489_3 (.CI(n35711), .I0(n16637[0]), .I1(n276_adj_3810), 
            .CO(n35712));
    SB_LUT4 add_3489_2_lut (.I0(GND_net), .I1(n86_adj_3796), .I2(n182_adj_3811), 
            .I3(GND_net), .O(n16629[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3489_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3489_2 (.CI(GND_net), .I0(n86_adj_3796), .I1(n182_adj_3811), 
            .CO(n35711));
    SB_LUT4 add_3404_16_lut (.I0(GND_net), .I1(n15850[13]), .I2(GND_net), 
            .I3(n35710), .O(n15640[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3404_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3404_15_lut (.I0(GND_net), .I1(n15850[12]), .I2(GND_net), 
            .I3(n35709), .O(n15640[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3404_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3404_15 (.CI(n35709), .I0(n15850[12]), .I1(GND_net), 
            .CO(n35710));
    SB_LUT4 add_3404_14_lut (.I0(GND_net), .I1(n15850[11]), .I2(GND_net), 
            .I3(n35708), .O(n15640[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3404_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3404_14 (.CI(n35708), .I0(n15850[11]), .I1(GND_net), 
            .CO(n35709));
    SB_LUT4 add_3404_13_lut (.I0(GND_net), .I1(n15850[10]), .I2(GND_net), 
            .I3(n35707), .O(n15640[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3404_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3404_13 (.CI(n35707), .I0(n15850[10]), .I1(GND_net), 
            .CO(n35708));
    SB_LUT4 add_3404_12_lut (.I0(GND_net), .I1(n15850[9]), .I2(GND_net), 
            .I3(n35706), .O(n15640[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3404_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_12_i205_2_lut (.I0(\Kd[3] ), .I1(n57[4]), .I2(GND_net), 
            .I3(GND_net), .O(n304));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i205_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_3404_12 (.CI(n35706), .I0(n15850[9]), .I1(GND_net), .CO(n35707));
    SB_LUT4 add_3404_11_lut (.I0(GND_net), .I1(n15850[8]), .I2(GND_net), 
            .I3(n35705), .O(n15640[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3404_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3404_11 (.CI(n35705), .I0(n15850[8]), .I1(GND_net), .CO(n35706));
    SB_LUT4 add_3404_10_lut (.I0(GND_net), .I1(n15850[7]), .I2(GND_net), 
            .I3(n35704), .O(n15640[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3404_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3404_10 (.CI(n35704), .I0(n15850[7]), .I1(GND_net), .CO(n35705));
    SB_LUT4 add_3404_9_lut (.I0(GND_net), .I1(n15850[6]), .I2(GND_net), 
            .I3(n35703), .O(n15640[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3404_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3404_9 (.CI(n35703), .I0(n15850[6]), .I1(GND_net), .CO(n35704));
    SB_LUT4 add_3404_8_lut (.I0(GND_net), .I1(n15850[5]), .I2(n728_adj_3812), 
            .I3(n35702), .O(n15640[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3404_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3404_8 (.CI(n35702), .I0(n15850[5]), .I1(n728_adj_3812), 
            .CO(n35703));
    SB_LUT4 add_3404_7_lut (.I0(GND_net), .I1(n15850[4]), .I2(n631_adj_3813), 
            .I3(n35701), .O(n15640[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3404_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3404_7 (.CI(n35701), .I0(n15850[4]), .I1(n631_adj_3813), 
            .CO(n35702));
    SB_LUT4 add_3404_6_lut (.I0(GND_net), .I1(n15850[3]), .I2(n534_adj_3814), 
            .I3(n35700), .O(n15640[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3404_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3404_6 (.CI(n35700), .I0(n15850[3]), .I1(n534_adj_3814), 
            .CO(n35701));
    SB_LUT4 add_3404_5_lut (.I0(GND_net), .I1(n15850[2]), .I2(n437_adj_3815), 
            .I3(n35699), .O(n15640[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3404_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3404_5 (.CI(n35699), .I0(n15850[2]), .I1(n437_adj_3815), 
            .CO(n35700));
    SB_LUT4 add_3404_4_lut (.I0(GND_net), .I1(n15850[1]), .I2(n340_adj_3816), 
            .I3(n35698), .O(n15640[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3404_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3404_4 (.CI(n35698), .I0(n15850[1]), .I1(n340_adj_3816), 
            .CO(n35699));
    SB_LUT4 add_3404_3_lut (.I0(GND_net), .I1(n15850[0]), .I2(n243_adj_3817), 
            .I3(n35697), .O(n15640[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3404_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3404_3 (.CI(n35697), .I0(n15850[0]), .I1(n243_adj_3817), 
            .CO(n35698));
    SB_LUT4 add_3404_2_lut (.I0(GND_net), .I1(n53_adj_3818), .I2(n146_adj_3819), 
            .I3(GND_net), .O(n15640[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3404_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3404_2 (.CI(GND_net), .I0(n53_adj_3818), .I1(n146_adj_3819), 
            .CO(n35697));
    SB_LUT4 add_3488_8_lut (.I0(GND_net), .I1(n16629[5]), .I2(n752_adj_3820), 
            .I3(n35696), .O(n16620[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3488_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3488_7_lut (.I0(GND_net), .I1(n16629[4]), .I2(n658_adj_3806), 
            .I3(n35695), .O(n16620[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3488_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3488_7 (.CI(n35695), .I0(n16629[4]), .I1(n658_adj_3806), 
            .CO(n35696));
    SB_LUT4 add_3488_6_lut (.I0(GND_net), .I1(n16629[3]), .I2(n558_adj_3807), 
            .I3(n35694), .O(n16620[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3488_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3488_6 (.CI(n35694), .I0(n16629[3]), .I1(n558_adj_3807), 
            .CO(n35695));
    SB_LUT4 state_23__I_0_add_2_20_lut (.I0(GND_net), .I1(\motor_state[18] ), 
            .I2(n58[18]), .I3(n34233), .O(\PID_CONTROLLER.err_31__N_2825 [18])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3231_10 (.CI(n35130), .I0(n12732[7]), .I1(GND_net), .CO(n35131));
    SB_CARRY add_13_add_1_20061_add_1_17 (.CI(n34870), .I0(n282[15]), .I1(n61[15]), 
            .CO(n34871));
    SB_LUT4 add_13_add_1_20061_add_1_16_lut (.I0(GND_net), .I1(n282[14]), 
            .I2(n61[14]), .I3(n34869), .O(n63[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_13_add_1_20061_add_1_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3301_5 (.CI(n34587), .I0(n14168[2]), .I1(n326), .CO(n34588));
    SB_CARRY add_3272_11 (.CI(n34398), .I0(n13594[8]), .I1(GND_net), .CO(n34399));
    SB_LUT4 add_3488_5_lut (.I0(GND_net), .I1(n16629[2]), .I2(n464_adj_3808), 
            .I3(n35693), .O(n16620[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3488_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3272_10_lut (.I0(GND_net), .I1(n13594[7]), .I2(GND_net), 
            .I3(n34397), .O(n13109[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3272_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3301_4_lut (.I0(GND_net), .I1(n14168[1]), .I2(n253), .I3(n34586), 
            .O(n13734[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3301_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3272_10 (.CI(n34397), .I0(n13594[7]), .I1(GND_net), .CO(n34398));
    SB_CARRY add_3301_4 (.CI(n34586), .I0(n14168[1]), .I1(n253), .CO(n34587));
    SB_CARRY state_23__I_0_add_2_20 (.CI(n34233), .I0(\motor_state[18] ), 
            .I1(n58[18]), .CO(n34234));
    SB_LUT4 add_3272_9_lut (.I0(GND_net), .I1(n13594[6]), .I2(GND_net), 
            .I3(n34396), .O(n13109[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3272_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3231_9_lut (.I0(GND_net), .I1(n12732[6]), .I2(GND_net), 
            .I3(n35129), .O(n12157[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3231_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3301_3_lut (.I0(GND_net), .I1(n14168[0]), .I2(n180), .I3(n34585), 
            .O(n13734[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3301_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3272_9 (.CI(n34396), .I0(n13594[6]), .I1(GND_net), .CO(n34397));
    SB_LUT4 add_3272_8_lut (.I0(GND_net), .I1(n13594[5]), .I2(n707_adj_3822), 
            .I3(n34395), .O(n13109[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3272_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3301_3 (.CI(n34585), .I0(n14168[0]), .I1(n180), .CO(n34586));
    SB_CARRY add_3488_5 (.CI(n35693), .I0(n16629[2]), .I1(n464_adj_3808), 
            .CO(n35694));
    SB_CARRY add_3272_8 (.CI(n34395), .I0(n13594[5]), .I1(n707_adj_3822), 
            .CO(n34396));
    SB_LUT4 add_3488_4_lut (.I0(GND_net), .I1(n16629[1]), .I2(n370_adj_3809), 
            .I3(n35692), .O(n16620[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3488_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3488_4 (.CI(n35692), .I0(n16629[1]), .I1(n370_adj_3809), 
            .CO(n35693));
    SB_LUT4 mult_10_i304_2_lut (.I0(\Kp[4] ), .I1(\PID_CONTROLLER.err[21] ), 
            .I2(GND_net), .I3(GND_net), .O(n452));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i304_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i471_2_lut (.I0(\Kp[7] ), .I1(\PID_CONTROLLER.err[7] ), 
            .I2(GND_net), .I3(GND_net), .O(n701_adj_3413));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i471_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 sub_11_inv_0_i16_1_lut (.I0(\PID_CONTROLLER.err[15] ), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n64[15]));   // verilog/motorControl.v(43[31:45])
    defparam sub_11_inv_0_i16_1_lut.LUT_INIT = 16'h5555;
    SB_DFF Kd_delay_counter_1015__i2 (.Q(Kd_delay_counter[2]), .C(clk32MHz), 
           .D(n69[2]));   // verilog/motorControl.v(55[27:47])
    SB_LUT4 add_3301_2_lut (.I0(GND_net), .I1(n35), .I2(n107), .I3(GND_net), 
            .O(n13734[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3301_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3488_3_lut (.I0(GND_net), .I1(n16629[0]), .I2(n276_adj_3810), 
            .I3(n35691), .O(n16620[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3488_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3488_3 (.CI(n35691), .I0(n16629[0]), .I1(n276_adj_3810), 
            .CO(n35692));
    SB_LUT4 add_3488_2_lut (.I0(GND_net), .I1(n86_adj_3796), .I2(n182_adj_3811), 
            .I3(GND_net), .O(n16620[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3488_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3488_2 (.CI(GND_net), .I0(n86_adj_3796), .I1(n182_adj_3811), 
            .CO(n35691));
    SB_LUT4 add_3418_15_lut (.I0(GND_net), .I1(n16031[12]), .I2(GND_net), 
            .I3(n35690), .O(n15850[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3418_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3418_14_lut (.I0(GND_net), .I1(n16031[11]), .I2(GND_net), 
            .I3(n35689), .O(n15850[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3418_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3418_14 (.CI(n35689), .I0(n16031[11]), .I1(GND_net), 
            .CO(n35690));
    SB_LUT4 add_3418_13_lut (.I0(GND_net), .I1(n16031[10]), .I2(GND_net), 
            .I3(n35688), .O(n15850[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3418_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3418_13 (.CI(n35688), .I0(n16031[10]), .I1(GND_net), 
            .CO(n35689));
    SB_LUT4 add_3418_12_lut (.I0(GND_net), .I1(n16031[9]), .I2(GND_net), 
            .I3(n35687), .O(n15850[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3418_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3418_12 (.CI(n35687), .I0(n16031[9]), .I1(GND_net), .CO(n35688));
    SB_LUT4 add_3418_11_lut (.I0(GND_net), .I1(n16031[8]), .I2(GND_net), 
            .I3(n35686), .O(n15850[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3418_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3418_11 (.CI(n35686), .I0(n16031[8]), .I1(GND_net), .CO(n35687));
    SB_LUT4 add_3418_10_lut (.I0(GND_net), .I1(n16031[7]), .I2(GND_net), 
            .I3(n35685), .O(n15850[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3418_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3272_7_lut (.I0(GND_net), .I1(n13594[4]), .I2(n610_adj_3823), 
            .I3(n34394), .O(n13109[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3272_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3418_10 (.CI(n35685), .I0(n16031[7]), .I1(GND_net), .CO(n35686));
    SB_DFF Kd_delay_counter_1015__i3 (.Q(Kd_delay_counter[3]), .C(clk32MHz), 
           .D(n69[3]));   // verilog/motorControl.v(55[27:47])
    SB_DFF Kd_delay_counter_1015__i4 (.Q(Kd_delay_counter[4]), .C(clk32MHz), 
           .D(n69[4]));   // verilog/motorControl.v(55[27:47])
    SB_DFF Kd_delay_counter_1015__i5 (.Q(Kd_delay_counter[5]), .C(clk32MHz), 
           .D(n69[5]));   // verilog/motorControl.v(55[27:47])
    SB_DFF Kd_delay_counter_1015__i6 (.Q(Kd_delay_counter[6]), .C(clk32MHz), 
           .D(n69[6]));   // verilog/motorControl.v(55[27:47])
    SB_DFF pwm_count_1016__i1 (.Q(pwm_count[1]), .C(clk32MHz), .D(n67[1]));   // verilog/motorControl.v(110[18:29])
    SB_LUT4 add_3067_12_lut (.I0(GND_net), .I1(n8274[9]), .I2(GND_net), 
            .I3(n35487), .O(n8253[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3067_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3418_9_lut (.I0(GND_net), .I1(n16031[6]), .I2(GND_net), 
            .I3(n35684), .O(n15850[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3418_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 state_23__I_0_add_2_19_lut (.I0(GND_net), .I1(\motor_state[17] ), 
            .I2(n58[17]), .I3(n34232), .O(\PID_CONTROLLER.err_31__N_2825 [17])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3059_6_lut (.I0(GND_net), .I1(n8078[3]), .I2(n498_adj_3825), 
            .I3(n35301), .O(n8049[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3059_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3272_7 (.CI(n34394), .I0(n13594[4]), .I1(n610_adj_3823), 
            .CO(n34395));
    SB_CARRY add_3231_9 (.CI(n35129), .I0(n12732[6]), .I1(GND_net), .CO(n35130));
    SB_CARRY add_3301_2 (.CI(GND_net), .I0(n35), .I1(n107), .CO(n34585));
    SB_LUT4 add_3272_6_lut (.I0(GND_net), .I1(n13594[3]), .I2(n513_adj_3826), 
            .I3(n34393), .O(n13109[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3272_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3231_8_lut (.I0(GND_net), .I1(n12732[5]), .I2(n545), .I3(n35128), 
            .O(n12157[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3231_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3272_6 (.CI(n34393), .I0(n13594[3]), .I1(n513_adj_3826), 
            .CO(n34394));
    SB_LUT4 add_3142_28_lut (.I0(GND_net), .I1(n10671[25]), .I2(GND_net), 
            .I3(n34584), .O(n9929[26])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3142_28_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3272_5_lut (.I0(GND_net), .I1(n13594[2]), .I2(n416_adj_3827), 
            .I3(n34392), .O(n13109[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3272_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_13_add_1_20061_add_1_16 (.CI(n34869), .I0(n282[14]), .I1(n61[14]), 
            .CO(n34870));
    SB_CARRY add_3272_5 (.CI(n34392), .I0(n13594[2]), .I1(n416_adj_3827), 
            .CO(n34393));
    SB_CARRY add_3063_4 (.CI(n35397), .I0(n8184[1]), .I1(n316_adj_3742), 
            .CO(n35398));
    SB_CARRY add_3059_6 (.CI(n35301), .I0(n8078[3]), .I1(n498_adj_3825), 
            .CO(n35302));
    SB_LUT4 add_3142_27_lut (.I0(GND_net), .I1(n10671[24]), .I2(GND_net), 
            .I3(n34583), .O(n9929[25])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3142_27_lut.LUT_INIT = 16'hC33C;
    SB_CARRY state_23__I_0_add_2_19 (.CI(n34232), .I0(\motor_state[17] ), 
            .I1(n58[17]), .CO(n34233));
    SB_CARRY add_3231_8 (.CI(n35128), .I0(n12732[5]), .I1(n545), .CO(n35129));
    SB_LUT4 add_13_add_1_20061_add_1_15_lut (.I0(GND_net), .I1(n282[13]), 
            .I2(n61[13]), .I3(n34868), .O(n63[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_13_add_1_20061_add_1_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3142_27 (.CI(n34583), .I0(n10671[24]), .I1(GND_net), 
            .CO(n34584));
    SB_LUT4 add_3142_26_lut (.I0(GND_net), .I1(n10671[23]), .I2(GND_net), 
            .I3(n34582), .O(n9929[24])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3142_26_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3272_4_lut (.I0(GND_net), .I1(n13594[1]), .I2(n319_adj_3828), 
            .I3(n34391), .O(n13109[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3272_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_13_add_1_20061_add_1_15 (.CI(n34868), .I0(n282[13]), .I1(n61[13]), 
            .CO(n34869));
    SB_CARRY add_3142_26 (.CI(n34582), .I0(n10671[23]), .I1(GND_net), 
            .CO(n34583));
    SB_LUT4 add_3142_25_lut (.I0(GND_net), .I1(n10671[22]), .I2(GND_net), 
            .I3(n34581), .O(n9929[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3142_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3272_4 (.CI(n34391), .I0(n13594[1]), .I1(n319_adj_3828), 
            .CO(n34392));
    SB_LUT4 add_3272_3_lut (.I0(GND_net), .I1(n13594[0]), .I2(n222_adj_3829), 
            .I3(n34390), .O(n13109[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3272_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3231_7_lut (.I0(GND_net), .I1(n12732[4]), .I2(n472), .I3(n35127), 
            .O(n12157[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3231_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_13_add_1_20061_add_1_14_lut (.I0(GND_net), .I1(n282[12]), 
            .I2(n61[12]), .I3(n34867), .O(n63[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_13_add_1_20061_add_1_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3418_9 (.CI(n35684), .I0(n16031[6]), .I1(GND_net), .CO(n35685));
    SB_CARRY add_3142_25 (.CI(n34581), .I0(n10671[22]), .I1(GND_net), 
            .CO(n34582));
    SB_LUT4 add_3142_24_lut (.I0(GND_net), .I1(n10671[21]), .I2(GND_net), 
            .I3(n34580), .O(n9929[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3142_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3418_8_lut (.I0(GND_net), .I1(n16031[5]), .I2(n731_adj_3830), 
            .I3(n35683), .O(n15850[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3418_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3074_8_lut (.I0(GND_net), .I1(n8393[5]), .I2(n737_adj_3831), 
            .I3(n35588), .O(n8379[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3074_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3418_8 (.CI(n35683), .I0(n16031[5]), .I1(n731_adj_3830), 
            .CO(n35684));
    SB_CARRY add_3272_3 (.CI(n34390), .I0(n13594[0]), .I1(n222_adj_3829), 
            .CO(n34391));
    SB_LUT4 add_3418_7_lut (.I0(GND_net), .I1(n16031[4]), .I2(n634_adj_3832), 
            .I3(n35682), .O(n15850[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3418_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3418_7 (.CI(n35682), .I0(n16031[4]), .I1(n634_adj_3832), 
            .CO(n35683));
    SB_CARRY add_3231_7 (.CI(n35127), .I0(n12732[4]), .I1(n472), .CO(n35128));
    SB_LUT4 add_3418_6_lut (.I0(GND_net), .I1(n16031[3]), .I2(n537_adj_3833), 
            .I3(n35681), .O(n15850[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3418_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3074_8 (.CI(n35588), .I0(n8393[5]), .I1(n737_adj_3831), 
            .CO(n35589));
    SB_LUT4 add_3272_2_lut (.I0(GND_net), .I1(n32_adj_3834), .I2(n125_adj_3835), 
            .I3(GND_net), .O(n13109[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3272_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3418_6 (.CI(n35681), .I0(n16031[3]), .I1(n537_adj_3833), 
            .CO(n35682));
    SB_CARRY add_13_add_1_20061_add_1_14 (.CI(n34867), .I0(n282[12]), .I1(n61[12]), 
            .CO(n34868));
    SB_CARRY add_3142_24 (.CI(n34580), .I0(n10671[21]), .I1(GND_net), 
            .CO(n34581));
    SB_LUT4 add_3074_7_lut (.I0(GND_net), .I1(n8393[4]), .I2(n640_adj_3836), 
            .I3(n35587), .O(n8379[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3074_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3418_5_lut (.I0(GND_net), .I1(n16031[2]), .I2(n440_adj_3837), 
            .I3(n35680), .O(n15850[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3418_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3142_23_lut (.I0(GND_net), .I1(n10671[20]), .I2(GND_net), 
            .I3(n34579), .O(n9929[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3142_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3418_5 (.CI(n35680), .I0(n16031[2]), .I1(n440_adj_3837), 
            .CO(n35681));
    SB_LUT4 state_23__I_0_add_2_18_lut (.I0(GND_net), .I1(\motor_state[16] ), 
            .I2(n58[16]), .I3(n34231), .O(\PID_CONTROLLER.err_31__N_2825 [16])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3418_4_lut (.I0(GND_net), .I1(n16031[1]), .I2(n343_adj_3839), 
            .I3(n35679), .O(n15850[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3418_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3074_7 (.CI(n35587), .I0(n8393[4]), .I1(n640_adj_3836), 
            .CO(n35588));
    SB_CARRY add_3272_2 (.CI(GND_net), .I0(n32_adj_3834), .I1(n125_adj_3835), 
            .CO(n34390));
    SB_CARRY add_3418_4 (.CI(n35679), .I0(n16031[1]), .I1(n343_adj_3839), 
            .CO(n35680));
    SB_LUT4 add_3294_22_lut (.I0(GND_net), .I1(n14035[19]), .I2(GND_net), 
            .I3(n34389), .O(n13594[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3294_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3418_3_lut (.I0(GND_net), .I1(n16031[0]), .I2(n246_adj_3840), 
            .I3(n35678), .O(n15850[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3418_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3059_5_lut (.I0(GND_net), .I1(n8078[2]), .I2(n401_adj_3841), 
            .I3(n35300), .O(n8049[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3059_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3074_6_lut (.I0(GND_net), .I1(n8393[3]), .I2(n543_adj_3842), 
            .I3(n35586), .O(n8379[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3074_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3231_6_lut (.I0(GND_net), .I1(n12732[3]), .I2(n399), .I3(n35126), 
            .O(n12157[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3231_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_13_add_1_20061_add_1_13_lut (.I0(GND_net), .I1(n282[11]), 
            .I2(n61[11]), .I3(n34866), .O(n63[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_13_add_1_20061_add_1_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_13_add_1_20061_add_1_13 (.CI(n34866), .I0(n282[11]), .I1(n61[11]), 
            .CO(n34867));
    SB_CARRY add_3418_3 (.CI(n35678), .I0(n16031[0]), .I1(n246_adj_3840), 
            .CO(n35679));
    SB_CARRY add_3142_23 (.CI(n34579), .I0(n10671[20]), .I1(GND_net), 
            .CO(n34580));
    SB_LUT4 add_3142_22_lut (.I0(GND_net), .I1(n10671[19]), .I2(GND_net), 
            .I3(n34578), .O(n9929[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3142_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3074_6 (.CI(n35586), .I0(n8393[3]), .I1(n543_adj_3842), 
            .CO(n35587));
    SB_CARRY add_3142_22 (.CI(n34578), .I0(n10671[19]), .I1(GND_net), 
            .CO(n34579));
    SB_CARRY state_23__I_0_add_2_18 (.CI(n34231), .I0(\motor_state[16] ), 
            .I1(n58[16]), .CO(n34232));
    SB_LUT4 add_3294_21_lut (.I0(GND_net), .I1(n14035[18]), .I2(GND_net), 
            .I3(n34388), .O(n13594[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3294_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3418_2_lut (.I0(GND_net), .I1(n56_adj_3843), .I2(n149_adj_3844), 
            .I3(GND_net), .O(n15850[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3418_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3294_21 (.CI(n34388), .I0(n14035[18]), .I1(GND_net), 
            .CO(n34389));
    SB_LUT4 add_3074_5_lut (.I0(GND_net), .I1(n8393[2]), .I2(n446), .I3(n35585), 
            .O(n8379[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3074_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_13_add_1_20061_add_1_12_lut (.I0(GND_net), .I1(n282[10]), 
            .I2(n61[10]), .I3(n34865), .O(n63[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_13_add_1_20061_add_1_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3142_21_lut (.I0(GND_net), .I1(n10671[18]), .I2(GND_net), 
            .I3(n34577), .O(n9929[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3142_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3142_21 (.CI(n34577), .I0(n10671[18]), .I1(GND_net), 
            .CO(n34578));
    SB_LUT4 add_3294_20_lut (.I0(GND_net), .I1(n14035[17]), .I2(GND_net), 
            .I3(n34387), .O(n13594[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3294_20_lut.LUT_INIT = 16'hC33C;
    SB_DFF pwm_count_1016__i2 (.Q(pwm_count[2]), .C(clk32MHz), .D(n67[2]));   // verilog/motorControl.v(110[18:29])
    SB_CARRY add_3294_20 (.CI(n34387), .I0(n14035[17]), .I1(GND_net), 
            .CO(n34388));
    SB_DFF pwm_count_1016__i3 (.Q(pwm_count[3]), .C(clk32MHz), .D(n67[3]));   // verilog/motorControl.v(110[18:29])
    SB_DFF pwm_count_1016__i4 (.Q(pwm_count[4]), .C(clk32MHz), .D(n67[4]));   // verilog/motorControl.v(110[18:29])
    SB_DFF pwm_count_1016__i5 (.Q(pwm_count[5]), .C(clk32MHz), .D(n67[5]));   // verilog/motorControl.v(110[18:29])
    SB_DFF pwm_count_1016__i6 (.Q(pwm_count[6]), .C(clk32MHz), .D(n67[6]));   // verilog/motorControl.v(110[18:29])
    SB_DFF pwm_count_1016__i7 (.Q(pwm_count[7]), .C(clk32MHz), .D(n67[7]));   // verilog/motorControl.v(110[18:29])
    SB_DFF pwm_count_1016__i8 (.Q(pwm_count[8]), .C(clk32MHz), .D(n67[8]));   // verilog/motorControl.v(110[18:29])
    SB_DFFE \PID_CONTROLLER.integral_1017__i1  (.Q(\PID_CONTROLLER.integral [1]), 
            .C(clk32MHz), .E(n55_adj_3594), .D(n66[1]));   // verilog/motorControl.v(41[21:33])
    SB_DFF \PID_CONTROLLER.err_prev__i1  (.Q(\PID_CONTROLLER.err_prev[0] ), 
           .C(clk32MHz), .D(n23589));   // verilog/motorControl.v(38[14] 59[8])
    SB_DFFE \PID_CONTROLLER.integral_1017__i2  (.Q(\PID_CONTROLLER.integral [2]), 
            .C(clk32MHz), .E(n55_adj_3594), .D(n66[2]));   // verilog/motorControl.v(41[21:33])
    SB_DFFE \PID_CONTROLLER.integral_1017__i3  (.Q(\PID_CONTROLLER.integral [3]), 
            .C(clk32MHz), .E(n55_adj_3594), .D(n66[3]));   // verilog/motorControl.v(41[21:33])
    SB_DFFE \PID_CONTROLLER.integral_1017__i4  (.Q(\PID_CONTROLLER.integral [4]), 
            .C(clk32MHz), .E(n55_adj_3594), .D(n66[4]));   // verilog/motorControl.v(41[21:33])
    SB_DFFE \PID_CONTROLLER.integral_1017__i5  (.Q(\PID_CONTROLLER.integral [5]), 
            .C(clk32MHz), .E(n55_adj_3594), .D(n66[5]));   // verilog/motorControl.v(41[21:33])
    SB_DFFE \PID_CONTROLLER.integral_1017__i6  (.Q(\PID_CONTROLLER.integral [6]), 
            .C(clk32MHz), .E(n55_adj_3594), .D(n66[6]));   // verilog/motorControl.v(41[21:33])
    SB_DFFE \PID_CONTROLLER.integral_1017__i7  (.Q(\PID_CONTROLLER.integral [7]), 
            .C(clk32MHz), .E(n55_adj_3594), .D(n66[7]));   // verilog/motorControl.v(41[21:33])
    SB_DFFE \PID_CONTROLLER.integral_1017__i8  (.Q(\PID_CONTROLLER.integral [8]), 
            .C(clk32MHz), .E(n55_adj_3594), .D(n66[8]));   // verilog/motorControl.v(41[21:33])
    SB_DFFE \PID_CONTROLLER.integral_1017__i9  (.Q(\PID_CONTROLLER.integral [9]), 
            .C(clk32MHz), .E(n55_adj_3594), .D(n66[9]));   // verilog/motorControl.v(41[21:33])
    SB_LUT4 add_3294_19_lut (.I0(GND_net), .I1(n14035[16]), .I2(GND_net), 
            .I3(n34386), .O(n13594[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3294_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 state_23__I_0_add_2_17_lut (.I0(GND_net), .I1(\motor_state[15] ), 
            .I2(n58[15]), .I3(n34230), .O(\PID_CONTROLLER.err_31__N_2825 [15])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3294_19 (.CI(n34386), .I0(n14035[16]), .I1(GND_net), 
            .CO(n34387));
    SB_LUT4 add_3063_3_lut (.I0(GND_net), .I1(n8184[0]), .I2(n219), .I3(n35396), 
            .O(n8159[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3063_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_13_add_1_20061_add_1_12 (.CI(n34865), .I0(n282[10]), .I1(n61[10]), 
            .CO(n34866));
    SB_CARRY add_3059_5 (.CI(n35300), .I0(n8078[2]), .I1(n401_adj_3841), 
            .CO(n35301));
    SB_CARRY add_3231_6 (.CI(n35126), .I0(n12732[3]), .I1(n399), .CO(n35127));
    SB_LUT4 add_13_add_1_20061_add_1_11_lut (.I0(GND_net), .I1(n282[9]), 
            .I2(n61[9]), .I3(n34864), .O(n63[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_13_add_1_20061_add_1_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3142_20_lut (.I0(GND_net), .I1(n10671[17]), .I2(GND_net), 
            .I3(n34576), .O(n9929[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3142_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3418_2 (.CI(GND_net), .I0(n56_adj_3843), .I1(n149_adj_3844), 
            .CO(n35678));
    SB_LUT4 mux_24_i1_3_lut (.I0(\PID_CONTROLLER.result [0]), .I1(n70[0]), 
            .I2(n421), .I3(GND_net), .O(n471));   // verilog/motorControl.v(49[18] 51[12])
    defparam mux_24_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_10_i101_2_lut (.I0(\Kp[1] ), .I1(\PID_CONTROLLER.err[17] ), 
            .I2(GND_net), .I3(GND_net), .O(n149_adj_3844));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i101_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i38_2_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err[18] ), 
            .I2(GND_net), .I3(GND_net), .O(n56_adj_3843));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i38_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i365_2_lut (.I0(\Kd[5] ), .I1(n57[19]), .I2(GND_net), 
            .I3(GND_net), .O(n543_adj_3842));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i365_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i270_2_lut (.I0(\Kd[4] ), .I1(n57[4]), .I2(GND_net), 
            .I3(GND_net), .O(n401_adj_3841));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i270_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i166_2_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err[17] ), 
            .I2(GND_net), .I3(GND_net), .O(n246_adj_3840));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i166_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i231_2_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err[17] ), 
            .I2(GND_net), .I3(GND_net), .O(n343_adj_3839));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i231_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 state_23__I_0_inv_0_i17_1_lut (.I0(setpoint[16]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n58[16]));   // verilog/motorControl.v(39[14:30])
    defparam state_23__I_0_inv_0_i17_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mux_24_i2_3_lut (.I0(\PID_CONTROLLER.result [1]), .I1(n70[1]), 
            .I2(n421), .I3(GND_net), .O(n470));   // verilog/motorControl.v(49[18] 51[12])
    defparam mux_24_i2_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_10_i296_2_lut (.I0(\Kp[4] ), .I1(\PID_CONTROLLER.err[17] ), 
            .I2(GND_net), .I3(GND_net), .O(n440_adj_3837));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i296_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i430_2_lut (.I0(\Kd[6] ), .I1(n57[19]), .I2(GND_net), 
            .I3(GND_net), .O(n640_adj_3836));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i430_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_24_i3_3_lut (.I0(\PID_CONTROLLER.result [2]), .I1(n70[2]), 
            .I2(n421), .I3(GND_net), .O(n469));   // verilog/motorControl.v(49[18] 51[12])
    defparam mux_24_i3_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_10_i85_2_lut (.I0(\Kp[1] ), .I1(\PID_CONTROLLER.err[9] ), 
            .I2(GND_net), .I3(GND_net), .O(n125_adj_3835));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i85_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i22_2_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err[10] ), 
            .I2(GND_net), .I3(GND_net), .O(n32_adj_3834));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i22_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i361_2_lut (.I0(\Kp[5] ), .I1(\PID_CONTROLLER.err[17] ), 
            .I2(GND_net), .I3(GND_net), .O(n537_adj_3833));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i361_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i426_2_lut (.I0(\Kp[6] ), .I1(\PID_CONTROLLER.err[17] ), 
            .I2(GND_net), .I3(GND_net), .O(n634_adj_3832));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i426_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i495_2_lut (.I0(\Kd[7] ), .I1(n57[19]), .I2(GND_net), 
            .I3(GND_net), .O(n737_adj_3831));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i495_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_24_i4_3_lut (.I0(\PID_CONTROLLER.result [3]), .I1(n70[3]), 
            .I2(n421), .I3(GND_net), .O(n468));   // verilog/motorControl.v(49[18] 51[12])
    defparam mux_24_i4_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_10_i491_2_lut (.I0(\Kp[7] ), .I1(\PID_CONTROLLER.err[17] ), 
            .I2(GND_net), .I3(GND_net), .O(n731_adj_3830));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i491_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i150_2_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err[9] ), 
            .I2(GND_net), .I3(GND_net), .O(n222_adj_3829));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i150_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i215_2_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err[9] ), 
            .I2(GND_net), .I3(GND_net), .O(n319_adj_3828));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i215_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i280_2_lut (.I0(\Kp[4] ), .I1(\PID_CONTROLLER.err[9] ), 
            .I2(GND_net), .I3(GND_net), .O(n416_adj_3827));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i280_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i345_2_lut (.I0(\Kp[5] ), .I1(\PID_CONTROLLER.err[9] ), 
            .I2(GND_net), .I3(GND_net), .O(n513_adj_3826));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i345_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_24_i5_3_lut (.I0(\PID_CONTROLLER.result [4]), .I1(n70[4]), 
            .I2(n421), .I3(GND_net), .O(n467));   // verilog/motorControl.v(49[18] 51[12])
    defparam mux_24_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_12_i335_2_lut (.I0(\Kd[5] ), .I1(n57[4]), .I2(GND_net), 
            .I3(GND_net), .O(n498_adj_3825));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i335_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 state_23__I_0_inv_0_i18_1_lut (.I0(setpoint[17]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n58[17]));   // verilog/motorControl.v(39[14:30])
    defparam state_23__I_0_inv_0_i18_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i410_2_lut (.I0(\Kp[6] ), .I1(\PID_CONTROLLER.err[9] ), 
            .I2(GND_net), .I3(GND_net), .O(n610_adj_3823));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i410_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1_4_lut_adj_1403 (.I0(pwm_23__N_2957), .I1(n1), .I2(\PWMLimit[5] ), 
            .I3(n387), .O(n24209));   // verilog/motorControl.v(44[10:51])
    defparam i1_4_lut_adj_1403.LUT_INIT = 16'ha088;
    SB_LUT4 mult_10_i475_2_lut (.I0(\Kp[7] ), .I1(\PID_CONTROLLER.err[9] ), 
            .I2(GND_net), .I3(GND_net), .O(n707_adj_3822));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i475_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1_4_lut_adj_1404 (.I0(pwm_23__N_2957), .I1(n27212), .I2(\PWMLimit[6] ), 
            .I3(n387), .O(n24210));   // verilog/motorControl.v(44[10:51])
    defparam i1_4_lut_adj_1404.LUT_INIT = 16'ha088;
    SB_LUT4 state_23__I_0_inv_0_i19_1_lut (.I0(setpoint[18]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n58[18]));   // verilog/motorControl.v(39[14:30])
    defparam state_23__I_0_inv_0_i19_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mux_24_i8_3_lut (.I0(\PID_CONTROLLER.result [7]), .I1(n70[7]), 
            .I2(n421), .I3(GND_net), .O(n464));   // verilog/motorControl.v(49[18] 51[12])
    defparam mux_24_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_10_i505_2_lut (.I0(\Kp[7] ), .I1(\PID_CONTROLLER.err[31] ), 
            .I2(GND_net), .I3(GND_net), .O(n752_adj_3820));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i505_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i99_2_lut (.I0(\Kp[1] ), .I1(\PID_CONTROLLER.err[16] ), 
            .I2(GND_net), .I3(GND_net), .O(n146_adj_3819));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i99_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i36_2_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err[17] ), 
            .I2(GND_net), .I3(GND_net), .O(n53_adj_3818));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i36_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_24_i9_3_lut (.I0(\PID_CONTROLLER.result [8]), .I1(n70[8]), 
            .I2(n421), .I3(GND_net), .O(n463));   // verilog/motorControl.v(49[18] 51[12])
    defparam mux_24_i9_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_10_i164_2_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err[16] ), 
            .I2(GND_net), .I3(GND_net), .O(n243_adj_3817));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i164_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i229_2_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err[16] ), 
            .I2(GND_net), .I3(GND_net), .O(n340_adj_3816));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i229_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i294_2_lut (.I0(\Kp[4] ), .I1(\PID_CONTROLLER.err[16] ), 
            .I2(GND_net), .I3(GND_net), .O(n437_adj_3815));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i294_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i359_2_lut (.I0(\Kp[5] ), .I1(\PID_CONTROLLER.err[16] ), 
            .I2(GND_net), .I3(GND_net), .O(n534_adj_3814));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i359_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i424_2_lut (.I0(\Kp[6] ), .I1(\PID_CONTROLLER.err[16] ), 
            .I2(GND_net), .I3(GND_net), .O(n631_adj_3813));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i424_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_24_i10_3_lut (.I0(\PID_CONTROLLER.result [9]), .I1(n70[9]), 
            .I2(n421), .I3(GND_net), .O(n462));   // verilog/motorControl.v(49[18] 51[12])
    defparam mux_24_i10_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_10_i489_2_lut (.I0(\Kp[7] ), .I1(\PID_CONTROLLER.err[16] ), 
            .I2(GND_net), .I3(GND_net), .O(n728_adj_3812));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i489_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i115_2_lut (.I0(\Kp[1] ), .I1(\PID_CONTROLLER.err[31] ), 
            .I2(GND_net), .I3(GND_net), .O(n182_adj_3811));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i115_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i375_2_lut (.I0(\Kp[5] ), .I1(\PID_CONTROLLER.err[31] ), 
            .I2(GND_net), .I3(GND_net), .O(n558_adj_3807));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i375_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_24_i11_3_lut (.I0(\PID_CONTROLLER.result [10]), .I1(n70[10]), 
            .I2(n421), .I3(GND_net), .O(n461));   // verilog/motorControl.v(49[18] 51[12])
    defparam mux_24_i11_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_24_i12_3_lut (.I0(\PID_CONTROLLER.result [11]), .I1(n70[10]), 
            .I2(n421), .I3(GND_net), .O(n460));   // verilog/motorControl.v(49[18] 51[12])
    defparam mux_24_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_10_i180_2_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err[31] ), 
            .I2(GND_net), .I3(GND_net), .O(n276_adj_3810));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i180_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i245_2_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err[31] ), 
            .I2(GND_net), .I3(GND_net), .O(n370_adj_3809));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i245_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i20072_3_lut (.I0(\PID_CONTROLLER.err[31] ), .I1(n33546), .I2(n35990), 
            .I3(GND_net), .O(n16644[1]));   // verilog/motorControl.v(43[17:23])
    defparam i20072_3_lut.LUT_INIT = 16'h6c6c;
    SB_LUT4 mux_24_i13_3_lut (.I0(\PID_CONTROLLER.result [12]), .I1(n70[10]), 
            .I2(n421), .I3(GND_net), .O(n459));   // verilog/motorControl.v(49[18] 51[12])
    defparam mux_24_i13_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_10_i310_2_lut (.I0(\Kp[4] ), .I1(\PID_CONTROLLER.err[31] ), 
            .I2(GND_net), .I3(GND_net), .O(n464_adj_3808));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i310_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i442_2_lut (.I0(\Kp[6] ), .I1(\PID_CONTROLLER.err[31] ), 
            .I2(GND_net), .I3(GND_net), .O(n658_adj_3806));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i442_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_24_i14_3_lut (.I0(\PID_CONTROLLER.result [13]), .I1(n70[10]), 
            .I2(n421), .I3(GND_net), .O(n458));   // verilog/motorControl.v(49[18] 51[12])
    defparam mux_24_i14_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i5_4_lut_adj_1405 (.I0(n33546), .I1(n7_adj_3851), .I2(n8_adj_3852), 
            .I3(n8_adj_3853), .O(n41719));   // verilog/motorControl.v(43[17:23])
    defparam i5_4_lut_adj_1405.LUT_INIT = 16'h6996;
    SB_LUT4 mult_10_i97_2_lut (.I0(\Kp[1] ), .I1(\PID_CONTROLLER.err[15] ), 
            .I2(GND_net), .I3(GND_net), .O(n143_adj_3805));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i97_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_24_i15_3_lut (.I0(\PID_CONTROLLER.result [14]), .I1(n70[10]), 
            .I2(n421), .I3(GND_net), .O(n457));   // verilog/motorControl.v(49[18] 51[12])
    defparam mux_24_i15_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_10_i34_2_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err[16] ), 
            .I2(GND_net), .I3(GND_net), .O(n50_adj_3804));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i34_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i162_2_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err[15] ), 
            .I2(GND_net), .I3(GND_net), .O(n240_adj_3803));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i162_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i227_2_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err[15] ), 
            .I2(GND_net), .I3(GND_net), .O(n337_adj_3802));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i227_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i292_2_lut (.I0(\Kp[4] ), .I1(\PID_CONTROLLER.err[15] ), 
            .I2(GND_net), .I3(GND_net), .O(n434_adj_3801));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i292_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i357_2_lut (.I0(\Kp[5] ), .I1(\PID_CONTROLLER.err[15] ), 
            .I2(GND_net), .I3(GND_net), .O(n531_adj_3800));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i357_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_24_i16_3_lut (.I0(\PID_CONTROLLER.result [15]), .I1(n70[10]), 
            .I2(n421), .I3(GND_net), .O(n456));   // verilog/motorControl.v(49[18] 51[12])
    defparam mux_24_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_10_i422_2_lut (.I0(\Kp[6] ), .I1(\PID_CONTROLLER.err[15] ), 
            .I2(GND_net), .I3(GND_net), .O(n628_adj_3799));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i422_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i487_2_lut (.I0(\Kp[7] ), .I1(\PID_CONTROLLER.err[15] ), 
            .I2(GND_net), .I3(GND_net), .O(n725_adj_3798));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i487_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i113_2_lut (.I0(\Kp[1] ), .I1(\PID_CONTROLLER.err[23] ), 
            .I2(GND_net), .I3(GND_net), .O(n167_adj_3797));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i113_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i50_2_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err[31] ), 
            .I2(GND_net), .I3(GND_net), .O(n86_adj_3796));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i50_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i178_2_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err[23] ), 
            .I2(GND_net), .I3(GND_net), .O(n264_adj_3795));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i178_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i243_2_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err[23] ), 
            .I2(GND_net), .I3(GND_net), .O(n361_adj_3794));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i243_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_24_i17_3_lut (.I0(\PID_CONTROLLER.result [16]), .I1(n70[10]), 
            .I2(n421), .I3(GND_net), .O(n455));   // verilog/motorControl.v(49[18] 51[12])
    defparam mux_24_i17_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_10_i308_2_lut (.I0(\Kp[4] ), .I1(\PID_CONTROLLER.err[23] ), 
            .I2(GND_net), .I3(GND_net), .O(n458_adj_3793));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i308_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i373_2_lut (.I0(\Kp[5] ), .I1(\PID_CONTROLLER.err[23] ), 
            .I2(GND_net), .I3(GND_net), .O(n555_adj_3792));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i373_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i400_2_lut (.I0(\Kd[6] ), .I1(n57[4]), .I2(GND_net), 
            .I3(GND_net), .O(n595_adj_3791));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i400_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i438_2_lut (.I0(\Kp[6] ), .I1(\PID_CONTROLLER.err[23] ), 
            .I2(GND_net), .I3(GND_net), .O(n652_adj_3790));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i438_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i503_2_lut (.I0(\Kp[7] ), .I1(\PID_CONTROLLER.err[23] ), 
            .I2(GND_net), .I3(GND_net), .O(n749_adj_3789));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i503_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i95_2_lut (.I0(\Kp[1] ), .I1(\PID_CONTROLLER.err[14] ), 
            .I2(GND_net), .I3(GND_net), .O(n140_adj_3788));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i95_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i32_2_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err[15] ), 
            .I2(GND_net), .I3(GND_net), .O(n47_adj_3787));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i32_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i160_2_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err[14] ), 
            .I2(GND_net), .I3(GND_net), .O(n237_adj_3786));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i160_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i225_2_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err[14] ), 
            .I2(GND_net), .I3(GND_net), .O(n334_adj_3785));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i225_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i290_2_lut (.I0(\Kp[4] ), .I1(\PID_CONTROLLER.err[14] ), 
            .I2(GND_net), .I3(GND_net), .O(n431_adj_3784));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i290_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1_4_lut_adj_1406 (.I0(pwm_23__N_2957), .I1(n44151), .I2(\PWMLimit[9] ), 
            .I3(n387), .O(n39108));
    defparam i1_4_lut_adj_1406.LUT_INIT = 16'ha088;
    SB_LUT4 mult_10_i355_2_lut (.I0(\Kp[5] ), .I1(\PID_CONTROLLER.err[14] ), 
            .I2(GND_net), .I3(GND_net), .O(n528_adj_3783));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i355_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i420_2_lut (.I0(\Kp[6] ), .I1(\PID_CONTROLLER.err[14] ), 
            .I2(GND_net), .I3(GND_net), .O(n625_adj_3782));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i420_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i485_2_lut (.I0(\Kp[7] ), .I1(\PID_CONTROLLER.err[14] ), 
            .I2(GND_net), .I3(GND_net), .O(n722_adj_3781));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i485_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_14_i51_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral [0]), 
            .I2(GND_net), .I3(GND_net), .O(n74_adj_3780));   // verilog/motorControl.v(43[48:59])
    defparam mult_14_i51_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_14_i4_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral [1]), 
            .I2(GND_net), .I3(GND_net), .O(n5_adj_3779));   // verilog/motorControl.v(43[48:59])
    defparam mult_14_i4_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_14_i100_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral [0]), 
            .I2(GND_net), .I3(GND_net), .O(n147_adj_3778));   // verilog/motorControl.v(43[48:59])
    defparam mult_14_i100_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_14_i149_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral [0]), 
            .I2(GND_net), .I3(GND_net), .O(n220_adj_3777));   // verilog/motorControl.v(43[48:59])
    defparam mult_14_i149_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_14_i198_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral [0]), 
            .I2(GND_net), .I3(GND_net), .O(n293));   // verilog/motorControl.v(43[48:59])
    defparam mult_14_i198_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_14_i247_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral [0]), 
            .I2(GND_net), .I3(GND_net), .O(n366));   // verilog/motorControl.v(43[48:59])
    defparam mult_14_i247_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i20344_2_lut_3_lut (.I0(\Kd[0] ), .I1(\Kd[1] ), .I2(\Kd[2] ), 
            .I3(GND_net), .O(n33872));   // verilog/motorControl.v(43[26:45])
    defparam i20344_2_lut_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 mult_14_i296_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral [0]), 
            .I2(GND_net), .I3(GND_net), .O(n439));   // verilog/motorControl.v(43[48:59])
    defparam mult_14_i296_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_14_i345_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral [0]), 
            .I2(GND_net), .I3(GND_net), .O(n512));   // verilog/motorControl.v(43[48:59])
    defparam mult_14_i345_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i20376_2_lut_3_lut (.I0(\Kd[0] ), .I1(\Kd[1] ), .I2(n57[25]), 
            .I3(GND_net), .O(n10111[0]));   // verilog/motorControl.v(43[26:45])
    defparam i20376_2_lut_3_lut.LUT_INIT = 16'h6060;
    SB_LUT4 mult_14_i53_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral [1]), 
            .I2(GND_net), .I3(GND_net), .O(n77));   // verilog/motorControl.v(43[48:59])
    defparam mult_14_i53_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_14_i6_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral [2]), 
            .I2(GND_net), .I3(GND_net), .O(n8_adj_3771));   // verilog/motorControl.v(43[48:59])
    defparam mult_14_i6_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_14_i102_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral [1]), 
            .I2(GND_net), .I3(GND_net), .O(n150_adj_3770));   // verilog/motorControl.v(43[48:59])
    defparam mult_14_i102_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_14_i151_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral [1]), 
            .I2(GND_net), .I3(GND_net), .O(n223_adj_3768));   // verilog/motorControl.v(43[48:59])
    defparam mult_14_i151_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_14_i200_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral [1]), 
            .I2(GND_net), .I3(GND_net), .O(n296_adj_3766));   // verilog/motorControl.v(43[48:59])
    defparam mult_14_i200_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_14_i249_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral [1]), 
            .I2(GND_net), .I3(GND_net), .O(n369));   // verilog/motorControl.v(43[48:59])
    defparam mult_14_i249_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_14_i298_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral [1]), 
            .I2(GND_net), .I3(GND_net), .O(n442));   // verilog/motorControl.v(43[48:59])
    defparam mult_14_i298_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_14_i347_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral [1]), 
            .I2(GND_net), .I3(GND_net), .O(n515));   // verilog/motorControl.v(43[48:59])
    defparam mult_14_i347_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1_3_lut_4_lut (.I0(n370), .I1(n4_adj_3856), .I2(n33872), 
            .I3(n57[25]), .O(n7_adj_3857));   // verilog/motorControl.v(43[26:45])
    defparam i1_3_lut_4_lut.LUT_INIT = 16'h6966;
    SB_LUT4 mult_14_i55_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral [2]), 
            .I2(GND_net), .I3(GND_net), .O(n80));   // verilog/motorControl.v(43[48:59])
    defparam mult_14_i55_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_14_i8_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral [3]), 
            .I2(GND_net), .I3(GND_net), .O(n11_adj_3760));   // verilog/motorControl.v(43[48:59])
    defparam mult_14_i8_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_14_i104_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral [2]), 
            .I2(GND_net), .I3(GND_net), .O(n153_adj_3759));   // verilog/motorControl.v(43[48:59])
    defparam mult_14_i104_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_22_i19_2_lut (.I0(\PID_CONTROLLER.result [9]), .I1(n70[9]), 
            .I2(GND_net), .I3(GND_net), .O(n19_adj_3858));   // verilog/motorControl.v(47[21:37])
    defparam LessThan_22_i19_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_14_i153_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral [2]), 
            .I2(GND_net), .I3(GND_net), .O(n226_adj_3757));   // verilog/motorControl.v(43[48:59])
    defparam mult_14_i153_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_22_i15_2_lut (.I0(\PID_CONTROLLER.result [7]), .I1(n70[7]), 
            .I2(GND_net), .I3(GND_net), .O(n15_adj_3859));   // verilog/motorControl.v(47[21:37])
    defparam LessThan_22_i15_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_14_i202_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral [2]), 
            .I2(GND_net), .I3(GND_net), .O(n299_adj_3755));   // verilog/motorControl.v(43[48:59])
    defparam mult_14_i202_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_22_i17_2_lut (.I0(\PID_CONTROLLER.result [8]), .I1(n70[8]), 
            .I2(GND_net), .I3(GND_net), .O(n17_adj_3860));   // verilog/motorControl.v(47[21:37])
    defparam LessThan_22_i17_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_14_i251_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral [2]), 
            .I2(GND_net), .I3(GND_net), .O(n372));   // verilog/motorControl.v(43[48:59])
    defparam mult_14_i251_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_22_i7_2_lut (.I0(\PID_CONTROLLER.result [3]), .I1(n70[3]), 
            .I2(GND_net), .I3(GND_net), .O(n7_adj_3861));   // verilog/motorControl.v(47[21:37])
    defparam LessThan_22_i7_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_22_i9_2_lut (.I0(\PID_CONTROLLER.result [4]), .I1(n70[4]), 
            .I2(GND_net), .I3(GND_net), .O(n9_adj_3862));   // verilog/motorControl.v(47[21:37])
    defparam LessThan_22_i9_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_14_i300_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral [2]), 
            .I2(GND_net), .I3(GND_net), .O(n445));   // verilog/motorControl.v(43[48:59])
    defparam mult_14_i300_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_14_i349_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral [2]), 
            .I2(GND_net), .I3(GND_net), .O(n518));   // verilog/motorControl.v(43[48:59])
    defparam mult_14_i349_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i4_2_lut (.I0(\PID_CONTROLLER.result [14]), .I1(\PID_CONTROLLER.result [16]), 
            .I2(GND_net), .I3(GND_net), .O(n18_adj_3863));
    defparam i4_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i10_4_lut (.I0(\PID_CONTROLLER.result [11]), .I1(\PID_CONTROLLER.result [27]), 
            .I2(\PID_CONTROLLER.result [15]), .I3(\PID_CONTROLLER.result [10]), 
            .O(n24_adj_3864));
    defparam i10_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 LessThan_22_i5_2_lut (.I0(\PID_CONTROLLER.result [2]), .I1(n70[2]), 
            .I2(GND_net), .I3(GND_net), .O(n5_adj_3865));   // verilog/motorControl.v(47[21:37])
    defparam LessThan_22_i5_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_12_i97_2_lut (.I0(\Kd[1] ), .I1(n57[15]), .I2(GND_net), 
            .I3(GND_net), .O(n143_adj_3750));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i97_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i34_2_lut (.I0(\Kd[0] ), .I1(n57[16]), .I2(GND_net), 
            .I3(GND_net), .O(n50_adj_3749));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i34_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i29019_4_lut (.I0(n11), .I1(n9_adj_3862), .I2(n7_adj_3861), 
            .I3(n5_adj_3865), .O(n44539));
    defparam i29019_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 mult_12_i162_2_lut (.I0(\Kd[2] ), .I1(n57[15]), .I2(GND_net), 
            .I3(GND_net), .O(n240_adj_3748));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i162_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i227_2_lut (.I0(\Kd[3] ), .I1(n57[15]), .I2(GND_net), 
            .I3(GND_net), .O(n337));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i227_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_22_i4_4_lut (.I0(n70[0]), .I1(n70[1]), .I2(\PID_CONTROLLER.result [1]), 
            .I3(\PID_CONTROLLER.result [0]), .O(n4_adj_3867));   // verilog/motorControl.v(47[21:37])
    defparam LessThan_22_i4_4_lut.LUT_INIT = 16'h0c8e;
    SB_LUT4 i30135_3_lut (.I0(n4_adj_3867), .I1(n415), .I2(n11), .I3(GND_net), 
            .O(n45656));   // verilog/motorControl.v(47[21:37])
    defparam i30135_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i30136_3_lut (.I0(n45656), .I1(n414), .I2(n13), .I3(GND_net), 
            .O(n45657));   // verilog/motorControl.v(47[21:37])
    defparam i30136_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_3_lut (.I0(\PID_CONTROLLER.result [27]), .I1(\PID_CONTROLLER.result [14]), 
            .I2(\PID_CONTROLLER.result [15]), .I3(GND_net), .O(n10_adj_3869));   // verilog/motorControl.v(38[14] 59[8])
    defparam i1_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 i8_4_lut (.I0(\PID_CONTROLLER.result [30]), .I1(n49_adj_3870), 
            .I2(\PID_CONTROLLER.result [12]), .I3(\PID_CONTROLLER.result [28]), 
            .O(n22_adj_3871));
    defparam i8_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i3_3_lut (.I0(\PID_CONTROLLER.result [16]), .I1(\PID_CONTROLLER.result [10]), 
            .I2(\PID_CONTROLLER.result [11]), .I3(GND_net), .O(n12_adj_3872));   // verilog/motorControl.v(38[14] 59[8])
    defparam i3_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 i7_4_lut (.I0(n70[10]), .I1(\PID_CONTROLLER.result [12]), .I2(\PID_CONTROLLER.result [26]), 
            .I3(n10_adj_3869), .O(n16_adj_3873));   // verilog/motorControl.v(38[14] 59[8])
    defparam i7_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i12_4_lut (.I0(\PID_CONTROLLER.result [29]), .I1(n24_adj_3864), 
            .I2(n18_adj_3863), .I3(n62_adj_3874), .O(n26_adj_3875));
    defparam i12_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i29320_4_lut (.I0(n40200), .I1(n16_adj_3873), .I2(n12_adj_3872), 
            .I3(n40124), .O(n44166));   // verilog/motorControl.v(38[14] 59[8])
    defparam i29320_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i11_3_lut (.I0(\PID_CONTROLLER.result [26]), .I1(n22_adj_3871), 
            .I2(n70[10]), .I3(GND_net), .O(n25_adj_3876));
    defparam i11_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 LessThan_22_i6_3_lut (.I0(n70[2]), .I1(n70[3]), .I2(n7_adj_3861), 
            .I3(GND_net), .O(n6_adj_3877));   // verilog/motorControl.v(47[21:37])
    defparam LessThan_22_i6_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i30287_3_lut (.I0(n6_adj_3877), .I1(n70[4]), .I2(n9_adj_3862), 
            .I3(GND_net), .O(n45808));   // verilog/motorControl.v(47[21:37])
    defparam i30287_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i30288_3_lut (.I0(n45808), .I1(n70[8]), .I2(n17_adj_3860), 
            .I3(GND_net), .O(n45809));   // verilog/motorControl.v(47[21:37])
    defparam i30288_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i29010_4_lut (.I0(n17_adj_3860), .I1(n15_adj_3859), .I2(n13), 
            .I3(n44539), .O(n44530));
    defparam i29010_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i29577_3_lut (.I0(n45657), .I1(n70[7]), .I2(n15_adj_3859), 
            .I3(GND_net), .O(n45098));   // verilog/motorControl.v(47[21:37])
    defparam i29577_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_14_i193_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral [9]), 
            .I2(GND_net), .I3(GND_net), .O(n253));   // verilog/motorControl.v(43[48:59])
    defparam mult_14_i193_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i30106_3_lut (.I0(n45809), .I1(n70[9]), .I2(n19_adj_3858), 
            .I3(GND_net), .O(n45627));   // verilog/motorControl.v(47[21:37])
    defparam i30106_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i28_4_lut (.I0(n25_adj_3876), .I1(n44166), .I2(\PID_CONTROLLER.result [13]), 
            .I3(n26_adj_3875), .O(n20_adj_3878));   // verilog/motorControl.v(38[14] 59[8])
    defparam i28_4_lut.LUT_INIT = 16'hc0c5;
    SB_LUT4 mult_10_i2_2_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err[0] ), 
            .I2(GND_net), .I3(GND_net), .O(n61[0]));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i2_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i30191_4_lut (.I0(n45627), .I1(n45098), .I2(n19_adj_3858), 
            .I3(n44530), .O(n45712));   // verilog/motorControl.v(47[21:37])
    defparam i30191_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 mult_14_i2_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral [0]), 
            .I2(GND_net), .I3(GND_net), .O(n282[0]));   // verilog/motorControl.v(43[48:59])
    defparam mult_14_i2_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 state_23__I_0_inv_0_i13_1_lut (.I0(setpoint[12]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n58[12]));   // verilog/motorControl.v(39[14:30])
    defparam state_23__I_0_inv_0_i13_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i29974_4_lut (.I0(n45712), .I1(\PID_CONTROLLER.result [31]), 
            .I2(n70[10]), .I3(n20_adj_3878), .O(n421));   // verilog/motorControl.v(47[21:37])
    defparam i29974_4_lut.LUT_INIT = 16'h8ecc;
    SB_LUT4 state_23__I_0_inv_0_i14_1_lut (.I0(setpoint[13]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n58[13]));   // verilog/motorControl.v(39[14:30])
    defparam state_23__I_0_inv_0_i14_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 \PID_CONTROLLER.result_31__I_0_i7_2_lut  (.I0(\deadband[3] ), 
            .I1(\PID_CONTROLLER.result [3]), .I2(GND_net), .I3(GND_net), 
            .O(n7_adj_3879));   // verilog/motorControl.v(44[10:27])
    defparam \PID_CONTROLLER.result_31__I_0_i7_2_lut .LUT_INIT = 16'h6666;
    SB_LUT4 \PID_CONTROLLER.result_31__I_0_i15_2_lut  (.I0(\deadband[7] ), 
            .I1(\PID_CONTROLLER.result [7]), .I2(GND_net), .I3(GND_net), 
            .O(n15_adj_3880));   // verilog/motorControl.v(44[10:27])
    defparam \PID_CONTROLLER.result_31__I_0_i15_2_lut .LUT_INIT = 16'h6666;
    SB_LUT4 \PID_CONTROLLER.result_31__I_0_i9_2_lut  (.I0(\deadband[4] ), 
            .I1(\PID_CONTROLLER.result [4]), .I2(GND_net), .I3(GND_net), 
            .O(n9_adj_3881));   // verilog/motorControl.v(44[10:27])
    defparam \PID_CONTROLLER.result_31__I_0_i9_2_lut .LUT_INIT = 16'h6666;
    SB_LUT4 \PID_CONTROLLER.result_31__I_0_i17_2_lut  (.I0(\deadband[8] ), 
            .I1(\PID_CONTROLLER.result [8]), .I2(GND_net), .I3(GND_net), 
            .O(n17_adj_3882));   // verilog/motorControl.v(44[10:27])
    defparam \PID_CONTROLLER.result_31__I_0_i17_2_lut .LUT_INIT = 16'h6666;
    SB_LUT4 state_23__I_0_inv_0_i15_1_lut (.I0(setpoint[14]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n58[14]));   // verilog/motorControl.v(39[14:30])
    defparam state_23__I_0_inv_0_i15_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i29784_4_lut (.I0(\deadband[9] ), .I1(n17_adj_3882), .I2(\PID_CONTROLLER.result [9]), 
            .I3(n9_adj_3881), .O(n45305));
    defparam i29784_4_lut.LUT_INIT = 16'hffde;
    SB_LUT4 i29778_4_lut (.I0(\deadband[9] ), .I1(\PID_CONTROLLER.result [10]), 
            .I2(\PID_CONTROLLER.result [11]), .I3(n45305), .O(n45299));
    defparam i29778_4_lut.LUT_INIT = 16'h7eff;
    SB_LUT4 i29792_3_lut (.I0(n15_adj_3880), .I1(n13_adj_10), .I2(n11_adj_11), 
            .I3(GND_net), .O(n45313));
    defparam i29792_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i29762_4_lut (.I0(\deadband[9] ), .I1(\PID_CONTROLLER.result [13]), 
            .I2(\PID_CONTROLLER.result [14]), .I3(n45313), .O(n45283));
    defparam i29762_4_lut.LUT_INIT = 16'h7eff;
    SB_LUT4 i29742_4_lut (.I0(\PID_CONTROLLER.result [17]), .I1(\PID_CONTROLLER.result [16]), 
            .I2(\deadband[9] ), .I3(n15_adj_3880), .O(n45263));
    defparam i29742_4_lut.LUT_INIT = 16'hff7e;
    SB_LUT4 \PID_CONTROLLER.result_31__I_0_i30_4_lut  (.I0(\PID_CONTROLLER.result [7]), 
            .I1(\PID_CONTROLLER.result [17]), .I2(\deadband[9] ), .I3(\PID_CONTROLLER.result [16]), 
            .O(n30_adj_3885));   // verilog/motorControl.v(44[10:27])
    defparam \PID_CONTROLLER.result_31__I_0_i30_4_lut .LUT_INIT = 16'h8f0e;
    SB_LUT4 i29804_4_lut (.I0(n9_adj_3881), .I1(n7_adj_3879), .I2(\deadband[2] ), 
            .I3(\PID_CONTROLLER.result [2]), .O(n45325));
    defparam i29804_4_lut.LUT_INIT = 16'heffe;
    SB_LUT4 i30061_4_lut (.I0(n15_adj_3880), .I1(n13_adj_10), .I2(n11_adj_11), 
            .I3(n45325), .O(n45582));
    defparam i30061_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i29788_4_lut (.I0(\deadband[9] ), .I1(n17_adj_3882), .I2(\PID_CONTROLLER.result [9]), 
            .I3(n45582), .O(n45309));
    defparam i29788_4_lut.LUT_INIT = 16'hdeff;
    SB_LUT4 state_23__I_0_inv_0_i20_1_lut (.I0(setpoint[19]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n58[19]));   // verilog/motorControl.v(39[14:30])
    defparam state_23__I_0_inv_0_i20_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i30307_4_lut (.I0(\deadband[9] ), .I1(\PID_CONTROLLER.result [10]), 
            .I2(\PID_CONTROLLER.result [11]), .I3(n45309), .O(n45828));
    defparam i30307_4_lut.LUT_INIT = 16'hff7e;
    SB_LUT4 i29155_4_lut (.I0(\deadband[9] ), .I1(\PID_CONTROLLER.result [12]), 
            .I2(\PID_CONTROLLER.result [13]), .I3(n45828), .O(n44676));
    defparam i29155_4_lut.LUT_INIT = 16'h5adb;
    SB_LUT4 i30045_4_lut (.I0(\deadband[9] ), .I1(\PID_CONTROLLER.result [14]), 
            .I2(\PID_CONTROLLER.result [15]), .I3(n44676), .O(n45566));
    defparam i30045_4_lut.LUT_INIT = 16'hff7e;
    SB_LUT4 i30467_4_lut (.I0(\PID_CONTROLLER.result [17]), .I1(\PID_CONTROLLER.result [16]), 
            .I2(\deadband[9] ), .I3(n45566), .O(n45988));
    defparam i30467_4_lut.LUT_INIT = 16'hff7e;
    SB_LUT4 i30619_4_lut (.I0(\PID_CONTROLLER.result [19]), .I1(\PID_CONTROLLER.result [18]), 
            .I2(\deadband[9] ), .I3(n45988), .O(n46140));
    defparam i30619_4_lut.LUT_INIT = 16'hff7e;
    SB_LUT4 state_23__I_0_inv_0_i21_1_lut (.I0(setpoint[20]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n58[20]));   // verilog/motorControl.v(39[14:30])
    defparam state_23__I_0_inv_0_i21_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 state_23__I_0_inv_0_i22_1_lut (.I0(setpoint[21]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n58[21]));   // verilog/motorControl.v(39[14:30])
    defparam state_23__I_0_inv_0_i22_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i30149_3_lut (.I0(n6_adj_3886), .I1(\PID_CONTROLLER.result [10]), 
            .I2(\deadband[9] ), .I3(GND_net), .O(n45670));   // verilog/motorControl.v(44[10:27])
    defparam i30149_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i29708_4_lut (.I0(\PID_CONTROLLER.result [22]), .I1(\PID_CONTROLLER.result [21]), 
            .I2(\deadband[9] ), .I3(\PID_CONTROLLER.result [9]), .O(n45229));
    defparam i29708_4_lut.LUT_INIT = 16'h7ffe;
    SB_LUT4 \PID_CONTROLLER.result_31__I_0_i24_4_lut  (.I0(\PID_CONTROLLER.result [9]), 
            .I1(\PID_CONTROLLER.result [22]), .I2(\deadband[9] ), .I3(\PID_CONTROLLER.result [21]), 
            .O(n24_adj_3887));   // verilog/motorControl.v(44[10:27])
    defparam \PID_CONTROLLER.result_31__I_0_i24_4_lut .LUT_INIT = 16'h8f0e;
    SB_LUT4 i29111_4_lut (.I0(\PID_CONTROLLER.result [21]), .I1(\PID_CONTROLLER.result [12]), 
            .I2(\deadband[9] ), .I3(n45299), .O(n44632));
    defparam i29111_4_lut.LUT_INIT = 16'h5adb;
    SB_LUT4 i17_rep_263_2_lut (.I0(\PID_CONTROLLER.result [22]), .I1(\deadband[9] ), 
            .I2(GND_net), .I3(GND_net), .O(n47290));   // verilog/TinyFPGA_B.v(65[22:30])
    defparam i17_rep_263_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i30403_3_lut (.I0(n24_adj_3887), .I1(n8_adj_3888), .I2(n45229), 
            .I3(GND_net), .O(n45924));   // verilog/motorControl.v(44[10:27])
    defparam i30403_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i29555_4_lut (.I0(n45670), .I1(\PID_CONTROLLER.result [12]), 
            .I2(\deadband[9] ), .I3(\PID_CONTROLLER.result [11]), .O(n45076));   // verilog/motorControl.v(44[10:27])
    defparam i29555_4_lut.LUT_INIT = 16'h8f0e;
    SB_LUT4 \PID_CONTROLLER.result_31__I_0_i4_4_lut  (.I0(\deadband[0] ), 
            .I1(\PID_CONTROLLER.result [1]), .I2(\deadband[1] ), .I3(\PID_CONTROLLER.result [0]), 
            .O(n4_adj_3889));   // verilog/motorControl.v(44[10:27])
    defparam \PID_CONTROLLER.result_31__I_0_i4_4_lut .LUT_INIT = 16'h4d0c;
    SB_LUT4 i30147_3_lut (.I0(n4_adj_3889), .I1(\PID_CONTROLLER.result [13]), 
            .I2(\deadband[9] ), .I3(GND_net), .O(n45668));   // verilog/motorControl.v(44[10:27])
    defparam i30147_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i29143_4_lut (.I0(\deadband[9] ), .I1(\PID_CONTROLLER.result [15]), 
            .I2(\PID_CONTROLLER.result [16]), .I3(n45283), .O(n44664));
    defparam i29143_4_lut.LUT_INIT = 16'h5adb;
    SB_LUT4 i19_rep_240_2_lut (.I0(\PID_CONTROLLER.result [17]), .I1(\deadband[9] ), 
            .I2(GND_net), .I3(GND_net), .O(n47267));   // verilog/TinyFPGA_B.v(65[22:30])
    defparam i19_rep_240_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_12_i465_2_lut (.I0(\Kd[7] ), .I1(n57[4]), .I2(GND_net), 
            .I3(GND_net), .O(n692_adj_3743));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i465_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i213_2_lut (.I0(\Kd[3] ), .I1(n57[8]), .I2(GND_net), 
            .I3(GND_net), .O(n316_adj_3742));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i213_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i30513_3_lut (.I0(n30_adj_3885), .I1(n10_adj_3890), .I2(n45263), 
            .I3(GND_net), .O(n46034));   // verilog/motorControl.v(44[10:27])
    defparam i30513_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i29557_4_lut (.I0(n45668), .I1(\PID_CONTROLLER.result [15]), 
            .I2(\deadband[9] ), .I3(\PID_CONTROLLER.result [14]), .O(n45078));   // verilog/motorControl.v(44[10:27])
    defparam i29557_4_lut.LUT_INIT = 16'h8f0e;
    SB_LUT4 i30641_4_lut (.I0(n45078), .I1(n46034), .I2(n47267), .I3(n44664), 
            .O(n46162));   // verilog/motorControl.v(44[10:27])
    defparam i30641_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i30642_3_lut (.I0(n46162), .I1(\PID_CONTROLLER.result [18]), 
            .I2(\deadband[9] ), .I3(GND_net), .O(n46163));   // verilog/motorControl.v(44[10:27])
    defparam i30642_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 mult_12_i292_2_lut (.I0(\Kd[4] ), .I1(n57[15]), .I2(GND_net), 
            .I3(GND_net), .O(n434));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i292_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i29117_4_lut (.I0(\PID_CONTROLLER.result [21]), .I1(\PID_CONTROLLER.result [20]), 
            .I2(\deadband[9] ), .I3(n46140), .O(n44638));
    defparam i29117_4_lut.LUT_INIT = 16'h5adb;
    SB_LUT4 i30596_4_lut (.I0(n45076), .I1(n45924), .I2(n47290), .I3(n44632), 
            .O(n46117));   // verilog/motorControl.v(44[10:27])
    defparam i30596_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 mult_12_i278_2_lut (.I0(\Kd[4] ), .I1(n57[8]), .I2(GND_net), 
            .I3(GND_net), .O(n413_adj_3740));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i278_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 state_23__I_0_inv_0_i23_1_lut (.I0(setpoint[22]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n58[22]));   // verilog/motorControl.v(39[14:30])
    defparam state_23__I_0_inv_0_i23_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i29563_4_lut (.I0(n46163), .I1(\PID_CONTROLLER.result [20]), 
            .I2(\deadband[9] ), .I3(\PID_CONTROLLER.result [19]), .O(n45084));   // verilog/motorControl.v(44[10:27])
    defparam i29563_4_lut.LUT_INIT = 16'h8f0e;
    SB_LUT4 i30637_4_lut (.I0(n45084), .I1(n46117), .I2(n47290), .I3(n44638), 
            .O(n46158));   // verilog/motorControl.v(44[10:27])
    defparam i30637_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i30603_4_lut (.I0(n46158), .I1(\PID_CONTROLLER.result [24]), 
            .I2(\deadband[9] ), .I3(\PID_CONTROLLER.result [23]), .O(n50_adj_3891));   // verilog/motorControl.v(44[10:27])
    defparam i30603_4_lut.LUT_INIT = 16'h8f0e;
    SB_LUT4 i24_4_lut (.I0(GATES_5__N_3048[4]), .I1(GATES_5__N_3048[5]), 
            .I2(n17_adj_3456), .I3(n878), .O(GATES_5__N_2788[5]));   // verilog/motorControl.v(86[14] 109[8])
    defparam i24_4_lut.LUT_INIT = 16'hac0c;
    SB_LUT4 i2_4_lut (.I0(hall1), .I1(GATES_5__N_3048[5]), .I2(hall2), 
            .I3(hall3), .O(GATES_5__N_3048[4]));   // verilog/motorControl.v(70[16] 85[10])
    defparam i2_4_lut.LUT_INIT = 16'h1050;
    SB_LUT4 GATES_5__I_0_i5_4_lut (.I0(n878), .I1(GATES_5__N_3048[4]), .I2(n17_adj_3456), 
            .I3(GATES_5__N_3048[5]), .O(GATES_5__N_2788[4]));   // verilog/motorControl.v(86[14] 109[8])
    defparam GATES_5__I_0_i5_4_lut.LUT_INIT = 16'hac0c;
    SB_LUT4 i3_4_lut (.I0(pwm_count[8]), .I1(n865), .I2(n868), .I3(n16), 
            .O(n19_adj_3893));
    defparam i3_4_lut.LUT_INIT = 16'h0223;
    SB_LUT4 i26666_3_lut (.I0(n866), .I1(n21), .I2(n853), .I3(GND_net), 
            .O(n42185));
    defparam i26666_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i26662_4_lut (.I0(n862), .I1(n864), .I2(n859), .I3(n861), 
            .O(n42181));
    defparam i26662_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i26664_4_lut (.I0(n856), .I1(n867), .I2(n863), .I3(n860), 
            .O(n42183));
    defparam i26664_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i13_4_lut_adj_1407 (.I0(n42185), .I1(n19_adj_3893), .I2(n855), 
            .I3(n857), .O(n29_adj_3894));
    defparam i13_4_lut_adj_1407.LUT_INIT = 16'h0004;
    SB_LUT4 i2_4_lut_adj_1408 (.I0(n29_adj_3894), .I1(hall3), .I2(n42183), 
            .I3(n42181), .O(n6_adj_3895));
    defparam i2_4_lut_adj_1408.LUT_INIT = 16'h333b;
    SB_LUT4 GATES_5__I_0_i4_4_lut (.I0(n5_adj_3441), .I1(GATES_5__N_3048[3]), 
            .I2(n17_adj_3456), .I3(n6_adj_3895), .O(GATES_5__N_2788[3]));   // verilog/motorControl.v(86[14] 109[8])
    defparam GATES_5__I_0_i4_4_lut.LUT_INIT = 16'h0c5c;
    SB_LUT4 i2_3_lut (.I0(hall2), .I1(GATES_5__N_3048[5]), .I2(hall3), 
            .I3(GND_net), .O(GATES_5__N_3048[3]));   // verilog/motorControl.v(70[16] 85[10])
    defparam i2_3_lut.LUT_INIT = 16'h0202;
    SB_LUT4 GATES_5__I_0_i3_4_lut (.I0(n44119), .I1(hall2), .I2(n17_adj_3456), 
            .I3(hall3), .O(GATES_5__N_2788[2]));   // verilog/motorControl.v(86[14] 109[8])
    defparam GATES_5__I_0_i3_4_lut.LUT_INIT = 16'ha3a0;
    SB_LUT4 mult_14_i57_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral [3]), 
            .I2(GND_net), .I3(GND_net), .O(n83));   // verilog/motorControl.v(43[48:59])
    defparam mult_14_i57_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_14_i10_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral [4]), 
            .I2(GND_net), .I3(GND_net), .O(n14_adj_3738));   // verilog/motorControl.v(43[48:59])
    defparam mult_14_i10_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 state_23__I_0_inv_0_i24_1_lut (.I0(setpoint[23]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n58[23]));   // verilog/motorControl.v(39[14:30])
    defparam state_23__I_0_inv_0_i24_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_14_i106_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral [3]), 
            .I2(GND_net), .I3(GND_net), .O(n156_adj_3735));   // verilog/motorControl.v(43[48:59])
    defparam mult_14_i106_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_14_i155_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral [3]), 
            .I2(GND_net), .I3(GND_net), .O(n229_adj_3733));   // verilog/motorControl.v(43[48:59])
    defparam mult_14_i155_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_14_i204_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral [3]), 
            .I2(GND_net), .I3(GND_net), .O(n302));   // verilog/motorControl.v(43[48:59])
    defparam mult_14_i204_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_14_i253_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral [3]), 
            .I2(GND_net), .I3(GND_net), .O(n375));   // verilog/motorControl.v(43[48:59])
    defparam mult_14_i253_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i343_2_lut (.I0(\Kd[5] ), .I1(n57[8]), .I2(GND_net), 
            .I3(GND_net), .O(n510_adj_3731));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i343_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_14_i302_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral [3]), 
            .I2(GND_net), .I3(GND_net), .O(n448));   // verilog/motorControl.v(43[48:59])
    defparam mult_14_i302_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 pwm_23__I_819_i17_2_lut (.I0(\PID_CONTROLLER.result [8]), .I1(pwm_23__N_2960[8]), 
            .I2(GND_net), .I3(GND_net), .O(n17_adj_3896));   // verilog/motorControl.v(44[31:51])
    defparam pwm_23__I_819_i17_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 pwm_23__I_819_i7_2_lut (.I0(\PID_CONTROLLER.result [3]), .I1(pwm_23__N_2960[3]), 
            .I2(GND_net), .I3(GND_net), .O(n7_adj_3897));   // verilog/motorControl.v(44[31:51])
    defparam pwm_23__I_819_i7_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 pwm_23__I_819_i9_2_lut (.I0(\PID_CONTROLLER.result [4]), .I1(pwm_23__N_2960[4]), 
            .I2(GND_net), .I3(GND_net), .O(n9_adj_3898));   // verilog/motorControl.v(44[31:51])
    defparam pwm_23__I_819_i9_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_14_i351_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral [3]), 
            .I2(GND_net), .I3(GND_net), .O(n521));   // verilog/motorControl.v(43[48:59])
    defparam mult_14_i351_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i2_3_lut_adj_1409 (.I0(\PID_CONTROLLER.result [28]), .I1(\PID_CONTROLLER.result [30]), 
            .I2(\PID_CONTROLLER.result [29]), .I3(GND_net), .O(n40124));   // verilog/motorControl.v(45[12:27])
    defparam i2_3_lut_adj_1409.LUT_INIT = 16'h8080;
    SB_LUT4 pwm_23__I_819_i15_2_lut (.I0(\PID_CONTROLLER.result [7]), .I1(pwm_23__N_2960[7]), 
            .I2(GND_net), .I3(GND_net), .O(n15_adj_3899));   // verilog/motorControl.v(44[31:51])
    defparam pwm_23__I_819_i15_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_12_i408_2_lut (.I0(\Kd[6] ), .I1(n57[8]), .I2(GND_net), 
            .I3(GND_net), .O(n607_adj_3728));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i408_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 pwm_23__I_819_i19_2_lut (.I0(\PID_CONTROLLER.result [9]), .I1(pwm_23__N_2960[9]), 
            .I2(GND_net), .I3(GND_net), .O(n19_adj_3900));   // verilog/motorControl.v(44[31:51])
    defparam pwm_23__I_819_i19_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i5_3_lut (.I0(\PID_CONTROLLER.result [25]), .I1(\PID_CONTROLLER.result [22]), 
            .I2(\PID_CONTROLLER.result [18]), .I3(GND_net), .O(n14_adj_3901));   // verilog/motorControl.v(38[14] 59[8])
    defparam i5_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 i6_4_lut (.I0(\PID_CONTROLLER.result [23]), .I1(\PID_CONTROLLER.result [21]), 
            .I2(\PID_CONTROLLER.result [19]), .I3(\PID_CONTROLLER.result [17]), 
            .O(n15_adj_3902));   // verilog/motorControl.v(38[14] 59[8])
    defparam i6_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i8_4_lut_adj_1410 (.I0(n15_adj_3902), .I1(\PID_CONTROLLER.result [20]), 
            .I2(n14_adj_3901), .I3(\PID_CONTROLLER.result [24]), .O(n40200));   // verilog/motorControl.v(38[14] 59[8])
    defparam i8_4_lut_adj_1410.LUT_INIT = 16'h8000;
    SB_LUT4 mult_12_i357_2_lut (.I0(\Kd[5] ), .I1(n57[15]), .I2(GND_net), 
            .I3(GND_net), .O(n531_adj_3726));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i357_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_20_i15_2_lut (.I0(\PWMLimit[7] ), .I1(\PID_CONTROLLER.result [7]), 
            .I2(GND_net), .I3(GND_net), .O(n15_adj_3903));   // verilog/motorControl.v(45[12:27])
    defparam LessThan_20_i15_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_20_i9_2_lut (.I0(\PWMLimit[4] ), .I1(\PID_CONTROLLER.result [4]), 
            .I2(GND_net), .I3(GND_net), .O(n9_adj_3904));   // verilog/motorControl.v(45[12:27])
    defparam LessThan_20_i9_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_4_lut_adj_1411 (.I0(Kd_delay_counter[1]), .I1(Kd_delay_counter[0]), 
            .I2(Kd_delay_counter[2]), .I3(Kd_delay_counter[6]), .O(n6_adj_3905));   // verilog/motorControl.v(56[10:29])
    defparam i1_4_lut_adj_1411.LUT_INIT = 16'hfffe;
    SB_LUT4 i4_4_lut (.I0(Kd_delay_counter[5]), .I1(Kd_delay_counter[4]), 
            .I2(Kd_delay_counter[3]), .I3(n6_adj_3905), .O(n41887));   // verilog/motorControl.v(56[10:29])
    defparam i4_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 mult_10_i73_2_lut (.I0(\Kp[1] ), .I1(\PID_CONTROLLER.err[3] ), 
            .I2(GND_net), .I3(GND_net), .O(n107_adj_3725));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i73_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_20_i4_4_lut (.I0(\PWMLimit[0] ), .I1(\PID_CONTROLLER.result [1]), 
            .I2(\PWMLimit[1] ), .I3(\PID_CONTROLLER.result [0]), .O(n4_adj_3906));   // verilog/motorControl.v(45[12:27])
    defparam LessThan_20_i4_4_lut.LUT_INIT = 16'h4d0c;
    SB_LUT4 mult_10_i10_2_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err[4] ), 
            .I2(GND_net), .I3(GND_net), .O(n14_adj_3724));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i10_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i30139_3_lut (.I0(n4_adj_3906), .I1(\PID_CONTROLLER.result[5] ), 
            .I2(n11_adj_12), .I3(GND_net), .O(n45660));   // verilog/motorControl.v(45[12:27])
    defparam i30139_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_10_i138_2_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err[3] ), 
            .I2(GND_net), .I3(GND_net), .O(n204_adj_3723));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i138_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i30140_3_lut (.I0(n45660), .I1(\PID_CONTROLLER.result[6] ), 
            .I2(n13_adj_13), .I3(GND_net), .O(n45661));   // verilog/motorControl.v(45[12:27])
    defparam i30140_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_12_i422_2_lut (.I0(\Kd[6] ), .I1(n57[15]), .I2(GND_net), 
            .I3(GND_net), .O(n628));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i422_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i29676_4_lut (.I0(n13_adj_13), .I1(n11_adj_12), .I2(n9_adj_3904), 
            .I3(n44552), .O(n45197));
    defparam i29676_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 mult_10_i203_2_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err[3] ), 
            .I2(GND_net), .I3(GND_net), .O(n301_adj_3722));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i203_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i473_2_lut (.I0(\Kd[7] ), .I1(n57[8]), .I2(GND_net), 
            .I3(GND_net), .O(n704_adj_3721));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i473_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_20_i8_3_lut (.I0(n6), .I1(\PID_CONTROLLER.result [4]), 
            .I2(n9_adj_3904), .I3(GND_net), .O(n8_adj_3909));   // verilog/motorControl.v(45[12:27])
    defparam LessThan_20_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i29567_3_lut (.I0(n45661), .I1(\PID_CONTROLLER.result [7]), 
            .I2(n15_adj_3903), .I3(GND_net), .O(n45088));   // verilog/motorControl.v(45[12:27])
    defparam i29567_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i30189_4_lut (.I0(n45088), .I1(n8_adj_3909), .I2(n15_adj_3903), 
            .I3(n45197), .O(n45710));   // verilog/motorControl.v(45[12:27])
    defparam i30189_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i30190_3_lut (.I0(n45710), .I1(\PID_CONTROLLER.result [8]), 
            .I2(\PWMLimit[8] ), .I3(GND_net), .O(n18_adj_3910));   // verilog/motorControl.v(45[12:27])
    defparam i30190_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 mult_14_i59_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral [4]), 
            .I2(GND_net), .I3(GND_net), .O(n86_adj_3720));   // verilog/motorControl.v(43[48:59])
    defparam mult_14_i59_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_14_i12_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral [5]), 
            .I2(GND_net), .I3(GND_net), .O(n17_adj_3719));   // verilog/motorControl.v(43[48:59])
    defparam mult_14_i12_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_14_i108_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral [4]), 
            .I2(GND_net), .I3(GND_net), .O(n159));   // verilog/motorControl.v(43[48:59])
    defparam mult_14_i108_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_14_i157_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral [4]), 
            .I2(GND_net), .I3(GND_net), .O(n232_adj_3718));   // verilog/motorControl.v(43[48:59])
    defparam mult_14_i157_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i3_4_lut_adj_1412 (.I0(\PID_CONTROLLER.result [11]), .I1(n18_adj_3910), 
            .I2(\PID_CONTROLLER.result [9]), .I3(\PID_CONTROLLER.result [10]), 
            .O(n41755));   // verilog/motorControl.v(45[12:27])
    defparam i3_4_lut_adj_1412.LUT_INIT = 16'hfffe;
    SB_LUT4 mult_14_i206_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral [4]), 
            .I2(GND_net), .I3(GND_net), .O(n305));   // verilog/motorControl.v(43[48:59])
    defparam mult_14_i206_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_14_i255_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral [4]), 
            .I2(GND_net), .I3(GND_net), .O(n378));   // verilog/motorControl.v(43[48:59])
    defparam mult_14_i255_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i2_4_lut_adj_1413 (.I0(n18_adj_3910), .I1(\PID_CONTROLLER.result [10]), 
            .I2(\PID_CONTROLLER.result [9]), .I3(\PID_CONTROLLER.result [11]), 
            .O(n41486));   // verilog/motorControl.v(45[12:27])
    defparam i2_4_lut_adj_1413.LUT_INIT = 16'h8000;
    SB_LUT4 mult_14_i304_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral [4]), 
            .I2(GND_net), .I3(GND_net), .O(n451));   // verilog/motorControl.v(43[48:59])
    defparam mult_14_i304_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_14_i353_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral [4]), 
            .I2(GND_net), .I3(GND_net), .O(n524));   // verilog/motorControl.v(43[48:59])
    defparam mult_14_i353_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i268_2_lut (.I0(\Kp[4] ), .I1(\PID_CONTROLLER.err[3] ), 
            .I2(GND_net), .I3(GND_net), .O(n398_adj_3713));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i268_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i333_2_lut (.I0(\Kp[5] ), .I1(\PID_CONTROLLER.err[3] ), 
            .I2(GND_net), .I3(GND_net), .O(n495_adj_3712));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i333_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1_4_lut_adj_1414 (.I0(\PID_CONTROLLER.result [12]), .I1(\PWMLimit[9] ), 
            .I2(n41486), .I3(n41755), .O(n26_adj_3911));   // verilog/motorControl.v(45[12:27])
    defparam i1_4_lut_adj_1414.LUT_INIT = 16'hb3a2;
    SB_LUT4 mult_10_i398_2_lut (.I0(\Kp[6] ), .I1(\PID_CONTROLLER.err[3] ), 
            .I2(GND_net), .I3(GND_net), .O(n592_adj_3711));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i398_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i463_2_lut (.I0(\Kp[7] ), .I1(\PID_CONTROLLER.err[3] ), 
            .I2(GND_net), .I3(GND_net), .O(n689_adj_3710));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i463_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i3_4_lut_adj_1415 (.I0(\PID_CONTROLLER.result [23]), .I1(\PID_CONTROLLER.result [24]), 
            .I2(\PID_CONTROLLER.result [22]), .I3(\PID_CONTROLLER.result [25]), 
            .O(n62_adj_3874));   // verilog/motorControl.v(38[14] 59[8])
    defparam i3_4_lut_adj_1415.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_adj_1416 (.I0(\PID_CONTROLLER.result [21]), .I1(\PID_CONTROLLER.result [19]), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_3912));   // verilog/motorControl.v(38[14] 59[8])
    defparam i1_2_lut_adj_1416.LUT_INIT = 16'heeee;
    SB_LUT4 i4_4_lut_adj_1417 (.I0(\PID_CONTROLLER.result [20]), .I1(\PID_CONTROLLER.result [17]), 
            .I2(\PID_CONTROLLER.result [18]), .I3(n6_adj_3912), .O(n49_adj_3870));   // verilog/motorControl.v(38[14] 59[8])
    defparam i4_4_lut_adj_1417.LUT_INIT = 16'hfffe;
    SB_LUT4 i3_4_lut_adj_1418 (.I0(\PID_CONTROLLER.result [15]), .I1(n26_adj_3911), 
            .I2(\PID_CONTROLLER.result [13]), .I3(\PID_CONTROLLER.result [14]), 
            .O(n41766));   // verilog/motorControl.v(45[12:27])
    defparam i3_4_lut_adj_1418.LUT_INIT = 16'hfffe;
    SB_LUT4 i2_4_lut_adj_1419 (.I0(n26_adj_3911), .I1(\PID_CONTROLLER.result [14]), 
            .I2(\PID_CONTROLLER.result [13]), .I3(\PID_CONTROLLER.result [15]), 
            .O(n41485));   // verilog/motorControl.v(45[12:27])
    defparam i2_4_lut_adj_1419.LUT_INIT = 16'h8000;
    SB_LUT4 i1_4_lut_adj_1420 (.I0(\PID_CONTROLLER.result [16]), .I1(\PWMLimit[9] ), 
            .I2(n41485), .I3(n41766), .O(n34_adj_3913));   // verilog/motorControl.v(45[12:27])
    defparam i1_4_lut_adj_1420.LUT_INIT = 16'hb3a2;
    SB_LUT4 i3_4_lut_adj_1421 (.I0(\PID_CONTROLLER.result [26]), .I1(n34_adj_3913), 
            .I2(n49_adj_3870), .I3(n62_adj_3874), .O(n41915));   // verilog/motorControl.v(38[14] 59[8])
    defparam i3_4_lut_adj_1421.LUT_INIT = 16'hfffe;
    SB_LUT4 i2_3_lut_adj_1422 (.I0(n40200), .I1(\PID_CONTROLLER.result [26]), 
            .I2(n34_adj_3913), .I3(GND_net), .O(n41828));
    defparam i2_3_lut_adj_1422.LUT_INIT = 16'h8080;
    SB_LUT4 i1_4_lut_adj_1423 (.I0(\PID_CONTROLLER.result [27]), .I1(\PWMLimit[9] ), 
            .I2(n41828), .I3(n41915), .O(n56_adj_3914));   // verilog/motorControl.v(45[12:27])
    defparam i1_4_lut_adj_1423.LUT_INIT = 16'hb3a2;
    SB_LUT4 i3_4_lut_adj_1424 (.I0(\PID_CONTROLLER.result [30]), .I1(n56_adj_3914), 
            .I2(\PID_CONTROLLER.result [28]), .I3(\PID_CONTROLLER.result [29]), 
            .O(n41769));   // verilog/motorControl.v(45[12:27])
    defparam i3_4_lut_adj_1424.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1425 (.I0(\PWMLimit[9] ), .I1(\PID_CONTROLLER.result [31]), 
            .I2(n40126), .I3(n41769), .O(n387));   // verilog/motorControl.v(45[12:27])
    defparam i1_4_lut_adj_1425.LUT_INIT = 16'hb3a2;
    SB_LUT4 i1_3_lut_adj_1426 (.I0(\PID_CONTROLLER.result [22]), .I1(\PID_CONTROLLER.result [21]), 
            .I2(pwm_23__N_2960[10]), .I3(GND_net), .O(n4_adj_3915));   // verilog/motorControl.v(44[31:51])
    defparam i1_3_lut_adj_1426.LUT_INIT = 16'h7e7e;
    SB_LUT4 i2_4_lut_adj_1427 (.I0(\PID_CONTROLLER.result [13]), .I1(\PID_CONTROLLER.result [30]), 
            .I2(n4_adj_3915), .I3(pwm_23__N_2960[10]), .O(n13_adj_3916));   // verilog/motorControl.v(44[31:51])
    defparam i2_4_lut_adj_1427.LUT_INIT = 16'hf7fe;
    SB_LUT4 mult_14_i61_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral [5]), 
            .I2(GND_net), .I3(GND_net), .O(n89));   // verilog/motorControl.v(43[48:59])
    defparam mult_14_i61_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i7_4_lut_adj_1428 (.I0(n13_adj_3916), .I1(\PID_CONTROLLER.result [11]), 
            .I2(\PID_CONTROLLER.result [20]), .I3(pwm_23__N_2960[10]), .O(n18_adj_3917));   // verilog/motorControl.v(44[31:51])
    defparam i7_4_lut_adj_1428.LUT_INIT = 16'hbffe;
    SB_LUT4 mult_14_i14_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral [6]), 
            .I2(GND_net), .I3(GND_net), .O(n20_adj_3709));   // verilog/motorControl.v(43[48:59])
    defparam mult_14_i14_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_14_i110_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral [5]), 
            .I2(GND_net), .I3(GND_net), .O(n162));   // verilog/motorControl.v(43[48:59])
    defparam mult_14_i110_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i5_3_lut_adj_1429 (.I0(\PID_CONTROLLER.result [15]), .I1(\PID_CONTROLLER.result [16]), 
            .I2(pwm_23__N_2960[10]), .I3(GND_net), .O(n16_adj_3918));   // verilog/motorControl.v(44[31:51])
    defparam i5_3_lut_adj_1429.LUT_INIT = 16'h7e7e;
    SB_LUT4 mult_12_i487_2_lut (.I0(\Kd[7] ), .I1(n57[15]), .I2(GND_net), 
            .I3(GND_net), .O(n725));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i487_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_14_i159_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral [5]), 
            .I2(GND_net), .I3(GND_net), .O(n235_adj_3708));   // verilog/motorControl.v(43[48:59])
    defparam mult_14_i159_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_14_i208_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral [5]), 
            .I2(GND_net), .I3(GND_net), .O(n308_adj_3706));   // verilog/motorControl.v(43[48:59])
    defparam mult_14_i208_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_14_i257_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral [5]), 
            .I2(GND_net), .I3(GND_net), .O(n381));   // verilog/motorControl.v(43[48:59])
    defparam mult_14_i257_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_14_i306_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral [5]), 
            .I2(GND_net), .I3(GND_net), .O(n454));   // verilog/motorControl.v(43[48:59])
    defparam mult_14_i306_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i6_4_lut_adj_1430 (.I0(\PID_CONTROLLER.result [12]), .I1(\PID_CONTROLLER.result [26]), 
            .I2(pwm_23__N_2960[10]), .I3(\PID_CONTROLLER.result [17]), .O(n17_adj_3919));   // verilog/motorControl.v(44[31:51])
    defparam i6_4_lut_adj_1430.LUT_INIT = 16'h7ffe;
    SB_LUT4 mult_14_i355_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral [5]), 
            .I2(GND_net), .I3(GND_net), .O(n527));   // verilog/motorControl.v(43[48:59])
    defparam mult_14_i355_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i4_3_lut (.I0(\PID_CONTROLLER.result [29]), .I1(\PID_CONTROLLER.result [19]), 
            .I2(pwm_23__N_2960[10]), .I3(GND_net), .O(n15_adj_3920));   // verilog/motorControl.v(44[31:51])
    defparam i4_3_lut.LUT_INIT = 16'h7e7e;
    SB_LUT4 i10_4_lut_adj_1431 (.I0(n15_adj_3920), .I1(n17_adj_3919), .I2(n16_adj_3918), 
            .I3(n18_adj_3917), .O(n41951));   // verilog/motorControl.v(44[31:51])
    defparam i10_4_lut_adj_1431.LUT_INIT = 16'hfffe;
    SB_LUT4 i14794_1_lut (.I0(\PID_CONTROLLER.result [0]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n28200));   // verilog/motorControl.v(38[14] 59[8])
    defparam i14794_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_17_inv_0_i1_1_lut (.I0(\deadband[0] ), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n82[0]));   // verilog/motorControl.v(44[41:50])
    defparam unary_minus_17_inv_0_i1_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 pwm_23__I_819_i5_2_lut (.I0(\PID_CONTROLLER.result [2]), .I1(pwm_23__N_2960[2]), 
            .I2(GND_net), .I3(GND_net), .O(n5_adj_3921));   // verilog/motorControl.v(44[31:51])
    defparam pwm_23__I_819_i5_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_12_i107_2_lut (.I0(\Kd[1] ), .I1(n57[20]), .I2(GND_net), 
            .I3(GND_net), .O(n158_adj_3700));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i107_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i29081_4_lut (.I0(n11_adj_14), .I1(n9_adj_3898), .I2(n7_adj_3897), 
            .I3(n5_adj_3921), .O(n44602));
    defparam i29081_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 mult_12_i44_2_lut (.I0(\Kd[0] ), .I1(n57[21]), .I2(GND_net), 
            .I3(GND_net), .O(n65_adj_3699));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i44_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 pwm_23__I_819_i8_3_lut (.I0(pwm_23__N_2960[4]), .I1(pwm_23__N_2960[8]), 
            .I2(n17_adj_3896), .I3(GND_net), .O(n8_adj_3923));   // verilog/motorControl.v(44[31:51])
    defparam pwm_23__I_819_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 pwm_23__I_819_i6_3_lut (.I0(pwm_23__N_2960[2]), .I1(pwm_23__N_2960[3]), 
            .I2(n7_adj_3897), .I3(GND_net), .O(n6_adj_3924));   // verilog/motorControl.v(44[31:51])
    defparam pwm_23__I_819_i6_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 pwm_23__I_819_i16_3_lut (.I0(n8_adj_3923), .I1(pwm_23__N_2960[9]), 
            .I2(n19_adj_3900), .I3(GND_net), .O(n16_adj_3925));   // verilog/motorControl.v(44[31:51])
    defparam pwm_23__I_819_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_12_i77_2_lut (.I0(\Kd[1] ), .I1(n57[5]), .I2(GND_net), 
            .I3(GND_net), .O(n113_adj_3698));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i77_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i14_2_lut (.I0(\Kd[0] ), .I1(n57[6]), .I2(GND_net), 
            .I3(GND_net), .O(n20_adj_3697));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i14_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i28891_4_lut (.I0(n50_adj_3891), .I1(\PID_CONTROLLER.result [26]), 
            .I2(\deadband[9] ), .I3(\PID_CONTROLLER.result [25]), .O(n44041));   // verilog/motorControl.v(44[10:27])
    defparam i28891_4_lut.LUT_INIT = 16'h8f0e;
    SB_LUT4 pwm_23__I_819_i4_3_lut (.I0(n44044), .I1(pwm_23__N_2960[1]), 
            .I2(\PID_CONTROLLER.result [1]), .I3(GND_net), .O(n4_adj_3926));   // verilog/motorControl.v(44[31:51])
    defparam pwm_23__I_819_i4_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 unary_minus_17_inv_0_i2_1_lut (.I0(\deadband[1] ), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n82[1]));   // verilog/motorControl.v(44[41:50])
    defparam unary_minus_17_inv_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i30141_3_lut (.I0(n4_adj_3926), .I1(\pwm_23__N_2960[5] ), .I2(n11_adj_14), 
            .I3(GND_net), .O(n45662));   // verilog/motorControl.v(44[31:51])
    defparam i30141_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_12_i172_2_lut (.I0(\Kd[2] ), .I1(n57[20]), .I2(GND_net), 
            .I3(GND_net), .O(n255_adj_3695));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i172_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i142_2_lut (.I0(\Kd[2] ), .I1(n57[5]), .I2(GND_net), 
            .I3(GND_net), .O(n210_adj_3694));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i142_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i207_2_lut (.I0(\Kd[3] ), .I1(n57[5]), .I2(GND_net), 
            .I3(GND_net), .O(n307_adj_3693));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i207_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i272_2_lut (.I0(\Kd[4] ), .I1(n57[5]), .I2(GND_net), 
            .I3(GND_net), .O(n404_adj_3692));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i272_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i30142_3_lut (.I0(n45662), .I1(\pwm_23__N_2960[6] ), .I2(n13_adj_15), 
            .I3(GND_net), .O(n45663));   // verilog/motorControl.v(44[31:51])
    defparam i30142_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i5_4_lut_adj_1432 (.I0(\PID_CONTROLLER.result [25]), .I1(\PID_CONTROLLER.result [18]), 
            .I2(pwm_23__N_2960[10]), .I3(n41951), .O(n14_adj_3928));   // verilog/motorControl.v(44[31:51])
    defparam i5_4_lut_adj_1432.LUT_INIT = 16'hff7e;
    SB_LUT4 i3_3_lut_adj_1433 (.I0(\PID_CONTROLLER.result [14]), .I1(\PID_CONTROLLER.result [24]), 
            .I2(pwm_23__N_2960[10]), .I3(GND_net), .O(n12_adj_3929));   // verilog/motorControl.v(44[31:51])
    defparam i3_3_lut_adj_1433.LUT_INIT = 16'h7e7e;
    SB_LUT4 i4_3_lut_adj_1434 (.I0(\PID_CONTROLLER.result [27]), .I1(\PID_CONTROLLER.result [28]), 
            .I2(pwm_23__N_2960[10]), .I3(GND_net), .O(n13_adj_3930));   // verilog/motorControl.v(44[31:51])
    defparam i4_3_lut_adj_1434.LUT_INIT = 16'h7e7e;
    SB_LUT4 i2_3_lut_adj_1435 (.I0(\PID_CONTROLLER.result [10]), .I1(\PID_CONTROLLER.result [23]), 
            .I2(pwm_23__N_2960[10]), .I3(GND_net), .O(n11_adj_3931));   // verilog/motorControl.v(44[31:51])
    defparam i2_3_lut_adj_1435.LUT_INIT = 16'h7e7e;
    SB_LUT4 i29071_4_lut (.I0(n17_adj_3896), .I1(n15_adj_3899), .I2(n13_adj_15), 
            .I3(n44602), .O(n44592));
    defparam i29071_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i30487_4_lut (.I0(n16_adj_3925), .I1(n6_adj_3924), .I2(n19_adj_3900), 
            .I3(n44590), .O(n46008));   // verilog/motorControl.v(44[31:51])
    defparam i30487_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i29565_3_lut (.I0(n45663), .I1(pwm_23__N_2960[7]), .I2(n15_adj_3899), 
            .I3(GND_net), .O(n45086));   // verilog/motorControl.v(44[31:51])
    defparam i29565_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8_4_lut_adj_1436 (.I0(n11_adj_3931), .I1(n13_adj_3930), .I2(n12_adj_3929), 
            .I3(n14_adj_3928), .O(n41904));   // verilog/motorControl.v(44[31:51])
    defparam i8_4_lut_adj_1436.LUT_INIT = 16'hfffe;
    SB_LUT4 i30635_4_lut (.I0(n45086), .I1(n46008), .I2(n19_adj_3900), 
            .I3(n44592), .O(n46156));   // verilog/motorControl.v(44[31:51])
    defparam i30635_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i29706_4_lut (.I0(\deadband[9] ), .I1(\PID_CONTROLLER.result [29]), 
            .I2(\PID_CONTROLLER.result [30]), .I3(\PID_CONTROLLER.result [28]), 
            .O(n45227));
    defparam i29706_4_lut.LUT_INIT = 16'h7ffe;
    SB_LUT4 \PID_CONTROLLER.result_31__I_0_i56_3_lut  (.I0(n44041), .I1(\PID_CONTROLLER.result [27]), 
            .I2(\deadband[9] ), .I3(GND_net), .O(n56_adj_3932));   // verilog/motorControl.v(44[10:27])
    defparam \PID_CONTROLLER.result_31__I_0_i56_3_lut .LUT_INIT = 16'h8e8e;
    SB_LUT4 \PID_CONTROLLER.result_31__I_0_i60_4_lut  (.I0(\PID_CONTROLLER.result [28]), 
            .I1(\PID_CONTROLLER.result [30]), .I2(\deadband[9] ), .I3(\PID_CONTROLLER.result [29]), 
            .O(n60));   // verilog/motorControl.v(44[10:27])
    defparam \PID_CONTROLLER.result_31__I_0_i60_4_lut .LUT_INIT = 16'h8f0e;
    SB_LUT4 i30605_4_lut (.I0(n46156), .I1(\PID_CONTROLLER.result [31]), 
            .I2(pwm_23__N_2960[10]), .I3(n41904), .O(pwm_23__N_2959));   // verilog/motorControl.v(44[31:51])
    defparam i30605_4_lut.LUT_INIT = 16'hcc8e;
    SB_LUT4 i30185_3_lut (.I0(n60), .I1(n56_adj_3932), .I2(n45227), .I3(GND_net), 
            .O(n45706));   // verilog/motorControl.v(44[10:27])
    defparam i30185_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 pwm_23__I_818_4_lut (.I0(n45706), .I1(pwm_23__N_2959), .I2(\deadband[9] ), 
            .I3(\PID_CONTROLLER.result [31]), .O(pwm_23__N_2957));   // verilog/motorControl.v(44[10:51])
    defparam pwm_23__I_818_4_lut.LUT_INIT = 16'hecfe;
    SB_LUT4 unary_minus_17_inv_0_i3_1_lut (.I0(\deadband[2] ), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n82[2]));   // verilog/motorControl.v(44[41:50])
    defparam unary_minus_17_inv_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_12_i237_2_lut (.I0(\Kd[3] ), .I1(n57[20]), .I2(GND_net), 
            .I3(GND_net), .O(n352_adj_3690));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i237_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i302_2_lut (.I0(\Kd[4] ), .I1(n57[20]), .I2(GND_net), 
            .I3(GND_net), .O(n449_adj_3689));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i302_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_14_i63_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral [6]), 
            .I2(GND_net), .I3(GND_net), .O(n92));   // verilog/motorControl.v(43[48:59])
    defparam mult_14_i63_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_14_i16_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral [7]), 
            .I2(GND_net), .I3(GND_net), .O(n23_adj_3688));   // verilog/motorControl.v(43[48:59])
    defparam mult_14_i16_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_14_i112_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral [6]), 
            .I2(GND_net), .I3(GND_net), .O(n165_adj_3687));   // verilog/motorControl.v(43[48:59])
    defparam mult_14_i112_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_14_i161_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral [6]), 
            .I2(GND_net), .I3(GND_net), .O(n238_adj_3685));   // verilog/motorControl.v(43[48:59])
    defparam mult_14_i161_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i337_2_lut (.I0(\Kd[5] ), .I1(n57[5]), .I2(GND_net), 
            .I3(GND_net), .O(n501_adj_3683));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i337_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i402_2_lut (.I0(\Kd[6] ), .I1(n57[5]), .I2(GND_net), 
            .I3(GND_net), .O(n598_adj_3682));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i402_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_14_i210_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral [6]), 
            .I2(GND_net), .I3(GND_net), .O(n311_adj_3681));   // verilog/motorControl.v(43[48:59])
    defparam mult_14_i210_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_17_inv_0_i4_1_lut (.I0(\deadband[3] ), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n82[3]));   // verilog/motorControl.v(44[41:50])
    defparam unary_minus_17_inv_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_14_i259_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral [6]), 
            .I2(GND_net), .I3(GND_net), .O(n384));   // verilog/motorControl.v(43[48:59])
    defparam mult_14_i259_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_14_i308_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral [6]), 
            .I2(GND_net), .I3(GND_net), .O(n457_c));   // verilog/motorControl.v(43[48:59])
    defparam mult_14_i308_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i467_2_lut (.I0(\Kd[7] ), .I1(n57[5]), .I2(GND_net), 
            .I3(GND_net), .O(n695_adj_3677));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i467_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_17_inv_0_i5_1_lut (.I0(\deadband[4] ), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n82[4]));   // verilog/motorControl.v(44[41:50])
    defparam unary_minus_17_inv_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_17_inv_0_i6_1_lut (.I0(\deadband[5] ), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n82[5]));   // verilog/motorControl.v(44[41:50])
    defparam unary_minus_17_inv_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_17_inv_0_i7_1_lut (.I0(\deadband[6] ), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n82[6]));   // verilog/motorControl.v(44[41:50])
    defparam unary_minus_17_inv_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_14_i357_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral [6]), 
            .I2(GND_net), .I3(GND_net), .O(n530));   // verilog/motorControl.v(43[48:59])
    defparam mult_14_i357_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_17_inv_0_i8_1_lut (.I0(\deadband[7] ), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n82[7]));   // verilog/motorControl.v(44[41:50])
    defparam unary_minus_17_inv_0_i8_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i93_2_lut (.I0(\Kp[1] ), .I1(\PID_CONTROLLER.err[13] ), 
            .I2(GND_net), .I3(GND_net), .O(n137_adj_3672));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i93_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i30_2_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err[14] ), 
            .I2(GND_net), .I3(GND_net), .O(n44_adj_3671));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i30_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i158_2_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err[13] ), 
            .I2(GND_net), .I3(GND_net), .O(n234_adj_3670));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i158_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 state_23__I_0_inv_0_i16_1_lut (.I0(setpoint[15]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n58[15]));   // verilog/motorControl.v(39[14:30])
    defparam state_23__I_0_inv_0_i16_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i223_2_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err[13] ), 
            .I2(GND_net), .I3(GND_net), .O(n331_adj_3669));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i223_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i288_2_lut (.I0(\Kp[4] ), .I1(\PID_CONTROLLER.err[13] ), 
            .I2(GND_net), .I3(GND_net), .O(n428_adj_3668));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i288_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_17_inv_0_i9_1_lut (.I0(\deadband[8] ), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n82[8]));   // verilog/motorControl.v(44[41:50])
    defparam unary_minus_17_inv_0_i9_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_17_inv_0_i32_1_lut (.I0(\deadband[9] ), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n82[31]));   // verilog/motorControl.v(44[41:50])
    defparam unary_minus_17_inv_0_i32_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i353_2_lut (.I0(\Kp[5] ), .I1(\PID_CONTROLLER.err[13] ), 
            .I2(GND_net), .I3(GND_net), .O(n525_adj_3664));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i353_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_inv_0_i1_1_lut (.I0(IntegralLimit[0]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n79[0]));   // verilog/motorControl.v(40[48:62])
    defparam unary_minus_5_inv_0_i1_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i418_2_lut (.I0(\Kp[6] ), .I1(\PID_CONTROLLER.err[13] ), 
            .I2(GND_net), .I3(GND_net), .O(n622_adj_3661));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i418_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i483_2_lut (.I0(\Kp[7] ), .I1(\PID_CONTROLLER.err[13] ), 
            .I2(GND_net), .I3(GND_net), .O(n719_adj_3660));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i483_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_inv_0_i2_1_lut (.I0(IntegralLimit[1]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n79[1]));   // verilog/motorControl.v(40[48:62])
    defparam unary_minus_5_inv_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_12_i93_2_lut (.I0(\Kd[1] ), .I1(n57[13]), .I2(GND_net), 
            .I3(GND_net), .O(n137_adj_3657));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i93_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i30_2_lut (.I0(\Kd[0] ), .I1(n57[14]), .I2(GND_net), 
            .I3(GND_net), .O(n44_adj_3656));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i30_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_inv_0_i3_1_lut (.I0(IntegralLimit[2]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n79[2]));   // verilog/motorControl.v(40[48:62])
    defparam unary_minus_5_inv_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_5_inv_0_i4_1_lut (.I0(IntegralLimit[3]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n79[3]));   // verilog/motorControl.v(40[48:62])
    defparam unary_minus_5_inv_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_5_inv_0_i5_1_lut (.I0(IntegralLimit[4]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n79[4]));   // verilog/motorControl.v(40[48:62])
    defparam unary_minus_5_inv_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_5_inv_0_i6_1_lut (.I0(IntegralLimit[5]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n79[5]));   // verilog/motorControl.v(40[48:62])
    defparam unary_minus_5_inv_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_5_inv_0_i7_1_lut (.I0(IntegralLimit[6]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n79[6]));   // verilog/motorControl.v(40[48:62])
    defparam unary_minus_5_inv_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_5_inv_0_i8_1_lut (.I0(IntegralLimit[7]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n79[7]));   // verilog/motorControl.v(40[48:62])
    defparam unary_minus_5_inv_0_i8_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_12_i158_2_lut (.I0(\Kd[2] ), .I1(n57[13]), .I2(GND_net), 
            .I3(GND_net), .O(n234_adj_3643));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i158_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i89_2_lut (.I0(\Kd[1] ), .I1(n57[11]), .I2(GND_net), 
            .I3(GND_net), .O(n131_adj_3642));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i89_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i26_2_lut (.I0(\Kd[0] ), .I1(n57[12]), .I2(GND_net), 
            .I3(GND_net), .O(n38_adj_3641));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i26_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i117_2_lut (.I0(\Kd[1] ), .I1(n57[25]), .I2(GND_net), 
            .I3(GND_net), .O(n182_adj_3640));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i117_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_inv_0_i9_1_lut (.I0(IntegralLimit[8]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n79[8]));   // verilog/motorControl.v(40[48:62])
    defparam unary_minus_5_inv_0_i9_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_12_i182_2_lut (.I0(\Kd[2] ), .I1(n57[25]), .I2(GND_net), 
            .I3(GND_net), .O(n276));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i182_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_inv_0_i10_1_lut (.I0(IntegralLimit[9]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n79[9]));   // verilog/motorControl.v(40[48:62])
    defparam unary_minus_5_inv_0_i10_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_12_i367_2_lut (.I0(\Kd[5] ), .I1(n57[20]), .I2(GND_net), 
            .I3(GND_net), .O(n546_adj_3635));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i367_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_inv_0_i11_1_lut (.I0(IntegralLimit[10]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n79[10]));   // verilog/motorControl.v(40[48:62])
    defparam unary_minus_5_inv_0_i11_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_5_inv_0_i12_1_lut (.I0(IntegralLimit[11]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n79[11]));   // verilog/motorControl.v(40[48:62])
    defparam unary_minus_5_inv_0_i12_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_5_inv_0_i13_1_lut (.I0(IntegralLimit[12]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n79[12]));   // verilog/motorControl.v(40[48:62])
    defparam unary_minus_5_inv_0_i13_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_12_i432_2_lut (.I0(\Kd[6] ), .I1(n57[20]), .I2(GND_net), 
            .I3(GND_net), .O(n643_adj_3627));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i432_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i154_2_lut (.I0(\Kd[2] ), .I1(n57[11]), .I2(GND_net), 
            .I3(GND_net), .O(n228_adj_3626));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i154_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i497_2_lut (.I0(\Kd[7] ), .I1(n57[20]), .I2(GND_net), 
            .I3(GND_net), .O(n740_adj_3625));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i497_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i223_2_lut (.I0(\Kd[3] ), .I1(n57[13]), .I2(GND_net), 
            .I3(GND_net), .O(n331));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i223_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i2_4_lut_adj_1437 (.I0(\Kd[2] ), .I1(\Kd[0] ), .I2(n57[25]), 
            .I3(\Kd[1] ), .O(n4_adj_3856));   // verilog/motorControl.v(43[26:45])
    defparam i2_4_lut_adj_1437.LUT_INIT = 16'ha080;
    SB_LUT4 mult_12_i247_2_lut (.I0(\Kd[3] ), .I1(n57[25]), .I2(GND_net), 
            .I3(GND_net), .O(n370));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i247_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i20345_3_lut (.I0(n57[25]), .I1(n33897), .I2(n33872), .I3(GND_net), 
            .O(n10111[1]));   // verilog/motorControl.v(43[26:45])
    defparam i20345_3_lut.LUT_INIT = 16'h6c6c;
    SB_LUT4 mult_12_i312_2_lut (.I0(\Kd[4] ), .I1(n57[25]), .I2(GND_net), 
            .I3(GND_net), .O(n464_adj_3628));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i312_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i379_2_lut (.I0(\Kd[5] ), .I1(n57[25]), .I2(GND_net), 
            .I3(GND_net), .O(n564));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i379_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i442_2_lut (.I0(\Kd[6] ), .I1(n57[25]), .I2(GND_net), 
            .I3(GND_net), .O(n658));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i442_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i5_4_lut_adj_1438 (.I0(n33897), .I1(n7_adj_3857), .I2(n8_adj_3933), 
            .I3(n8_adj_3934), .O(n41372));   // verilog/motorControl.v(43[26:45])
    defparam i5_4_lut_adj_1438.LUT_INIT = 16'h6996;
    SB_LUT4 unary_minus_5_inv_0_i14_1_lut (.I0(IntegralLimit[13]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n79[13]));   // verilog/motorControl.v(40[48:62])
    defparam unary_minus_5_inv_0_i14_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_12_i2_2_lut (.I0(\Kd[0] ), .I1(n57[0]), .I2(GND_net), 
            .I3(GND_net), .O(n191[0]));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i2_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_inv_0_i15_1_lut (.I0(IntegralLimit[14]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n79[14]));   // verilog/motorControl.v(40[48:62])
    defparam unary_minus_5_inv_0_i15_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_14_i65_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral [7]), 
            .I2(GND_net), .I3(GND_net), .O(n95));   // verilog/motorControl.v(43[48:59])
    defparam mult_14_i65_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_14_i18_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral [8]), 
            .I2(GND_net), .I3(GND_net), .O(n26_adj_3620));   // verilog/motorControl.v(43[48:59])
    defparam mult_14_i18_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_14_i114_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral [7]), 
            .I2(GND_net), .I3(GND_net), .O(n168_adj_3619));   // verilog/motorControl.v(43[48:59])
    defparam mult_14_i114_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_14_i163_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral [7]), 
            .I2(GND_net), .I3(GND_net), .O(n241_adj_3617));   // verilog/motorControl.v(43[48:59])
    defparam mult_14_i163_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_14_i212_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral [7]), 
            .I2(GND_net), .I3(GND_net), .O(n314_adj_3615));   // verilog/motorControl.v(43[48:59])
    defparam mult_14_i212_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i219_2_lut (.I0(\Kd[3] ), .I1(n57[11]), .I2(GND_net), 
            .I3(GND_net), .O(n325_adj_3613));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i219_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i288_2_lut (.I0(\Kd[4] ), .I1(n57[13]), .I2(GND_net), 
            .I3(GND_net), .O(n428));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i288_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_14_i261_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral [7]), 
            .I2(GND_net), .I3(GND_net), .O(n387_c));   // verilog/motorControl.v(43[48:59])
    defparam mult_14_i261_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_inv_0_i16_1_lut (.I0(IntegralLimit[15]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n79[15]));   // verilog/motorControl.v(40[48:62])
    defparam unary_minus_5_inv_0_i16_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_14_i310_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral [7]), 
            .I2(GND_net), .I3(GND_net), .O(n460_c));   // verilog/motorControl.v(43[48:59])
    defparam mult_14_i310_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_inv_0_i17_1_lut (.I0(IntegralLimit[16]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n79[16]));   // verilog/motorControl.v(40[48:62])
    defparam unary_minus_5_inv_0_i17_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_14_i359_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral [7]), 
            .I2(GND_net), .I3(GND_net), .O(n533));   // verilog/motorControl.v(43[48:59])
    defparam mult_14_i359_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_inv_0_i18_1_lut (.I0(IntegralLimit[17]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n79[17]));   // verilog/motorControl.v(40[48:62])
    defparam unary_minus_5_inv_0_i18_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_5_inv_0_i19_1_lut (.I0(IntegralLimit[18]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n79[18]));   // verilog/motorControl.v(40[48:62])
    defparam unary_minus_5_inv_0_i19_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_12_i353_2_lut (.I0(\Kd[5] ), .I1(n57[13]), .I2(GND_net), 
            .I3(GND_net), .O(n525));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i353_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i99_2_lut (.I0(\Kd[1] ), .I1(n57[16]), .I2(GND_net), 
            .I3(GND_net), .O(n146_adj_3600));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i99_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i36_2_lut (.I0(\Kd[0] ), .I1(n57[17]), .I2(GND_net), 
            .I3(GND_net), .O(n53_adj_3599));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i36_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_inv_0_i20_1_lut (.I0(IntegralLimit[19]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n79[19]));   // verilog/motorControl.v(40[48:62])
    defparam unary_minus_5_inv_0_i20_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i4_2_lut_adj_1439 (.I0(n19_adj_3636), .I1(n25_adj_3629), .I2(GND_net), 
            .I3(GND_net), .O(n18_adj_3935));   // verilog/motorControl.v(40[38:63])
    defparam i4_2_lut_adj_1439.LUT_INIT = 16'heeee;
    SB_LUT4 i10_4_lut_adj_1440 (.I0(n33_adj_3608), .I1(n43_adj_3575), .I2(n27_adj_3623), 
            .I3(n35_adj_3604), .O(n24_adj_3936));   // verilog/motorControl.v(40[38:63])
    defparam i10_4_lut_adj_1440.LUT_INIT = 16'hfffe;
    SB_LUT4 i8_4_lut_adj_1441 (.I0(n41_adj_3592), .I1(n45_adj_3573), .I2(n31_adj_3611), 
            .I3(n23_adj_3631), .O(n22_adj_3937));   // verilog/motorControl.v(40[38:63])
    defparam i8_4_lut_adj_1441.LUT_INIT = 16'hfffe;
    SB_LUT4 i12_4_lut_adj_1442 (.I0(n29_adj_3621), .I1(n24_adj_3936), .I2(n18_adj_3935), 
            .I3(n37_adj_3601), .O(n26_adj_3938));   // verilog/motorControl.v(40[38:63])
    defparam i12_4_lut_adj_1442.LUT_INIT = 16'hfffe;
    SB_LUT4 i13_4_lut_adj_1443 (.I0(n21_adj_3633), .I1(n26_adj_3938), .I2(n22_adj_3937), 
            .I3(n39_adj_3597), .O(n41724));   // verilog/motorControl.v(40[38:63])
    defparam i13_4_lut_adj_1443.LUT_INIT = 16'hfffe;
    SB_LUT4 LessThan_4_i11_2_lut (.I0(\PID_CONTROLLER.integral [5]), .I1(IntegralLimit[5]), 
            .I2(GND_net), .I3(GND_net), .O(n11_adj_3939));   // verilog/motorControl.v(40[10:34])
    defparam LessThan_4_i11_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_4_i9_2_lut (.I0(\PID_CONTROLLER.integral [4]), .I1(IntegralLimit[4]), 
            .I2(GND_net), .I3(GND_net), .O(n9_adj_3940));   // verilog/motorControl.v(40[10:34])
    defparam LessThan_4_i9_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_4_i17_2_lut (.I0(\PID_CONTROLLER.integral [8]), .I1(IntegralLimit[8]), 
            .I2(GND_net), .I3(GND_net), .O(n17_adj_3941));   // verilog/motorControl.v(40[10:34])
    defparam LessThan_4_i17_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i29874_4_lut (.I0(\PID_CONTROLLER.integral [9]), .I1(n17_adj_3941), 
            .I2(IntegralLimit[9]), .I3(n9_adj_3940), .O(n45395));
    defparam i29874_4_lut.LUT_INIT = 16'hffde;
    SB_LUT4 i29872_4_lut (.I0(\PID_CONTROLLER.integral [9]), .I1(IntegralLimit[10]), 
            .I2(IntegralLimit[11]), .I3(n45395), .O(n45393));
    defparam i29872_4_lut.LUT_INIT = 16'h7eff;
    SB_LUT4 i29224_4_lut (.I0(n11_adj_3648), .I1(n9_adj_3650), .I2(n7_adj_3652), 
            .I3(n5_adj_3654), .O(n44745));
    defparam i29224_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 LessThan_4_i13_rep_450_2_lut (.I0(\PID_CONTROLLER.integral [6]), 
            .I1(IntegralLimit[6]), .I2(GND_net), .I3(GND_net), .O(n47477));   // verilog/motorControl.v(40[10:34])
    defparam LessThan_4_i13_rep_450_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i29878_4_lut (.I0(\PID_CONTROLLER.integral [7]), .I1(n47477), 
            .I2(IntegralLimit[7]), .I3(n11_adj_3939), .O(n45399));
    defparam i29878_4_lut.LUT_INIT = 16'hffde;
    SB_LUT4 i29866_4_lut (.I0(\PID_CONTROLLER.integral [9]), .I1(IntegralLimit[13]), 
            .I2(IntegralLimit[14]), .I3(n45399), .O(n45387));
    defparam i29866_4_lut.LUT_INIT = 16'h7eff;
    SB_LUT4 i29266_4_lut (.I0(\PID_CONTROLLER.integral [9]), .I1(\PID_CONTROLLER.integral [7]), 
            .I2(IntegralLimit[16]), .I3(IntegralLimit[7]), .O(n44787));
    defparam i29266_4_lut.LUT_INIT = 16'h7bde;
    SB_LUT4 LessThan_4_i35_rep_438_2_lut (.I0(\PID_CONTROLLER.integral [9]), 
            .I1(IntegralLimit[17]), .I2(GND_net), .I3(GND_net), .O(n47465));   // verilog/motorControl.v(40[10:34])
    defparam LessThan_4_i35_rep_438_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_4_i10_3_lut (.I0(IntegralLimit[5]), .I1(IntegralLimit[6]), 
            .I2(\PID_CONTROLLER.integral [6]), .I3(GND_net), .O(n10_adj_3942));   // verilog/motorControl.v(40[10:34])
    defparam LessThan_4_i10_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 LessThan_4_i30_4_lut (.I0(IntegralLimit[7]), .I1(IntegralLimit[17]), 
            .I2(\PID_CONTROLLER.integral [9]), .I3(IntegralLimit[16]), .O(n30_adj_3943));   // verilog/motorControl.v(40[10:34])
    defparam LessThan_4_i30_4_lut.LUT_INIT = 16'h8f0e;
    SB_LUT4 LessThan_4_i5_2_lut (.I0(\PID_CONTROLLER.integral [2]), .I1(IntegralLimit[2]), 
            .I2(GND_net), .I3(GND_net), .O(n5_adj_3944));   // verilog/motorControl.v(40[10:34])
    defparam LessThan_4_i5_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i29882_4_lut (.I0(n9_adj_3940), .I1(\PID_CONTROLLER.integral [3]), 
            .I2(n5_adj_3944), .I3(IntegralLimit[3]), .O(n45403));
    defparam i29882_4_lut.LUT_INIT = 16'hfbfe;
    SB_LUT4 i29880_4_lut (.I0(\PID_CONTROLLER.integral [6]), .I1(n11_adj_3939), 
            .I2(IntegralLimit[6]), .I3(n45403), .O(n45401));
    defparam i29880_4_lut.LUT_INIT = 16'hdeff;
    SB_LUT4 i29290_4_lut (.I0(n17_adj_3941), .I1(\PID_CONTROLLER.integral [7]), 
            .I2(n45401), .I3(IntegralLimit[7]), .O(n44811));
    defparam i29290_4_lut.LUT_INIT = 16'haeab;
    SB_LUT4 i30099_4_lut (.I0(\PID_CONTROLLER.integral [9]), .I1(IntegralLimit[9]), 
            .I2(IntegralLimit[10]), .I3(n44811), .O(n45620));
    defparam i30099_4_lut.LUT_INIT = 16'hff7e;
    SB_LUT4 i30485_4_lut (.I0(\PID_CONTROLLER.integral [9]), .I1(IntegralLimit[11]), 
            .I2(IntegralLimit[12]), .I3(n45620), .O(n46006));
    defparam i30485_4_lut.LUT_INIT = 16'hff7e;
    SB_LUT4 i29868_4_lut (.I0(\PID_CONTROLLER.integral [9]), .I1(IntegralLimit[13]), 
            .I2(IntegralLimit[14]), .I3(n46006), .O(n45389));
    defparam i29868_4_lut.LUT_INIT = 16'h7eff;
    SB_LUT4 i30319_4_lut (.I0(\PID_CONTROLLER.integral [9]), .I1(IntegralLimit[15]), 
            .I2(IntegralLimit[16]), .I3(n45389), .O(n45840));
    defparam i30319_4_lut.LUT_INIT = 16'hff7e;
    SB_LUT4 i30558_4_lut (.I0(\PID_CONTROLLER.integral [9]), .I1(IntegralLimit[17]), 
            .I2(IntegralLimit[18]), .I3(n45840), .O(n46079));
    defparam i30558_4_lut.LUT_INIT = 16'hff7e;
    SB_LUT4 i30661_4_lut (.I0(\PID_CONTROLLER.integral [9]), .I1(IntegralLimit[19]), 
            .I2(IntegralLimit[20]), .I3(n46079), .O(n46182));
    defparam i30661_4_lut.LUT_INIT = 16'hff7e;
    SB_LUT4 LessThan_4_i6_3_lut (.I0(IntegralLimit[2]), .I1(IntegralLimit[3]), 
            .I2(\PID_CONTROLLER.integral [3]), .I3(GND_net), .O(n6_adj_3945));   // verilog/motorControl.v(40[10:34])
    defparam LessThan_4_i6_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i29367_4_lut (.I0(\PID_CONTROLLER.integral [9]), .I1(IntegralLimit[21]), 
            .I2(IntegralLimit[22]), .I3(IntegralLimit[9]), .O(n44888));
    defparam i29367_4_lut.LUT_INIT = 16'h7ffe;
    SB_LUT4 LessThan_4_i24_4_lut (.I0(IntegralLimit[9]), .I1(IntegralLimit[22]), 
            .I2(\PID_CONTROLLER.integral [9]), .I3(IntegralLimit[21]), .O(n24_adj_3946));   // verilog/motorControl.v(40[10:34])
    defparam LessThan_4_i24_4_lut.LUT_INIT = 16'h8f0e;
    SB_LUT4 i30177_3_lut (.I0(n6_adj_3945), .I1(IntegralLimit[10]), .I2(\PID_CONTROLLER.integral [9]), 
            .I3(GND_net), .O(n45698));   // verilog/motorControl.v(40[10:34])
    defparam i30177_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i29242_4_lut (.I0(\PID_CONTROLLER.integral [9]), .I1(IntegralLimit[12]), 
            .I2(IntegralLimit[21]), .I3(n45393), .O(n44763));
    defparam i29242_4_lut.LUT_INIT = 16'h5adb;
    SB_LUT4 LessThan_4_i45_rep_403_2_lut (.I0(\PID_CONTROLLER.integral [9]), 
            .I1(IntegralLimit[22]), .I2(GND_net), .I3(GND_net), .O(n47430));   // verilog/motorControl.v(40[10:34])
    defparam LessThan_4_i45_rep_403_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i30179_3_lut (.I0(n24_adj_3946), .I1(n8_adj_3947), .I2(n44888), 
            .I3(GND_net), .O(n45700));   // verilog/motorControl.v(40[10:34])
    defparam i30179_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i29543_4_lut (.I0(n45698), .I1(IntegralLimit[12]), .I2(\PID_CONTROLLER.integral [9]), 
            .I3(IntegralLimit[11]), .O(n45064));   // verilog/motorControl.v(40[10:34])
    defparam i29543_4_lut.LUT_INIT = 16'h8f0e;
    SB_LUT4 LessThan_6_i4_4_lut (.I0(n76[0]), .I1(\PID_CONTROLLER.integral [1]), 
            .I2(n3_adj_3658), .I3(\PID_CONTROLLER.integral [0]), .O(n4_adj_3948));   // verilog/motorControl.v(40[38:63])
    defparam LessThan_6_i4_4_lut.LUT_INIT = 16'hc5c0;
    SB_LUT4 i30151_3_lut (.I0(n4_adj_3948), .I1(\PID_CONTROLLER.integral [5]), 
            .I2(n11_adj_3648), .I3(GND_net), .O(n45672));   // verilog/motorControl.v(40[38:63])
    defparam i30151_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i30152_3_lut (.I0(n45672), .I1(\PID_CONTROLLER.integral [6]), 
            .I2(n13_adj_3646), .I3(GND_net), .O(n45673));   // verilog/motorControl.v(40[38:63])
    defparam i30152_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_6_i8_3_lut (.I0(\PID_CONTROLLER.integral [4]), .I1(\PID_CONTROLLER.integral [8]), 
            .I2(n17_adj_3638), .I3(GND_net), .O(n8_adj_3949));   // verilog/motorControl.v(40[38:63])
    defparam LessThan_6_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i29214_2_lut (.I0(n17_adj_3638), .I1(n9_adj_3650), .I2(GND_net), 
            .I3(GND_net), .O(n44735));
    defparam i29214_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 LessThan_6_i6_3_lut (.I0(\PID_CONTROLLER.integral [2]), .I1(\PID_CONTROLLER.integral [3]), 
            .I2(n7_adj_3652), .I3(GND_net), .O(n6_adj_3950));   // verilog/motorControl.v(40[38:63])
    defparam LessThan_6_i6_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_6_i16_3_lut (.I0(n8_adj_3949), .I1(\PID_CONTROLLER.integral [9]), 
            .I2(n41724), .I3(GND_net), .O(n16_adj_3951));   // verilog/motorControl.v(40[38:63])
    defparam LessThan_6_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i29218_4_lut (.I0(n17_adj_3638), .I1(n15_adj_3644), .I2(n13_adj_3646), 
            .I3(n44745), .O(n44739));
    defparam i29218_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i30277_4_lut (.I0(n16_adj_3951), .I1(n6_adj_3950), .I2(n41724), 
            .I3(n44735), .O(n45798));   // verilog/motorControl.v(40[38:63])
    defparam i30277_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i29553_3_lut (.I0(n45673), .I1(\PID_CONTROLLER.integral [7]), 
            .I2(n15_adj_3644), .I3(GND_net), .O(n45074));   // verilog/motorControl.v(40[38:63])
    defparam i29553_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i30535_4_lut (.I0(n45074), .I1(n45798), .I2(n41724), .I3(n44739), 
            .O(n46056));   // verilog/motorControl.v(40[38:63])
    defparam i30535_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 LessThan_4_i4_4_lut (.I0(\PID_CONTROLLER.integral [0]), .I1(IntegralLimit[1]), 
            .I2(\PID_CONTROLLER.integral [1]), .I3(IntegralLimit[0]), .O(n4_adj_3952));   // verilog/motorControl.v(40[10:34])
    defparam LessThan_4_i4_4_lut.LUT_INIT = 16'h4d0c;
    SB_LUT4 i30157_3_lut (.I0(n4_adj_3952), .I1(IntegralLimit[13]), .I2(\PID_CONTROLLER.integral [9]), 
            .I3(GND_net), .O(n45678));   // verilog/motorControl.v(40[10:34])
    defparam i30157_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i29268_4_lut (.I0(\PID_CONTROLLER.integral [9]), .I1(IntegralLimit[15]), 
            .I2(IntegralLimit[16]), .I3(n45387), .O(n44789));
    defparam i29268_4_lut.LUT_INIT = 16'h5adb;
    SB_LUT4 i30511_4_lut (.I0(n30_adj_3943), .I1(n10_adj_3942), .I2(n47465), 
            .I3(n44787), .O(n46032));   // verilog/motorControl.v(40[10:34])
    defparam i30511_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i29545_4_lut (.I0(n45678), .I1(IntegralLimit[15]), .I2(\PID_CONTROLLER.integral [9]), 
            .I3(IntegralLimit[14]), .O(n45066));   // verilog/motorControl.v(40[10:34])
    defparam i29545_4_lut.LUT_INIT = 16'h8f0e;
    SB_LUT4 i30639_4_lut (.I0(n45066), .I1(n46032), .I2(n47465), .I3(n44789), 
            .O(n46160));   // verilog/motorControl.v(40[10:34])
    defparam i30639_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i30640_3_lut (.I0(n46160), .I1(IntegralLimit[18]), .I2(\PID_CONTROLLER.integral [9]), 
            .I3(GND_net), .O(n46161));   // verilog/motorControl.v(40[10:34])
    defparam i30640_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i29844_4_lut (.I0(\PID_CONTROLLER.integral [9]), .I1(IntegralLimit[21]), 
            .I2(IntegralLimit[22]), .I3(n46182), .O(n45365));
    defparam i29844_4_lut.LUT_INIT = 16'h7eff;
    SB_LUT4 i30415_4_lut (.I0(n45064), .I1(n45700), .I2(n47430), .I3(n44763), 
            .O(n45936));   // verilog/motorControl.v(40[10:34])
    defparam i30415_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i29551_4_lut (.I0(n46161), .I1(IntegralLimit[20]), .I2(\PID_CONTROLLER.integral [9]), 
            .I3(IntegralLimit[19]), .O(n45072));   // verilog/motorControl.v(40[10:34])
    defparam i29551_4_lut.LUT_INIT = 16'h8f0e;
    SB_LUT4 i30536_3_lut (.I0(n46056), .I1(n76[23]), .I2(\PID_CONTROLLER.integral [9]), 
            .I3(GND_net), .O(n46057));   // verilog/motorControl.v(40[38:63])
    defparam i30536_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i30533_3_lut (.I0(n45072), .I1(n45936), .I2(n45365), .I3(GND_net), 
            .O(n46054));   // verilog/motorControl.v(40[10:34])
    defparam i30533_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8_4_lut_adj_1444 (.I0(n46054), .I1(n46057), .I2(\PID_CONTROLLER.integral [9]), 
            .I3(IntegralLimit[23]), .O(n55_adj_3594));   // verilog/motorControl.v(40[10:63])
    defparam i8_4_lut_adj_1444.LUT_INIT = 16'h80c8;
    SB_LUT4 unary_minus_5_inv_0_i21_1_lut (.I0(IntegralLimit[20]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n79[20]));   // verilog/motorControl.v(40[48:62])
    defparam unary_minus_5_inv_0_i21_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_12_i164_2_lut (.I0(\Kd[2] ), .I1(n57[16]), .I2(GND_net), 
            .I3(GND_net), .O(n243_adj_3590));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i164_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i229_2_lut (.I0(\Kd[3] ), .I1(n57[16]), .I2(GND_net), 
            .I3(GND_net), .O(n340));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i229_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i418_2_lut (.I0(\Kd[6] ), .I1(n57[13]), .I2(GND_net), 
            .I3(GND_net), .O(n622));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i418_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i109_2_lut (.I0(\Kd[1] ), .I1(n57[21]), .I2(GND_net), 
            .I3(GND_net), .O(n161_adj_3589));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i109_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i46_2_lut (.I0(\Kd[0] ), .I1(n57[22]), .I2(GND_net), 
            .I3(GND_net), .O(n68_adj_3588));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i46_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i174_2_lut (.I0(\Kd[2] ), .I1(n57[21]), .I2(GND_net), 
            .I3(GND_net), .O(n258_adj_3587));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i174_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i239_2_lut (.I0(\Kd[3] ), .I1(n57[21]), .I2(GND_net), 
            .I3(GND_net), .O(n355_adj_3586));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i239_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i304_2_lut (.I0(\Kd[4] ), .I1(n57[21]), .I2(GND_net), 
            .I3(GND_net), .O(n452_adj_3585));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i304_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i369_2_lut (.I0(\Kd[5] ), .I1(n57[21]), .I2(GND_net), 
            .I3(GND_net), .O(n549_adj_3584));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i369_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i434_2_lut (.I0(\Kd[6] ), .I1(n57[21]), .I2(GND_net), 
            .I3(GND_net), .O(n646_adj_3583));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i434_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i499_2_lut (.I0(\Kd[7] ), .I1(n57[21]), .I2(GND_net), 
            .I3(GND_net), .O(n743_adj_3582));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i499_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i294_2_lut (.I0(\Kd[4] ), .I1(n57[16]), .I2(GND_net), 
            .I3(GND_net), .O(n437_adj_3581));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i294_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_14_i67_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral [8]), 
            .I2(GND_net), .I3(GND_net), .O(n98_adj_3580));   // verilog/motorControl.v(43[48:59])
    defparam mult_14_i67_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_14_i116_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral [8]), 
            .I2(GND_net), .I3(GND_net), .O(n171_adj_3579));   // verilog/motorControl.v(43[48:59])
    defparam mult_14_i116_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_inv_0_i22_1_lut (.I0(IntegralLimit[21]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n79[21]));   // verilog/motorControl.v(40[48:62])
    defparam unary_minus_5_inv_0_i22_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_5_inv_0_i23_1_lut (.I0(IntegralLimit[22]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n79[22]));   // verilog/motorControl.v(40[48:62])
    defparam unary_minus_5_inv_0_i23_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_5_inv_0_i24_1_lut (.I0(IntegralLimit[23]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n79[23]));   // verilog/motorControl.v(40[48:62])
    defparam unary_minus_5_inv_0_i24_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_14_i165_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral [8]), 
            .I2(GND_net), .I3(GND_net), .O(n244_adj_3571));   // verilog/motorControl.v(43[48:59])
    defparam mult_14_i165_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_21_inv_0_i1_1_lut (.I0(\PWMLimit[0] ), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n75[0]));   // verilog/motorControl.v(47[28:37])
    defparam unary_minus_21_inv_0_i1_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_14_i214_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral [8]), 
            .I2(GND_net), .I3(GND_net), .O(n317));   // verilog/motorControl.v(43[48:59])
    defparam mult_14_i214_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i111_2_lut (.I0(\Kd[1] ), .I1(n57[22]), .I2(GND_net), 
            .I3(GND_net), .O(n164_adj_3568));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i111_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i48_2_lut (.I0(\Kd[0] ), .I1(n57[23]), .I2(GND_net), 
            .I3(GND_net), .O(n71_adj_3567));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i48_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i284_2_lut (.I0(\Kd[4] ), .I1(n57[11]), .I2(GND_net), 
            .I3(GND_net), .O(n422_adj_3566));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i284_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i359_2_lut (.I0(\Kd[5] ), .I1(n57[16]), .I2(GND_net), 
            .I3(GND_net), .O(n534));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i359_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_14_i263_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral [8]), 
            .I2(GND_net), .I3(GND_net), .O(n390));   // verilog/motorControl.v(43[48:59])
    defparam mult_14_i263_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_14_i312_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral [8]), 
            .I2(GND_net), .I3(GND_net), .O(n463_c));   // verilog/motorControl.v(43[48:59])
    defparam mult_14_i312_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_14_i361_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral [8]), 
            .I2(GND_net), .I3(GND_net), .O(n536));   // verilog/motorControl.v(43[48:59])
    defparam mult_14_i361_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i85_2_lut (.I0(\Kd[1] ), .I1(n57[9]), .I2(GND_net), 
            .I3(GND_net), .O(n125));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i85_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i22_2_lut (.I0(\Kd[0] ), .I1(n57[10]), .I2(GND_net), 
            .I3(GND_net), .O(n32_adj_3562));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i22_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_21_inv_0_i2_1_lut (.I0(\PWMLimit[1] ), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n75[1]));   // verilog/motorControl.v(47[28:37])
    defparam unary_minus_21_inv_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_12_i150_2_lut (.I0(\Kd[2] ), .I1(n57[9]), .I2(GND_net), 
            .I3(GND_net), .O(n222_adj_3558));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i150_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i424_2_lut (.I0(\Kd[6] ), .I1(n57[16]), .I2(GND_net), 
            .I3(GND_net), .O(n631));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i424_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_21_inv_0_i3_1_lut (.I0(\PWMLimit[2] ), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n75[2]));   // verilog/motorControl.v(47[28:37])
    defparam unary_minus_21_inv_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_12_i176_2_lut (.I0(\Kd[2] ), .I1(n57[22]), .I2(GND_net), 
            .I3(GND_net), .O(n261_adj_3556));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i176_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_21_inv_0_i4_1_lut (.I0(\PWMLimit[3] ), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n75[3]));   // verilog/motorControl.v(47[28:37])
    defparam unary_minus_21_inv_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_21_inv_0_i5_1_lut (.I0(\PWMLimit[4] ), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n75[4]));   // verilog/motorControl.v(47[28:37])
    defparam unary_minus_21_inv_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_12_i349_2_lut (.I0(\Kd[5] ), .I1(n57[11]), .I2(GND_net), 
            .I3(GND_net), .O(n519_adj_3551));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i349_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i483_2_lut (.I0(\Kd[7] ), .I1(n57[13]), .I2(GND_net), 
            .I3(GND_net), .O(n719));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i483_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i241_2_lut (.I0(\Kd[3] ), .I1(n57[22]), .I2(GND_net), 
            .I3(GND_net), .O(n358_adj_3550));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i241_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i306_2_lut (.I0(\Kd[4] ), .I1(n57[22]), .I2(GND_net), 
            .I3(GND_net), .O(n455_adj_3549));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i306_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i489_2_lut (.I0(\Kd[7] ), .I1(n57[16]), .I2(GND_net), 
            .I3(GND_net), .O(n728));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i489_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i371_2_lut (.I0(\Kd[5] ), .I1(n57[22]), .I2(GND_net), 
            .I3(GND_net), .O(n552_adj_3548));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i371_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i414_2_lut (.I0(\Kd[6] ), .I1(n57[11]), .I2(GND_net), 
            .I3(GND_net), .O(n616_adj_3547));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i414_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_21_inv_0_i6_1_lut (.I0(\PWMLimit[5] ), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n75[5]));   // verilog/motorControl.v(47[28:37])
    defparam unary_minus_21_inv_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_21_inv_0_i7_1_lut (.I0(\PWMLimit[6] ), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n75[6]));   // verilog/motorControl.v(47[28:37])
    defparam unary_minus_21_inv_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 LessThan_4_i8_3_lut_3_lut (.I0(IntegralLimit[4]), .I1(IntegralLimit[8]), 
            .I2(\PID_CONTROLLER.integral [8]), .I3(GND_net), .O(n8_adj_3947));   // verilog/motorControl.v(40[10:34])
    defparam LessThan_4_i8_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i20400_3_lut_4_lut (.I0(n10111[2]), .I1(\Kd[4] ), .I2(n57[25]), 
            .I3(n6_adj_3953), .O(n8_adj_3933));   // verilog/motorControl.v(43[26:45])
    defparam i20400_3_lut_4_lut.LUT_INIT = 16'hea80;
    SB_LUT4 i2_3_lut_4_lut (.I0(\Kd[5] ), .I1(n57[25]), .I2(\Kd[4] ), 
            .I3(n6_adj_3953), .O(n8_adj_3934));   // verilog/motorControl.v(43[26:45])
    defparam i2_3_lut_4_lut.LUT_INIT = 16'hb748;
    SB_LUT4 i20392_3_lut_4_lut (.I0(n10111[1]), .I1(\Kd[3] ), .I2(n57[25]), 
            .I3(n4_adj_3856), .O(n6_adj_3953));   // verilog/motorControl.v(43[26:45])
    defparam i20392_3_lut_4_lut.LUT_INIT = 16'hea80;
    SB_LUT4 i20296_2_lut_3_lut (.I0(\Kd[0] ), .I1(n57[25]), .I2(\Kd[1] ), 
            .I3(GND_net), .O(n33897));   // verilog/motorControl.v(43[26:45])
    defparam i20296_2_lut_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 i1_3_lut_4_lut_adj_1445 (.I0(n10111[2]), .I1(\Kd[4] ), .I2(n57[25]), 
            .I3(n6_adj_3953), .O(n10111[3]));   // verilog/motorControl.v(43[26:45])
    defparam i1_3_lut_4_lut_adj_1445.LUT_INIT = 16'h956a;
    SB_LUT4 mult_12_i436_2_lut (.I0(\Kd[6] ), .I1(n57[22]), .I2(GND_net), 
            .I3(GND_net), .O(n649_adj_3544));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i436_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i215_2_lut (.I0(\Kd[3] ), .I1(n57[9]), .I2(GND_net), 
            .I3(GND_net), .O(n319));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i215_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i501_2_lut (.I0(\Kd[7] ), .I1(n57[22]), .I2(GND_net), 
            .I3(GND_net), .O(n746_adj_3543));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i501_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i29069_2_lut_4_lut (.I0(\PID_CONTROLLER.result [8]), .I1(pwm_23__N_2960[8]), 
            .I2(\PID_CONTROLLER.result [4]), .I3(pwm_23__N_2960[4]), .O(n44590));
    defparam i29069_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 i1_2_lut_4_lut (.I0(\PID_CONTROLLER.result [28]), .I1(\PID_CONTROLLER.result [30]), 
            .I2(\PID_CONTROLLER.result [29]), .I3(n56_adj_3914), .O(n40126));   // verilog/motorControl.v(45[12:27])
    defparam i1_2_lut_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 mult_12_i113_2_lut (.I0(\Kd[1] ), .I1(n57[23]), .I2(GND_net), 
            .I3(GND_net), .O(n167_adj_3542));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i113_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i50_2_lut (.I0(\Kd[0] ), .I1(n57[24]), .I2(GND_net), 
            .I3(GND_net), .O(n74));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i50_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i28843_2_lut_4_lut (.I0(hall2), .I1(GATES_5__N_3048[5]), .I2(hall3), 
            .I3(n878), .O(n44119));   // verilog/motorControl.v(86[14] 109[8])
    defparam i28843_2_lut_4_lut.LUT_INIT = 16'h0200;
    SB_LUT4 \PID_CONTROLLER.result_31__I_0_i8_3_lut_3_lut  (.I0(\PID_CONTROLLER.result [4]), 
            .I1(\PID_CONTROLLER.result [8]), .I2(\deadband[8] ), .I3(GND_net), 
            .O(n8_adj_3888));   // verilog/motorControl.v(44[10:27])
    defparam \PID_CONTROLLER.result_31__I_0_i8_3_lut_3_lut .LUT_INIT = 16'h8e8e;
    SB_LUT4 \PID_CONTROLLER.result_31__I_0_i6_3_lut_3_lut  (.I0(\PID_CONTROLLER.result [2]), 
            .I1(\PID_CONTROLLER.result [3]), .I2(\deadband[3] ), .I3(GND_net), 
            .O(n6_adj_3886));   // verilog/motorControl.v(44[10:27])
    defparam \PID_CONTROLLER.result_31__I_0_i6_3_lut_3_lut .LUT_INIT = 16'h8e8e;
    SB_LUT4 \PID_CONTROLLER.result_31__I_0_i10_3_lut_3_lut  (.I0(\PID_CONTROLLER.result[5] ), 
            .I1(\PID_CONTROLLER.result[6] ), .I2(\deadband[6] ), .I3(GND_net), 
            .O(n10_adj_3890));   // verilog/motorControl.v(44[10:27])
    defparam \PID_CONTROLLER.result_31__I_0_i10_3_lut_3_lut .LUT_INIT = 16'h8e8e;
    SB_LUT4 mult_12_i178_2_lut (.I0(\Kd[2] ), .I1(n57[23]), .I2(GND_net), 
            .I3(GND_net), .O(n264));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i178_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i243_2_lut (.I0(\Kd[3] ), .I1(n57[23]), .I2(GND_net), 
            .I3(GND_net), .O(n361));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i243_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_21_inv_0_i8_1_lut (.I0(\PWMLimit[7] ), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n75[7]));   // verilog/motorControl.v(47[28:37])
    defparam unary_minus_21_inv_0_i8_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1_2_lut_3_lut_4_lut (.I0(\Kd[3] ), .I1(n57[25]), .I2(n4_adj_3856), 
            .I3(n10111[1]), .O(n10111[2]));   // verilog/motorControl.v(43[26:45])
    defparam i1_2_lut_3_lut_4_lut.LUT_INIT = 16'h8778;
    SB_LUT4 i20093_3_lut_4_lut (.I0(n16637[2]), .I1(\Kp[4] ), .I2(\PID_CONTROLLER.err[31] ), 
            .I3(n6_adj_3954), .O(n8_adj_3852));   // verilog/motorControl.v(43[17:23])
    defparam i20093_3_lut_4_lut.LUT_INIT = 16'hea80;
    SB_LUT4 i2_3_lut_4_lut_adj_1446 (.I0(\Kp[5] ), .I1(\PID_CONTROLLER.err[31] ), 
            .I2(\Kp[4] ), .I3(n6_adj_3954), .O(n8_adj_3853));   // verilog/motorControl.v(43[17:23])
    defparam i2_3_lut_4_lut_adj_1446.LUT_INIT = 16'hb748;
    SB_LUT4 i20085_3_lut_4_lut (.I0(n16644[1]), .I1(\Kp[3] ), .I2(\PID_CONTROLLER.err[31] ), 
            .I3(n4_adj_3955), .O(n6_adj_3954));   // verilog/motorControl.v(43[17:23])
    defparam i20085_3_lut_4_lut.LUT_INIT = 16'hea80;
    SB_LUT4 i20244_4_lut_4_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err[31] ), 
            .I2(n16637[0]), .I3(n33546), .O(n4_adj_3955));   // verilog/motorControl.v(43[17:23])
    defparam i20244_4_lut_4_lut.LUT_INIT = 16'hf8a0;
    SB_LUT4 i20232_2_lut_3_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err[31] ), 
            .I2(\Kp[1] ), .I3(GND_net), .O(n33546));   // verilog/motorControl.v(43[17:23])
    defparam i20232_2_lut_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 i1_3_lut_4_lut_adj_1447 (.I0(n16637[2]), .I1(\Kp[4] ), .I2(\PID_CONTROLLER.err[31] ), 
            .I3(n6_adj_3954), .O(n16637[3]));   // verilog/motorControl.v(43[17:23])
    defparam i1_3_lut_4_lut_adj_1447.LUT_INIT = 16'h956a;
    SB_LUT4 mult_12_i308_2_lut (.I0(\Kd[4] ), .I1(n57[23]), .I2(GND_net), 
            .I3(GND_net), .O(n458_c));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i308_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i373_2_lut (.I0(\Kd[5] ), .I1(n57[23]), .I2(GND_net), 
            .I3(GND_net), .O(n555));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i373_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_21_inv_0_i9_1_lut (.I0(\PWMLimit[8] ), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n75[8]));   // verilog/motorControl.v(47[28:37])
    defparam unary_minus_21_inv_0_i9_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i71_2_lut (.I0(\Kp[1] ), .I1(\PID_CONTROLLER.err[2] ), 
            .I2(GND_net), .I3(GND_net), .O(n104_adj_3538));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i71_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i8_2_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err[3] ), 
            .I2(GND_net), .I3(GND_net), .O(n11_adj_3537));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i8_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_21_inv_0_i32_1_lut (.I0(\PWMLimit[9] ), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_3536));   // verilog/motorControl.v(47[28:37])
    defparam unary_minus_21_inv_0_i32_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i12058_1_lut (.I0(pwm_count[0]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n25474));   // verilog/motorControl.v(110[18:29])
    defparam i12058_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_70_inv_0_i1_1_lut (.I0(pwm[0]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n73[0]));   // verilog/motorControl.v(86[38:44])
    defparam unary_minus_70_inv_0_i1_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_70_inv_0_i2_1_lut (.I0(pwm[1]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n73[1]));   // verilog/motorControl.v(86[38:44])
    defparam unary_minus_70_inv_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i136_2_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err[2] ), 
            .I2(GND_net), .I3(GND_net), .O(n201_adj_3533));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i136_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i67_2_lut (.I0(\Kd[1] ), .I1(n57[0]), .I2(GND_net), 
            .I3(GND_net), .O(n98_adj_3532));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i67_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i4_2_lut (.I0(\Kd[0] ), .I1(n57[1]), .I2(GND_net), 
            .I3(GND_net), .O(n5_adj_3531));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i4_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i479_2_lut (.I0(\Kd[7] ), .I1(n57[11]), .I2(GND_net), 
            .I3(GND_net), .O(n713_adj_3529));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i479_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i438_2_lut (.I0(\Kd[6] ), .I1(n57[23]), .I2(GND_net), 
            .I3(GND_net), .O(n652));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i438_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_70_inv_0_i3_1_lut (.I0(pwm[2]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n73[2]));   // verilog/motorControl.v(86[38:44])
    defparam unary_minus_70_inv_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_70_inv_0_i4_1_lut (.I0(pwm[3]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n73[3]));   // verilog/motorControl.v(86[38:44])
    defparam unary_minus_70_inv_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i201_2_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err[2] ), 
            .I2(GND_net), .I3(GND_net), .O(n298_adj_3526));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i201_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i132_2_lut (.I0(\Kd[2] ), .I1(n57[0]), .I2(GND_net), 
            .I3(GND_net), .O(n195_adj_3525));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i132_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_70_inv_0_i5_1_lut (.I0(pwm[4]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n73[4]));   // verilog/motorControl.v(86[38:44])
    defparam unary_minus_70_inv_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_70_inv_0_i6_1_lut (.I0(pwm[5]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n73[5]));   // verilog/motorControl.v(86[38:44])
    defparam unary_minus_70_inv_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_70_inv_0_i7_1_lut (.I0(pwm[6]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n73[6]));   // verilog/motorControl.v(86[38:44])
    defparam unary_minus_70_inv_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_12_i503_2_lut (.I0(\Kd[7] ), .I1(n57[23]), .I2(GND_net), 
            .I3(GND_net), .O(n749));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i503_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i115_2_lut (.I0(\Kd[1] ), .I1(n57[24]), .I2(GND_net), 
            .I3(GND_net), .O(n170_adj_3521));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i115_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i52_2_lut (.I0(\Kd[0] ), .I1(n57[25]), .I2(GND_net), 
            .I3(GND_net), .O(n86));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i52_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i266_2_lut (.I0(\Kp[4] ), .I1(\PID_CONTROLLER.err[2] ), 
            .I2(GND_net), .I3(GND_net), .O(n395_adj_3520));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i266_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_70_inv_0_i8_1_lut (.I0(pwm[7]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n73[7]));   // verilog/motorControl.v(86[38:44])
    defparam unary_minus_70_inv_0_i8_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_70_inv_0_i9_1_lut (.I0(pwm[8]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n73[8]));   // verilog/motorControl.v(86[38:44])
    defparam unary_minus_70_inv_0_i9_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_70_inv_0_i10_1_lut (.I0(pwm[9]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n73[9]));   // verilog/motorControl.v(86[38:44])
    defparam unary_minus_70_inv_0_i10_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_70_inv_0_i11_1_lut (.I0(pwm[10]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n73[10]));   // verilog/motorControl.v(86[38:44])
    defparam unary_minus_70_inv_0_i11_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i331_2_lut (.I0(\Kp[5] ), .I1(\PID_CONTROLLER.err[2] ), 
            .I2(GND_net), .I3(GND_net), .O(n492_adj_3515));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i331_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_70_inv_0_i12_1_lut (.I0(pwm[11]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n73[11]));   // verilog/motorControl.v(86[38:44])
    defparam unary_minus_70_inv_0_i12_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i396_2_lut (.I0(\Kp[6] ), .I1(\PID_CONTROLLER.err[2] ), 
            .I2(GND_net), .I3(GND_net), .O(n589_adj_3513));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i396_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i197_2_lut (.I0(\Kd[3] ), .I1(n57[0]), .I2(GND_net), 
            .I3(GND_net), .O(n292_adj_3512));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i197_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i79_2_lut (.I0(\Kd[1] ), .I1(n57[6]), .I2(GND_net), 
            .I3(GND_net), .O(n116_adj_3511));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i79_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i16_2_lut (.I0(\Kd[0] ), .I1(n57[7]), .I2(GND_net), 
            .I3(GND_net), .O(n23_adj_3510));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i16_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_70_inv_0_i13_1_lut (.I0(pwm[12]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n73[12]));   // verilog/motorControl.v(86[38:44])
    defparam unary_minus_70_inv_0_i13_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_70_inv_0_i14_1_lut (.I0(pwm[13]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n73[13]));   // verilog/motorControl.v(86[38:44])
    defparam unary_minus_70_inv_0_i14_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_12_i180_2_lut (.I0(\Kd[2] ), .I1(n57[24]), .I2(GND_net), 
            .I3(GND_net), .O(n267));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i180_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i245_2_lut (.I0(\Kd[3] ), .I1(n57[24]), .I2(GND_net), 
            .I3(GND_net), .O(n364_adj_3507));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i245_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i461_2_lut (.I0(\Kp[7] ), .I1(\PID_CONTROLLER.err[2] ), 
            .I2(GND_net), .I3(GND_net), .O(n686_adj_3506));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i461_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_70_inv_0_i15_1_lut (.I0(pwm[14]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n73[14]));   // verilog/motorControl.v(86[38:44])
    defparam unary_minus_70_inv_0_i15_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_12_i262_2_lut (.I0(\Kd[4] ), .I1(n57[0]), .I2(GND_net), 
            .I3(GND_net), .O(n389_adj_3504));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i262_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i280_2_lut (.I0(\Kd[4] ), .I1(n57[9]), .I2(GND_net), 
            .I3(GND_net), .O(n416));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i280_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_70_inv_0_i16_1_lut (.I0(pwm[15]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n73[15]));   // verilog/motorControl.v(86[38:44])
    defparam unary_minus_70_inv_0_i16_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_70_inv_0_i17_1_lut (.I0(pwm[16]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n73[16]));   // verilog/motorControl.v(86[38:44])
    defparam unary_minus_70_inv_0_i17_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_12_i144_2_lut (.I0(\Kd[2] ), .I1(n57[6]), .I2(GND_net), 
            .I3(GND_net), .O(n213_adj_3502));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i144_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_70_inv_0_i18_1_lut (.I0(pwm[17]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n73[17]));   // verilog/motorControl.v(86[38:44])
    defparam unary_minus_70_inv_0_i18_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_70_inv_0_i19_1_lut (.I0(pwm[18]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n73[18]));   // verilog/motorControl.v(86[38:44])
    defparam unary_minus_70_inv_0_i19_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_70_inv_0_i20_1_lut (.I0(pwm[19]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n73[19]));   // verilog/motorControl.v(86[38:44])
    defparam unary_minus_70_inv_0_i20_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_12_i310_2_lut (.I0(\Kd[4] ), .I1(n57[24]), .I2(GND_net), 
            .I3(GND_net), .O(n461_c));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i310_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i375_2_lut (.I0(\Kd[5] ), .I1(n57[24]), .I2(GND_net), 
            .I3(GND_net), .O(n558));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i375_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_70_inv_0_i21_1_lut (.I0(pwm[20]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n73[20]));   // verilog/motorControl.v(86[38:44])
    defparam unary_minus_70_inv_0_i21_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_12_i327_2_lut (.I0(\Kd[5] ), .I1(n57[0]), .I2(GND_net), 
            .I3(GND_net), .O(n486_adj_3497));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i327_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_70_inv_0_i22_1_lut (.I0(pwm[21]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n73[21]));   // verilog/motorControl.v(86[38:44])
    defparam unary_minus_70_inv_0_i22_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i111_2_lut (.I0(\Kp[1] ), .I1(\PID_CONTROLLER.err[22] ), 
            .I2(GND_net), .I3(GND_net), .O(n164));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i111_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i48_2_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err[23] ), 
            .I2(GND_net), .I3(GND_net), .O(n71));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i48_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i392_2_lut (.I0(\Kd[6] ), .I1(n57[0]), .I2(GND_net), 
            .I3(GND_net), .O(n583_adj_3496));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i392_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i176_2_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err[22] ), 
            .I2(GND_net), .I3(GND_net), .O(n261));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i176_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i241_2_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err[22] ), 
            .I2(GND_net), .I3(GND_net), .O(n358));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i241_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i306_2_lut (.I0(\Kp[4] ), .I1(\PID_CONTROLLER.err[22] ), 
            .I2(GND_net), .I3(GND_net), .O(n455_c));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i306_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i457_2_lut (.I0(\Kd[7] ), .I1(n57[0]), .I2(GND_net), 
            .I3(GND_net), .O(n680_adj_3495));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i457_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i209_2_lut (.I0(\Kd[3] ), .I1(n57[6]), .I2(GND_net), 
            .I3(GND_net), .O(n310_adj_3494));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i209_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i371_2_lut (.I0(\Kp[5] ), .I1(\PID_CONTROLLER.err[22] ), 
            .I2(GND_net), .I3(GND_net), .O(n552));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i371_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_70_inv_0_i23_1_lut (.I0(pwm[22]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n73[22]));   // verilog/motorControl.v(86[38:44])
    defparam unary_minus_70_inv_0_i23_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_70_inv_0_i24_1_lut (.I0(pwm[23]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(GATES_5__N_3055));   // verilog/motorControl.v(86[38:44])
    defparam unary_minus_70_inv_0_i24_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i436_2_lut (.I0(\Kp[6] ), .I1(\PID_CONTROLLER.err[22] ), 
            .I2(GND_net), .I3(GND_net), .O(n649));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i436_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i345_2_lut (.I0(\Kd[5] ), .I1(n57[9]), .I2(GND_net), 
            .I3(GND_net), .O(n513));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i345_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i501_2_lut (.I0(\Kp[7] ), .I1(\PID_CONTROLLER.err[22] ), 
            .I2(GND_net), .I3(GND_net), .O(n746));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i501_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i91_2_lut (.I0(\Kp[1] ), .I1(\PID_CONTROLLER.err[12] ), 
            .I2(GND_net), .I3(GND_net), .O(n134_adj_3489));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i91_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i28_2_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err[13] ), 
            .I2(GND_net), .I3(GND_net), .O(n41_adj_3488));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i28_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i440_2_lut (.I0(\Kd[6] ), .I1(n57[24]), .I2(GND_net), 
            .I3(GND_net), .O(n655));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i440_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i156_2_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err[12] ), 
            .I2(GND_net), .I3(GND_net), .O(n231_adj_3487));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i156_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i410_2_lut (.I0(\Kd[6] ), .I1(n57[9]), .I2(GND_net), 
            .I3(GND_net), .O(n610));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i410_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i221_2_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err[12] ), 
            .I2(GND_net), .I3(GND_net), .O(n328_adj_3486));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i221_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i286_2_lut (.I0(\Kp[4] ), .I1(\PID_CONTROLLER.err[12] ), 
            .I2(GND_net), .I3(GND_net), .O(n425_adj_3485));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i286_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i505_2_lut (.I0(\Kd[7] ), .I1(n57[24]), .I2(GND_net), 
            .I3(GND_net), .O(n752));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i505_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i351_2_lut (.I0(\Kp[5] ), .I1(\PID_CONTROLLER.err[12] ), 
            .I2(GND_net), .I3(GND_net), .O(n522_adj_3484));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i351_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i101_2_lut (.I0(\Kd[1] ), .I1(n57[17]), .I2(GND_net), 
            .I3(GND_net), .O(n149_adj_3483));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i101_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i38_2_lut (.I0(\Kd[0] ), .I1(n57[18]), .I2(GND_net), 
            .I3(GND_net), .O(n56));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i38_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i274_2_lut (.I0(\Kd[4] ), .I1(n57[6]), .I2(GND_net), 
            .I3(GND_net), .O(n407_adj_3482));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i274_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i416_2_lut (.I0(\Kp[6] ), .I1(\PID_CONTROLLER.err[12] ), 
            .I2(GND_net), .I3(GND_net), .O(n619_adj_3480));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i416_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i339_2_lut (.I0(\Kd[5] ), .I1(n57[6]), .I2(GND_net), 
            .I3(GND_net), .O(n504_adj_3479));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i339_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i166_2_lut (.I0(\Kd[2] ), .I1(n57[17]), .I2(GND_net), 
            .I3(GND_net), .O(n246));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i166_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i231_2_lut (.I0(\Kd[3] ), .I1(n57[17]), .I2(GND_net), 
            .I3(GND_net), .O(n343));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i231_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i296_2_lut (.I0(\Kd[4] ), .I1(n57[17]), .I2(GND_net), 
            .I3(GND_net), .O(n440));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i296_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i361_2_lut (.I0(\Kd[5] ), .I1(n57[17]), .I2(GND_net), 
            .I3(GND_net), .O(n537));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i361_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i426_2_lut (.I0(\Kd[6] ), .I1(n57[17]), .I2(GND_net), 
            .I3(GND_net), .O(n634));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i426_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i475_2_lut (.I0(\Kd[7] ), .I1(n57[9]), .I2(GND_net), 
            .I3(GND_net), .O(n707));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i475_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i481_2_lut (.I0(\Kp[7] ), .I1(\PID_CONTROLLER.err[12] ), 
            .I2(GND_net), .I3(GND_net), .O(n716_adj_3477));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i481_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i404_2_lut (.I0(\Kd[6] ), .I1(n57[6]), .I2(GND_net), 
            .I3(GND_net), .O(n601_adj_3476));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i404_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i491_2_lut (.I0(\Kd[7] ), .I1(n57[17]), .I2(GND_net), 
            .I3(GND_net), .O(n731));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i491_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i95_2_lut (.I0(\Kd[1] ), .I1(n57[14]), .I2(GND_net), 
            .I3(GND_net), .O(n140_adj_3474));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i95_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i32_2_lut (.I0(\Kd[0] ), .I1(n57[15]), .I2(GND_net), 
            .I3(GND_net), .O(n47_adj_3473));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i32_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i469_2_lut (.I0(\Kd[7] ), .I1(n57[6]), .I2(GND_net), 
            .I3(GND_net), .O(n698_adj_3472));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i469_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i69_2_lut (.I0(\Kp[1] ), .I1(\PID_CONTROLLER.err[1] ), 
            .I2(GND_net), .I3(GND_net), .O(n101_adj_3471));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i69_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i6_2_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err[2] ), 
            .I2(GND_net), .I3(GND_net), .O(n8_adj_3470));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i6_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i134_2_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err[1] ), 
            .I2(GND_net), .I3(GND_net), .O(n198_adj_3469));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i134_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i105_2_lut (.I0(\Kp[1] ), .I1(\PID_CONTROLLER.err[19] ), 
            .I2(GND_net), .I3(GND_net), .O(n155_adj_3468));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i105_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i42_2_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err[20] ), 
            .I2(GND_net), .I3(GND_net), .O(n62_adj_3467));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i42_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i103_2_lut (.I0(\Kd[1] ), .I1(n57[18]), .I2(GND_net), 
            .I3(GND_net), .O(n152_adj_3466));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i103_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i40_2_lut (.I0(\Kd[0] ), .I1(n57[19]), .I2(GND_net), 
            .I3(GND_net), .O(n59_adj_3465));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i40_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i89_2_lut (.I0(\Kp[1] ), .I1(\PID_CONTROLLER.err[11] ), 
            .I2(GND_net), .I3(GND_net), .O(n131_adj_3463));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i89_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i26_2_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err[12] ), 
            .I2(GND_net), .I3(GND_net), .O(n38));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i26_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i160_2_lut (.I0(\Kd[2] ), .I1(n57[14]), .I2(GND_net), 
            .I3(GND_net), .O(n237));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i160_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i154_2_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err[11] ), 
            .I2(GND_net), .I3(GND_net), .O(n228_adj_3462));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i154_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i199_2_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err[1] ), 
            .I2(GND_net), .I3(GND_net), .O(n295_adj_3461));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i199_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i219_2_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err[11] ), 
            .I2(GND_net), .I3(GND_net), .O(n325));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i219_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i284_2_lut (.I0(\Kp[4] ), .I1(\PID_CONTROLLER.err[11] ), 
            .I2(GND_net), .I3(GND_net), .O(n422));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i284_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i170_2_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err[19] ), 
            .I2(GND_net), .I3(GND_net), .O(n252_adj_3460));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i170_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i168_2_lut (.I0(\Kd[2] ), .I1(n57[18]), .I2(GND_net), 
            .I3(GND_net), .O(n249_adj_3459));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i168_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i264_2_lut (.I0(\Kp[4] ), .I1(\PID_CONTROLLER.err[1] ), 
            .I2(GND_net), .I3(GND_net), .O(n392_adj_3458));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i264_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i349_2_lut (.I0(\Kp[5] ), .I1(\PID_CONTROLLER.err[11] ), 
            .I2(GND_net), .I3(GND_net), .O(n519));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i349_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i329_2_lut (.I0(\Kp[5] ), .I1(\PID_CONTROLLER.err[1] ), 
            .I2(GND_net), .I3(GND_net), .O(n489_adj_3457));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i329_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i394_2_lut (.I0(\Kp[6] ), .I1(\PID_CONTROLLER.err[1] ), 
            .I2(GND_net), .I3(GND_net), .O(n586_adj_3455));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i394_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i459_2_lut (.I0(\Kp[7] ), .I1(\PID_CONTROLLER.err[1] ), 
            .I2(GND_net), .I3(GND_net), .O(n683_adj_3454));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i459_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i414_2_lut (.I0(\Kp[6] ), .I1(\PID_CONTROLLER.err[11] ), 
            .I2(GND_net), .I3(GND_net), .O(n616));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i414_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 sub_11_inv_0_i1_1_lut (.I0(\PID_CONTROLLER.err[0] ), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n64[0]));   // verilog/motorControl.v(43[31:45])
    defparam sub_11_inv_0_i1_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i479_2_lut (.I0(\Kp[7] ), .I1(\PID_CONTROLLER.err[11] ), 
            .I2(GND_net), .I3(GND_net), .O(n713));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i479_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i235_2_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err[19] ), 
            .I2(GND_net), .I3(GND_net), .O(n349_adj_3453));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i235_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i107_2_lut (.I0(\Kp[1] ), .I1(\PID_CONTROLLER.err[20] ), 
            .I2(GND_net), .I3(GND_net), .O(n158));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i107_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i44_2_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err[21] ), 
            .I2(GND_net), .I3(GND_net), .O(n65));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i44_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i172_2_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err[20] ), 
            .I2(GND_net), .I3(GND_net), .O(n255));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i172_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i237_2_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err[20] ), 
            .I2(GND_net), .I3(GND_net), .O(n352));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i237_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 sub_11_inv_0_i2_1_lut (.I0(\PID_CONTROLLER.err[1] ), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n64[1]));   // verilog/motorControl.v(43[31:45])
    defparam sub_11_inv_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i302_2_lut (.I0(\Kp[4] ), .I1(\PID_CONTROLLER.err[20] ), 
            .I2(GND_net), .I3(GND_net), .O(n449));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i302_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i367_2_lut (.I0(\Kp[5] ), .I1(\PID_CONTROLLER.err[20] ), 
            .I2(GND_net), .I3(GND_net), .O(n546));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i367_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i432_2_lut (.I0(\Kp[6] ), .I1(\PID_CONTROLLER.err[20] ), 
            .I2(GND_net), .I3(GND_net), .O(n643));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i432_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i497_2_lut (.I0(\Kp[7] ), .I1(\PID_CONTROLLER.err[20] ), 
            .I2(GND_net), .I3(GND_net), .O(n740));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i497_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i83_2_lut (.I0(\Kp[1] ), .I1(\PID_CONTROLLER.err[8] ), 
            .I2(GND_net), .I3(GND_net), .O(n122_adj_3450));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i83_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i20_2_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err[9] ), 
            .I2(GND_net), .I3(GND_net), .O(n29_adj_3449));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i20_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i148_2_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err[8] ), 
            .I2(GND_net), .I3(GND_net), .O(n219_adj_3448));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i148_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i213_2_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err[8] ), 
            .I2(GND_net), .I3(GND_net), .O(n316_adj_3447));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i213_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i300_2_lut (.I0(\Kp[4] ), .I1(\PID_CONTROLLER.err[19] ), 
            .I2(GND_net), .I3(GND_net), .O(n446_adj_3446));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i300_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 sub_11_inv_0_i3_1_lut (.I0(\PID_CONTROLLER.err[2] ), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n64[2]));   // verilog/motorControl.v(43[31:45])
    defparam sub_11_inv_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_12_i225_2_lut (.I0(\Kd[3] ), .I1(n57[14]), .I2(GND_net), 
            .I3(GND_net), .O(n334));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i225_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i365_2_lut (.I0(\Kp[5] ), .I1(\PID_CONTROLLER.err[19] ), 
            .I2(GND_net), .I3(GND_net), .O(n543));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i365_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i430_2_lut (.I0(\Kp[6] ), .I1(\PID_CONTROLLER.err[19] ), 
            .I2(GND_net), .I3(GND_net), .O(n640));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i430_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i233_2_lut (.I0(\Kd[3] ), .I1(n57[18]), .I2(GND_net), 
            .I3(GND_net), .O(n346_adj_3445));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i233_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i290_2_lut (.I0(\Kd[4] ), .I1(n57[14]), .I2(GND_net), 
            .I3(GND_net), .O(n431));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i290_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i69_2_lut (.I0(\Kd[1] ), .I1(n57[1]), .I2(GND_net), 
            .I3(GND_net), .O(n101));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i69_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i6_2_lut (.I0(\Kd[0] ), .I1(n57[2]), .I2(GND_net), 
            .I3(GND_net), .O(n8));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i6_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i278_2_lut (.I0(\Kp[4] ), .I1(\PID_CONTROLLER.err[8] ), 
            .I2(GND_net), .I3(GND_net), .O(n413));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i278_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i495_2_lut (.I0(\Kp[7] ), .I1(\PID_CONTROLLER.err[19] ), 
            .I2(GND_net), .I3(GND_net), .O(n737));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i495_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i298_2_lut (.I0(\Kd[4] ), .I1(n57[18]), .I2(GND_net), 
            .I3(GND_net), .O(n443_adj_3443));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i298_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i355_2_lut (.I0(\Kd[5] ), .I1(n57[14]), .I2(GND_net), 
            .I3(GND_net), .O(n528));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i355_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i343_2_lut (.I0(\Kp[5] ), .I1(\PID_CONTROLLER.err[8] ), 
            .I2(GND_net), .I3(GND_net), .O(n510_adj_3442));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i343_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i408_2_lut (.I0(\Kp[6] ), .I1(\PID_CONTROLLER.err[8] ), 
            .I2(GND_net), .I3(GND_net), .O(n607));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i408_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i134_2_lut (.I0(\Kd[2] ), .I1(n57[1]), .I2(GND_net), 
            .I3(GND_net), .O(n198));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i134_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i420_2_lut (.I0(\Kd[6] ), .I1(n57[14]), .I2(GND_net), 
            .I3(GND_net), .O(n625));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i420_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i363_2_lut (.I0(\Kd[5] ), .I1(n57[18]), .I2(GND_net), 
            .I3(GND_net), .O(n540_adj_3439));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i363_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i199_2_lut (.I0(\Kd[3] ), .I1(n57[1]), .I2(GND_net), 
            .I3(GND_net), .O(n295));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i199_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i473_2_lut (.I0(\Kp[7] ), .I1(\PID_CONTROLLER.err[8] ), 
            .I2(GND_net), .I3(GND_net), .O(n704));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i473_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i485_2_lut (.I0(\Kd[7] ), .I1(n57[14]), .I2(GND_net), 
            .I3(GND_net), .O(n722));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i485_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1_3_lut_4_lut_4_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err[31] ), 
            .I2(n4_adj_3955), .I3(n35990), .O(n7_adj_3851));   // verilog/motorControl.v(43[17:23])
    defparam i1_3_lut_4_lut_4_lut.LUT_INIT = 16'h78b4;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1448 (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err[31] ), 
            .I2(n4_adj_3955), .I3(n16644[1]), .O(n16637[2]));   // verilog/motorControl.v(43[17:23])
    defparam i1_2_lut_3_lut_4_lut_adj_1448.LUT_INIT = 16'h8778;
    SB_LUT4 mult_12_i71_2_lut (.I0(\Kd[1] ), .I1(n57[2]), .I2(GND_net), 
            .I3(GND_net), .O(n104));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i71_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i8_2_lut (.I0(\Kd[0] ), .I1(n57[3]), .I2(GND_net), 
            .I3(GND_net), .O(n11_adj_3438));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i8_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i428_2_lut (.I0(\Kd[6] ), .I1(n57[18]), .I2(GND_net), 
            .I3(GND_net), .O(n637_adj_3437));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i428_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i493_2_lut (.I0(\Kd[7] ), .I1(n57[18]), .I2(GND_net), 
            .I3(GND_net), .O(n734_adj_3436));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i493_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i264_2_lut (.I0(\Kd[4] ), .I1(n57[1]), .I2(GND_net), 
            .I3(GND_net), .O(n392));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i264_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i329_2_lut (.I0(\Kd[5] ), .I1(n57[1]), .I2(GND_net), 
            .I3(GND_net), .O(n489));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i329_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i136_2_lut (.I0(\Kd[2] ), .I1(n57[2]), .I2(GND_net), 
            .I3(GND_net), .O(n201));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i136_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i103_2_lut (.I0(\Kp[1] ), .I1(\PID_CONTROLLER.err[18] ), 
            .I2(GND_net), .I3(GND_net), .O(n152_adj_3435));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i103_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i40_2_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err[19] ), 
            .I2(GND_net), .I3(GND_net), .O(n59));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i40_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i394_2_lut (.I0(\Kd[6] ), .I1(n57[1]), .I2(GND_net), 
            .I3(GND_net), .O(n586));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i394_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i168_2_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err[18] ), 
            .I2(GND_net), .I3(GND_net), .O(n249));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i168_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i459_2_lut (.I0(\Kd[7] ), .I1(n57[1]), .I2(GND_net), 
            .I3(GND_net), .O(n683));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i459_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 sub_11_inv_0_i4_1_lut (.I0(\PID_CONTROLLER.err[3] ), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n64[3]));   // verilog/motorControl.v(43[31:45])
    defparam sub_11_inv_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i233_2_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err[18] ), 
            .I2(GND_net), .I3(GND_net), .O(n346));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i233_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i298_2_lut (.I0(\Kp[4] ), .I1(\PID_CONTROLLER.err[18] ), 
            .I2(GND_net), .I3(GND_net), .O(n443));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i298_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i363_2_lut (.I0(\Kp[5] ), .I1(\PID_CONTROLLER.err[18] ), 
            .I2(GND_net), .I3(GND_net), .O(n540));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i363_2_lut.LUT_INIT = 16'h8888;
    
endmodule
//
// Verilog Description of module pll32MHz
//

module pll32MHz (GND_net, CLK_c, VCC_net, clk32MHz) /* synthesis lattice_noprune=1, syn_preserve=0, syn_module_defined=1, syn_noprune=0 */ ;
    input GND_net;
    input CLK_c;
    input VCC_net;
    output clk32MHz;
    
    wire clk32MHz /* synthesis SET_AS_NETWORK=clk32MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(34[8:16])
    
    SB_PLL40_CORE pll32MHz_inst (.REFERENCECLK(CLK_c), .PLLOUTGLOBAL(clk32MHz), 
            .BYPASS(GND_net), .RESETB(VCC_net)) /* synthesis lattice_noprune=1, syn_instantiated=1, LSE_LINE_FILE_ID=47, LSE_LCOL=12, LSE_RCOL=39, LSE_LLINE=35, LSE_RLINE=38, syn_preserve=0 */ ;   // verilog/TinyFPGA_B.v(35[12] 38[39])
    defparam pll32MHz_inst.FEEDBACK_PATH = "PHASE_AND_DELAY";
    defparam pll32MHz_inst.DELAY_ADJUSTMENT_MODE_FEEDBACK = "FIXED";
    defparam pll32MHz_inst.DELAY_ADJUSTMENT_MODE_RELATIVE = "FIXED";
    defparam pll32MHz_inst.SHIFTREG_DIV_MODE = 2'b00;
    defparam pll32MHz_inst.FDA_FEEDBACK = 4'b0000;
    defparam pll32MHz_inst.FDA_RELATIVE = 4'b0000;
    defparam pll32MHz_inst.PLLOUT_SELECT = "SHIFTREG_0deg";
    defparam pll32MHz_inst.DIVR = 4'b0000;
    defparam pll32MHz_inst.DIVF = 7'b0000001;
    defparam pll32MHz_inst.DIVQ = 3'b011;
    defparam pll32MHz_inst.FILTER_RANGE = 3'b001;
    defparam pll32MHz_inst.ENABLE_ICEGATE = 1'b0;
    defparam pll32MHz_inst.TEST_MODE = 1'b0;
    defparam pll32MHz_inst.EXTERNAL_DIVIDE_FACTOR = 1;
    
endmodule
//
// Verilog Description of module coms
//

module coms (clk32MHz, n24165, IntegralLimit, GND_net, n24164, n24163, 
            n24117, gearBoxRatio, n24116, n24115, n24114, n24113, 
            n24112, n24111, n24110, \data_in_frame[5] , \data_in_frame[3] , 
            n22338, pwm, n24109, n24108, n24107, n24106, n24105, 
            encoder0_position, n24104, n24103, n24102, n24101, n24100, 
            n24099, \data_in[0] , n24098, n24097, n24096, n24095, 
            n24094, n24093, n24092, \data_in[1] , n24091, encoder1_position, 
            n24269, \deadband[9] , n24268, \deadband[8] , n24267, 
            \deadband[7] , n24266, \deadband[6] , n24265, \deadband[5] , 
            n24264, \deadband[4] , n24263, \deadband[3] , n24262, 
            \deadband[2] , n24260, \deadband[1] , n24259, setpoint, 
            n24258, n24257, n24256, n24255, n24254, n24253, n24252, 
            n24251, n24250, n24249, n24248, n24247, n24246, n24245, 
            n24244, n24243, n24242, n24241, n24240, n24239, n24238, 
            n24237, VCC_net, byte_transmit_counter, n24169, n24168, 
            n24167, n24166, n24079, \data_in[2] , n24078, n24077, 
            n24076, \data_in[3] , n24075, n24074, n24073, n24072, 
            n24071, n24070, n24069, n24068, \data_out_frame[0][2] , 
            n24067, \data_out_frame[0][3] , n24066, \data_out_frame[0][4] , 
            n24063, \data_out_frame[5][2] , n24132, \Ki[5] , n24131, 
            \Ki[6] , n24130, \Ki[7] , n24129, \Kd[1] , n24128, \Kd[2] , 
            n24127, \Kd[3] , n24126, \Kd[4] , \data_in_frame[9] , 
            \data_in_frame[7] , n24125, \Kd[5] , n24090, n24089, n24088, 
            n24087, n40207, rx_data_ready, displacement, n24086, n24137, 
            \Kp[7] , n24136, \Ki[1] , n24124, \Kd[6] , n24085, n24162, 
            n24161, n24160, n24159, n24158, \data_out_frame[18][3] , 
            \data_in_frame[8] , rx_data, \data_out_frame[19][3] , n24157, 
            \data_out_frame[20][7] , n24156, n23930, \data_in_frame[1] , 
            n23929, n23928, n23927, n23926, \data_in_frame[6][1] , 
            \data_in_frame[6][0] , n23925, n23924, n23923, \data_in_frame[13] , 
            \data_in_frame[2] , n23914, n24155, n23913, n23912, n23911, 
            n23910, n23909, n23908, n23907, \data_in_frame[4] , n23898, 
            n23897, n23896, \data_in_frame[10] , n23895, n23894, n23893, 
            n23892, n23891, \data_in_frame[12][1] , \data_in_frame[12][0] , 
            n24151, n23866, n23865, n23864, n23863, n23862, n23861, 
            n23860, n23859, n23850, \data_in_frame[11] , n23849, n23848, 
            n23847, n23846, n23845, n23844, n23843, n24150, n24149, 
            n17, \data_in_frame[19] , n40227, n24148, n24147, n23834, 
            \data_in_frame[18] , n23833, n23832, n23831, n23830, n23829, 
            n23828, n23827, \data_in_frame[21] , \data_in_frame[17] , 
            n23802, n24084, n23801, n23800, n23799, n23798, n23797, 
            n23796, n23795, n23786, \data_out_frame[22][7] , \data_out_frame[21][7] , 
            n23785, n23784, n23783, n24135, \Ki[2] , n23782, n24134, 
            \Ki[3] , n23781, n24133, \Ki[4] , n23780, n23779, n23770, 
            n23769, n23768, n23767, n23766, n23765, n23764, n23763, 
            n23762, control_mode, n23761, n23760, n23759, n23758, 
            n23757, n23756, n23755, \PWMLimit[1] , n23754, \PWMLimit[2] , 
            n23753, \PWMLimit[3] , n23752, \PWMLimit[4] , n23751, 
            \PWMLimit[5] , n27220, \PWMLimit[6] , n23749, \PWMLimit[7] , 
            n23748, \PWMLimit[8] , n23747, \PWMLimit[9] , n24083, 
            n24082, n24123, \Kd[7] , n24081, n24080, n24122, n24146, 
            n24145, n24144, n24143, \Kp[1] , n24142, \Kp[2] , n24141, 
            \Kp[3] , n24140, \Kp[4] , n24139, \Kp[5] , n24138, \Kp[6] , 
            LED_c, n24121, n24120, n24119, n24118, n23600, \deadband[0] , 
            n23599, n23588, \PWMLimit[0] , n23587, n23585, n23584, 
            n23583, \Kd[0] , n23582, \Ki[0] , n23581, \Kp[0] , n23580, 
            n5019, n23458, n40218, n21, Kp_23__N_516, n22, n3792, 
            n3793, n23430, n3794, n3795, n3796, n3797, n3798, 
            n3799, n3800, n3801, n3802, n3803, n3804, n3805, n3806, 
            n3807, n3808, n3809, n3810, n3811, n3812, n3813, n3815, 
            n3814, n40209, n40222, n40213, n23399, n40216, n40225, 
            n40211, n313, \r_Clock_Count[8] , n314, \r_Clock_Count[7] , 
            n23624, n23627, n23630, \r_Clock_Count[6] , n23633, \r_Clock_Count[5] , 
            n23636, \r_Clock_Count[4] , n23639, \r_Clock_Count[3] , 
            n23642, \r_Clock_Count[2] , n23645, \r_Clock_Count[1] , 
            n23649, r_Bit_Index, n23652, n23695, n315, n316, n317, 
            n318, n319, n320, n23644, \r_SM_Main[2] , tx_o, tx_enable, 
            n23477, n23562, n4034, r_Rx_Data, \r_SM_Main[2]_adj_3 , 
            \r_SM_Main[1] , n23655, r_Bit_Index_adj_9, n23658, n28263, 
            n23698, n24171, PIN_13_N_26, n23665, n23664, n23663, 
            n23662, n23661, n23660, n23659, n23594, n22466, n4, 
            n28231, n1, n27725, n4_adj_7, n4_adj_8, n22471, n44134, 
            n44133, n23471, n23560, n4012) /* synthesis lattice_noprune=1, syn_preserve=0, syn_module_defined=1, syn_noprune=0 */ ;
    input clk32MHz;
    input n24165;
    output [23:0]IntegralLimit;
    input GND_net;
    input n24164;
    input n24163;
    input n24117;
    output [23:0]gearBoxRatio;
    input n24116;
    input n24115;
    input n24114;
    input n24113;
    input n24112;
    input n24111;
    input n24110;
    output [7:0]\data_in_frame[5] ;
    output [7:0]\data_in_frame[3] ;
    output n22338;
    input [23:0]pwm;
    input n24109;
    input n24108;
    input n24107;
    input n24106;
    input n24105;
    input [23:0]encoder0_position;
    input n24104;
    input n24103;
    input n24102;
    input n24101;
    input n24100;
    input n24099;
    output [7:0]\data_in[0] ;
    input n24098;
    input n24097;
    input n24096;
    input n24095;
    input n24094;
    input n24093;
    input n24092;
    output [7:0]\data_in[1] ;
    input n24091;
    input [23:0]encoder1_position;
    input n24269;
    output \deadband[9] ;
    input n24268;
    output \deadband[8] ;
    input n24267;
    output \deadband[7] ;
    input n24266;
    output \deadband[6] ;
    input n24265;
    output \deadband[5] ;
    input n24264;
    output \deadband[4] ;
    input n24263;
    output \deadband[3] ;
    input n24262;
    output \deadband[2] ;
    input n24260;
    output \deadband[1] ;
    input n24259;
    output [23:0]setpoint;
    input n24258;
    input n24257;
    input n24256;
    input n24255;
    input n24254;
    input n24253;
    input n24252;
    input n24251;
    input n24250;
    input n24249;
    input n24248;
    input n24247;
    input n24246;
    input n24245;
    input n24244;
    input n24243;
    input n24242;
    input n24241;
    input n24240;
    input n24239;
    input n24238;
    input n24237;
    input VCC_net;
    output [7:0]byte_transmit_counter;
    input n24169;
    input n24168;
    input n24167;
    input n24166;
    input n24079;
    output [7:0]\data_in[2] ;
    input n24078;
    input n24077;
    input n24076;
    output [7:0]\data_in[3] ;
    input n24075;
    input n24074;
    input n24073;
    input n24072;
    input n24071;
    input n24070;
    input n24069;
    input n24068;
    output \data_out_frame[0][2] ;
    input n24067;
    output \data_out_frame[0][3] ;
    input n24066;
    output \data_out_frame[0][4] ;
    input n24063;
    output \data_out_frame[5][2] ;
    input n24132;
    output \Ki[5] ;
    input n24131;
    output \Ki[6] ;
    input n24130;
    output \Ki[7] ;
    input n24129;
    output \Kd[1] ;
    input n24128;
    output \Kd[2] ;
    input n24127;
    output \Kd[3] ;
    input n24126;
    output \Kd[4] ;
    output [7:0]\data_in_frame[9] ;
    output [7:0]\data_in_frame[7] ;
    input n24125;
    output \Kd[5] ;
    input n24090;
    input n24089;
    input n24088;
    input n24087;
    output n40207;
    output rx_data_ready;
    input [23:0]displacement;
    input n24086;
    input n24137;
    output \Kp[7] ;
    input n24136;
    output \Ki[1] ;
    input n24124;
    output \Kd[6] ;
    input n24085;
    input n24162;
    input n24161;
    input n24160;
    input n24159;
    input n24158;
    output \data_out_frame[18][3] ;
    output [7:0]\data_in_frame[8] ;
    output [7:0]rx_data;
    output \data_out_frame[19][3] ;
    input n24157;
    output \data_out_frame[20][7] ;
    input n24156;
    input n23930;
    output [7:0]\data_in_frame[1] ;
    input n23929;
    input n23928;
    input n23927;
    input n23926;
    output \data_in_frame[6][1] ;
    output \data_in_frame[6][0] ;
    input n23925;
    input n23924;
    input n23923;
    output [7:0]\data_in_frame[13] ;
    output [7:0]\data_in_frame[2] ;
    input n23914;
    input n24155;
    input n23913;
    input n23912;
    input n23911;
    input n23910;
    input n23909;
    input n23908;
    input n23907;
    output [7:0]\data_in_frame[4] ;
    input n23898;
    input n23897;
    input n23896;
    output [7:0]\data_in_frame[10] ;
    input n23895;
    input n23894;
    input n23893;
    input n23892;
    input n23891;
    output \data_in_frame[12][1] ;
    output \data_in_frame[12][0] ;
    input n24151;
    input n23866;
    input n23865;
    input n23864;
    input n23863;
    input n23862;
    input n23861;
    input n23860;
    input n23859;
    input n23850;
    output [7:0]\data_in_frame[11] ;
    input n23849;
    input n23848;
    input n23847;
    input n23846;
    input n23845;
    input n23844;
    input n23843;
    input n24150;
    input n24149;
    input n17;
    output [7:0]\data_in_frame[19] ;
    output n40227;
    input n24148;
    input n24147;
    input n23834;
    output [7:0]\data_in_frame[18] ;
    input n23833;
    input n23832;
    input n23831;
    input n23830;
    input n23829;
    input n23828;
    input n23827;
    output [7:0]\data_in_frame[21] ;
    output [7:0]\data_in_frame[17] ;
    input n23802;
    input n24084;
    input n23801;
    input n23800;
    input n23799;
    input n23798;
    input n23797;
    input n23796;
    input n23795;
    input n23786;
    output \data_out_frame[22][7] ;
    output \data_out_frame[21][7] ;
    input n23785;
    input n23784;
    input n23783;
    input n24135;
    output \Ki[2] ;
    input n23782;
    input n24134;
    output \Ki[3] ;
    input n23781;
    input n24133;
    output \Ki[4] ;
    input n23780;
    input n23779;
    input n23770;
    input n23769;
    input n23768;
    input n23767;
    input n23766;
    input n23765;
    input n23764;
    input n23763;
    input n23762;
    output [7:0]control_mode;
    input n23761;
    input n23760;
    input n23759;
    input n23758;
    input n23757;
    input n23756;
    input n23755;
    output \PWMLimit[1] ;
    input n23754;
    output \PWMLimit[2] ;
    input n23753;
    output \PWMLimit[3] ;
    input n23752;
    output \PWMLimit[4] ;
    input n23751;
    output \PWMLimit[5] ;
    input n27220;
    output \PWMLimit[6] ;
    input n23749;
    output \PWMLimit[7] ;
    input n23748;
    output \PWMLimit[8] ;
    input n23747;
    output \PWMLimit[9] ;
    input n24083;
    input n24082;
    input n24123;
    output \Kd[7] ;
    input n24081;
    input n24080;
    input n24122;
    input n24146;
    input n24145;
    input n24144;
    input n24143;
    output \Kp[1] ;
    input n24142;
    output \Kp[2] ;
    input n24141;
    output \Kp[3] ;
    input n24140;
    output \Kp[4] ;
    input n24139;
    output \Kp[5] ;
    input n24138;
    output \Kp[6] ;
    output LED_c;
    input n24121;
    input n24120;
    input n24119;
    input n24118;
    input n23600;
    output \deadband[0] ;
    input n23599;
    input n23588;
    output \PWMLimit[0] ;
    input n23587;
    input n23585;
    input n23584;
    input n23583;
    output \Kd[0] ;
    input n23582;
    output \Ki[0] ;
    input n23581;
    output \Kp[0] ;
    input n23580;
    output n5019;
    output n23458;
    output n40218;
    input n21;
    input Kp_23__N_516;
    input n22;
    output n3792;
    output n3793;
    output n23430;
    output n3794;
    output n3795;
    output n3796;
    output n3797;
    output n3798;
    output n3799;
    output n3800;
    output n3801;
    output n3802;
    output n3803;
    output n3804;
    output n3805;
    output n3806;
    output n3807;
    output n3808;
    output n3809;
    output n3810;
    output n3811;
    output n3812;
    output n3813;
    output n3815;
    output n3814;
    output n40209;
    output n40222;
    output n40213;
    output n23399;
    output n40216;
    output n40225;
    output n40211;
    output n313;
    output \r_Clock_Count[8] ;
    output n314;
    output \r_Clock_Count[7] ;
    input n23624;
    input n23627;
    input n23630;
    output \r_Clock_Count[6] ;
    input n23633;
    output \r_Clock_Count[5] ;
    input n23636;
    output \r_Clock_Count[4] ;
    input n23639;
    output \r_Clock_Count[3] ;
    input n23642;
    output \r_Clock_Count[2] ;
    input n23645;
    output \r_Clock_Count[1] ;
    input n23649;
    output [2:0]r_Bit_Index;
    input n23652;
    input n23695;
    output n315;
    output n316;
    output n317;
    output n318;
    output n319;
    output n320;
    output n23644;
    output \r_SM_Main[2] ;
    output tx_o;
    output tx_enable;
    output n23477;
    output n23562;
    output n4034;
    output r_Rx_Data;
    output \r_SM_Main[2]_adj_3 ;
    output \r_SM_Main[1] ;
    input n23655;
    output [2:0]r_Bit_Index_adj_9;
    input n23658;
    input n28263;
    input n23698;
    input n24171;
    input PIN_13_N_26;
    input n23665;
    input n23664;
    input n23663;
    input n23662;
    input n23661;
    input n23660;
    input n23659;
    input n23594;
    output n22466;
    output n4;
    output n28231;
    output n1;
    output n27725;
    output n4_adj_7;
    output n4_adj_8;
    output n22471;
    output n44134;
    output n44133;
    output n23471;
    output n23560;
    output n4012;
    
    wire clk32MHz /* synthesis SET_AS_NETWORK=clk32MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(34[8:16])
    
    wire n24043;
    wire [7:0]\data_out_frame[7] ;   // verilog/coms.v(95[12:26])
    
    wire n24042, n24041;
    wire [7:0]\data_out_frame[8] ;   // verilog/coms.v(95[12:26])
    
    wire n24040, n34041;
    wire [31:0]\FRAME_MATCHER.i ;   // verilog/coms.v(113[11:12])
    
    wire n34042, n2, n34040, n1498, n34029, n34030, n24039, n2_adj_3119, 
        n34039, n40371, n22873;
    wire [31:0]\FRAME_MATCHER.state ;   // verilog/coms.v(110[11:16])
    wire [7:0]\data_out_frame[17] ;   // verilog/coms.v(95[12:26])
    
    wire n23963;
    wire [7:0]\data_out_frame[15] ;   // verilog/coms.v(95[12:26])
    
    wire n23980, n24038, n24037, n24036, n24035, n24034, n24033;
    wire [7:0]\data_out_frame[9] ;   // verilog/coms.v(95[12:26])
    
    wire n24047, n24032;
    wire [7:0]\data_out_frame[11] ;   // verilog/coms.v(95[12:26])
    
    wire n24012, n24234, n23668, n2_adj_3120, n34028, n23671;
    wire [7:0]byte_transmit_counter_c;   // verilog/coms.v(100[12:33])
    
    wire n23674, n23677, n23680, n24178, n24177, n24031, n24030, 
        n24029, n24028, n24027, n24026, n24025;
    wire [7:0]\data_out_frame[10] ;   // verilog/coms.v(95[12:26])
    
    wire n24024, n24023, n24022, n24021, n24020, n24019, n24018, 
        n24017, n24065;
    wire [7:0]\data_out_frame[5] ;   // verilog/coms.v(95[12:26])
    
    wire n24064, n24062, n24061, n24060, n24059, n24058, n24057;
    wire [7:0]\data_out_frame[6] ;   // verilog/coms.v(95[12:26])
    
    wire n24056, n24055, n24054, n24053, n24052, n24051, n24050, 
        n24049, n24016;
    wire [7:0]\data_out_frame[12] ;   // verilog/coms.v(95[12:26])
    
    wire n24007, n24015, n24048, n40591, n24014, n24013, n8, n24011, 
        n24010, n24009, n24008, n24006, n24005, n24004, n24003, 
        n24002, n24001;
    wire [7:0]\data_out_frame[13] ;   // verilog/coms.v(95[12:26])
    
    wire n24000, n23999, n23998, n23997, n23996, n40205, n23995, 
        n24046, n23994, n23993;
    wire [7:0]\data_out_frame[14] ;   // verilog/coms.v(95[12:26])
    
    wire n23992, \FRAME_MATCHER.rx_data_ready_prev , n2_adj_3121, n34038, 
        n23991, n23990, n23989;
    wire [7:0]\data_out_frame[20] ;   // verilog/coms.v(95[12:26])
    
    wire n23943, n23988, n23987, n23986, n23985, n23984, n23983, 
        n23982, n23981, n23979, n23978, n23977;
    wire [7:0]\data_out_frame[16] ;   // verilog/coms.v(95[12:26])
    
    wire n23976, n23975, n23974, n23973, n23972, n23971, n23970, 
        n23969, n23968, n23967, n23966, n23965, n23964, n23962, 
        n23961;
    wire [7:0]\data_out_frame[18] ;   // verilog/coms.v(95[12:26])
    
    wire n23960, n23959, n23958;
    wire [7:0]\data_in_frame[6] ;   // verilog/coms.v(94[12:25])
    
    wire n40619;
    wire [7:0]\data_in_frame[20] ;   // verilog/coms.v(94[12:25])
    
    wire n23771, n23772, n23773, n23774, n23957, n23956, n23955, 
        n23954, n164, n23953;
    wire [7:0]\data_out_frame[19] ;   // verilog/coms.v(95[12:26])
    
    wire n9, n8_adj_3122, n40212, n23883, n23884, n23952, n23885, 
        n23951, n23950, n23949, n23948, n23886, n23947, n23887, 
        n23946, n23775, n23945, n23944, n23942, n23941, n23940, 
        n23939, n23938, n23937;
    wire [7:0]\data_in_frame[0] ;   // verilog/coms.v(94[12:25])
    
    wire n23936, n23935, n23776, n23934, n24045, n23933, n23777, 
        n23932, n23931, n23888, n23889, n23890, n27747, n23875, 
        n23876, n23877, n23878, n23879, n41901, n23880, n23922, 
        n23921, n23881, n23920, n23919, n23918, n23778, n23882, 
        n23917, n8_adj_3123, n40221, n23867, n23916, n23915, n23868, 
        n23869, n23870, n23871, n23872, n23906, n23905, n23904, 
        n102, n23903, n23902, n23901, n23900, n23873, n23899, 
        n23874, n8_adj_3124, n23851, n23852;
    wire [7:0]\data_in_frame[16] ;   // verilog/coms.v(94[12:25])
    
    wire n40515, n37274, n23853, n2_adj_3125, n34037, n23854, n23855, 
        n23856, n23857, n23858;
    wire [7:0]\data_in_frame[12] ;   // verilog/coms.v(94[12:25])
    
    wire n23835, n23836, n23837, n23838, n23839, n23840, n23841, 
        n23842, Kp_23__N_908;
    wire [7:0]\data_in_frame[15] ;   // verilog/coms.v(94[12:25])
    
    wire n37237, n6, n22648, n15, n23101, n40831, n40773, n10;
    wire [7:0]\data_in_frame[14] ;   // verilog/coms.v(94[12:25])
    
    wire n40570, n36853, n37336;
    wire [7:0]\data_out_frame[21] ;   // verilog/coms.v(95[12:26])
    
    wire n19, n44438, n5;
    wire [7:0]\data_out_frame[22] ;   // verilog/coms.v(95[12:26])
    
    wire n42234, n46934, n42235, n42206, n42208, n46988, n47018, 
        n42207, n47003, n47006, n2_adj_3126, n34027, n2_adj_3127, 
        n34036, n40782, n40644, n37268, n40858, n40318, n40503, 
        n23275, Kp_23__N_379, n40481, n8_adj_3128, n40779, n40584, 
        n22842, n40752, n14, n10_adj_3129, n23157, n37248, n40478, 
        n40261, n40708, n40463, n40432, n40255, n4_c, n6_adj_3130, 
        Kp_23__N_329, n16, n10_adj_3131, n40834, n40308, n40383, 
        n18, n10_adj_3132, n20, Kp_23__N_326, n19_adj_3133, n9_adj_3134, 
        n40674, n40437, n23290, Kp_23__N_459, n40846, n5_adj_3135, 
        n40705, n40531, n40728, n40460, n40417, n23045, n2_adj_3136, 
        n34035, n10_adj_3137, n14_adj_3138, n37239, n40864, n40647, 
        n41875, n19_adj_3139, n44182, n47021, n16_adj_3140, n47024, 
        n40258, n23301, n47015, n14_adj_3141, n47009, n47012, n44143, 
        n5_adj_3142, n13, n42272, n42273, n46997, n42270, n42269, 
        n47000, n44012, n34061, n19614;
    wire [7:0]n2236;
    
    wire n34060, n34059, n34058, n13_adj_3143, n14_adj_3144, n27691, 
        n42278, n42279, n46991, n42276, n42275, n46994, n12, n46985, 
        n40420, n40487, n10_adj_3145, n46979, n46982, n40398, n41720, 
        n46973, n23826, n46976, n23825, n22997, n40746, n40554, 
        n41390, n23824, n46967, n23823, n46970, n23822, n41776, 
        n23821, n46961, n23820, n46964, n23819, n37284, n41583, 
        n23818, n46955, n23817, n46958, n23816, n47038, n23815, 
        n46949, n23814, n46952, n23813, n40567, n4_adj_3146, n23812, 
        n46943, n23811, n46946, n23810, n37241, n10_adj_3147, n23809, 
        n46937, n23808, n46940, n23807, n40362, n37310, n41687, 
        n23806, n2_adj_3148, n34034, n23805, n2_adj_3149, n34026, 
        n34057, n2_adj_3150, n34033, n34056, n2_adj_3151, n34025, 
        n23804, n23803, n46931, n39646, n39508, n2_adj_3152, n34024, 
        n34055, n39642, n39518, n39640, n39510, n27682, n39514, 
        n39638, n39550, n2_adj_3153, n34032, n39636, n39516, tx_transmit_N_2648, 
        n39634, n39496, n39632, n39492, n39744, n39494, n39686, 
        n39552, n39684, n39554, n39676, n35999, n39674, n39556, 
        n39672, n39512, n39670, n39522, n39668, n39436, n39666, 
        n39558, n39664, n39560, n39662, n39562, n39660, n39564, 
        n39658, n39566, n39656, n39568, n39654, n39570, n39652, 
        n39402, n39650, n39572, n39584, n28159, n27700, n28157, 
        n39648, n39406, n39506, n39742, n39504, n47026, n2_adj_3154, 
        n34054, n23794, n23793, n23792, n23791, n23790, n23789, 
        n23788, n23787, n41574, n23452, n41743, n40703, n40448, 
        n40449, n40375, n40513, n40514, n41732, n41124, n41129, 
        n41339, n41672, n41758, n41498, n41847, n3, n2_adj_3155, 
        n34053, n3_adj_3156, n2_adj_3157, n3_adj_3158, n2_adj_3159, 
        n3_adj_3160, n2_adj_3161, n3_adj_3162, n2_adj_3163, n3_adj_3164, 
        n2_adj_3165, n3_adj_3166, n2_adj_3167, n3_adj_3168, n2_adj_3169, 
        n3_adj_3170, n2_adj_3171, n3_adj_3172, n2_adj_3173, n3_adj_3174, 
        n2_adj_3175, n3_adj_3176, n2_adj_3177, n3_adj_3178, n2_adj_3179, 
        n3_adj_3180, n3_adj_3181, n3_adj_3182, n3_adj_3183, n3_adj_3184, 
        n3_adj_3185, n3_adj_3186, n3_adj_3187, n3_adj_3188, n3_adj_3189, 
        n2_adj_3190, n3_adj_3191, n2_adj_3192, n3_adj_3193, n2_adj_3194, 
        n3_adj_3195, n3_adj_3196, n3_adj_3197, n3_adj_3198, n3_adj_3199, 
        n3_adj_3200, n34052, n40352, n40564, n10_adj_3201, n34051, 
        n34050, n47027, n34049, n34031, n14_adj_3202, n11, n12_adj_3203, 
        n46919, n9_adj_3204, n8_adj_3205, n46922, n39256;
    wire [2:0]r_SM_Main_2__N_2756;
    
    wire n28289, n41389, n42155, n34048, n19_adj_3206, n40886, n46913, 
        n2_adj_3207, n31577, n40110, n20_adj_3208, n19_adj_3209, n34047, 
        n21_c, n40247, n10_adj_3210, n14_adj_3211, n40573, n47033, 
        n40106, n28279, n41005, n9_adj_3212, n18_adj_3213, n10_adj_3214, 
        n14_adj_3215, n46916, n34046, n41262, n30, n40668, n41134, 
        n28, n34045, n42187, n37295, n41676, n27, n11_adj_3216, 
        n34044, n3_adj_3217, n34043, n39520, n23586, n24044, n5021, 
        n28145;
    wire [31:0]\FRAME_MATCHER.state_31__N_1925 ;
    
    wire n41462, n10_adj_3218, n40840, n46907, n5_adj_3219, \FRAME_MATCHER.i_31__N_1825 , 
        n40163, n2857, n41799, \FRAME_MATCHER.i_31__N_1823 , n20075, 
        n46910, n47, n2_adj_3220, n6_adj_3221, n44587, n5_adj_3222, 
        n22_c, n43966, n42230, n42232, n19_adj_3224, n42201, n44581, 
        n5_adj_3225, n42202, n42227, n42229, n19_adj_3226, n44575, 
        n5_adj_3227, n42198, n46904, n42199, n42224, n42226, n46892, 
        n42225;
    wire [7:0]tx_data;   // verilog/coms.v(103[13:20])
    
    wire n19_adj_3228, n42195, n46898, n42196, n45804, n44129, n6_adj_3229, 
        n5_adj_3230, n42215, n42217, n42216, n44126, n19_adj_3231, 
        n6_adj_3232, n5_adj_3233, n42240, n42241, n42212, n42214, 
        n42213, n19_adj_3234, n44556, n5_adj_3235, n42237, n42238, 
        n42209, n42211, n4_adj_3236, n40828, n42210, n12_adj_3237, 
        n5_adj_3238, n43, n40791, n40662, n40339, n6_adj_3239, n40776, 
        n10_adj_3240, n40843, n40737, n14_adj_3241, n40653, n40359, 
        n22641, n6_adj_3242, n40495, n40637, n105, n27701, n28285, 
        n28293, n40173, n40867, n22816, n6_adj_3243, n40365, n40671, 
        n22716, n40699, n40450, n40392, n14_adj_3244, n10_adj_3245, 
        n23120, n22794, n40693, n40466, n40285, n41155, n11_adj_3246, 
        \FRAME_MATCHER.i_31__N_1821 , n52, n40788, n40755, n50, n40731, 
        n51, Kp_23__N_839, n49, n40876, n40734, n46, n40650, n48, 
        n40800, n40595, n47_adj_3247, n58, \FRAME_MATCHER.i_31__N_1827 , 
        n53, n37228, n63, n63_adj_3248, n63_adj_3249, n40193, n740, 
        n5_adj_3250, n40598, Kp_23__N_786, n40797, n41003, n15_adj_3251, 
        n41586, n37304, n3761, n6_adj_3252, n22250, n41620, n12_adj_3253, 
        n41987, n40377, n12_adj_3254, n23257, n6_adj_3255, n40540, 
        n16_adj_3256, n21050, n41706, n15_adj_3257, n36562, n40794, 
        n23094, n17_adj_3258, n18_adj_3259, n40332, n20_adj_3260, 
        n41807, n1_c, n36591, n22721, n40849, n40855, n46901, 
        n6_adj_3261, n6_adj_3262, n40677, n10_adj_3263, n23224, n23098, 
        n40322, n10_adj_3264, n40616, n6_adj_3265, n10_adj_3266, n22670, 
        n23350, n40326, n14_adj_3268, n10_adj_3269, n14_adj_3270, 
        n22_adj_3271, n40819, n21_adj_3272, n23, \FRAME_MATCHER.i_31__N_1824 , 
        n12_adj_3273, n36582, n40528, n12_adj_3274, n4_adj_3275, n10_adj_3276, 
        n40659, n6_adj_3277, n13_adj_3278, n15_adj_3279;
    wire [31:0]n7;
    
    wire tx_active, n28275, Kp_23__N_152, n736, n22347, n22400, 
        n4_adj_3280, n12_adj_3281, n27743, n41992, n40758, n6_adj_3282, 
        n27693, n44105, n8_adj_3283, n23400, n41662, n40279, n40612, 
        n40761, n12_adj_3284, n40628, n40292, n23166, n41642, n40401, 
        n10_adj_3285, n40282, n40380, n37253, n40822, n41673, n41806, 
        n36572, n8_adj_3286, n36494, n22729, n40690, n40415, n40810, 
        n10_adj_3287, n36991, n40490, n40329, n23285, n36529, n40535, 
        n36532, n10_adj_3288, n40356, n22132, n14_adj_3289, n40551, 
        n1695, n40561, n40641, n40785, n40656, n23316, n40311, 
        n36597, n12_adj_3290, n40767, n40837, n40631, n12_adj_3291, 
        n40861, n40723, n40665, n40349, n22047, n36629, n10_adj_3292, 
        n41402, n36837, n40506, n40474, n37234, n18_adj_3293, n30_adj_3294, 
        n40714, n28_adj_3295, n22635, n40764, n40609, n23383, n40588, 
        n29, n40622, n40870, n40581, n40368, n27_adj_3296, n37246, 
        n36588, n1787, n40558, n41416, n22840, n40813, n40576, 
        n42020, n40825, n40577, n40770, n6_adj_3297, n40298, n22666, 
        n40453, n37308, n10_adj_3298, n41192, n22071, n28_adj_3299, 
        n22134, n40429, n30_adj_3300, n40408, n31, n23169, n29_adj_3301, 
        n32, n37255, n10_adj_3302, n40343, n22515, n40423, n1595, 
        n6_adj_3303, n41850, n23107, n12_adj_3304, n40749, n40496, 
        n22095, n10_adj_3305, n31_adj_3306, n19864, n40414, n6_adj_3307, 
        n41802, n23038, n22_adj_3308, n23000, n40335, n20_adj_3309, 
        n16_adj_3310, n24, n23248, n40518, n48_adj_3311, n40604, 
        n54, n23004, n52_adj_3312, n22630, n53_adj_3313, n51_adj_3314, 
        n93, n40386, n50_adj_3315, n36, n56, n60, n40499, n55, 
        n37341, n1664, n40852, n40720, n16_adj_3316, n40806, n40873, 
        n17_adj_3317, n1515, n30_adj_3318, n22511, n41479, n40443, 
        n34, n40471, n32_adj_3319, n22051, n1716, n40711, n33, 
        n31_adj_3320, n40717, n6_adj_3321, n37264, n40634, n40249, 
        n1506, n37222, n40684, n23218, n40548, n18_adj_3322, n16_adj_3323, 
        n20_adj_3324, n40740, n40521, n6_adj_3325, n40816, n4_adj_3326, 
        n23323, n6_adj_3327, n40381, n40456, n40803, n18_adj_3328, 
        n20_adj_3329, n16_adj_3330, n6_adj_3331, n40696, n23029, n14_adj_3332, 
        n15_adj_3333, n40440, n46895, n40681, n40295, n6_adj_3334, 
        n40625, n10_adj_3335, n40289, n14_adj_3336, n15_adj_3337, 
        n4_adj_3338, n10_adj_3339, n9_adj_3340, n40411, n5_adj_3341, 
        n1_adj_3342, n36044, n8_adj_3343, n44171, n44173, n36224, 
        n10_adj_3344, n17_adj_3345, n6_adj_3346, n6_adj_3347, n8_adj_3348, 
        n42018, n14_adj_3349, n13_adj_3350, n9_adj_3351, n11_adj_3352, 
        n10_adj_3353, n14_adj_3354, n22476, n15_adj_3355, n22256, 
        n16_adj_3356, n17_adj_3357, n22341, n10_adj_3358, n12_adj_3359, 
        n13_adj_3360, n22374, n18_adj_3361, n20_adj_3362, n15_adj_3363, 
        n16_adj_3364, n17_adj_3365, n20_adj_3366, n19_adj_3367, n42179, 
        n28265, n46889;
    
    SB_DFF data_out_frame_0___i63 (.Q(\data_out_frame[7] [6]), .C(clk32MHz), 
           .D(n24043));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i64 (.Q(\data_out_frame[7] [7]), .C(clk32MHz), 
           .D(n24042));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i65 (.Q(\data_out_frame[8] [0]), .C(clk32MHz), 
           .D(n24041));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i66 (.Q(\data_out_frame[8] [1]), .C(clk32MHz), 
           .D(n24040));   // verilog/coms.v(126[12] 289[6])
    SB_DFF IntegralLimit_i0_i5 (.Q(IntegralLimit[5]), .C(clk32MHz), .D(n24165));   // verilog/coms.v(126[12] 289[6])
    SB_CARRY add_44_20 (.CI(n34041), .I0(\FRAME_MATCHER.i [18]), .I1(GND_net), 
            .CO(n34042));
    SB_LUT4 add_44_19_lut (.I0(n1498), .I1(\FRAME_MATCHER.i [17]), .I2(GND_net), 
            .I3(n34040), .O(n2)) /* synthesis syn_instantiated=1 */ ;
    defparam add_44_19_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_44_8 (.CI(n34029), .I0(\FRAME_MATCHER.i [6]), .I1(GND_net), 
            .CO(n34030));
    SB_CARRY add_44_19 (.CI(n34040), .I0(\FRAME_MATCHER.i [17]), .I1(GND_net), 
            .CO(n34041));
    SB_DFF IntegralLimit_i0_i6 (.Q(IntegralLimit[6]), .C(clk32MHz), .D(n24164));   // verilog/coms.v(126[12] 289[6])
    SB_DFF IntegralLimit_i0_i7 (.Q(IntegralLimit[7]), .C(clk32MHz), .D(n24163));   // verilog/coms.v(126[12] 289[6])
    SB_DFF gearBoxRatio_i0_i6 (.Q(gearBoxRatio[6]), .C(clk32MHz), .D(n24117));   // verilog/coms.v(126[12] 289[6])
    SB_DFF gearBoxRatio_i0_i7 (.Q(gearBoxRatio[7]), .C(clk32MHz), .D(n24116));   // verilog/coms.v(126[12] 289[6])
    SB_DFF gearBoxRatio_i0_i8 (.Q(gearBoxRatio[8]), .C(clk32MHz), .D(n24115));   // verilog/coms.v(126[12] 289[6])
    SB_DFF gearBoxRatio_i0_i9 (.Q(gearBoxRatio[9]), .C(clk32MHz), .D(n24114));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i67 (.Q(\data_out_frame[8] [2]), .C(clk32MHz), 
           .D(n24039));   // verilog/coms.v(126[12] 289[6])
    SB_DFF gearBoxRatio_i0_i10 (.Q(gearBoxRatio[10]), .C(clk32MHz), .D(n24113));   // verilog/coms.v(126[12] 289[6])
    SB_DFF gearBoxRatio_i0_i11 (.Q(gearBoxRatio[11]), .C(clk32MHz), .D(n24112));   // verilog/coms.v(126[12] 289[6])
    SB_DFF gearBoxRatio_i0_i12 (.Q(gearBoxRatio[12]), .C(clk32MHz), .D(n24111));   // verilog/coms.v(126[12] 289[6])
    SB_DFF gearBoxRatio_i0_i13 (.Q(gearBoxRatio[13]), .C(clk32MHz), .D(n24110));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 add_44_18_lut (.I0(n1498), .I1(\FRAME_MATCHER.i [16]), .I2(GND_net), 
            .I3(n34039), .O(n2_adj_3119)) /* synthesis syn_instantiated=1 */ ;
    defparam add_44_18_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i1_4_lut (.I0(\data_in_frame[5] [3]), .I1(\data_in_frame[3] [2]), 
            .I2(n40371), .I3(\data_in_frame[3] [1]), .O(n22873));
    defparam i1_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i10545_3_lut_4_lut (.I0(\FRAME_MATCHER.state [2]), .I1(n22338), 
            .I2(pwm[6]), .I3(\data_out_frame[17] [6]), .O(n23963));
    defparam i10545_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i10562_3_lut_4_lut (.I0(\FRAME_MATCHER.state [2]), .I1(n22338), 
            .I2(pwm[21]), .I3(\data_out_frame[15] [5]), .O(n23980));
    defparam i10562_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_CARRY add_44_18 (.CI(n34039), .I0(\FRAME_MATCHER.i [16]), .I1(GND_net), 
            .CO(n34040));
    SB_DFF data_out_frame_0___i68 (.Q(\data_out_frame[8] [3]), .C(clk32MHz), 
           .D(n24038));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i69 (.Q(\data_out_frame[8] [4]), .C(clk32MHz), 
           .D(n24037));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i70 (.Q(\data_out_frame[8] [5]), .C(clk32MHz), 
           .D(n24036));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i71 (.Q(\data_out_frame[8] [6]), .C(clk32MHz), 
           .D(n24035));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i72 (.Q(\data_out_frame[8] [7]), .C(clk32MHz), 
           .D(n24034));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i73 (.Q(\data_out_frame[9] [0]), .C(clk32MHz), 
           .D(n24033));   // verilog/coms.v(126[12] 289[6])
    SB_DFF gearBoxRatio_i0_i14 (.Q(gearBoxRatio[14]), .C(clk32MHz), .D(n24109));   // verilog/coms.v(126[12] 289[6])
    SB_DFF gearBoxRatio_i0_i15 (.Q(gearBoxRatio[15]), .C(clk32MHz), .D(n24108));   // verilog/coms.v(126[12] 289[6])
    SB_DFF gearBoxRatio_i0_i16 (.Q(gearBoxRatio[16]), .C(clk32MHz), .D(n24107));   // verilog/coms.v(126[12] 289[6])
    SB_DFF gearBoxRatio_i0_i17 (.Q(gearBoxRatio[17]), .C(clk32MHz), .D(n24106));   // verilog/coms.v(126[12] 289[6])
    SB_DFF gearBoxRatio_i0_i18 (.Q(gearBoxRatio[18]), .C(clk32MHz), .D(n24105));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i10629_3_lut_4_lut (.I0(\FRAME_MATCHER.state [2]), .I1(n22338), 
            .I2(encoder0_position[10]), .I3(\data_out_frame[7] [2]), .O(n24047));
    defparam i10629_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_DFF gearBoxRatio_i0_i19 (.Q(gearBoxRatio[19]), .C(clk32MHz), .D(n24104));   // verilog/coms.v(126[12] 289[6])
    SB_DFF gearBoxRatio_i0_i20 (.Q(gearBoxRatio[20]), .C(clk32MHz), .D(n24103));   // verilog/coms.v(126[12] 289[6])
    SB_DFF gearBoxRatio_i0_i21 (.Q(gearBoxRatio[21]), .C(clk32MHz), .D(n24102));   // verilog/coms.v(126[12] 289[6])
    SB_DFF gearBoxRatio_i0_i22 (.Q(gearBoxRatio[22]), .C(clk32MHz), .D(n24101));   // verilog/coms.v(126[12] 289[6])
    SB_DFF gearBoxRatio_i0_i23 (.Q(gearBoxRatio[23]), .C(clk32MHz), .D(n24100));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_0___i2 (.Q(\data_in[0] [1]), .C(clk32MHz), .D(n24099));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_0___i3 (.Q(\data_in[0] [2]), .C(clk32MHz), .D(n24098));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_0___i4 (.Q(\data_in[0] [3]), .C(clk32MHz), .D(n24097));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_0___i5 (.Q(\data_in[0] [4]), .C(clk32MHz), .D(n24096));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_0___i6 (.Q(\data_in[0] [5]), .C(clk32MHz), .D(n24095));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_0___i7 (.Q(\data_in[0] [6]), .C(clk32MHz), .D(n24094));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_0___i8 (.Q(\data_in[0] [7]), .C(clk32MHz), .D(n24093));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_0___i9 (.Q(\data_in[1] [0]), .C(clk32MHz), .D(n24092));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_0___i10 (.Q(\data_in[1] [1]), .C(clk32MHz), .D(n24091));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i74 (.Q(\data_out_frame[9] [1]), .C(clk32MHz), 
           .D(n24032));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i10594_3_lut_4_lut (.I0(\FRAME_MATCHER.state [2]), .I1(n22338), 
            .I2(encoder1_position[5]), .I3(\data_out_frame[11] [5]), .O(n24012));
    defparam i10594_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_DFF deadband_i0_i9 (.Q(\deadband[9] ), .C(clk32MHz), .D(n24269));   // verilog/coms.v(126[12] 289[6])
    SB_DFF deadband_i0_i8 (.Q(\deadband[8] ), .C(clk32MHz), .D(n24268));   // verilog/coms.v(126[12] 289[6])
    SB_DFF deadband_i0_i7 (.Q(\deadband[7] ), .C(clk32MHz), .D(n24267));   // verilog/coms.v(126[12] 289[6])
    SB_DFF deadband_i0_i6 (.Q(\deadband[6] ), .C(clk32MHz), .D(n24266));   // verilog/coms.v(126[12] 289[6])
    SB_DFF deadband_i0_i5 (.Q(\deadband[5] ), .C(clk32MHz), .D(n24265));   // verilog/coms.v(126[12] 289[6])
    SB_DFF deadband_i0_i4 (.Q(\deadband[4] ), .C(clk32MHz), .D(n24264));   // verilog/coms.v(126[12] 289[6])
    SB_DFF deadband_i0_i3 (.Q(\deadband[3] ), .C(clk32MHz), .D(n24263));   // verilog/coms.v(126[12] 289[6])
    SB_DFF deadband_i0_i2 (.Q(\deadband[2] ), .C(clk32MHz), .D(n24262));   // verilog/coms.v(126[12] 289[6])
    SB_DFF deadband_i0_i1 (.Q(\deadband[1] ), .C(clk32MHz), .D(n24260));   // verilog/coms.v(126[12] 289[6])
    SB_DFF setpoint__i23 (.Q(setpoint[23]), .C(clk32MHz), .D(n24259));   // verilog/coms.v(126[12] 289[6])
    SB_DFF setpoint__i22 (.Q(setpoint[22]), .C(clk32MHz), .D(n24258));   // verilog/coms.v(126[12] 289[6])
    SB_DFF setpoint__i21 (.Q(setpoint[21]), .C(clk32MHz), .D(n24257));   // verilog/coms.v(126[12] 289[6])
    SB_DFF setpoint__i20 (.Q(setpoint[20]), .C(clk32MHz), .D(n24256));   // verilog/coms.v(126[12] 289[6])
    SB_DFF setpoint__i19 (.Q(setpoint[19]), .C(clk32MHz), .D(n24255));   // verilog/coms.v(126[12] 289[6])
    SB_DFF setpoint__i18 (.Q(setpoint[18]), .C(clk32MHz), .D(n24254));   // verilog/coms.v(126[12] 289[6])
    SB_DFF setpoint__i17 (.Q(setpoint[17]), .C(clk32MHz), .D(n24253));   // verilog/coms.v(126[12] 289[6])
    SB_DFF setpoint__i16 (.Q(setpoint[16]), .C(clk32MHz), .D(n24252));   // verilog/coms.v(126[12] 289[6])
    SB_DFF setpoint__i15 (.Q(setpoint[15]), .C(clk32MHz), .D(n24251));   // verilog/coms.v(126[12] 289[6])
    SB_DFF setpoint__i14 (.Q(setpoint[14]), .C(clk32MHz), .D(n24250));   // verilog/coms.v(126[12] 289[6])
    SB_DFF setpoint__i13 (.Q(setpoint[13]), .C(clk32MHz), .D(n24249));   // verilog/coms.v(126[12] 289[6])
    SB_DFF setpoint__i12 (.Q(setpoint[12]), .C(clk32MHz), .D(n24248));   // verilog/coms.v(126[12] 289[6])
    SB_DFF setpoint__i11 (.Q(setpoint[11]), .C(clk32MHz), .D(n24247));   // verilog/coms.v(126[12] 289[6])
    SB_DFF setpoint__i10 (.Q(setpoint[10]), .C(clk32MHz), .D(n24246));   // verilog/coms.v(126[12] 289[6])
    SB_DFF setpoint__i9 (.Q(setpoint[9]), .C(clk32MHz), .D(n24245));   // verilog/coms.v(126[12] 289[6])
    SB_DFF setpoint__i8 (.Q(setpoint[8]), .C(clk32MHz), .D(n24244));   // verilog/coms.v(126[12] 289[6])
    SB_DFF setpoint__i7 (.Q(setpoint[7]), .C(clk32MHz), .D(n24243));   // verilog/coms.v(126[12] 289[6])
    SB_DFF setpoint__i6 (.Q(setpoint[6]), .C(clk32MHz), .D(n24242));   // verilog/coms.v(126[12] 289[6])
    SB_DFF setpoint__i5 (.Q(setpoint[5]), .C(clk32MHz), .D(n24241));   // verilog/coms.v(126[12] 289[6])
    SB_DFF setpoint__i4 (.Q(setpoint[4]), .C(clk32MHz), .D(n24240));   // verilog/coms.v(126[12] 289[6])
    SB_DFF setpoint__i3 (.Q(setpoint[3]), .C(clk32MHz), .D(n24239));   // verilog/coms.v(126[12] 289[6])
    SB_DFF setpoint__i2 (.Q(setpoint[2]), .C(clk32MHz), .D(n24238));   // verilog/coms.v(126[12] 289[6])
    SB_DFF setpoint__i1 (.Q(setpoint[1]), .C(clk32MHz), .D(n24237));   // verilog/coms.v(126[12] 289[6])
    SB_DFFE byte_transmit_counter_i0_i0 (.Q(byte_transmit_counter[0]), .C(clk32MHz), 
            .E(VCC_net), .D(n24234));   // verilog/coms.v(126[12] 289[6])
    SB_DFF byte_transmit_counter_i0_i1 (.Q(byte_transmit_counter[1]), .C(clk32MHz), 
           .D(n23668));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 add_44_7_lut (.I0(n1498), .I1(\FRAME_MATCHER.i [5]), .I2(GND_net), 
            .I3(n34028), .O(n2_adj_3120)) /* synthesis syn_instantiated=1 */ ;
    defparam add_44_7_lut.LUT_INIT = 16'h8228;
    SB_DFF byte_transmit_counter_i0_i2 (.Q(byte_transmit_counter_c[2]), .C(clk32MHz), 
           .D(n23671));   // verilog/coms.v(126[12] 289[6])
    SB_DFF byte_transmit_counter_i0_i3 (.Q(byte_transmit_counter_c[3]), .C(clk32MHz), 
           .D(n23674));   // verilog/coms.v(126[12] 289[6])
    SB_DFF byte_transmit_counter_i0_i4 (.Q(byte_transmit_counter_c[4]), .C(clk32MHz), 
           .D(n23677));   // verilog/coms.v(126[12] 289[6])
    SB_DFF byte_transmit_counter_i0_i5 (.Q(byte_transmit_counter_c[5]), .C(clk32MHz), 
           .D(n23680));   // verilog/coms.v(126[12] 289[6])
    SB_DFF byte_transmit_counter_i0_i6 (.Q(byte_transmit_counter_c[6]), .C(clk32MHz), 
           .D(n24178));   // verilog/coms.v(126[12] 289[6])
    SB_DFF byte_transmit_counter_i0_i7 (.Q(byte_transmit_counter_c[7]), .C(clk32MHz), 
           .D(n24177));   // verilog/coms.v(126[12] 289[6])
    SB_DFF IntegralLimit_i0_i1 (.Q(IntegralLimit[1]), .C(clk32MHz), .D(n24169));   // verilog/coms.v(126[12] 289[6])
    SB_DFF IntegralLimit_i0_i2 (.Q(IntegralLimit[2]), .C(clk32MHz), .D(n24168));   // verilog/coms.v(126[12] 289[6])
    SB_DFF IntegralLimit_i0_i3 (.Q(IntegralLimit[3]), .C(clk32MHz), .D(n24167));   // verilog/coms.v(126[12] 289[6])
    SB_DFF IntegralLimit_i0_i4 (.Q(IntegralLimit[4]), .C(clk32MHz), .D(n24166));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i75 (.Q(\data_out_frame[9] [2]), .C(clk32MHz), 
           .D(n24031));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_0___i22 (.Q(\data_in[2] [5]), .C(clk32MHz), .D(n24079));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i76 (.Q(\data_out_frame[9] [3]), .C(clk32MHz), 
           .D(n24030));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_0___i23 (.Q(\data_in[2] [6]), .C(clk32MHz), .D(n24078));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i77 (.Q(\data_out_frame[9] [4]), .C(clk32MHz), 
           .D(n24029));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_0___i24 (.Q(\data_in[2] [7]), .C(clk32MHz), .D(n24077));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i78 (.Q(\data_out_frame[9] [5]), .C(clk32MHz), 
           .D(n24028));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_0___i25 (.Q(\data_in[3] [0]), .C(clk32MHz), .D(n24076));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i79 (.Q(\data_out_frame[9] [6]), .C(clk32MHz), 
           .D(n24027));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_0___i26 (.Q(\data_in[3] [1]), .C(clk32MHz), .D(n24075));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i80 (.Q(\data_out_frame[9] [7]), .C(clk32MHz), 
           .D(n24026));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_0___i27 (.Q(\data_in[3] [2]), .C(clk32MHz), .D(n24074));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i81 (.Q(\data_out_frame[10] [0]), .C(clk32MHz), 
           .D(n24025));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_0___i28 (.Q(\data_in[3] [3]), .C(clk32MHz), .D(n24073));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i82 (.Q(\data_out_frame[10] [1]), .C(clk32MHz), 
           .D(n24024));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_0___i29 (.Q(\data_in[3] [4]), .C(clk32MHz), .D(n24072));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i83 (.Q(\data_out_frame[10] [2]), .C(clk32MHz), 
           .D(n24023));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_0___i30 (.Q(\data_in[3] [5]), .C(clk32MHz), .D(n24071));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i84 (.Q(\data_out_frame[10] [3]), .C(clk32MHz), 
           .D(n24022));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_0___i31 (.Q(\data_in[3] [6]), .C(clk32MHz), .D(n24070));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i85 (.Q(\data_out_frame[10] [4]), .C(clk32MHz), 
           .D(n24021));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_0___i32 (.Q(\data_in[3] [7]), .C(clk32MHz), .D(n24069));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i86 (.Q(\data_out_frame[10] [5]), .C(clk32MHz), 
           .D(n24020));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i3 (.Q(\data_out_frame[0][2] ), .C(clk32MHz), 
           .D(n24068));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i87 (.Q(\data_out_frame[10] [6]), .C(clk32MHz), 
           .D(n24019));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i4 (.Q(\data_out_frame[0][3] ), .C(clk32MHz), 
           .D(n24067));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i88 (.Q(\data_out_frame[10] [7]), .C(clk32MHz), 
           .D(n24018));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i5 (.Q(\data_out_frame[0][4] ), .C(clk32MHz), 
           .D(n24066));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i89 (.Q(\data_out_frame[11] [0]), .C(clk32MHz), 
           .D(n24017));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i41 (.Q(\data_out_frame[5] [0]), .C(clk32MHz), 
           .D(n24065));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i42 (.Q(\data_out_frame[5] [1]), .C(clk32MHz), 
           .D(n24064));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i43 (.Q(\data_out_frame[5][2] ), .C(clk32MHz), 
           .D(n24063));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i44 (.Q(\data_out_frame[5] [3]), .C(clk32MHz), 
           .D(n24062));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i45 (.Q(\data_out_frame[5] [4]), .C(clk32MHz), 
           .D(n24061));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i46 (.Q(\data_out_frame[5] [5]), .C(clk32MHz), 
           .D(n24060));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i47 (.Q(\data_out_frame[5] [6]), .C(clk32MHz), 
           .D(n24059));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i48 (.Q(\data_out_frame[5] [7]), .C(clk32MHz), 
           .D(n24058));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i49 (.Q(\data_out_frame[6] [0]), .C(clk32MHz), 
           .D(n24057));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i50 (.Q(\data_out_frame[6] [1]), .C(clk32MHz), 
           .D(n24056));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i51 (.Q(\data_out_frame[6] [2]), .C(clk32MHz), 
           .D(n24055));   // verilog/coms.v(126[12] 289[6])
    SB_DFF Ki_i5 (.Q(\Ki[5] ), .C(clk32MHz), .D(n24132));   // verilog/coms.v(126[12] 289[6])
    SB_DFF Ki_i6 (.Q(\Ki[6] ), .C(clk32MHz), .D(n24131));   // verilog/coms.v(126[12] 289[6])
    SB_DFF Ki_i7 (.Q(\Ki[7] ), .C(clk32MHz), .D(n24130));   // verilog/coms.v(126[12] 289[6])
    SB_DFF Kd_i1 (.Q(\Kd[1] ), .C(clk32MHz), .D(n24129));   // verilog/coms.v(126[12] 289[6])
    SB_DFF Kd_i2 (.Q(\Kd[2] ), .C(clk32MHz), .D(n24128));   // verilog/coms.v(126[12] 289[6])
    SB_DFF Kd_i3 (.Q(\Kd[3] ), .C(clk32MHz), .D(n24127));   // verilog/coms.v(126[12] 289[6])
    SB_DFF Kd_i4 (.Q(\Kd[4] ), .C(clk32MHz), .D(n24126));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i52 (.Q(\data_out_frame[6] [3]), .C(clk32MHz), 
           .D(n24054));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i53 (.Q(\data_out_frame[6] [4]), .C(clk32MHz), 
           .D(n24053));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i54 (.Q(\data_out_frame[6] [5]), .C(clk32MHz), 
           .D(n24052));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i55 (.Q(\data_out_frame[6] [6]), .C(clk32MHz), 
           .D(n24051));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i56 (.Q(\data_out_frame[6] [7]), .C(clk32MHz), 
           .D(n24050));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i57 (.Q(\data_out_frame[7] [0]), .C(clk32MHz), 
           .D(n24049));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i90 (.Q(\data_out_frame[11] [1]), .C(clk32MHz), 
           .D(n24016));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i10589_3_lut_4_lut (.I0(\FRAME_MATCHER.state [2]), .I1(n22338), 
            .I2(setpoint[18]), .I3(\data_out_frame[12] [2]), .O(n24007));
    defparam i10589_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_DFF data_out_frame_0___i91 (.Q(\data_out_frame[11] [2]), .C(clk32MHz), 
           .D(n24015));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i58 (.Q(\data_out_frame[7] [1]), .C(clk32MHz), 
           .D(n24048));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i59 (.Q(\data_out_frame[7] [2]), .C(clk32MHz), 
           .D(n24047));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i2_3_lut (.I0(\data_in_frame[9] [5]), .I1(\data_in_frame[7] [4]), 
            .I2(n22873), .I3(GND_net), .O(n40591));
    defparam i2_3_lut.LUT_INIT = 16'h9696;
    SB_DFF data_out_frame_0___i92 (.Q(\data_out_frame[11] [3]), .C(clk32MHz), 
           .D(n24014));   // verilog/coms.v(126[12] 289[6])
    SB_DFF Kd_i5 (.Q(\Kd[5] ), .C(clk32MHz), .D(n24125));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i93 (.Q(\data_out_frame[11] [4]), .C(clk32MHz), 
           .D(n24013));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_0___i11 (.Q(\data_in[1] [2]), .C(clk32MHz), .D(n24090));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 equal_63_i8_2_lut_3_lut (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(\FRAME_MATCHER.i [0]), .I3(GND_net), .O(n8));   // verilog/coms.v(154[7:23])
    defparam equal_63_i8_2_lut_3_lut.LUT_INIT = 16'hfbfb;
    SB_DFF data_out_frame_0___i94 (.Q(\data_out_frame[11] [5]), .C(clk32MHz), 
           .D(n24012));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i95 (.Q(\data_out_frame[11] [6]), .C(clk32MHz), 
           .D(n24011));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i96 (.Q(\data_out_frame[11] [7]), .C(clk32MHz), 
           .D(n24010));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i97 (.Q(\data_out_frame[12] [0]), .C(clk32MHz), 
           .D(n24009));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i98 (.Q(\data_out_frame[12] [1]), .C(clk32MHz), 
           .D(n24008));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i99 (.Q(\data_out_frame[12] [2]), .C(clk32MHz), 
           .D(n24007));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i100 (.Q(\data_out_frame[12] [3]), .C(clk32MHz), 
           .D(n24006));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i101 (.Q(\data_out_frame[12] [4]), .C(clk32MHz), 
           .D(n24005));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i102 (.Q(\data_out_frame[12] [5]), .C(clk32MHz), 
           .D(n24004));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i103 (.Q(\data_out_frame[12] [6]), .C(clk32MHz), 
           .D(n24003));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_0___i12 (.Q(\data_in[1] [3]), .C(clk32MHz), .D(n24089));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i104 (.Q(\data_out_frame[12] [7]), .C(clk32MHz), 
           .D(n24002));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i105 (.Q(\data_out_frame[13] [0]), .C(clk32MHz), 
           .D(n24001));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i106 (.Q(\data_out_frame[13] [1]), .C(clk32MHz), 
           .D(n24000));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i107 (.Q(\data_out_frame[13] [2]), .C(clk32MHz), 
           .D(n23999));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_0___i13 (.Q(\data_in[1] [4]), .C(clk32MHz), .D(n24088));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_0___i14 (.Q(\data_in[1] [5]), .C(clk32MHz), .D(n24087));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i108 (.Q(\data_out_frame[13] [3]), .C(clk32MHz), 
           .D(n23998));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i109 (.Q(\data_out_frame[13] [4]), .C(clk32MHz), 
           .D(n23997));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i110 (.Q(\data_out_frame[13] [5]), .C(clk32MHz), 
           .D(n23996));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i1_2_lut_3_lut_4_lut (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(n40205), .I3(\FRAME_MATCHER.i [0]), .O(n40207));   // verilog/coms.v(154[7:23])
    defparam i1_2_lut_3_lut_4_lut.LUT_INIT = 16'hfbff;
    SB_DFF data_out_frame_0___i111 (.Q(\data_out_frame[13] [6]), .C(clk32MHz), 
           .D(n23995));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i60 (.Q(\data_out_frame[7] [3]), .C(clk32MHz), 
           .D(n24046));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i112 (.Q(\data_out_frame[13] [7]), .C(clk32MHz), 
           .D(n23994));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i113 (.Q(\data_out_frame[14] [0]), .C(clk32MHz), 
           .D(n23993));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i114 (.Q(\data_out_frame[14] [1]), .C(clk32MHz), 
           .D(n23992));   // verilog/coms.v(126[12] 289[6])
    SB_DFF \FRAME_MATCHER.rx_data_ready_prev_3228  (.Q(\FRAME_MATCHER.rx_data_ready_prev ), 
           .C(clk32MHz), .D(rx_data_ready));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 add_44_17_lut (.I0(n1498), .I1(\FRAME_MATCHER.i [15]), .I2(GND_net), 
            .I3(n34038), .O(n2_adj_3121)) /* synthesis syn_instantiated=1 */ ;
    defparam add_44_17_lut.LUT_INIT = 16'h8228;
    SB_DFF data_out_frame_0___i115 (.Q(\data_out_frame[14] [2]), .C(clk32MHz), 
           .D(n23991));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i116 (.Q(\data_out_frame[14] [3]), .C(clk32MHz), 
           .D(n23990));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i10625_3_lut_4_lut (.I0(\FRAME_MATCHER.state [2]), .I1(n22338), 
            .I2(encoder0_position[14]), .I3(\data_out_frame[7] [6]), .O(n24043));
    defparam i10625_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_DFF data_out_frame_0___i117 (.Q(\data_out_frame[14] [4]), .C(clk32MHz), 
           .D(n23989));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i10525_3_lut_4_lut (.I0(\FRAME_MATCHER.state [2]), .I1(n22338), 
            .I2(displacement[2]), .I3(\data_out_frame[20] [2]), .O(n23943));
    defparam i10525_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_DFF data_out_frame_0___i118 (.Q(\data_out_frame[14] [5]), .C(clk32MHz), 
           .D(n23988));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i119 (.Q(\data_out_frame[14] [6]), .C(clk32MHz), 
           .D(n23987));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_0___i15 (.Q(\data_in[1] [6]), .C(clk32MHz), .D(n24086));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i120 (.Q(\data_out_frame[14] [7]), .C(clk32MHz), 
           .D(n23986));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i121 (.Q(\data_out_frame[15] [0]), .C(clk32MHz), 
           .D(n23985));   // verilog/coms.v(126[12] 289[6])
    SB_DFF Kp_i7 (.Q(\Kp[7] ), .C(clk32MHz), .D(n24137));   // verilog/coms.v(126[12] 289[6])
    SB_DFF Ki_i1 (.Q(\Ki[1] ), .C(clk32MHz), .D(n24136));   // verilog/coms.v(126[12] 289[6])
    SB_DFF Kd_i6 (.Q(\Kd[6] ), .C(clk32MHz), .D(n24124));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i122 (.Q(\data_out_frame[15] [1]), .C(clk32MHz), 
           .D(n23984));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_0___i16 (.Q(\data_in[1] [7]), .C(clk32MHz), .D(n24085));   // verilog/coms.v(126[12] 289[6])
    SB_DFF IntegralLimit_i0_i8 (.Q(IntegralLimit[8]), .C(clk32MHz), .D(n24162));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i123 (.Q(\data_out_frame[15] [2]), .C(clk32MHz), 
           .D(n23983));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i124 (.Q(\data_out_frame[15] [3]), .C(clk32MHz), 
           .D(n23982));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i125 (.Q(\data_out_frame[15] [4]), .C(clk32MHz), 
           .D(n23981));   // verilog/coms.v(126[12] 289[6])
    SB_DFF IntegralLimit_i0_i9 (.Q(IntegralLimit[9]), .C(clk32MHz), .D(n24161));   // verilog/coms.v(126[12] 289[6])
    SB_DFF IntegralLimit_i0_i10 (.Q(IntegralLimit[10]), .C(clk32MHz), .D(n24160));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i126 (.Q(\data_out_frame[15] [5]), .C(clk32MHz), 
           .D(n23980));   // verilog/coms.v(126[12] 289[6])
    SB_DFF IntegralLimit_i0_i11 (.Q(IntegralLimit[11]), .C(clk32MHz), .D(n24159));   // verilog/coms.v(126[12] 289[6])
    SB_DFF IntegralLimit_i0_i12 (.Q(IntegralLimit[12]), .C(clk32MHz), .D(n24158));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i127 (.Q(\data_out_frame[15] [6]), .C(clk32MHz), 
           .D(n23979));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i128 (.Q(\data_out_frame[15] [7]), .C(clk32MHz), 
           .D(n23978));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i129 (.Q(\data_out_frame[16] [0]), .C(clk32MHz), 
           .D(n23977));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i130 (.Q(\data_out_frame[16] [1]), .C(clk32MHz), 
           .D(n23976));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i131 (.Q(\data_out_frame[16] [2]), .C(clk32MHz), 
           .D(n23975));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i132 (.Q(\data_out_frame[16] [3]), .C(clk32MHz), 
           .D(n23974));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i133 (.Q(\data_out_frame[16] [4]), .C(clk32MHz), 
           .D(n23973));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i134 (.Q(\data_out_frame[16] [5]), .C(clk32MHz), 
           .D(n23972));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i135 (.Q(\data_out_frame[16] [6]), .C(clk32MHz), 
           .D(n23971));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i136 (.Q(\data_out_frame[16] [7]), .C(clk32MHz), 
           .D(n23970));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i137 (.Q(\data_out_frame[17] [0]), .C(clk32MHz), 
           .D(n23969));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i138 (.Q(\data_out_frame[17] [1]), .C(clk32MHz), 
           .D(n23968));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i139 (.Q(\data_out_frame[17] [2]), .C(clk32MHz), 
           .D(n23967));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i140 (.Q(\data_out_frame[17] [3]), .C(clk32MHz), 
           .D(n23966));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i141 (.Q(\data_out_frame[17] [4]), .C(clk32MHz), 
           .D(n23965));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i142 (.Q(\data_out_frame[17] [5]), .C(clk32MHz), 
           .D(n23964));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i143 (.Q(\data_out_frame[17] [6]), .C(clk32MHz), 
           .D(n23963));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i144 (.Q(\data_out_frame[17] [7]), .C(clk32MHz), 
           .D(n23962));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i145 (.Q(\data_out_frame[18] [0]), .C(clk32MHz), 
           .D(n23961));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i146 (.Q(\data_out_frame[18] [1]), .C(clk32MHz), 
           .D(n23960));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i147 (.Q(\data_out_frame[18] [2]), .C(clk32MHz), 
           .D(n23959));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i148 (.Q(\data_out_frame[18][3] ), .C(clk32MHz), 
           .D(n23958));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i1_2_lut_3_lut (.I0(\data_in_frame[6] [5]), .I1(\data_in_frame[6] [4]), 
            .I2(\data_in_frame[8] [6]), .I3(GND_net), .O(n40619));   // verilog/coms.v(72[16:43])
    defparam i1_2_lut_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 i10353_3_lut_4_lut (.I0(n8), .I1(n40205), .I2(rx_data[7]), 
            .I3(\data_in_frame[20] [7]), .O(n23771));
    defparam i10353_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10354_3_lut_4_lut (.I0(n8), .I1(n40205), .I2(rx_data[6]), 
            .I3(\data_in_frame[20] [6]), .O(n23772));
    defparam i10354_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10355_3_lut_4_lut (.I0(n8), .I1(n40205), .I2(rx_data[5]), 
            .I3(\data_in_frame[20] [5]), .O(n23773));
    defparam i10355_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10356_3_lut_4_lut (.I0(n8), .I1(n40205), .I2(rx_data[4]), 
            .I3(\data_in_frame[20] [4]), .O(n23774));
    defparam i10356_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF data_out_frame_0___i149 (.Q(\data_out_frame[18] [4]), .C(clk32MHz), 
           .D(n23957));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i150 (.Q(\data_out_frame[18] [5]), .C(clk32MHz), 
           .D(n23956));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i151 (.Q(\data_out_frame[18] [6]), .C(clk32MHz), 
           .D(n23955));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i152 (.Q(\data_out_frame[18] [7]), .C(clk32MHz), 
           .D(n23954));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i17_2_lut (.I0(rx_data_ready), .I1(\FRAME_MATCHER.rx_data_ready_prev ), 
            .I2(GND_net), .I3(GND_net), .O(n164));   // verilog/coms.v(153[9:50])
    defparam i17_2_lut.LUT_INIT = 16'h2222;
    SB_DFF data_out_frame_0___i153 (.Q(\data_out_frame[19] [0]), .C(clk32MHz), 
           .D(n23953));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 equal_53_i9_2_lut (.I0(\FRAME_MATCHER.i [4]), .I1(\FRAME_MATCHER.i [5]), 
            .I2(GND_net), .I3(GND_net), .O(n9));   // verilog/coms.v(154[7:23])
    defparam equal_53_i9_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i10465_3_lut_4_lut (.I0(n8_adj_3122), .I1(n40212), .I2(rx_data[7]), 
            .I3(\data_in_frame[6] [7]), .O(n23883));
    defparam i10465_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10466_3_lut_4_lut (.I0(n8_adj_3122), .I1(n40212), .I2(rx_data[6]), 
            .I3(\data_in_frame[6] [6]), .O(n23884));
    defparam i10466_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF data_out_frame_0___i154 (.Q(\data_out_frame[19] [1]), .C(clk32MHz), 
           .D(n23952));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i10467_3_lut_4_lut (.I0(n8_adj_3122), .I1(n40212), .I2(rx_data[5]), 
            .I3(\data_in_frame[6] [5]), .O(n23885));
    defparam i10467_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF data_out_frame_0___i155 (.Q(\data_out_frame[19] [2]), .C(clk32MHz), 
           .D(n23951));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i156 (.Q(\data_out_frame[19][3] ), .C(clk32MHz), 
           .D(n23950));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i157 (.Q(\data_out_frame[19] [4]), .C(clk32MHz), 
           .D(n23949));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i158 (.Q(\data_out_frame[19] [5]), .C(clk32MHz), 
           .D(n23948));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i10468_3_lut_4_lut (.I0(n8_adj_3122), .I1(n40212), .I2(rx_data[4]), 
            .I3(\data_in_frame[6] [4]), .O(n23886));
    defparam i10468_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF data_out_frame_0___i159 (.Q(\data_out_frame[19] [6]), .C(clk32MHz), 
           .D(n23947));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i10469_3_lut_4_lut (.I0(n8_adj_3122), .I1(n40212), .I2(rx_data[3]), 
            .I3(\data_in_frame[6] [3]), .O(n23887));
    defparam i10469_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF data_out_frame_0___i160 (.Q(\data_out_frame[19] [7]), .C(clk32MHz), 
           .D(n23946));   // verilog/coms.v(126[12] 289[6])
    SB_DFF IntegralLimit_i0_i13 (.Q(IntegralLimit[13]), .C(clk32MHz), .D(n24157));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i10357_3_lut_4_lut (.I0(n8), .I1(n40205), .I2(rx_data[3]), 
            .I3(\data_in_frame[20] [3]), .O(n23775));
    defparam i10357_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF data_out_frame_0___i161 (.Q(\data_out_frame[20] [0]), .C(clk32MHz), 
           .D(n23945));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i162 (.Q(\data_out_frame[20] [1]), .C(clk32MHz), 
           .D(n23944));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i163 (.Q(\data_out_frame[20] [2]), .C(clk32MHz), 
           .D(n23943));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i164 (.Q(\data_out_frame[20] [3]), .C(clk32MHz), 
           .D(n23942));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i165 (.Q(\data_out_frame[20] [4]), .C(clk32MHz), 
           .D(n23941));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i166 (.Q(\data_out_frame[20] [5]), .C(clk32MHz), 
           .D(n23940));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i167 (.Q(\data_out_frame[20] [6]), .C(clk32MHz), 
           .D(n23939));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i168 (.Q(\data_out_frame[20][7] ), .C(clk32MHz), 
           .D(n23938));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i2 (.Q(\data_in_frame[0] [1]), .C(clk32MHz), 
           .D(n23937));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i3 (.Q(\data_in_frame[0] [2]), .C(clk32MHz), 
           .D(n23936));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i4 (.Q(\data_in_frame[0] [3]), .C(clk32MHz), 
           .D(n23935));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i10358_3_lut_4_lut (.I0(n8), .I1(n40205), .I2(rx_data[2]), 
            .I3(\data_in_frame[20] [2]), .O(n23776));
    defparam i10358_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF data_in_frame_0__i5 (.Q(\data_in_frame[0] [4]), .C(clk32MHz), 
           .D(n23934));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i61 (.Q(\data_out_frame[7] [4]), .C(clk32MHz), 
           .D(n24045));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i6 (.Q(\data_in_frame[0] [5]), .C(clk32MHz), 
           .D(n23933));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i10359_3_lut_4_lut (.I0(n8), .I1(n40205), .I2(rx_data[1]), 
            .I3(\data_in_frame[20] [1]), .O(n23777));
    defparam i10359_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF IntegralLimit_i0_i14 (.Q(IntegralLimit[14]), .C(clk32MHz), .D(n24156));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i7 (.Q(\data_in_frame[0] [6]), .C(clk32MHz), 
           .D(n23932));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i8 (.Q(\data_in_frame[0] [7]), .C(clk32MHz), 
           .D(n23931));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i9 (.Q(\data_in_frame[1] [0]), .C(clk32MHz), 
           .D(n23930));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i10470_3_lut_4_lut (.I0(n8_adj_3122), .I1(n40212), .I2(rx_data[2]), 
            .I3(\data_in_frame[6] [2]), .O(n23888));
    defparam i10470_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF data_in_frame_0__i10 (.Q(\data_in_frame[1] [1]), .C(clk32MHz), 
           .D(n23929));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i11 (.Q(\data_in_frame[1] [2]), .C(clk32MHz), 
           .D(n23928));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i12 (.Q(\data_in_frame[1] [3]), .C(clk32MHz), 
           .D(n23927));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i13 (.Q(\data_in_frame[1] [4]), .C(clk32MHz), 
           .D(n23926));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i10471_3_lut_4_lut (.I0(n8_adj_3122), .I1(n40212), .I2(rx_data[1]), 
            .I3(\data_in_frame[6][1] ), .O(n23889));
    defparam i10471_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10472_3_lut_4_lut (.I0(n8_adj_3122), .I1(n40212), .I2(rx_data[0]), 
            .I3(\data_in_frame[6][0] ), .O(n23890));
    defparam i10472_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13817_3_lut_4_lut (.I0(n27747), .I1(n40212), .I2(\data_in_frame[7] [7]), 
            .I3(rx_data[7]), .O(n23875));
    defparam i13817_3_lut_4_lut.LUT_INIT = 16'hf2d0;
    SB_LUT4 i10458_3_lut_4_lut (.I0(n27747), .I1(n40212), .I2(rx_data[6]), 
            .I3(\data_in_frame[7] [6]), .O(n23876));
    defparam i10458_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i10459_3_lut_4_lut (.I0(n27747), .I1(n40212), .I2(rx_data[5]), 
            .I3(\data_in_frame[7] [5]), .O(n23877));
    defparam i10459_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i10460_3_lut_4_lut (.I0(n27747), .I1(n40212), .I2(rx_data[4]), 
            .I3(\data_in_frame[7] [4]), .O(n23878));
    defparam i10460_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF data_in_frame_0__i14 (.Q(\data_in_frame[1] [5]), .C(clk32MHz), 
           .D(n23925));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i10461_3_lut_4_lut (.I0(n27747), .I1(n40212), .I2(rx_data[3]), 
            .I3(\data_in_frame[7] [3]), .O(n23879));
    defparam i10461_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF data_in_frame_0__i15 (.Q(\data_in_frame[1] [6]), .C(clk32MHz), 
           .D(n23924));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i16 (.Q(\data_in_frame[1] [7]), .C(clk32MHz), 
           .D(n23923));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i2_3_lut_adj_840 (.I0(\data_in_frame[13] [7]), .I1(n40591), 
            .I2(\data_in_frame[9] [3]), .I3(GND_net), .O(n41901));
    defparam i2_3_lut_adj_840.LUT_INIT = 16'h9696;
    SB_LUT4 i10462_3_lut_4_lut (.I0(n27747), .I1(n40212), .I2(rx_data[2]), 
            .I3(\data_in_frame[7] [2]), .O(n23880));
    defparam i10462_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF data_in_frame_0__i17 (.Q(\data_in_frame[2] [0]), .C(clk32MHz), 
           .D(n23922));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i18 (.Q(\data_in_frame[2] [1]), .C(clk32MHz), 
           .D(n23921));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i10463_3_lut_4_lut (.I0(n27747), .I1(n40212), .I2(rx_data[1]), 
            .I3(\data_in_frame[7] [1]), .O(n23881));
    defparam i10463_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF data_in_frame_0__i19 (.Q(\data_in_frame[2] [2]), .C(clk32MHz), 
           .D(n23920));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i20 (.Q(\data_in_frame[2] [3]), .C(clk32MHz), 
           .D(n23919));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i21 (.Q(\data_in_frame[2] [4]), .C(clk32MHz), 
           .D(n23918));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i10360_3_lut_4_lut (.I0(n8), .I1(n40205), .I2(rx_data[0]), 
            .I3(\data_in_frame[20] [0]), .O(n23778));
    defparam i10360_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10464_3_lut_4_lut (.I0(n27747), .I1(n40212), .I2(rx_data[0]), 
            .I3(\data_in_frame[7] [0]), .O(n23882));
    defparam i10464_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF data_in_frame_0__i22 (.Q(\data_in_frame[2] [5]), .C(clk32MHz), 
           .D(n23917));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i10449_3_lut_4_lut (.I0(n8_adj_3123), .I1(n40221), .I2(rx_data[7]), 
            .I3(\data_in_frame[8] [7]), .O(n23867));
    defparam i10449_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF data_in_frame_0__i23 (.Q(\data_in_frame[2] [6]), .C(clk32MHz), 
           .D(n23916));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i24 (.Q(\data_in_frame[2] [7]), .C(clk32MHz), 
           .D(n23915));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i25 (.Q(\data_in_frame[3] [0]), .C(clk32MHz), 
           .D(n23914));   // verilog/coms.v(126[12] 289[6])
    SB_DFF IntegralLimit_i0_i15 (.Q(IntegralLimit[15]), .C(clk32MHz), .D(n24155));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i26 (.Q(\data_in_frame[3] [1]), .C(clk32MHz), 
           .D(n23913));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i27 (.Q(\data_in_frame[3] [2]), .C(clk32MHz), 
           .D(n23912));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i10450_3_lut_4_lut (.I0(n8_adj_3123), .I1(n40221), .I2(rx_data[6]), 
            .I3(\data_in_frame[8] [6]), .O(n23868));
    defparam i10450_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10451_3_lut_4_lut (.I0(n8_adj_3123), .I1(n40221), .I2(rx_data[5]), 
            .I3(\data_in_frame[8] [5]), .O(n23869));
    defparam i10451_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10452_3_lut_4_lut (.I0(n8_adj_3123), .I1(n40221), .I2(rx_data[4]), 
            .I3(\data_in_frame[8] [4]), .O(n23870));
    defparam i10452_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10453_3_lut_4_lut (.I0(n8_adj_3123), .I1(n40221), .I2(rx_data[3]), 
            .I3(\data_in_frame[8] [3]), .O(n23871));
    defparam i10453_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF data_in_frame_0__i28 (.Q(\data_in_frame[3] [3]), .C(clk32MHz), 
           .D(n23911));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i29 (.Q(\data_in_frame[3] [4]), .C(clk32MHz), 
           .D(n23910));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i30 (.Q(\data_in_frame[3] [5]), .C(clk32MHz), 
           .D(n23909));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i31 (.Q(\data_in_frame[3] [6]), .C(clk32MHz), 
           .D(n23908));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i32 (.Q(\data_in_frame[3] [7]), .C(clk32MHz), 
           .D(n23907));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i10454_3_lut_4_lut (.I0(n8_adj_3123), .I1(n40221), .I2(rx_data[2]), 
            .I3(\data_in_frame[8] [2]), .O(n23872));
    defparam i10454_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF data_in_frame_0__i33 (.Q(\data_in_frame[4] [0]), .C(clk32MHz), 
           .D(n23906));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i34 (.Q(\data_in_frame[4] [1]), .C(clk32MHz), 
           .D(n23905));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i35 (.Q(\data_in_frame[4] [2]), .C(clk32MHz), 
           .D(n23904));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i1_2_lut (.I0(\FRAME_MATCHER.state [2]), .I1(\FRAME_MATCHER.state [3]), 
            .I2(GND_net), .I3(GND_net), .O(n102));   // verilog/coms.v(126[12] 289[6])
    defparam i1_2_lut.LUT_INIT = 16'h2222;
    SB_DFF data_in_frame_0__i36 (.Q(\data_in_frame[4] [3]), .C(clk32MHz), 
           .D(n23903));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i37 (.Q(\data_in_frame[4] [4]), .C(clk32MHz), 
           .D(n23902));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i38 (.Q(\data_in_frame[4] [5]), .C(clk32MHz), 
           .D(n23901));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i39 (.Q(\data_in_frame[4] [6]), .C(clk32MHz), 
           .D(n23900));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i10455_3_lut_4_lut (.I0(n8_adj_3123), .I1(n40221), .I2(rx_data[1]), 
            .I3(\data_in_frame[8] [1]), .O(n23873));
    defparam i10455_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF data_in_frame_0__i40 (.Q(\data_in_frame[4] [7]), .C(clk32MHz), 
           .D(n23899));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i41 (.Q(\data_in_frame[5] [0]), .C(clk32MHz), 
           .D(n23898));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i42 (.Q(\data_in_frame[5] [1]), .C(clk32MHz), 
           .D(n23897));   // verilog/coms.v(126[12] 289[6])
    SB_CARRY add_44_17 (.CI(n34038), .I0(\FRAME_MATCHER.i [15]), .I1(GND_net), 
            .CO(n34039));
    SB_DFF data_in_frame_0__i43 (.Q(\data_in_frame[5] [2]), .C(clk32MHz), 
           .D(n23896));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i10456_3_lut_4_lut (.I0(n8_adj_3123), .I1(n40221), .I2(rx_data[0]), 
            .I3(\data_in_frame[8] [0]), .O(n23874));
    defparam i10456_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_CARRY add_44_7 (.CI(n34028), .I0(\FRAME_MATCHER.i [5]), .I1(GND_net), 
            .CO(n34029));
    SB_LUT4 i10433_3_lut_4_lut (.I0(n8_adj_3124), .I1(n40221), .I2(rx_data[7]), 
            .I3(\data_in_frame[10] [7]), .O(n23851));
    defparam i10433_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF data_in_frame_0__i44 (.Q(\data_in_frame[5] [3]), .C(clk32MHz), 
           .D(n23895));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i10434_3_lut_4_lut (.I0(n8_adj_3124), .I1(n40221), .I2(rx_data[6]), 
            .I3(\data_in_frame[10] [6]), .O(n23852));
    defparam i10434_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_841 (.I0(\data_in_frame[16] [3]), .I1(n40515), 
            .I2(GND_net), .I3(GND_net), .O(n37274));
    defparam i1_2_lut_adj_841.LUT_INIT = 16'h6666;
    SB_LUT4 i10435_3_lut_4_lut (.I0(n8_adj_3124), .I1(n40221), .I2(rx_data[5]), 
            .I3(\data_in_frame[10] [5]), .O(n23853));
    defparam i10435_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF data_in_frame_0__i45 (.Q(\data_in_frame[5] [4]), .C(clk32MHz), 
           .D(n23894));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 add_44_16_lut (.I0(n1498), .I1(\FRAME_MATCHER.i [14]), .I2(GND_net), 
            .I3(n34037), .O(n2_adj_3125)) /* synthesis syn_instantiated=1 */ ;
    defparam add_44_16_lut.LUT_INIT = 16'h8228;
    SB_DFF data_in_frame_0__i46 (.Q(\data_in_frame[5] [5]), .C(clk32MHz), 
           .D(n23893));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i47 (.Q(\data_in_frame[5] [6]), .C(clk32MHz), 
           .D(n23892));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i48 (.Q(\data_in_frame[5] [7]), .C(clk32MHz), 
           .D(n23891));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i49 (.Q(\data_in_frame[6][0] ), .C(clk32MHz), 
           .D(n23890));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i50 (.Q(\data_in_frame[6][1] ), .C(clk32MHz), 
           .D(n23889));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i10436_3_lut_4_lut (.I0(n8_adj_3124), .I1(n40221), .I2(rx_data[4]), 
            .I3(\data_in_frame[10] [4]), .O(n23854));
    defparam i10436_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF data_in_frame_0__i51 (.Q(\data_in_frame[6] [2]), .C(clk32MHz), 
           .D(n23888));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i52 (.Q(\data_in_frame[6] [3]), .C(clk32MHz), 
           .D(n23887));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i53 (.Q(\data_in_frame[6] [4]), .C(clk32MHz), 
           .D(n23886));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i54 (.Q(\data_in_frame[6] [5]), .C(clk32MHz), 
           .D(n23885));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i10437_3_lut_4_lut (.I0(n8_adj_3124), .I1(n40221), .I2(rx_data[3]), 
            .I3(\data_in_frame[10] [3]), .O(n23855));
    defparam i10437_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF data_in_frame_0__i55 (.Q(\data_in_frame[6] [6]), .C(clk32MHz), 
           .D(n23884));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i10438_3_lut_4_lut (.I0(n8_adj_3124), .I1(n40221), .I2(rx_data[2]), 
            .I3(\data_in_frame[10] [2]), .O(n23856));
    defparam i10438_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF data_in_frame_0__i56 (.Q(\data_in_frame[6] [7]), .C(clk32MHz), 
           .D(n23883));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i10439_3_lut_4_lut (.I0(n8_adj_3124), .I1(n40221), .I2(rx_data[1]), 
            .I3(\data_in_frame[10] [1]), .O(n23857));
    defparam i10439_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF data_in_frame_0__i57 (.Q(\data_in_frame[7] [0]), .C(clk32MHz), 
           .D(n23882));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i58 (.Q(\data_in_frame[7] [1]), .C(clk32MHz), 
           .D(n23881));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i59 (.Q(\data_in_frame[7] [2]), .C(clk32MHz), 
           .D(n23880));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i10440_3_lut_4_lut (.I0(n8_adj_3124), .I1(n40221), .I2(rx_data[0]), 
            .I3(\data_in_frame[10] [0]), .O(n23858));
    defparam i10440_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF data_in_frame_0__i60 (.Q(\data_in_frame[7] [3]), .C(clk32MHz), 
           .D(n23879));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i61 (.Q(\data_in_frame[7] [4]), .C(clk32MHz), 
           .D(n23878));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i62 (.Q(\data_in_frame[7] [5]), .C(clk32MHz), 
           .D(n23877));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i63 (.Q(\data_in_frame[7] [6]), .C(clk32MHz), 
           .D(n23876));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i64 (.Q(\data_in_frame[7] [7]), .C(clk32MHz), 
           .D(n23875));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i65 (.Q(\data_in_frame[8] [0]), .C(clk32MHz), 
           .D(n23874));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i10417_3_lut_4_lut (.I0(n8), .I1(n40221), .I2(rx_data[7]), 
            .I3(\data_in_frame[12] [7]), .O(n23835));
    defparam i10417_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10418_3_lut_4_lut (.I0(n8), .I1(n40221), .I2(rx_data[6]), 
            .I3(\data_in_frame[12] [6]), .O(n23836));
    defparam i10418_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10419_3_lut_4_lut (.I0(n8), .I1(n40221), .I2(rx_data[5]), 
            .I3(\data_in_frame[12] [5]), .O(n23837));
    defparam i10419_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF data_in_frame_0__i66 (.Q(\data_in_frame[8] [1]), .C(clk32MHz), 
           .D(n23873));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i10420_3_lut_4_lut (.I0(n8), .I1(n40221), .I2(rx_data[4]), 
            .I3(\data_in_frame[12] [4]), .O(n23838));
    defparam i10420_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF data_in_frame_0__i67 (.Q(\data_in_frame[8] [2]), .C(clk32MHz), 
           .D(n23872));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i10421_3_lut_4_lut (.I0(n8), .I1(n40221), .I2(rx_data[3]), 
            .I3(\data_in_frame[12] [3]), .O(n23839));
    defparam i10421_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF data_in_frame_0__i68 (.Q(\data_in_frame[8] [3]), .C(clk32MHz), 
           .D(n23871));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i10422_3_lut_4_lut (.I0(n8), .I1(n40221), .I2(rx_data[2]), 
            .I3(\data_in_frame[12] [2]), .O(n23840));
    defparam i10422_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10423_3_lut_4_lut (.I0(n8), .I1(n40221), .I2(rx_data[1]), 
            .I3(\data_in_frame[12][1] ), .O(n23841));
    defparam i10423_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10424_3_lut_4_lut (.I0(n8), .I1(n40221), .I2(rx_data[0]), 
            .I3(\data_in_frame[12][0] ), .O(n23842));
    defparam i10424_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_4_lut (.I0(\data_in_frame[16] [0]), .I1(Kp_23__N_908), 
            .I2(\data_in_frame[15] [5]), .I3(n37237), .O(n6));
    defparam i1_2_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i4_2_lut_4_lut (.I0(\data_in_frame[16] [0]), .I1(Kp_23__N_908), 
            .I2(\data_in_frame[15] [5]), .I3(n22648), .O(n15));
    defparam i4_2_lut_4_lut.LUT_INIT = 16'h6996;
    SB_DFF data_in_frame_0__i69 (.Q(\data_in_frame[8] [4]), .C(clk32MHz), 
           .D(n23870));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i3_4_lut (.I0(\data_in_frame[6] [7]), .I1(\data_in_frame[7] [1]), 
            .I2(n41901), .I3(n23101), .O(n40831));
    defparam i3_4_lut.LUT_INIT = 16'h6996;
    SB_DFF data_in_frame_0__i70 (.Q(\data_in_frame[8] [5]), .C(clk32MHz), 
           .D(n23869));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i71 (.Q(\data_in_frame[8] [6]), .C(clk32MHz), 
           .D(n23868));   // verilog/coms.v(126[12] 289[6])
    SB_DFF IntegralLimit_i0_i16 (.Q(IntegralLimit[16]), .C(clk32MHz), .D(n24151));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i72 (.Q(\data_in_frame[8] [7]), .C(clk32MHz), 
           .D(n23867));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i1_2_lut_4_lut_adj_842 (.I0(n40773), .I1(n10), .I2(\data_in_frame[14] [4]), 
            .I3(\data_in_frame[16] [5]), .O(n40570));
    defparam i1_2_lut_4_lut_adj_842.LUT_INIT = 16'h6996;
    SB_DFF data_in_frame_0__i73 (.Q(\data_in_frame[9] [0]), .C(clk32MHz), 
           .D(n23866));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i1_2_lut_4_lut_adj_843 (.I0(n40773), .I1(n10), .I2(\data_in_frame[14] [4]), 
            .I3(n36853), .O(n37336));
    defparam i1_2_lut_4_lut_adj_843.LUT_INIT = 16'h6996;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_0_i19_3_lut (.I0(\data_out_frame[20] [0]), 
            .I1(\data_out_frame[21] [0]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n19));   // verilog/coms.v(104[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_0_i19_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i28918_4_lut (.I0(byte_transmit_counter[0]), .I1(\data_out_frame[5] [0]), 
            .I2(byte_transmit_counter[1]), .I3(byte_transmit_counter_c[2]), 
            .O(n44438));   // verilog/coms.v(104[34:55])
    defparam i28918_4_lut.LUT_INIT = 16'h880a;
    SB_DFF data_in_frame_0__i74 (.Q(\data_in_frame[9] [1]), .C(clk32MHz), 
           .D(n23865));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i75 (.Q(\data_in_frame[9] [2]), .C(clk32MHz), 
           .D(n23864));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i76 (.Q(\data_in_frame[9] [3]), .C(clk32MHz), 
           .D(n23863));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_0_i5_3_lut (.I0(\data_out_frame[6] [0]), 
            .I1(\data_out_frame[7] [0]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n5));   // verilog/coms.v(104[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_0_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i26715_4_lut (.I0(n19), .I1(\data_out_frame[22] [0]), .I2(byte_transmit_counter[1]), 
            .I3(byte_transmit_counter[0]), .O(n42234));
    defparam i26715_4_lut.LUT_INIT = 16'h0aca;
    SB_DFF data_in_frame_0__i77 (.Q(\data_in_frame[9] [4]), .C(clk32MHz), 
           .D(n23862));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i78 (.Q(\data_in_frame[9] [5]), .C(clk32MHz), 
           .D(n23861));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i26716_3_lut (.I0(n46934), .I1(n42234), .I2(byte_transmit_counter_c[2]), 
            .I3(GND_net), .O(n42235));
    defparam i26716_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i26687_4_lut (.I0(n5), .I1(n44438), .I2(byte_transmit_counter_c[2]), 
            .I3(byte_transmit_counter[1]), .O(n42206));
    defparam i26687_4_lut.LUT_INIT = 16'haccc;
    SB_LUT4 i26689_4_lut (.I0(n42206), .I1(n42235), .I2(byte_transmit_counter_c[4]), 
            .I3(byte_transmit_counter_c[3]), .O(n42208));
    defparam i26689_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i26688_3_lut (.I0(n46988), .I1(n47018), .I2(byte_transmit_counter_c[2]), 
            .I3(GND_net), .O(n42207));
    defparam i26688_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 n47003_bdd_4_lut_4_lut (.I0(\data_out_frame[0][4] ), .I1(byte_transmit_counter[0]), 
            .I2(byte_transmit_counter_c[2]), .I3(n47003), .O(n47006));
    defparam n47003_bdd_4_lut_4_lut.LUT_INIT = 16'hfc02;
    SB_DFF data_in_frame_0__i79 (.Q(\data_in_frame[9] [6]), .C(clk32MHz), 
           .D(n23860));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i80 (.Q(\data_in_frame[9] [7]), .C(clk32MHz), 
           .D(n23859));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i81 (.Q(\data_in_frame[10] [0]), .C(clk32MHz), 
           .D(n23858));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i82 (.Q(\data_in_frame[10] [1]), .C(clk32MHz), 
           .D(n23857));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i83 (.Q(\data_in_frame[10] [2]), .C(clk32MHz), 
           .D(n23856));   // verilog/coms.v(126[12] 289[6])
    SB_CARRY add_44_16 (.CI(n34037), .I0(\FRAME_MATCHER.i [14]), .I1(GND_net), 
            .CO(n34038));
    SB_DFF data_in_frame_0__i84 (.Q(\data_in_frame[10] [3]), .C(clk32MHz), 
           .D(n23855));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i85 (.Q(\data_in_frame[10] [4]), .C(clk32MHz), 
           .D(n23854));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i86 (.Q(\data_in_frame[10] [5]), .C(clk32MHz), 
           .D(n23853));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i87 (.Q(\data_in_frame[10] [6]), .C(clk32MHz), 
           .D(n23852));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i88 (.Q(\data_in_frame[10] [7]), .C(clk32MHz), 
           .D(n23851));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i89 (.Q(\data_in_frame[11] [0]), .C(clk32MHz), 
           .D(n23850));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i90 (.Q(\data_in_frame[11] [1]), .C(clk32MHz), 
           .D(n23849));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i91 (.Q(\data_in_frame[11] [2]), .C(clk32MHz), 
           .D(n23848));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i92 (.Q(\data_in_frame[11] [3]), .C(clk32MHz), 
           .D(n23847));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i93 (.Q(\data_in_frame[11] [4]), .C(clk32MHz), 
           .D(n23846));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i94 (.Q(\data_in_frame[11] [5]), .C(clk32MHz), 
           .D(n23845));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i95 (.Q(\data_in_frame[11] [6]), .C(clk32MHz), 
           .D(n23844));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 add_44_6_lut (.I0(n1498), .I1(\FRAME_MATCHER.i [4]), .I2(GND_net), 
            .I3(n34027), .O(n2_adj_3126)) /* synthesis syn_instantiated=1 */ ;
    defparam add_44_6_lut.LUT_INIT = 16'h8228;
    SB_LUT4 add_44_15_lut (.I0(n1498), .I1(\FRAME_MATCHER.i [13]), .I2(GND_net), 
            .I3(n34036), .O(n2_adj_3127)) /* synthesis syn_instantiated=1 */ ;
    defparam add_44_15_lut.LUT_INIT = 16'h8228;
    SB_DFF data_in_frame_0__i96 (.Q(\data_in_frame[11] [7]), .C(clk32MHz), 
           .D(n23843));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i97 (.Q(\data_in_frame[12][0] ), .C(clk32MHz), 
           .D(n23842));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i98 (.Q(\data_in_frame[12][1] ), .C(clk32MHz), 
           .D(n23841));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i99 (.Q(\data_in_frame[12] [2]), .C(clk32MHz), 
           .D(n23840));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i100 (.Q(\data_in_frame[12] [3]), .C(clk32MHz), 
           .D(n23839));   // verilog/coms.v(126[12] 289[6])
    SB_DFF IntegralLimit_i0_i17 (.Q(IntegralLimit[17]), .C(clk32MHz), .D(n24150));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i3_4_lut_adj_844 (.I0(\data_in_frame[11] [5]), .I1(n40831), 
            .I2(n40782), .I3(n40644), .O(n37268));
    defparam i3_4_lut_adj_844.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_845 (.I0(\data_in_frame[7] [2]), .I1(\data_in_frame[4] [6]), 
            .I2(\data_in_frame[7] [3]), .I3(GND_net), .O(n40858));
    defparam i2_3_lut_adj_845.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_adj_846 (.I0(\data_in_frame[11] [6]), .I1(n40858), 
            .I2(\data_in_frame[9] [4]), .I3(GND_net), .O(n40318));
    defparam i2_3_lut_adj_846.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_847 (.I0(\data_in_frame[3] [7]), .I1(\data_in_frame[3] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n40503));   // verilog/coms.v(83[17:28])
    defparam i1_2_lut_adj_847.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_848 (.I0(\data_in_frame[4] [0]), .I1(n40503), .I2(\data_in_frame[1] [6]), 
            .I3(\data_in_frame[1] [4]), .O(n23275));   // verilog/coms.v(83[17:28])
    defparam i3_4_lut_adj_848.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_849 (.I0(\data_in_frame[8] [2]), .I1(Kp_23__N_379), 
            .I2(n23275), .I3(GND_net), .O(n40481));   // verilog/coms.v(70[16:41])
    defparam i2_3_lut_adj_849.LUT_INIT = 16'h9696;
    SB_LUT4 i3_4_lut_adj_850 (.I0(\data_in_frame[1] [3]), .I1(\data_in_frame[1] [5]), 
            .I2(\data_in_frame[3] [6]), .I3(\data_in_frame[3] [5]), .O(Kp_23__N_379));   // verilog/coms.v(75[16:43])
    defparam i3_4_lut_adj_850.LUT_INIT = 16'h6996;
    SB_LUT4 equal_1013_i8_2_lut (.I0(Kp_23__N_379), .I1(\data_in_frame[5] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n8_adj_3128));   // verilog/coms.v(230[9:81])
    defparam equal_1013_i8_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_851 (.I0(\data_in_frame[14] [5]), .I1(n40779), 
            .I2(n40584), .I3(n22842), .O(n40752));
    defparam i3_4_lut_adj_851.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut (.I0(n40481), .I1(\data_in_frame[5] [7]), .I2(\data_in_frame[10] [3]), 
            .I3(\data_in_frame[8] [0]), .O(n14));
    defparam i6_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut (.I0(\data_in_frame[12] [4]), .I1(n14), .I2(n10_adj_3129), 
            .I3(n23157), .O(n22648));
    defparam i7_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_852 (.I0(n22648), .I1(n40752), .I2(GND_net), 
            .I3(GND_net), .O(n37248));
    defparam i1_2_lut_adj_852.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_853 (.I0(\data_in_frame[0] [5]), .I1(\data_in_frame[2] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n40478));   // verilog/coms.v(74[16:27])
    defparam i1_2_lut_adj_853.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_854 (.I0(\data_in_frame[0] [1]), .I1(\data_in_frame[2] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n40261));   // verilog/coms.v(166[9:87])
    defparam i1_2_lut_adj_854.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_855 (.I0(\data_in_frame[3] [5]), .I1(\data_in_frame[3] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n40708));   // verilog/coms.v(74[16:43])
    defparam i1_2_lut_adj_855.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_856 (.I0(\data_in_frame[1] [2]), .I1(\data_in_frame[1] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n40463));   // verilog/coms.v(74[16:43])
    defparam i1_2_lut_adj_856.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_857 (.I0(\data_in_frame[5] [4]), .I1(n40432), .I2(n40255), 
            .I3(\data_in_frame[1] [2]), .O(n23157));   // verilog/coms.v(76[16:27])
    defparam i3_4_lut_adj_857.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_858 (.I0(\data_in_frame[0] [6]), .I1(\data_in_frame[1] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n40432));   // verilog/coms.v(76[16:27])
    defparam i1_2_lut_adj_858.LUT_INIT = 16'h6666;
    SB_LUT4 i1_4_lut_adj_859 (.I0(\data_in_frame[5] [2]), .I1(n4_c), .I2(n6_adj_3130), 
            .I3(\data_in_frame[3] [1]), .O(n22842));
    defparam i1_4_lut_adj_859.LUT_INIT = 16'h6996;
    SB_LUT4 equal_1013_i16_2_lut (.I0(Kp_23__N_329), .I1(\data_in_frame[4] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n16));   // verilog/coms.v(230[9:81])
    defparam equal_1013_i16_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut (.I0(n16), .I1(\data_in_frame[7] [4]), .I2(n22842), 
            .I3(\data_in_frame[9] [6]), .O(n10_adj_3131));
    defparam i4_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i5_3_lut (.I0(n23157), .I1(n10_adj_3131), .I2(\data_in_frame[7] [5]), 
            .I3(GND_net), .O(n40834));
    defparam i5_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_adj_860 (.I0(\data_in_frame[1] [3]), .I1(\data_in_frame[1] [1]), 
            .I2(\data_in_frame[0] [7]), .I3(GND_net), .O(n40308));   // verilog/coms.v(71[16:34])
    defparam i2_3_lut_adj_860.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_adj_861 (.I0(\data_in_frame[3] [2]), .I1(\data_in_frame[3] [3]), 
            .I2(\data_in_frame[0] [7]), .I3(GND_net), .O(n40255));   // verilog/coms.v(71[16:34])
    defparam i2_3_lut_adj_861.LUT_INIT = 16'h9696;
    SB_LUT4 i7_4_lut_adj_862 (.I0(\data_in_frame[2] [7]), .I1(\data_in_frame[2] [3]), 
            .I2(n40383), .I3(n40478), .O(n18));   // verilog/coms.v(71[16:34])
    defparam i7_4_lut_adj_862.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_863 (.I0(n40503), .I1(\data_in_frame[1] [5]), .I2(\data_in_frame[1] [1]), 
            .I3(n40708), .O(n10_adj_3132));   // verilog/coms.v(71[16:34])
    defparam i4_4_lut_adj_863.LUT_INIT = 16'h6996;
    SB_LUT4 i9_4_lut (.I0(n40463), .I1(n18), .I2(n40261), .I3(n40432), 
            .O(n20));   // verilog/coms.v(71[16:34])
    defparam i9_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i8_4_lut (.I0(\data_in_frame[1] [7]), .I1(\data_in_frame[0] [3]), 
            .I2(n40308), .I3(Kp_23__N_326), .O(n19_adj_3133));   // verilog/coms.v(71[16:34])
    defparam i8_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_864 (.I0(n19_adj_3133), .I1(n9_adj_3134), .I2(n20), 
            .I3(n10_adj_3132), .O(n40674));
    defparam i1_4_lut_adj_864.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_865 (.I0(\data_in_frame[12][0] ), .I1(n40834), 
            .I2(\data_in_frame[11] [7]), .I3(GND_net), .O(n40644));
    defparam i2_3_lut_adj_865.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_adj_866 (.I0(n4_c), .I1(n40437), .I2(\data_in_frame[5] [0]), 
            .I3(GND_net), .O(n23290));
    defparam i2_3_lut_adj_866.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_adj_867 (.I0(\data_in_frame[9] [6]), .I1(\data_in_frame[12] [2]), 
            .I2(Kp_23__N_459), .I3(GND_net), .O(n40846));
    defparam i2_3_lut_adj_867.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_adj_868 (.I0(\data_in_frame[2] [4]), .I1(\data_in_frame[0] [2]), 
            .I2(\data_in_frame[0] [3]), .I3(GND_net), .O(n5_adj_3135));   // verilog/coms.v(166[9:87])
    defparam i2_3_lut_adj_868.LUT_INIT = 16'h9696;
    SB_DFF data_in_frame_0__i101 (.Q(\data_in_frame[12] [4]), .C(clk32MHz), 
           .D(n23838));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i2_3_lut_4_lut (.I0(\data_in_frame[8] [5]), .I1(\data_in_frame[6] [3]), 
            .I2(\data_in_frame[12] [7]), .I3(n40705), .O(n40531));   // verilog/coms.v(72[16:43])
    defparam i2_3_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_869 (.I0(\data_in_frame[8] [5]), .I1(\data_in_frame[6] [3]), 
            .I2(\data_in_frame[13] [4]), .I3(n40728), .O(n40460));   // verilog/coms.v(72[16:43])
    defparam i2_3_lut_4_lut_adj_869.LUT_INIT = 16'h6996;
    SB_DFF IntegralLimit_i0_i18 (.Q(IntegralLimit[18]), .C(clk32MHz), .D(n24149));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i3_4_lut_adj_870 (.I0(\data_in_frame[8] [0]), .I1(n40417), .I2(\data_in_frame[10] [1]), 
            .I3(n23045), .O(n40779));
    defparam i3_4_lut_adj_870.LUT_INIT = 16'h6996;
    SB_CARRY add_44_15 (.CI(n34036), .I0(\FRAME_MATCHER.i [13]), .I1(GND_net), 
            .CO(n34037));
    SB_CARRY add_44_6 (.CI(n34027), .I0(\FRAME_MATCHER.i [4]), .I1(GND_net), 
            .CO(n34028));
    SB_LUT4 add_44_14_lut (.I0(n1498), .I1(\FRAME_MATCHER.i [12]), .I2(GND_net), 
            .I3(n34035), .O(n2_adj_3136)) /* synthesis syn_instantiated=1 */ ;
    defparam add_44_14_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i2_2_lut (.I0(n40779), .I1(Kp_23__N_326), .I2(GND_net), .I3(GND_net), 
            .O(n10_adj_3137));
    defparam i2_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i6_4_lut_adj_871 (.I0(n40846), .I1(n23290), .I2(n40644), .I3(\data_in_frame[14] [2]), 
            .O(n14_adj_3138));
    defparam i6_4_lut_adj_871.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut_adj_872 (.I0(\data_in_frame[14] [3]), .I1(n14_adj_3138), 
            .I2(n10_adj_3137), .I3(n40318), .O(n37239));
    defparam i7_4_lut_adj_872.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_873 (.I0(\data_in_frame[12][0] ), .I1(n40864), 
            .I2(\data_in_frame[14] [2]), .I3(GND_net), .O(n40647));
    defparam i2_3_lut_adj_873.LUT_INIT = 16'h9696;
    SB_LUT4 i3_4_lut_adj_874 (.I0(n23045), .I1(n40647), .I2(\data_in_frame[7] [6]), 
            .I3(\data_in_frame[9] [7]), .O(n41875));
    defparam i3_4_lut_adj_874.LUT_INIT = 16'h6996;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut (.I0(byte_transmit_counter[1]), 
            .I1(n19_adj_3139), .I2(n44182), .I3(byte_transmit_counter_c[2]), 
            .O(n47021));
    defparam byte_transmit_counter_1__bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_LUT4 n47021_bdd_4_lut (.I0(n47021), .I1(n17), .I2(n16_adj_3140), 
            .I3(byte_transmit_counter_c[2]), .O(n47024));
    defparam n47021_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i3_4_lut_adj_875 (.I0(\data_in_frame[16] [4]), .I1(n40258), 
            .I2(n37239), .I3(\data_in_frame[19] [0]), .O(n23301));
    defparam i3_4_lut_adj_875.LUT_INIT = 16'h6996;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[14] [0]), .I2(\data_out_frame[15] [0]), 
            .I3(byte_transmit_counter[1]), .O(n47015));
    defparam byte_transmit_counter_0__bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_LUT4 n47015_bdd_4_lut (.I0(n47015), .I1(\data_out_frame[13] [0]), 
            .I2(\data_out_frame[12] [0]), .I3(byte_transmit_counter[1]), 
            .O(n47018));
    defparam n47015_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i6_4_lut_adj_876 (.I0(\data_in_frame[0] [7]), .I1(\data_in_frame[0] [4]), 
            .I2(\data_in_frame[0] [5]), .I3(\data_in_frame[0] [6]), .O(n14_adj_3141));
    defparam i6_4_lut_adj_876.LUT_INIT = 16'h8000;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_31475 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[18] [7]), .I2(\data_out_frame[19] [7]), 
            .I3(byte_transmit_counter[1]), .O(n47009));
    defparam byte_transmit_counter_0__bdd_4_lut_31475.LUT_INIT = 16'he4aa;
    SB_LUT4 n47009_bdd_4_lut (.I0(n47009), .I1(\data_out_frame[17] [7]), 
            .I2(\data_out_frame[16] [7]), .I3(byte_transmit_counter[1]), 
            .O(n47012));
    defparam n47009_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_31480 (.I0(byte_transmit_counter[1]), 
            .I1(n44143), .I2(n5_adj_3142), .I3(byte_transmit_counter_c[2]), 
            .O(n47003));
    defparam byte_transmit_counter_1__bdd_4_lut_31480.LUT_INIT = 16'he4aa;
    SB_LUT4 i5_4_lut (.I0(\data_in_frame[0] [0]), .I1(\data_in_frame[0] [1]), 
            .I2(\data_in_frame[0] [3]), .I3(\data_in_frame[0] [2]), .O(n13));
    defparam i5_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_31465 (.I0(byte_transmit_counter[1]), 
            .I1(n42272), .I2(n42273), .I3(byte_transmit_counter_c[2]), 
            .O(n46997));
    defparam byte_transmit_counter_1__bdd_4_lut_31465.LUT_INIT = 16'he4aa;
    SB_LUT4 n46997_bdd_4_lut (.I0(n46997), .I1(n42270), .I2(n42269), .I3(byte_transmit_counter_c[2]), 
            .O(n47000));
    defparam n46997_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_877 (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(n40221), .I3(\FRAME_MATCHER.i [0]), .O(n40227));   // verilog/coms.v(154[7:23])
    defparam i1_2_lut_3_lut_4_lut_adj_877.LUT_INIT = 16'hfbff;
    SB_DFF IntegralLimit_i0_i19 (.Q(IntegralLimit[19]), .C(clk32MHz), .D(n24148));   // verilog/coms.v(126[12] 289[6])
    SB_DFF IntegralLimit_i0_i20 (.Q(IntegralLimit[20]), .C(clk32MHz), .D(n24147));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 add_547_9_lut (.I0(n19614), .I1(byte_transmit_counter_c[7]), 
            .I2(GND_net), .I3(n34061), .O(n44012)) /* synthesis syn_instantiated=1 */ ;
    defparam add_547_9_lut.LUT_INIT = 16'h8228;
    SB_LUT4 add_547_8_lut (.I0(GND_net), .I1(byte_transmit_counter_c[6]), 
            .I2(GND_net), .I3(n34060), .O(n2236[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_547_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_547_8 (.CI(n34060), .I0(byte_transmit_counter_c[6]), .I1(GND_net), 
            .CO(n34061));
    SB_LUT4 add_547_7_lut (.I0(GND_net), .I1(byte_transmit_counter_c[5]), 
            .I2(GND_net), .I3(n34059), .O(n2236[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_547_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_547_7 (.CI(n34059), .I0(byte_transmit_counter_c[5]), .I1(GND_net), 
            .CO(n34060));
    SB_CARRY add_44_14 (.CI(n34035), .I0(\FRAME_MATCHER.i [12]), .I1(GND_net), 
            .CO(n34036));
    SB_LUT4 add_547_6_lut (.I0(GND_net), .I1(byte_transmit_counter_c[4]), 
            .I2(GND_net), .I3(n34058), .O(n2236[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_547_6_lut.LUT_INIT = 16'hC33C;
    SB_DFF data_in_frame_0__i102 (.Q(\data_in_frame[12] [5]), .C(clk32MHz), 
           .D(n23837));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i5_4_lut_adj_878 (.I0(\data_in_frame[0] [0]), .I1(\data_in_frame[0] [1]), 
            .I2(\data_in_frame[0] [3]), .I3(\data_in_frame[0] [2]), .O(n13_adj_3143));   // verilog/coms.v(232[13:35])
    defparam i5_4_lut_adj_878.LUT_INIT = 16'hfffe;
    SB_LUT4 i14290_4_lut (.I0(n13_adj_3143), .I1(n13), .I2(n14_adj_3144), 
            .I3(n14_adj_3141), .O(n27691));
    defparam i14290_4_lut.LUT_INIT = 16'h32fa;
    SB_DFF data_in_frame_0__i103 (.Q(\data_in_frame[12] [6]), .C(clk32MHz), 
           .D(n23836));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_31460 (.I0(byte_transmit_counter[1]), 
            .I1(n42278), .I2(n42279), .I3(byte_transmit_counter_c[2]), 
            .O(n46991));
    defparam byte_transmit_counter_1__bdd_4_lut_31460.LUT_INIT = 16'he4aa;
    SB_DFF data_in_frame_0__i104 (.Q(\data_in_frame[12] [7]), .C(clk32MHz), 
           .D(n23835));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 n46991_bdd_4_lut (.I0(n46991), .I1(n42276), .I2(n42275), .I3(byte_transmit_counter_c[2]), 
            .O(n46994));
    defparam n46991_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF data_in_frame_0__i105 (.Q(\data_in_frame[13] [0]), .C(clk32MHz), 
           .D(n23834));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i5_4_lut_adj_879 (.I0(\data_in_frame[18] [7]), .I1(n23301), 
            .I2(\data_in_frame[18] [5]), .I3(n37274), .O(n12));
    defparam i5_4_lut_adj_879.LUT_INIT = 16'h6996;
    SB_DFF data_in_frame_0__i106 (.Q(\data_in_frame[13] [1]), .C(clk32MHz), 
           .D(n23833));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_31470 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[10] [0]), .I2(\data_out_frame[11] [0]), 
            .I3(byte_transmit_counter[1]), .O(n46985));
    defparam byte_transmit_counter_0__bdd_4_lut_31470.LUT_INIT = 16'he4aa;
    SB_DFF data_in_frame_0__i107 (.Q(\data_in_frame[13] [2]), .C(clk32MHz), 
           .D(n23832));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 n46985_bdd_4_lut (.I0(n46985), .I1(\data_out_frame[9] [0]), 
            .I2(\data_out_frame[8] [0]), .I3(byte_transmit_counter[1]), 
            .O(n46988));
    defparam n46985_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF data_in_frame_0__i108 (.Q(\data_in_frame[13] [3]), .C(clk32MHz), 
           .D(n23831));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i4_4_lut_adj_880 (.I0(n40420), .I1(\data_in_frame[18] [3]), 
            .I2(\data_in_frame[20] [4]), .I3(n40487), .O(n10_adj_3145));
    defparam i4_4_lut_adj_880.LUT_INIT = 16'h6996;
    SB_DFF data_in_frame_0__i109 (.Q(\data_in_frame[13] [4]), .C(clk32MHz), 
           .D(n23830));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_31450 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[10] [1]), .I2(\data_out_frame[11] [1]), 
            .I3(byte_transmit_counter[1]), .O(n46979));
    defparam byte_transmit_counter_0__bdd_4_lut_31450.LUT_INIT = 16'he4aa;
    SB_DFF data_in_frame_0__i110 (.Q(\data_in_frame[13] [5]), .C(clk32MHz), 
           .D(n23829));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 n46979_bdd_4_lut (.I0(n46979), .I1(\data_out_frame[9] [1]), 
            .I2(\data_out_frame[8] [1]), .I3(byte_transmit_counter[1]), 
            .O(n46982));
    defparam n46979_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF data_in_frame_0__i111 (.Q(\data_in_frame[13] [6]), .C(clk32MHz), 
           .D(n23828));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i2_3_lut_adj_881 (.I0(\data_in_frame[18] [4]), .I1(n40398), 
            .I2(\data_in_frame[20] [6]), .I3(GND_net), .O(n41720));   // verilog/coms.v(83[17:63])
    defparam i2_3_lut_adj_881.LUT_INIT = 16'h9696;
    SB_DFF data_in_frame_0__i112 (.Q(\data_in_frame[13] [7]), .C(clk32MHz), 
           .D(n23827));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_31445 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[14] [1]), .I2(\data_out_frame[15] [1]), 
            .I3(byte_transmit_counter[1]), .O(n46973));
    defparam byte_transmit_counter_0__bdd_4_lut_31445.LUT_INIT = 16'he4aa;
    SB_DFF data_in_frame_0__i113 (.Q(\data_in_frame[14] [0]), .C(clk32MHz), 
           .D(n23826));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 n46973_bdd_4_lut (.I0(n46973), .I1(\data_out_frame[13] [1]), 
            .I2(\data_out_frame[12] [1]), .I3(byte_transmit_counter[1]), 
            .O(n46976));
    defparam n46973_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF data_in_frame_0__i114 (.Q(\data_in_frame[14] [1]), .C(clk32MHz), 
           .D(n23825));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i2_4_lut (.I0(n22997), .I1(n40746), .I2(n40554), .I3(\data_in_frame[21] [7]), 
            .O(n41390));
    defparam i2_4_lut.LUT_INIT = 16'h6996;
    SB_DFF data_in_frame_0__i115 (.Q(\data_in_frame[14] [2]), .C(clk32MHz), 
           .D(n23824));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_31440 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[10] [2]), .I2(\data_out_frame[11] [2]), 
            .I3(byte_transmit_counter[1]), .O(n46967));
    defparam byte_transmit_counter_0__bdd_4_lut_31440.LUT_INIT = 16'he4aa;
    SB_DFF data_in_frame_0__i116 (.Q(\data_in_frame[14] [3]), .C(clk32MHz), 
           .D(n23823));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 n46967_bdd_4_lut (.I0(n46967), .I1(\data_out_frame[9] [2]), 
            .I2(\data_out_frame[8] [2]), .I3(byte_transmit_counter[1]), 
            .O(n46970));
    defparam n46967_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF data_in_frame_0__i117 (.Q(\data_in_frame[14] [4]), .C(clk32MHz), 
           .D(n23822));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i5_3_lut_adj_882 (.I0(\data_in_frame[18] [2]), .I1(n10_adj_3145), 
            .I2(\data_in_frame[16] [2]), .I3(GND_net), .O(n41776));
    defparam i5_3_lut_adj_882.LUT_INIT = 16'h9696;
    SB_DFF data_in_frame_0__i118 (.Q(\data_in_frame[14] [5]), .C(clk32MHz), 
           .D(n23821));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_31435 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[14] [2]), .I2(\data_out_frame[15] [2]), 
            .I3(byte_transmit_counter[1]), .O(n46961));
    defparam byte_transmit_counter_0__bdd_4_lut_31435.LUT_INIT = 16'he4aa;
    SB_DFF data_in_frame_0__i119 (.Q(\data_in_frame[14] [6]), .C(clk32MHz), 
           .D(n23820));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 n46961_bdd_4_lut (.I0(n46961), .I1(\data_out_frame[13] [2]), 
            .I2(\data_out_frame[12] [2]), .I3(byte_transmit_counter[1]), 
            .O(n46964));
    defparam n46961_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF data_in_frame_0__i120 (.Q(\data_in_frame[14] [7]), .C(clk32MHz), 
           .D(n23819));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i6_4_lut_adj_883 (.I0(\data_in_frame[20] [7]), .I1(n12), .I2(n40570), 
            .I3(n37284), .O(n41583));
    defparam i6_4_lut_adj_883.LUT_INIT = 16'h6996;
    SB_DFF data_in_frame_0__i121 (.Q(\data_in_frame[15] [0]), .C(clk32MHz), 
           .D(n23818));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_31430 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[10] [3]), .I2(\data_out_frame[11] [3]), 
            .I3(byte_transmit_counter[1]), .O(n46955));
    defparam byte_transmit_counter_0__bdd_4_lut_31430.LUT_INIT = 16'he4aa;
    SB_DFF data_in_frame_0__i122 (.Q(\data_in_frame[15] [1]), .C(clk32MHz), 
           .D(n23817));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 n46955_bdd_4_lut (.I0(n46955), .I1(\data_out_frame[9] [3]), 
            .I2(\data_out_frame[8] [3]), .I3(byte_transmit_counter[1]), 
            .O(n46958));
    defparam n46955_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF data_in_frame_0__i123 (.Q(\data_in_frame[15] [2]), .C(clk32MHz), 
           .D(n23816));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i1_rep_11_2_lut (.I0(\data_in_frame[17] [7]), .I1(\data_in_frame[17] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n47038));
    defparam i1_rep_11_2_lut.LUT_INIT = 16'h6666;
    SB_DFF data_in_frame_0__i124 (.Q(\data_in_frame[15] [3]), .C(clk32MHz), 
           .D(n23815));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_31425 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[14] [3]), .I2(\data_out_frame[15] [3]), 
            .I3(byte_transmit_counter[1]), .O(n46949));
    defparam byte_transmit_counter_0__bdd_4_lut_31425.LUT_INIT = 16'he4aa;
    SB_DFF data_in_frame_0__i125 (.Q(\data_in_frame[15] [4]), .C(clk32MHz), 
           .D(n23814));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 n46949_bdd_4_lut (.I0(n46949), .I1(\data_out_frame[13] [3]), 
            .I2(\data_out_frame[12] [3]), .I3(byte_transmit_counter[1]), 
            .O(n46952));
    defparam n46949_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF data_in_frame_0__i126 (.Q(\data_in_frame[15] [5]), .C(clk32MHz), 
           .D(n23813));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i1_2_lut_adj_884 (.I0(n40567), .I1(\data_in_frame[20] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n4_adj_3146));
    defparam i1_2_lut_adj_884.LUT_INIT = 16'h6666;
    SB_DFF data_in_frame_0__i127 (.Q(\data_in_frame[15] [6]), .C(clk32MHz), 
           .D(n23812));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_31420 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[18] [2]), .I2(\data_out_frame[19] [2]), 
            .I3(byte_transmit_counter[1]), .O(n46943));
    defparam byte_transmit_counter_0__bdd_4_lut_31420.LUT_INIT = 16'he4aa;
    SB_DFF data_in_frame_0__i128 (.Q(\data_in_frame[15] [7]), .C(clk32MHz), 
           .D(n23811));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 n46943_bdd_4_lut (.I0(n46943), .I1(\data_out_frame[17] [2]), 
            .I2(\data_out_frame[16] [2]), .I3(byte_transmit_counter[1]), 
            .O(n46946));
    defparam n46943_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF data_in_frame_0__i129 (.Q(\data_in_frame[16] [0]), .C(clk32MHz), 
           .D(n23810));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i4_4_lut_adj_885 (.I0(\data_in_frame[20] [2]), .I1(n37241), 
            .I2(n22997), .I3(n47038), .O(n10_adj_3147));
    defparam i4_4_lut_adj_885.LUT_INIT = 16'h9669;
    SB_DFF data_in_frame_0__i130 (.Q(\data_in_frame[16] [1]), .C(clk32MHz), 
           .D(n23809));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_31415 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[18] [1]), .I2(\data_out_frame[19] [1]), 
            .I3(byte_transmit_counter[1]), .O(n46937));
    defparam byte_transmit_counter_0__bdd_4_lut_31415.LUT_INIT = 16'he4aa;
    SB_DFF data_in_frame_0__i131 (.Q(\data_in_frame[16] [2]), .C(clk32MHz), 
           .D(n23808));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 n46937_bdd_4_lut (.I0(n46937), .I1(\data_out_frame[17] [1]), 
            .I2(\data_out_frame[16] [1]), .I3(byte_transmit_counter[1]), 
            .O(n46940));
    defparam n46937_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF data_in_frame_0__i132 (.Q(\data_in_frame[16] [3]), .C(clk32MHz), 
           .D(n23807));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i3_4_lut_adj_886 (.I0(\data_in_frame[17] [7]), .I1(n40362), 
            .I2(n37310), .I3(\data_in_frame[20] [1]), .O(n41687));
    defparam i3_4_lut_adj_886.LUT_INIT = 16'h9669;
    SB_DFF data_in_frame_0__i133 (.Q(\data_in_frame[16] [4]), .C(clk32MHz), 
           .D(n23806));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 add_44_13_lut (.I0(n1498), .I1(\FRAME_MATCHER.i [11]), .I2(GND_net), 
            .I3(n34034), .O(n2_adj_3148)) /* synthesis syn_instantiated=1 */ ;
    defparam add_44_13_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_547_6 (.CI(n34058), .I0(byte_transmit_counter_c[4]), .I1(GND_net), 
            .CO(n34059));
    SB_DFF data_in_frame_0__i134 (.Q(\data_in_frame[16] [5]), .C(clk32MHz), 
           .D(n23805));   // verilog/coms.v(126[12] 289[6])
    SB_CARRY add_44_13 (.CI(n34034), .I0(\FRAME_MATCHER.i [11]), .I1(GND_net), 
            .CO(n34035));
    SB_LUT4 add_44_5_lut (.I0(n1498), .I1(\FRAME_MATCHER.i [3]), .I2(GND_net), 
            .I3(n34026), .O(n2_adj_3149)) /* synthesis syn_instantiated=1 */ ;
    defparam add_44_5_lut.LUT_INIT = 16'h8228;
    SB_LUT4 add_547_5_lut (.I0(GND_net), .I1(byte_transmit_counter_c[3]), 
            .I2(GND_net), .I3(n34057), .O(n2236[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_547_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_44_5 (.CI(n34026), .I0(\FRAME_MATCHER.i [3]), .I1(GND_net), 
            .CO(n34027));
    SB_LUT4 add_44_12_lut (.I0(n1498), .I1(\FRAME_MATCHER.i [10]), .I2(GND_net), 
            .I3(n34033), .O(n2_adj_3150)) /* synthesis syn_instantiated=1 */ ;
    defparam add_44_12_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_547_5 (.CI(n34057), .I0(byte_transmit_counter_c[3]), .I1(GND_net), 
            .CO(n34058));
    SB_LUT4 add_547_4_lut (.I0(GND_net), .I1(byte_transmit_counter_c[2]), 
            .I2(GND_net), .I3(n34056), .O(n2236[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_547_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_44_4_lut (.I0(n1498), .I1(\FRAME_MATCHER.i [2]), .I2(GND_net), 
            .I3(n34025), .O(n2_adj_3151)) /* synthesis syn_instantiated=1 */ ;
    defparam add_44_4_lut.LUT_INIT = 16'h8228;
    SB_DFF data_in_frame_0__i135 (.Q(\data_in_frame[16] [6]), .C(clk32MHz), 
           .D(n23804));   // verilog/coms.v(126[12] 289[6])
    SB_CARRY add_44_4 (.CI(n34025), .I0(\FRAME_MATCHER.i [2]), .I1(GND_net), 
            .CO(n34026));
    SB_DFF data_in_frame_0__i136 (.Q(\data_in_frame[16] [7]), .C(clk32MHz), 
           .D(n23803));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i137 (.Q(\data_in_frame[17] [0]), .C(clk32MHz), 
           .D(n23802));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_31410 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[18] [0]), .I2(\data_out_frame[19] [0]), 
            .I3(byte_transmit_counter[1]), .O(n46931));
    defparam byte_transmit_counter_0__bdd_4_lut_31410.LUT_INIT = 16'he4aa;
    SB_DFF data_in_0___i17 (.Q(\data_in[2] [0]), .C(clk32MHz), .D(n24084));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.state_i31  (.Q(\FRAME_MATCHER.state [31]), .C(clk32MHz), 
            .D(n39646), .S(n39508));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 add_44_3_lut (.I0(n1498), .I1(\FRAME_MATCHER.i [1]), .I2(GND_net), 
            .I3(n34024), .O(n2_adj_3152)) /* synthesis syn_instantiated=1 */ ;
    defparam add_44_3_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_44_12 (.CI(n34033), .I0(\FRAME_MATCHER.i [10]), .I1(GND_net), 
            .CO(n34034));
    SB_CARRY add_547_4 (.CI(n34056), .I0(byte_transmit_counter_c[2]), .I1(GND_net), 
            .CO(n34057));
    SB_LUT4 add_547_3_lut (.I0(GND_net), .I1(byte_transmit_counter[1]), 
            .I2(GND_net), .I3(n34055), .O(n2236[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_547_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_547_3 (.CI(n34055), .I0(byte_transmit_counter[1]), .I1(GND_net), 
            .CO(n34056));
    SB_DFFSS \FRAME_MATCHER.state_i30  (.Q(\FRAME_MATCHER.state [30]), .C(clk32MHz), 
            .D(n39642), .S(n39518));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.state_i29  (.Q(\FRAME_MATCHER.state [29]), .C(clk32MHz), 
            .D(n39640), .S(n39510));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.state_i28  (.Q(\FRAME_MATCHER.state [28]), .C(clk32MHz), 
            .D(n27682), .S(n39514));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.state_i27  (.Q(\FRAME_MATCHER.state [27]), .C(clk32MHz), 
            .D(n39638), .S(n39550));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 add_44_11_lut (.I0(n1498), .I1(\FRAME_MATCHER.i [9]), .I2(GND_net), 
            .I3(n34032), .O(n2_adj_3153)) /* synthesis syn_instantiated=1 */ ;
    defparam add_44_11_lut.LUT_INIT = 16'h8228;
    SB_DFFSS \FRAME_MATCHER.state_i26  (.Q(\FRAME_MATCHER.state [26]), .C(clk32MHz), 
            .D(n39636), .S(n39516));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 add_547_2_lut (.I0(GND_net), .I1(byte_transmit_counter[0]), 
            .I2(tx_transmit_N_2648), .I3(GND_net), .O(n2236[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_547_2_lut.LUT_INIT = 16'hC33C;
    SB_DFFSS \FRAME_MATCHER.state_i25  (.Q(\FRAME_MATCHER.state [25]), .C(clk32MHz), 
            .D(n39634), .S(n39496));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.state_i24  (.Q(\FRAME_MATCHER.state [24]), .C(clk32MHz), 
            .D(n39632), .S(n39492));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.state_i23  (.Q(\FRAME_MATCHER.state [23]), .C(clk32MHz), 
            .D(n39744), .S(n39494));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.state_i22  (.Q(\FRAME_MATCHER.state [22]), .C(clk32MHz), 
            .D(n39686), .S(n39552));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.state_i21  (.Q(\FRAME_MATCHER.state [21]), .C(clk32MHz), 
            .D(n39684), .S(n39554));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.state_i20  (.Q(\FRAME_MATCHER.state [20]), .C(clk32MHz), 
            .D(n39676), .S(n35999));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.state_i19  (.Q(\FRAME_MATCHER.state [19]), .C(clk32MHz), 
            .D(n39674), .S(n39556));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.state_i18  (.Q(\FRAME_MATCHER.state [18]), .C(clk32MHz), 
            .D(n39672), .S(n39512));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.state_i17  (.Q(\FRAME_MATCHER.state [17]), .C(clk32MHz), 
            .D(n39670), .S(n39522));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.state_i16  (.Q(\FRAME_MATCHER.state [16]), .C(clk32MHz), 
            .D(n39668), .S(n39436));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.state_i15  (.Q(\FRAME_MATCHER.state [15]), .C(clk32MHz), 
            .D(n39666), .S(n39558));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.state_i14  (.Q(\FRAME_MATCHER.state [14]), .C(clk32MHz), 
            .D(n39664), .S(n39560));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.state_i13  (.Q(\FRAME_MATCHER.state [13]), .C(clk32MHz), 
            .D(n39662), .S(n39562));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.state_i12  (.Q(\FRAME_MATCHER.state [12]), .C(clk32MHz), 
            .D(n39660), .S(n39564));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.state_i11  (.Q(\FRAME_MATCHER.state [11]), .C(clk32MHz), 
            .D(n39658), .S(n39566));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.state_i10  (.Q(\FRAME_MATCHER.state [10]), .C(clk32MHz), 
            .D(n39656), .S(n39568));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.state_i9  (.Q(\FRAME_MATCHER.state [9]), .C(clk32MHz), 
            .D(n39654), .S(n39570));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.state_i8  (.Q(\FRAME_MATCHER.state [8]), .C(clk32MHz), 
            .D(n39652), .S(n39402));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.state_i7  (.Q(\FRAME_MATCHER.state [7]), .C(clk32MHz), 
            .D(n39650), .S(n39572));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.state_i6  (.Q(\FRAME_MATCHER.state [6]), .C(clk32MHz), 
            .D(n39584), .S(n28159));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.state_i5  (.Q(\FRAME_MATCHER.state [5]), .C(clk32MHz), 
            .D(n27700), .S(n28157));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.state_i4  (.Q(\FRAME_MATCHER.state [4]), .C(clk32MHz), 
            .D(n39648), .S(n39406));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.state_i3  (.Q(\FRAME_MATCHER.state [3]), .C(clk32MHz), 
            .D(n39506), .S(n39742));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.state_i1  (.Q(\FRAME_MATCHER.state [1]), .C(clk32MHz), 
            .D(n39504), .S(n47026));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i138 (.Q(\data_in_frame[17] [1]), .C(clk32MHz), 
           .D(n23801));   // verilog/coms.v(126[12] 289[6])
    SB_CARRY add_44_3 (.CI(n34024), .I0(\FRAME_MATCHER.i [1]), .I1(GND_net), 
            .CO(n34025));
    SB_CARRY add_44_11 (.CI(n34032), .I0(\FRAME_MATCHER.i [9]), .I1(GND_net), 
            .CO(n34033));
    SB_CARRY add_547_2 (.CI(GND_net), .I0(byte_transmit_counter[0]), .I1(tx_transmit_N_2648), 
            .CO(n34055));
    SB_LUT4 add_44_33_lut (.I0(n1498), .I1(\FRAME_MATCHER.i [31]), .I2(GND_net), 
            .I3(n34054), .O(n2_adj_3154)) /* synthesis syn_instantiated=1 */ ;
    defparam add_44_33_lut.LUT_INIT = 16'h8228;
    SB_DFF data_in_frame_0__i139 (.Q(\data_in_frame[17] [2]), .C(clk32MHz), 
           .D(n23800));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i140 (.Q(\data_in_frame[17] [3]), .C(clk32MHz), 
           .D(n23799));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i141 (.Q(\data_in_frame[17] [4]), .C(clk32MHz), 
           .D(n23798));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i142 (.Q(\data_in_frame[17] [5]), .C(clk32MHz), 
           .D(n23797));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i143 (.Q(\data_in_frame[17] [6]), .C(clk32MHz), 
           .D(n23796));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i144 (.Q(\data_in_frame[17] [7]), .C(clk32MHz), 
           .D(n23795));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i145 (.Q(\data_in_frame[18] [0]), .C(clk32MHz), 
           .D(n23794));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i146 (.Q(\data_in_frame[18] [1]), .C(clk32MHz), 
           .D(n23793));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i147 (.Q(\data_in_frame[18] [2]), .C(clk32MHz), 
           .D(n23792));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i148 (.Q(\data_in_frame[18] [3]), .C(clk32MHz), 
           .D(n23791));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i149 (.Q(\data_in_frame[18] [4]), .C(clk32MHz), 
           .D(n23790));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i150 (.Q(\data_in_frame[18] [5]), .C(clk32MHz), 
           .D(n23789));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i151 (.Q(\data_in_frame[18] [6]), .C(clk32MHz), 
           .D(n23788));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i152 (.Q(\data_in_frame[18] [7]), .C(clk32MHz), 
           .D(n23787));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i153 (.Q(\data_in_frame[19] [0]), .C(clk32MHz), 
           .D(n23786));   // verilog/coms.v(126[12] 289[6])
    SB_DFFE data_out_frame_0___i184 (.Q(\data_out_frame[22][7] ), .C(clk32MHz), 
            .E(n23452), .D(n41574));   // verilog/coms.v(126[12] 289[6])
    SB_DFFE data_out_frame_0___i183 (.Q(\data_out_frame[22] [6]), .C(clk32MHz), 
            .E(n23452), .D(n41743));   // verilog/coms.v(126[12] 289[6])
    SB_DFFE data_out_frame_0___i182 (.Q(\data_out_frame[22] [5]), .C(clk32MHz), 
            .E(n23452), .D(n40703));   // verilog/coms.v(126[12] 289[6])
    SB_DFFE data_out_frame_0___i181 (.Q(\data_out_frame[22] [4]), .C(clk32MHz), 
            .E(n23452), .D(n40448));   // verilog/coms.v(126[12] 289[6])
    SB_DFFE data_out_frame_0___i180 (.Q(\data_out_frame[22] [3]), .C(clk32MHz), 
            .E(n23452), .D(n40449));   // verilog/coms.v(126[12] 289[6])
    SB_DFFE data_out_frame_0___i179 (.Q(\data_out_frame[22] [2]), .C(clk32MHz), 
            .E(n23452), .D(n40375));   // verilog/coms.v(126[12] 289[6])
    SB_DFFE data_out_frame_0___i178 (.Q(\data_out_frame[22] [1]), .C(clk32MHz), 
            .E(n23452), .D(n40513));   // verilog/coms.v(126[12] 289[6])
    SB_DFFE data_out_frame_0___i177 (.Q(\data_out_frame[22] [0]), .C(clk32MHz), 
            .E(n23452), .D(n40514));   // verilog/coms.v(126[12] 289[6])
    SB_DFFE data_out_frame_0___i176 (.Q(\data_out_frame[21][7] ), .C(clk32MHz), 
            .E(n23452), .D(n41732));   // verilog/coms.v(126[12] 289[6])
    SB_DFFE data_out_frame_0___i175 (.Q(\data_out_frame[21] [6]), .C(clk32MHz), 
            .E(n23452), .D(n41124));   // verilog/coms.v(126[12] 289[6])
    SB_DFFE data_out_frame_0___i174 (.Q(\data_out_frame[21] [5]), .C(clk32MHz), 
            .E(n23452), .D(n41129));   // verilog/coms.v(126[12] 289[6])
    SB_DFFE data_out_frame_0___i173 (.Q(\data_out_frame[21] [4]), .C(clk32MHz), 
            .E(n23452), .D(n41339));   // verilog/coms.v(126[12] 289[6])
    SB_DFFE data_out_frame_0___i172 (.Q(\data_out_frame[21] [3]), .C(clk32MHz), 
            .E(n23452), .D(n41672));   // verilog/coms.v(126[12] 289[6])
    SB_DFFE data_out_frame_0___i171 (.Q(\data_out_frame[21] [2]), .C(clk32MHz), 
            .E(n23452), .D(n41758));   // verilog/coms.v(126[12] 289[6])
    SB_DFFE data_out_frame_0___i170 (.Q(\data_out_frame[21] [1]), .C(clk32MHz), 
            .E(n23452), .D(n41498));   // verilog/coms.v(126[12] 289[6])
    SB_DFFE data_out_frame_0___i169 (.Q(\data_out_frame[21] [0]), .C(clk32MHz), 
            .E(n23452), .D(n41847));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i154 (.Q(\data_in_frame[19] [1]), .C(clk32MHz), 
           .D(n23785));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.i_i31  (.Q(\FRAME_MATCHER.i [31]), .C(clk32MHz), 
            .D(n2_adj_3154), .S(n3));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 add_44_32_lut (.I0(n1498), .I1(\FRAME_MATCHER.i [30]), .I2(GND_net), 
            .I3(n34053), .O(n2_adj_3155)) /* synthesis syn_instantiated=1 */ ;
    defparam add_44_32_lut.LUT_INIT = 16'h8228;
    SB_LUT4 n46931_bdd_4_lut (.I0(n46931), .I1(\data_out_frame[17] [0]), 
            .I2(\data_out_frame[16] [0]), .I3(byte_transmit_counter[1]), 
            .O(n46934));
    defparam n46931_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFFSS \FRAME_MATCHER.i_i30  (.Q(\FRAME_MATCHER.i [30]), .C(clk32MHz), 
            .D(n2_adj_3155), .S(n3_adj_3156));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.i_i29  (.Q(\FRAME_MATCHER.i [29]), .C(clk32MHz), 
            .D(n2_adj_3157), .S(n3_adj_3158));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.i_i28  (.Q(\FRAME_MATCHER.i [28]), .C(clk32MHz), 
            .D(n2_adj_3159), .S(n3_adj_3160));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.i_i27  (.Q(\FRAME_MATCHER.i [27]), .C(clk32MHz), 
            .D(n2_adj_3161), .S(n3_adj_3162));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.i_i26  (.Q(\FRAME_MATCHER.i [26]), .C(clk32MHz), 
            .D(n2_adj_3163), .S(n3_adj_3164));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.i_i25  (.Q(\FRAME_MATCHER.i [25]), .C(clk32MHz), 
            .D(n2_adj_3165), .S(n3_adj_3166));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.i_i24  (.Q(\FRAME_MATCHER.i [24]), .C(clk32MHz), 
            .D(n2_adj_3167), .S(n3_adj_3168));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.i_i23  (.Q(\FRAME_MATCHER.i [23]), .C(clk32MHz), 
            .D(n2_adj_3169), .S(n3_adj_3170));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.i_i22  (.Q(\FRAME_MATCHER.i [22]), .C(clk32MHz), 
            .D(n2_adj_3171), .S(n3_adj_3172));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.i_i21  (.Q(\FRAME_MATCHER.i [21]), .C(clk32MHz), 
            .D(n2_adj_3173), .S(n3_adj_3174));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.i_i20  (.Q(\FRAME_MATCHER.i [20]), .C(clk32MHz), 
            .D(n2_adj_3175), .S(n3_adj_3176));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.i_i19  (.Q(\FRAME_MATCHER.i [19]), .C(clk32MHz), 
            .D(n2_adj_3177), .S(n3_adj_3178));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.i_i18  (.Q(\FRAME_MATCHER.i [18]), .C(clk32MHz), 
            .D(n2_adj_3179), .S(n3_adj_3180));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.i_i17  (.Q(\FRAME_MATCHER.i [17]), .C(clk32MHz), 
            .D(n2), .S(n3_adj_3181));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.i_i16  (.Q(\FRAME_MATCHER.i [16]), .C(clk32MHz), 
            .D(n2_adj_3119), .S(n3_adj_3182));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.i_i15  (.Q(\FRAME_MATCHER.i [15]), .C(clk32MHz), 
            .D(n2_adj_3121), .S(n3_adj_3183));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.i_i14  (.Q(\FRAME_MATCHER.i [14]), .C(clk32MHz), 
            .D(n2_adj_3125), .S(n3_adj_3184));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.i_i13  (.Q(\FRAME_MATCHER.i [13]), .C(clk32MHz), 
            .D(n2_adj_3127), .S(n3_adj_3185));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.i_i12  (.Q(\FRAME_MATCHER.i [12]), .C(clk32MHz), 
            .D(n2_adj_3136), .S(n3_adj_3186));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.i_i11  (.Q(\FRAME_MATCHER.i [11]), .C(clk32MHz), 
            .D(n2_adj_3148), .S(n3_adj_3187));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.i_i10  (.Q(\FRAME_MATCHER.i [10]), .C(clk32MHz), 
            .D(n2_adj_3150), .S(n3_adj_3188));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.i_i9  (.Q(\FRAME_MATCHER.i [9]), .C(clk32MHz), 
            .D(n2_adj_3153), .S(n3_adj_3189));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.i_i8  (.Q(\FRAME_MATCHER.i [8]), .C(clk32MHz), 
            .D(n2_adj_3190), .S(n3_adj_3191));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.i_i7  (.Q(\FRAME_MATCHER.i [7]), .C(clk32MHz), 
            .D(n2_adj_3192), .S(n3_adj_3193));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.i_i6  (.Q(\FRAME_MATCHER.i [6]), .C(clk32MHz), 
            .D(n2_adj_3194), .S(n3_adj_3195));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.i_i5  (.Q(\FRAME_MATCHER.i [5]), .C(clk32MHz), 
            .D(n2_adj_3120), .S(n3_adj_3196));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.i_i4  (.Q(\FRAME_MATCHER.i [4]), .C(clk32MHz), 
            .D(n2_adj_3126), .S(n3_adj_3197));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.i_i3  (.Q(\FRAME_MATCHER.i [3]), .C(clk32MHz), 
            .D(n2_adj_3149), .S(n3_adj_3198));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.i_i2  (.Q(\FRAME_MATCHER.i [2]), .C(clk32MHz), 
            .D(n2_adj_3151), .S(n3_adj_3199));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.i_i1  (.Q(\FRAME_MATCHER.i [1]), .C(clk32MHz), 
            .D(n2_adj_3152), .S(n3_adj_3200));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i155 (.Q(\data_in_frame[19] [2]), .C(clk32MHz), 
           .D(n23784));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i156 (.Q(\data_in_frame[19] [3]), .C(clk32MHz), 
           .D(n23783));   // verilog/coms.v(126[12] 289[6])
    SB_DFF Ki_i2 (.Q(\Ki[2] ), .C(clk32MHz), .D(n24135));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i157 (.Q(\data_in_frame[19] [4]), .C(clk32MHz), 
           .D(n23782));   // verilog/coms.v(126[12] 289[6])
    SB_DFF Ki_i3 (.Q(\Ki[3] ), .C(clk32MHz), .D(n24134));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i158 (.Q(\data_in_frame[19] [5]), .C(clk32MHz), 
           .D(n23781));   // verilog/coms.v(126[12] 289[6])
    SB_DFF Ki_i4 (.Q(\Ki[4] ), .C(clk32MHz), .D(n24133));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i159 (.Q(\data_in_frame[19] [6]), .C(clk32MHz), 
           .D(n23780));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i160 (.Q(\data_in_frame[19] [7]), .C(clk32MHz), 
           .D(n23779));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i161 (.Q(\data_in_frame[20] [0]), .C(clk32MHz), 
           .D(n23778));   // verilog/coms.v(126[12] 289[6])
    SB_CARRY add_44_32 (.CI(n34053), .I0(\FRAME_MATCHER.i [30]), .I1(GND_net), 
            .CO(n34054));
    SB_LUT4 add_44_31_lut (.I0(n1498), .I1(\FRAME_MATCHER.i [29]), .I2(GND_net), 
            .I3(n34052), .O(n2_adj_3157)) /* synthesis syn_instantiated=1 */ ;
    defparam add_44_31_lut.LUT_INIT = 16'h8228;
    SB_DFF data_in_frame_0__i162 (.Q(\data_in_frame[20] [1]), .C(clk32MHz), 
           .D(n23777));   // verilog/coms.v(126[12] 289[6])
    SB_CARRY add_44_31 (.CI(n34052), .I0(\FRAME_MATCHER.i [29]), .I1(GND_net), 
            .CO(n34053));
    SB_DFF data_in_frame_0__i163 (.Q(\data_in_frame[20] [2]), .C(clk32MHz), 
           .D(n23776));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i164 (.Q(\data_in_frame[20] [3]), .C(clk32MHz), 
           .D(n23775));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i165 (.Q(\data_in_frame[20] [4]), .C(clk32MHz), 
           .D(n23774));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i166 (.Q(\data_in_frame[20] [5]), .C(clk32MHz), 
           .D(n23773));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i167 (.Q(\data_in_frame[20] [6]), .C(clk32MHz), 
           .D(n23772));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i168 (.Q(\data_in_frame[20] [7]), .C(clk32MHz), 
           .D(n23771));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i169 (.Q(\data_in_frame[21] [0]), .C(clk32MHz), 
           .D(n23770));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i170 (.Q(\data_in_frame[21] [1]), .C(clk32MHz), 
           .D(n23769));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i171 (.Q(\data_in_frame[21] [2]), .C(clk32MHz), 
           .D(n23768));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i172 (.Q(\data_in_frame[21] [3]), .C(clk32MHz), 
           .D(n23767));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i173 (.Q(\data_in_frame[21] [4]), .C(clk32MHz), 
           .D(n23766));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i174 (.Q(\data_in_frame[21] [5]), .C(clk32MHz), 
           .D(n23765));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i175 (.Q(\data_in_frame[21] [6]), .C(clk32MHz), 
           .D(n23764));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i176 (.Q(\data_in_frame[21] [7]), .C(clk32MHz), 
           .D(n23763));   // verilog/coms.v(126[12] 289[6])
    SB_DFF control_mode_i0_i1 (.Q(control_mode[1]), .C(clk32MHz), .D(n23762));   // verilog/coms.v(126[12] 289[6])
    SB_DFF control_mode_i0_i2 (.Q(control_mode[2]), .C(clk32MHz), .D(n23761));   // verilog/coms.v(126[12] 289[6])
    SB_DFF control_mode_i0_i3 (.Q(control_mode[3]), .C(clk32MHz), .D(n23760));   // verilog/coms.v(126[12] 289[6])
    SB_DFF control_mode_i0_i4 (.Q(control_mode[4]), .C(clk32MHz), .D(n23759));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i2_4_lut_adj_887 (.I0(n41687), .I1(n40352), .I2(n40564), .I3(\data_in_frame[21] [2]), 
            .O(n10_adj_3201));
    defparam i2_4_lut_adj_887.LUT_INIT = 16'h8228;
    SB_LUT4 add_44_30_lut (.I0(n1498), .I1(\FRAME_MATCHER.i [28]), .I2(GND_net), 
            .I3(n34051), .O(n2_adj_3159)) /* synthesis syn_instantiated=1 */ ;
    defparam add_44_30_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_44_30 (.CI(n34051), .I0(\FRAME_MATCHER.i [28]), .I1(GND_net), 
            .CO(n34052));
    SB_DFF control_mode_i0_i5 (.Q(control_mode[5]), .C(clk32MHz), .D(n23758));   // verilog/coms.v(126[12] 289[6])
    SB_DFF control_mode_i0_i6 (.Q(control_mode[6]), .C(clk32MHz), .D(n23757));   // verilog/coms.v(126[12] 289[6])
    SB_DFF control_mode_i0_i7 (.Q(control_mode[7]), .C(clk32MHz), .D(n23756));   // verilog/coms.v(126[12] 289[6])
    SB_DFF PWMLimit_i0_i1 (.Q(\PWMLimit[1] ), .C(clk32MHz), .D(n23755));   // verilog/coms.v(126[12] 289[6])
    SB_DFF PWMLimit_i0_i2 (.Q(\PWMLimit[2] ), .C(clk32MHz), .D(n23754));   // verilog/coms.v(126[12] 289[6])
    SB_DFF PWMLimit_i0_i3 (.Q(\PWMLimit[3] ), .C(clk32MHz), .D(n23753));   // verilog/coms.v(126[12] 289[6])
    SB_DFF PWMLimit_i0_i4 (.Q(\PWMLimit[4] ), .C(clk32MHz), .D(n23752));   // verilog/coms.v(126[12] 289[6])
    SB_DFF PWMLimit_i0_i5 (.Q(\PWMLimit[5] ), .C(clk32MHz), .D(n23751));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 add_44_29_lut (.I0(n1498), .I1(\FRAME_MATCHER.i [27]), .I2(GND_net), 
            .I3(n34050), .O(n2_adj_3161)) /* synthesis syn_instantiated=1 */ ;
    defparam add_44_29_lut.LUT_INIT = 16'h8228;
    SB_DFF PWMLimit_i0_i6 (.Q(\PWMLimit[6] ), .C(clk32MHz), .D(n27220));   // verilog/coms.v(126[12] 289[6])
    SB_DFF PWMLimit_i0_i7 (.Q(\PWMLimit[7] ), .C(clk32MHz), .D(n23749));   // verilog/coms.v(126[12] 289[6])
    SB_DFF PWMLimit_i0_i8 (.Q(\PWMLimit[8] ), .C(clk32MHz), .D(n23748));   // verilog/coms.v(126[12] 289[6])
    SB_DFF PWMLimit_i0_i9 (.Q(\PWMLimit[9] ), .C(clk32MHz), .D(n23747));   // verilog/coms.v(126[12] 289[6])
    SB_CARRY add_44_29 (.CI(n34050), .I0(\FRAME_MATCHER.i [27]), .I1(GND_net), 
            .CO(n34051));
    SB_DFF \FRAME_MATCHER.state_i2  (.Q(\FRAME_MATCHER.state [2]), .C(clk32MHz), 
           .D(n47027));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 add_44_28_lut (.I0(n1498), .I1(\FRAME_MATCHER.i [26]), .I2(GND_net), 
            .I3(n34049), .O(n2_adj_3163)) /* synthesis syn_instantiated=1 */ ;
    defparam add_44_28_lut.LUT_INIT = 16'h8228;
    SB_LUT4 add_44_10_lut (.I0(n1498), .I1(\FRAME_MATCHER.i [8]), .I2(GND_net), 
            .I3(n34031), .O(n2_adj_3190)) /* synthesis syn_instantiated=1 */ ;
    defparam add_44_10_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i6_4_lut_adj_888 (.I0(n41583), .I1(n41776), .I2(n41390), .I3(n41720), 
            .O(n14_adj_3202));
    defparam i6_4_lut_adj_888.LUT_INIT = 16'h0080;
    SB_DFF data_in_0___i18 (.Q(\data_in[2] [1]), .C(clk32MHz), .D(n24083));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_31455 (.I0(byte_transmit_counter[1]), 
            .I1(n11), .I2(n12_adj_3203), .I3(byte_transmit_counter_c[2]), 
            .O(n46919));
    defparam byte_transmit_counter_1__bdd_4_lut_31455.LUT_INIT = 16'he4aa;
    SB_LUT4 n46919_bdd_4_lut (.I0(n46919), .I1(n9_adj_3204), .I2(n8_adj_3205), 
            .I3(byte_transmit_counter_c[2]), .O(n46922));
    defparam n46919_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF data_in_0___i19 (.Q(\data_in[2] [2]), .C(clk32MHz), .D(n24082));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSR tx_transmit_3227 (.Q(r_SM_Main_2__N_2756[0]), .C(clk32MHz), 
            .D(n39256), .R(n28289));   // verilog/coms.v(126[12] 289[6])
    SB_DFF Kd_i7 (.Q(\Kd[7] ), .C(clk32MHz), .D(n24123));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_0___i20 (.Q(\data_in[2] [3]), .C(clk32MHz), .D(n24081));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i10401_3_lut_4_lut (.I0(n8_adj_3122), .I1(n40221), .I2(rx_data[7]), 
            .I3(\data_in_frame[14] [7]), .O(n23819));
    defparam i10401_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF data_in_0___i21 (.Q(\data_in[2] [4]), .C(clk32MHz), .D(n24080));   // verilog/coms.v(126[12] 289[6])
    SB_DFF gearBoxRatio_i0_i1 (.Q(gearBoxRatio[1]), .C(clk32MHz), .D(n24122));   // verilog/coms.v(126[12] 289[6])
    SB_CARRY add_44_28 (.CI(n34049), .I0(\FRAME_MATCHER.i [26]), .I1(GND_net), 
            .CO(n34050));
    SB_DFF IntegralLimit_i0_i21 (.Q(IntegralLimit[21]), .C(clk32MHz), .D(n24146));   // verilog/coms.v(126[12] 289[6])
    SB_CARRY add_44_10 (.CI(n34031), .I0(\FRAME_MATCHER.i [8]), .I1(GND_net), 
            .CO(n34032));
    SB_LUT4 add_44_9_lut (.I0(n1498), .I1(\FRAME_MATCHER.i [7]), .I2(GND_net), 
            .I3(n34030), .O(n2_adj_3192)) /* synthesis syn_instantiated=1 */ ;
    defparam add_44_9_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i26636_4_lut (.I0(n41389), .I1(n10_adj_3147), .I2(\data_in_frame[18] [1]), 
            .I3(n4_adj_3146), .O(n42155));
    defparam i26636_4_lut.LUT_INIT = 16'heb7d;
    SB_LUT4 add_44_27_lut (.I0(n1498), .I1(\FRAME_MATCHER.i [25]), .I2(GND_net), 
            .I3(n34048), .O(n2_adj_3165)) /* synthesis syn_instantiated=1 */ ;
    defparam add_44_27_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i10402_3_lut_4_lut (.I0(n8_adj_3122), .I1(n40221), .I2(rx_data[6]), 
            .I3(\data_in_frame[14] [6]), .O(n23820));
    defparam i10402_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF IntegralLimit_i0_i22 (.Q(IntegralLimit[22]), .C(clk32MHz), .D(n24145));   // verilog/coms.v(126[12] 289[6])
    SB_DFF IntegralLimit_i0_i23 (.Q(IntegralLimit[23]), .C(clk32MHz), .D(n24144));   // verilog/coms.v(126[12] 289[6])
    SB_DFF Kp_i1 (.Q(\Kp[1] ), .C(clk32MHz), .D(n24143));   // verilog/coms.v(126[12] 289[6])
    SB_DFF Kp_i2 (.Q(\Kp[2] ), .C(clk32MHz), .D(n24142));   // verilog/coms.v(126[12] 289[6])
    SB_DFF Kp_i3 (.Q(\Kp[3] ), .C(clk32MHz), .D(n24141));   // verilog/coms.v(126[12] 289[6])
    SB_DFF Kp_i4 (.Q(\Kp[4] ), .C(clk32MHz), .D(n24140));   // verilog/coms.v(126[12] 289[6])
    SB_DFF Kp_i5 (.Q(\Kp[5] ), .C(clk32MHz), .D(n24139));   // verilog/coms.v(126[12] 289[6])
    SB_DFF Kp_i6 (.Q(\Kp[6] ), .C(clk32MHz), .D(n24138));   // verilog/coms.v(126[12] 289[6])
    SB_DFFE LED_3230 (.Q(LED_c), .C(clk32MHz), .E(n40886), .D(n19_adj_3206));   // verilog/coms.v(126[12] 289[6])
    SB_CARRY add_44_27 (.CI(n34048), .I0(\FRAME_MATCHER.i [25]), .I1(GND_net), 
            .CO(n34049));
    SB_LUT4 i10403_3_lut_4_lut (.I0(n8_adj_3122), .I1(n40221), .I2(rx_data[5]), 
            .I3(\data_in_frame[14] [5]), .O(n23821));
    defparam i10403_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_31405 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[10] [5]), .I2(\data_out_frame[11] [5]), 
            .I3(byte_transmit_counter[1]), .O(n46913));
    defparam byte_transmit_counter_0__bdd_4_lut_31405.LUT_INIT = 16'he4aa;
    SB_LUT4 add_44_2_lut (.I0(n1498), .I1(\FRAME_MATCHER.i [0]), .I2(n164), 
            .I3(GND_net), .O(n2_adj_3207)) /* synthesis syn_instantiated=1 */ ;
    defparam add_44_2_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i3_4_lut_adj_889 (.I0(\FRAME_MATCHER.state [18]), .I1(\FRAME_MATCHER.state [16]), 
            .I2(\FRAME_MATCHER.state [20]), .I3(\FRAME_MATCHER.state [24]), 
            .O(n31577));   // verilog/coms.v(126[12] 289[6])
    defparam i3_4_lut_adj_889.LUT_INIT = 16'hfffe;
    SB_LUT4 i3_4_lut_adj_890 (.I0(\FRAME_MATCHER.state [4]), .I1(\FRAME_MATCHER.state [7]), 
            .I2(\FRAME_MATCHER.state [5]), .I3(\FRAME_MATCHER.state [6]), 
            .O(n40110));
    defparam i3_4_lut_adj_890.LUT_INIT = 16'hfffe;
    SB_LUT4 i8_4_lut_adj_891 (.I0(\FRAME_MATCHER.state [19]), .I1(\FRAME_MATCHER.state [29]), 
            .I2(\FRAME_MATCHER.state [26]), .I3(\FRAME_MATCHER.state [30]), 
            .O(n20_adj_3208));
    defparam i8_4_lut_adj_891.LUT_INIT = 16'hfffe;
    SB_LUT4 i7_4_lut_adj_892 (.I0(\FRAME_MATCHER.state [17]), .I1(\FRAME_MATCHER.state [21]), 
            .I2(\FRAME_MATCHER.state [31]), .I3(\FRAME_MATCHER.state [28]), 
            .O(n19_adj_3209));
    defparam i7_4_lut_adj_892.LUT_INIT = 16'hfffe;
    SB_LUT4 add_44_26_lut (.I0(n1498), .I1(\FRAME_MATCHER.i [24]), .I2(GND_net), 
            .I3(n34047), .O(n2_adj_3167)) /* synthesis syn_instantiated=1 */ ;
    defparam add_44_26_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i10404_3_lut_4_lut (.I0(n8_adj_3122), .I1(n40221), .I2(rx_data[4]), 
            .I3(\data_in_frame[14] [4]), .O(n23822));
    defparam i10404_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10405_3_lut_4_lut (.I0(n8_adj_3122), .I1(n40221), .I2(rx_data[3]), 
            .I3(\data_in_frame[14] [3]), .O(n23823));
    defparam i10405_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i9_4_lut_adj_893 (.I0(\FRAME_MATCHER.state [22]), .I1(\FRAME_MATCHER.state [23]), 
            .I2(\FRAME_MATCHER.state [25]), .I3(\FRAME_MATCHER.state [27]), 
            .O(n21_c));
    defparam i9_4_lut_adj_893.LUT_INIT = 16'hfffe;
    SB_LUT4 i11_3_lut (.I0(n21_c), .I1(n19_adj_3209), .I2(n20_adj_3208), 
            .I3(GND_net), .O(n40247));
    defparam i11_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i2_2_lut_adj_894 (.I0(\FRAME_MATCHER.state [13]), .I1(\FRAME_MATCHER.state [8]), 
            .I2(GND_net), .I3(GND_net), .O(n10_adj_3210));
    defparam i2_2_lut_adj_894.LUT_INIT = 16'heeee;
    SB_LUT4 i6_4_lut_adj_895 (.I0(\FRAME_MATCHER.state [10]), .I1(\FRAME_MATCHER.state [11]), 
            .I2(\FRAME_MATCHER.state [12]), .I3(\FRAME_MATCHER.state [9]), 
            .O(n14_adj_3211));
    defparam i6_4_lut_adj_895.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_rep_6_2_lut (.I0(n40573), .I1(n40746), .I2(GND_net), .I3(GND_net), 
            .O(n47033));
    defparam i1_rep_6_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i7_4_lut_adj_896 (.I0(\FRAME_MATCHER.state [15]), .I1(n14_adj_3211), 
            .I2(n10_adj_3210), .I3(\FRAME_MATCHER.state [14]), .O(n40106));
    defparam i7_4_lut_adj_896.LUT_INIT = 16'hfffe;
    SB_LUT4 i3_4_lut_adj_897 (.I0(n40106), .I1(n40247), .I2(n40110), .I3(n31577), 
            .O(n28279));
    defparam i3_4_lut_adj_897.LUT_INIT = 16'hfffe;
    SB_LUT4 i25487_2_lut (.I0(n28279), .I1(\FRAME_MATCHER.state [0]), .I2(GND_net), 
            .I3(GND_net), .O(n41005));
    defparam i25487_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i1_2_lut_adj_898 (.I0(\data_in_frame[0] [5]), .I1(\data_in_frame[0] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n9_adj_3212));
    defparam i1_2_lut_adj_898.LUT_INIT = 16'heeee;
    SB_LUT4 i1_2_lut_adj_899 (.I0(\data_in_frame[1] [6]), .I1(\data_in_frame[1] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n18_adj_3213));
    defparam i1_2_lut_adj_899.LUT_INIT = 16'h8888;
    SB_LUT4 i4_4_lut_adj_900 (.I0(n40362), .I1(n37241), .I2(n37310), .I3(n40554), 
            .O(n10_adj_3214));
    defparam i4_4_lut_adj_900.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_901 (.I0(\data_in_frame[0] [2]), .I1(\data_in_frame[1] [1]), 
            .I2(\data_in_frame[2] [0]), .I3(\data_in_frame[2] [5]), .O(n14_adj_3215));
    defparam i6_4_lut_adj_901.LUT_INIT = 16'hfffe;
    SB_CARRY add_44_26 (.CI(n34047), .I0(\FRAME_MATCHER.i [24]), .I1(GND_net), 
            .CO(n34048));
    SB_LUT4 n46913_bdd_4_lut (.I0(n46913), .I1(\data_out_frame[9] [5]), 
            .I2(\data_out_frame[8] [5]), .I3(byte_transmit_counter[1]), 
            .O(n46916));
    defparam n46913_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 add_44_25_lut (.I0(n1498), .I1(\FRAME_MATCHER.i [23]), .I2(GND_net), 
            .I3(n34046), .O(n2_adj_3169)) /* synthesis syn_instantiated=1 */ ;
    defparam add_44_25_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_44_9 (.CI(n34030), .I0(\FRAME_MATCHER.i [7]), .I1(GND_net), 
            .CO(n34031));
    SB_CARRY add_44_25 (.CI(n34046), .I0(\FRAME_MATCHER.i [23]), .I1(GND_net), 
            .CO(n34047));
    SB_LUT4 i10406_3_lut_4_lut (.I0(n8_adj_3122), .I1(n40221), .I2(rx_data[2]), 
            .I3(\data_in_frame[14] [2]), .O(n23824));
    defparam i10406_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i7_4_lut_adj_902 (.I0(n9_adj_3212), .I1(n14_adj_3215), .I2(\data_in_frame[2] [4]), 
            .I3(\data_in_frame[2] [3]), .O(n41262));
    defparam i7_4_lut_adj_902.LUT_INIT = 16'hfffe;
    SB_LUT4 i13_4_lut (.I0(\data_in_frame[0] [3]), .I1(\data_in_frame[0] [1]), 
            .I2(\data_in_frame[0] [4]), .I3(n18_adj_3213), .O(n30));
    defparam i13_4_lut.LUT_INIT = 16'h0100;
    SB_LUT4 i2_3_lut_adj_903 (.I0(n40352), .I1(n40668), .I2(\data_in_frame[21] [3]), 
            .I3(GND_net), .O(n41134));
    defparam i2_3_lut_adj_903.LUT_INIT = 16'h9696;
    SB_LUT4 i11_4_lut (.I0(\data_in_frame[2] [1]), .I1(\data_in_frame[1] [5]), 
            .I2(\data_in_frame[1] [4]), .I3(\data_in_frame[2] [7]), .O(n28));
    defparam i11_4_lut.LUT_INIT = 16'h0080;
    SB_LUT4 add_44_24_lut (.I0(n1498), .I1(\FRAME_MATCHER.i [22]), .I2(GND_net), 
            .I3(n34045), .O(n2_adj_3171)) /* synthesis syn_instantiated=1 */ ;
    defparam add_44_24_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i26668_4_lut (.I0(\data_in_frame[2] [6]), .I1(\data_in_frame[2] [2]), 
            .I2(\data_in_frame[0] [0]), .I3(\data_in_frame[0] [6]), .O(n42187));
    defparam i26668_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i3_4_lut_adj_904 (.I0(\data_in_frame[19] [3]), .I1(n40573), 
            .I2(n37295), .I3(\data_in_frame[21] [5]), .O(n41676));
    defparam i3_4_lut_adj_904.LUT_INIT = 16'h6996;
    SB_LUT4 i10_4_lut (.I0(n41262), .I1(\data_in_frame[1] [2]), .I2(\data_in_frame[1] [3]), 
            .I3(\data_in_frame[1] [0]), .O(n27));
    defparam i10_4_lut.LUT_INIT = 16'h4000;
    SB_LUT4 i2_4_lut_adj_905 (.I0(\data_in_frame[17] [6]), .I1(n41134), 
            .I2(n10_adj_3214), .I3(\data_in_frame[20] [0]), .O(n11_adj_3216));
    defparam i2_4_lut_adj_905.LUT_INIT = 16'h4884;
    SB_LUT4 i10407_3_lut_4_lut (.I0(n8_adj_3122), .I1(n40221), .I2(rx_data[1]), 
            .I3(\data_in_frame[14] [1]), .O(n23825));
    defparam i10407_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_CARRY add_44_24 (.CI(n34045), .I0(\FRAME_MATCHER.i [22]), .I1(GND_net), 
            .CO(n34046));
    SB_LUT4 add_44_8_lut (.I0(n1498), .I1(\FRAME_MATCHER.i [6]), .I2(GND_net), 
            .I3(n34029), .O(n2_adj_3194)) /* synthesis syn_instantiated=1 */ ;
    defparam add_44_8_lut.LUT_INIT = 16'h8228;
    SB_DFF gearBoxRatio_i0_i2 (.Q(gearBoxRatio[2]), .C(clk32MHz), .D(n24121));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i10408_3_lut_4_lut (.I0(n8_adj_3122), .I1(n40221), .I2(rx_data[0]), 
            .I3(\data_in_frame[14] [0]), .O(n23826));
    defparam i10408_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10393_3_lut_4_lut (.I0(n27747), .I1(n40221), .I2(rx_data[7]), 
            .I3(\data_in_frame[15] [7]), .O(n23811));
    defparam i10393_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 add_44_23_lut (.I0(n1498), .I1(\FRAME_MATCHER.i [21]), .I2(GND_net), 
            .I3(n34044), .O(n2_adj_3173)) /* synthesis syn_instantiated=1 */ ;
    defparam add_44_23_lut.LUT_INIT = 16'h8228;
    SB_DFF gearBoxRatio_i0_i3 (.Q(gearBoxRatio[3]), .C(clk32MHz), .D(n24120));   // verilog/coms.v(126[12] 289[6])
    SB_DFF gearBoxRatio_i0_i4 (.Q(gearBoxRatio[4]), .C(clk32MHz), .D(n24119));   // verilog/coms.v(126[12] 289[6])
    SB_DFF gearBoxRatio_i0_i5 (.Q(gearBoxRatio[5]), .C(clk32MHz), .D(n24118));   // verilog/coms.v(126[12] 289[6])
    SB_DFF deadband_i0_i0 (.Q(\deadband[0] ), .C(clk32MHz), .D(n23600));   // verilog/coms.v(126[12] 289[6])
    SB_CARRY add_44_23 (.CI(n34044), .I0(\FRAME_MATCHER.i [21]), .I1(GND_net), 
            .CO(n34045));
    SB_DFFSS \FRAME_MATCHER.i_i0  (.Q(\FRAME_MATCHER.i [0]), .C(clk32MHz), 
            .D(n2_adj_3207), .S(n3_adj_3217));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 add_44_22_lut (.I0(n1498), .I1(\FRAME_MATCHER.i [20]), .I2(GND_net), 
            .I3(n34043), .O(n2_adj_3175)) /* synthesis syn_instantiated=1 */ ;
    defparam add_44_22_lut.LUT_INIT = 16'h8228;
    SB_DFF setpoint__i0 (.Q(setpoint[0]), .C(clk32MHz), .D(n23599));   // verilog/coms.v(126[12] 289[6])
    SB_CARRY add_44_22 (.CI(n34043), .I0(\FRAME_MATCHER.i [20]), .I1(GND_net), 
            .CO(n34044));
    SB_LUT4 add_44_21_lut (.I0(n1498), .I1(\FRAME_MATCHER.i [19]), .I2(GND_net), 
            .I3(n34042), .O(n2_adj_3177)) /* synthesis syn_instantiated=1 */ ;
    defparam add_44_21_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_44_21 (.CI(n34042), .I0(\FRAME_MATCHER.i [19]), .I1(GND_net), 
            .CO(n34043));
    SB_DFF \FRAME_MATCHER.state_i0  (.Q(\FRAME_MATCHER.state [0]), .C(clk32MHz), 
           .D(n39520));   // verilog/coms.v(126[12] 289[6])
    SB_DFF PWMLimit_i0_i0 (.Q(\PWMLimit[0] ), .C(clk32MHz), .D(n23588));   // verilog/coms.v(126[12] 289[6])
    SB_DFF control_mode_i0_i0 (.Q(control_mode[0]), .C(clk32MHz), .D(n23587));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i1 (.Q(\data_in_frame[0] [0]), .C(clk32MHz), 
           .D(n23586));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_0___i1 (.Q(\data_in[0] [0]), .C(clk32MHz), .D(n23585));   // verilog/coms.v(126[12] 289[6])
    SB_DFF gearBoxRatio_i0_i0 (.Q(gearBoxRatio[0]), .C(clk32MHz), .D(n23584));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i62 (.Q(\data_out_frame[7] [5]), .C(clk32MHz), 
           .D(n24044));   // verilog/coms.v(126[12] 289[6])
    SB_DFF Kd_i0 (.Q(\Kd[0] ), .C(clk32MHz), .D(n23583));   // verilog/coms.v(126[12] 289[6])
    SB_CARRY add_44_2 (.CI(GND_net), .I0(\FRAME_MATCHER.i [0]), .I1(n164), 
            .CO(n34024));
    SB_DFF Ki_i0 (.Q(\Ki[0] ), .C(clk32MHz), .D(n23582));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 add_44_20_lut (.I0(n1498), .I1(\FRAME_MATCHER.i [18]), .I2(GND_net), 
            .I3(n34041), .O(n2_adj_3179)) /* synthesis syn_instantiated=1 */ ;
    defparam add_44_20_lut.LUT_INIT = 16'h8228;
    SB_DFF Kp_i0 (.Q(\Kp[0] ), .C(clk32MHz), .D(n23581));   // verilog/coms.v(126[12] 289[6])
    SB_DFF IntegralLimit_i0_i0 (.Q(IntegralLimit[0]), .C(clk32MHz), .D(n23580));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i10394_3_lut_4_lut (.I0(n27747), .I1(n40221), .I2(rx_data[6]), 
            .I3(\data_in_frame[15] [6]), .O(n23812));
    defparam i10394_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1_2_lut_3_lut_adj_906 (.I0(\data_in_frame[7] [4]), .I1(\data_in_frame[10] [0]), 
            .I2(\data_in_frame[7] [5]), .I3(GND_net), .O(n23045));
    defparam i1_2_lut_3_lut_adj_906.LUT_INIT = 16'h9696;
    SB_LUT4 i10395_3_lut_4_lut (.I0(n27747), .I1(n40221), .I2(rx_data[5]), 
            .I3(\data_in_frame[15] [5]), .O(n23813));
    defparam i10395_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i10396_3_lut_4_lut (.I0(n27747), .I1(n40221), .I2(rx_data[4]), 
            .I3(\data_in_frame[15] [4]), .O(n23814));
    defparam i10396_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1_4_lut_adj_907 (.I0(n5021), .I1(n28145), .I2(\FRAME_MATCHER.state_31__N_1925 [3]), 
            .I3(n5019), .O(n23458));
    defparam i1_4_lut_adj_907.LUT_INIT = 16'ha022;
    SB_LUT4 i10397_3_lut_4_lut (.I0(n27747), .I1(n40221), .I2(rx_data[3]), 
            .I3(\data_in_frame[15] [3]), .O(n23815));
    defparam i10397_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i2_4_lut_adj_908 (.I0(\FRAME_MATCHER.state [3]), .I1(n41005), 
            .I2(\FRAME_MATCHER.state [1]), .I3(\FRAME_MATCHER.state [2]), 
            .O(n5019));
    defparam i2_4_lut_adj_908.LUT_INIT = 16'h0012;
    SB_LUT4 i1_4_lut_adj_909 (.I0(n41462), .I1(n42155), .I2(n14_adj_3202), 
            .I3(n10_adj_3201), .O(n10_adj_3218));
    defparam i1_4_lut_adj_909.LUT_INIT = 16'h1000;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_910 (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(n40212), .I3(\FRAME_MATCHER.i [0]), .O(n40218));   // verilog/coms.v(154[7:23])
    defparam i1_2_lut_3_lut_4_lut_adj_910.LUT_INIT = 16'hfbff;
    SB_LUT4 i2_3_lut_4_lut_adj_911 (.I0(\data_in_frame[7] [4]), .I1(\data_in_frame[10] [0]), 
            .I2(\data_in_frame[11] [7]), .I3(\data_in_frame[14] [3]), .O(n40840));
    defparam i2_3_lut_4_lut_adj_911.LUT_INIT = 16'h6996;
    SB_LUT4 i10398_3_lut_4_lut (.I0(n27747), .I1(n40221), .I2(rx_data[2]), 
            .I3(\data_in_frame[15] [2]), .O(n23816));
    defparam i10398_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i10399_3_lut_4_lut (.I0(n27747), .I1(n40221), .I2(rx_data[1]), 
            .I3(\data_in_frame[15] [1]), .O(n23817));
    defparam i10399_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_31392 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[18] [6]), .I2(\data_out_frame[19] [6]), 
            .I3(byte_transmit_counter[1]), .O(n46907));
    defparam byte_transmit_counter_0__bdd_4_lut_31392.LUT_INIT = 16'he4aa;
    SB_LUT4 i10400_3_lut_4_lut (.I0(n27747), .I1(n40221), .I2(rx_data[0]), 
            .I3(\data_in_frame[15] [0]), .O(n23818));
    defparam i10400_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i10385_3_lut_4_lut (.I0(n8_adj_3123), .I1(n40205), .I2(rx_data[7]), 
            .I3(\data_in_frame[16] [7]), .O(n23803));
    defparam i10385_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10386_3_lut_4_lut (.I0(n8_adj_3123), .I1(n40205), .I2(rx_data[6]), 
            .I3(\data_in_frame[16] [6]), .O(n23804));
    defparam i10386_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_4_lut_adj_912 (.I0(\data_in_frame[0] [4]), .I1(\data_in_frame[2] [5]), 
            .I2(\data_in_frame[0] [3]), .I3(n40437), .O(Kp_23__N_329));   // verilog/coms.v(74[16:43])
    defparam i1_2_lut_4_lut_adj_912.LUT_INIT = 16'h6996;
    SB_LUT4 i10387_3_lut_4_lut (.I0(n8_adj_3123), .I1(n40205), .I2(rx_data[5]), 
            .I3(\data_in_frame[16] [5]), .O(n23805));
    defparam i10387_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i3_4_lut_adj_913 (.I0(n5_adj_3219), .I1(\FRAME_MATCHER.i_31__N_1825 ), 
            .I2(n40163), .I3(n2857), .O(n41799));
    defparam i3_4_lut_adj_913.LUT_INIT = 16'hfafe;
    SB_LUT4 i1_2_lut_4_lut_adj_914 (.I0(\data_in_frame[0] [4]), .I1(\data_in_frame[2] [5]), 
            .I2(\data_in_frame[0] [3]), .I3(n5_adj_3135), .O(Kp_23__N_326));   // verilog/coms.v(74[16:43])
    defparam i1_2_lut_4_lut_adj_914.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_915 (.I0(\FRAME_MATCHER.i_31__N_1823 ), .I1(n20075), 
            .I2(n41799), .I3(\FRAME_MATCHER.state [0]), .O(n39520));
    defparam i1_4_lut_adj_915.LUT_INIT = 16'hfaba;
    SB_LUT4 n46907_bdd_4_lut (.I0(n46907), .I1(\data_out_frame[17] [6]), 
            .I2(\data_out_frame[16] [6]), .I3(byte_transmit_counter[1]), 
            .O(n46910));
    defparam n46907_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i2_3_lut_4_lut_adj_916 (.I0(\data_in_frame[3] [0]), .I1(\data_in_frame[0] [7]), 
            .I2(\data_in_frame[1] [1]), .I3(n40674), .O(n40437));   // verilog/coms.v(69[16:69])
    defparam i2_3_lut_4_lut_adj_916.LUT_INIT = 16'h6996;
    SB_LUT4 i10388_3_lut_4_lut (.I0(n8_adj_3123), .I1(n40205), .I2(rx_data[4]), 
            .I3(\data_in_frame[16] [4]), .O(n23806));
    defparam i10388_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10389_3_lut_4_lut (.I0(n8_adj_3123), .I1(n40205), .I2(rx_data[3]), 
            .I3(\data_in_frame[16] [3]), .O(n23807));
    defparam i10389_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10390_3_lut_4_lut (.I0(n8_adj_3123), .I1(n40205), .I2(rx_data[2]), 
            .I3(\data_in_frame[16] [2]), .O(n23808));
    defparam i10390_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10391_3_lut_4_lut (.I0(n8_adj_3123), .I1(n40205), .I2(rx_data[1]), 
            .I3(\data_in_frame[16] [1]), .O(n23809));
    defparam i10391_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10392_3_lut_4_lut (.I0(n8_adj_3123), .I1(n40205), .I2(rx_data[0]), 
            .I3(\data_in_frame[16] [0]), .O(n23810));
    defparam i10392_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_4_lut_adj_917 (.I0(n47), .I1(n2_adj_3220), .I2(n6_adj_3221), 
            .I3(\FRAME_MATCHER.state [7]), .O(n39572));
    defparam i1_2_lut_4_lut_adj_917.LUT_INIT = 16'hfe00;
    SB_LUT4 i1_2_lut_4_lut_adj_918 (.I0(n47), .I1(n2_adj_3220), .I2(n6_adj_3221), 
            .I3(\FRAME_MATCHER.state [9]), .O(n39570));
    defparam i1_2_lut_4_lut_adj_918.LUT_INIT = 16'hfe00;
    SB_LUT4 i29066_2_lut (.I0(byte_transmit_counter_c[2]), .I1(\data_out_frame[5] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n44587));   // verilog/coms.v(104[34:55])
    defparam i29066_2_lut.LUT_INIT = 16'hdddd;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_7_i5_3_lut (.I0(\data_out_frame[6] [7]), 
            .I1(\data_out_frame[7] [7]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n5_adj_3222));   // verilog/coms.v(104[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_7_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_7_i22_3_lut (.I0(n47012), .I1(n21), 
            .I2(byte_transmit_counter_c[2]), .I3(GND_net), .O(n22_c));   // verilog/coms.v(104[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_7_i22_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i26711_4_lut (.I0(n5_adj_3222), .I1(n44587), .I2(n43966), 
            .I3(byte_transmit_counter[0]), .O(n42230));
    defparam i26711_4_lut.LUT_INIT = 16'haca0;
    SB_LUT4 i26713_4_lut (.I0(n42230), .I1(n22_c), .I2(byte_transmit_counter_c[4]), 
            .I3(byte_transmit_counter_c[3]), .O(n42232));
    defparam i26713_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_6_i19_3_lut (.I0(\data_out_frame[20] [6]), 
            .I1(\data_out_frame[21] [6]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n19_adj_3224));   // verilog/coms.v(104[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_6_i19_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i26682_4_lut (.I0(n19_adj_3224), .I1(\data_out_frame[22] [6]), 
            .I2(byte_transmit_counter[1]), .I3(byte_transmit_counter[0]), 
            .O(n42201));
    defparam i26682_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i29060_2_lut (.I0(byte_transmit_counter_c[2]), .I1(\data_out_frame[5] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n44581));   // verilog/coms.v(104[34:55])
    defparam i29060_2_lut.LUT_INIT = 16'hdddd;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_6_i5_3_lut (.I0(\data_out_frame[6] [6]), 
            .I1(\data_out_frame[7] [6]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n5_adj_3225));   // verilog/coms.v(104[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_6_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i26683_3_lut (.I0(n46910), .I1(n42201), .I2(byte_transmit_counter_c[2]), 
            .I3(GND_net), .O(n42202));
    defparam i26683_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i26708_4_lut (.I0(n5_adj_3225), .I1(n44581), .I2(n43966), 
            .I3(byte_transmit_counter[0]), .O(n42227));
    defparam i26708_4_lut.LUT_INIT = 16'haca0;
    SB_LUT4 i26710_4_lut (.I0(n42227), .I1(n42202), .I2(byte_transmit_counter_c[4]), 
            .I3(byte_transmit_counter_c[3]), .O(n42229));
    defparam i26710_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i1_2_lut_4_lut_adj_919 (.I0(n47), .I1(n2_adj_3220), .I2(n6_adj_3221), 
            .I3(\FRAME_MATCHER.state [10]), .O(n39568));
    defparam i1_2_lut_4_lut_adj_919.LUT_INIT = 16'hfe00;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_5_i19_3_lut (.I0(\data_out_frame[20] [5]), 
            .I1(\data_out_frame[21] [5]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n19_adj_3226));   // verilog/coms.v(104[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_5_i19_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_5_i6_3_lut (.I0(\data_out_frame[5] [5]), 
            .I1(byte_transmit_counter[1]), .I2(byte_transmit_counter_c[2]), 
            .I3(GND_net), .O(n44575));   // verilog/coms.v(104[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_5_i6_3_lut.LUT_INIT = 16'ha3a3;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_5_i5_3_lut (.I0(\data_out_frame[6] [5]), 
            .I1(\data_out_frame[7] [5]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n5_adj_3227));   // verilog/coms.v(104[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_5_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i26679_4_lut (.I0(n19_adj_3226), .I1(\data_out_frame[22] [5]), 
            .I2(byte_transmit_counter[1]), .I3(byte_transmit_counter[0]), 
            .O(n42198));
    defparam i26679_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i26680_3_lut (.I0(n46904), .I1(n42198), .I2(byte_transmit_counter_c[2]), 
            .I3(GND_net), .O(n42199));
    defparam i26680_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i26705_4_lut (.I0(n5_adj_3227), .I1(byte_transmit_counter[0]), 
            .I2(n43966), .I3(n44575), .O(n42224));
    defparam i26705_4_lut.LUT_INIT = 16'haca0;
    SB_LUT4 i26707_4_lut (.I0(n42224), .I1(n42199), .I2(byte_transmit_counter_c[4]), 
            .I3(byte_transmit_counter_c[3]), .O(n42226));
    defparam i26707_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i26706_3_lut (.I0(n46916), .I1(n46892), .I2(byte_transmit_counter_c[2]), 
            .I3(GND_net), .O(n42225));
    defparam i26706_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_4_lut_adj_920 (.I0(n47), .I1(n2_adj_3220), .I2(n6_adj_3221), 
            .I3(\FRAME_MATCHER.state [11]), .O(n39566));
    defparam i1_2_lut_4_lut_adj_920.LUT_INIT = 16'hfe00;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_7_i31_3_lut_4_lut (.I0(byte_transmit_counter_c[4]), 
            .I1(byte_transmit_counter_c[3]), .I2(n42232), .I3(n46994), 
            .O(tx_data[7]));   // verilog/coms.v(104[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_7_i31_3_lut_4_lut.LUT_INIT = 16'hf4b0;
    SB_LUT4 i1_2_lut_4_lut_adj_921 (.I0(n47), .I1(n2_adj_3220), .I2(n6_adj_3221), 
            .I3(\FRAME_MATCHER.state [12]), .O(n39564));
    defparam i1_2_lut_4_lut_adj_921.LUT_INIT = 16'hfe00;
    SB_LUT4 i1_2_lut_4_lut_adj_922 (.I0(n47), .I1(n2_adj_3220), .I2(n6_adj_3221), 
            .I3(\FRAME_MATCHER.state [13]), .O(n39562));
    defparam i1_2_lut_4_lut_adj_922.LUT_INIT = 16'hfe00;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_4_i19_3_lut (.I0(\data_out_frame[20] [4]), 
            .I1(\data_out_frame[21] [4]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n19_adj_3228));   // verilog/coms.v(104[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_4_i19_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_6_i31_3_lut_4_lut (.I0(byte_transmit_counter_c[4]), 
            .I1(byte_transmit_counter_c[3]), .I2(n42229), .I3(n47000), 
            .O(tx_data[6]));   // verilog/coms.v(104[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_6_i31_3_lut_4_lut.LUT_INIT = 16'hf4b0;
    SB_LUT4 i26676_4_lut (.I0(n19_adj_3228), .I1(\data_out_frame[22] [4]), 
            .I2(byte_transmit_counter[1]), .I3(byte_transmit_counter[0]), 
            .O(n42195));
    defparam i26676_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i26677_3_lut (.I0(n46898), .I1(n42195), .I2(byte_transmit_counter_c[2]), 
            .I3(GND_net), .O(n42196));
    defparam i26677_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i30283_3_lut (.I0(n47006), .I1(n46922), .I2(byte_transmit_counter_c[3]), 
            .I3(GND_net), .O(n45804));   // verilog/coms.v(104[34:55])
    defparam i30283_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i30284_4_lut (.I0(n45804), .I1(n42196), .I2(byte_transmit_counter_c[4]), 
            .I3(byte_transmit_counter_c[3]), .O(tx_data[4]));   // verilog/coms.v(104[34:55])
    defparam i30284_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i1_2_lut_4_lut_adj_923 (.I0(n47), .I1(n2_adj_3220), .I2(n6_adj_3221), 
            .I3(\FRAME_MATCHER.state [14]), .O(n39560));
    defparam i1_2_lut_4_lut_adj_923.LUT_INIT = 16'hfe00;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_5_i31_3_lut_4_lut (.I0(byte_transmit_counter_c[4]), 
            .I1(byte_transmit_counter_c[3]), .I2(n42226), .I3(n42225), 
            .O(tx_data[5]));   // verilog/coms.v(104[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_5_i31_3_lut_4_lut.LUT_INIT = 16'hf4b0;
    SB_LUT4 i1_2_lut_4_lut_adj_924 (.I0(n47), .I1(n2_adj_3220), .I2(n6_adj_3221), 
            .I3(\FRAME_MATCHER.state [15]), .O(n39558));
    defparam i1_2_lut_4_lut_adj_924.LUT_INIT = 16'hfe00;
    SB_LUT4 i29041_2_lut (.I0(\data_out_frame[0][3] ), .I1(byte_transmit_counter[1]), 
            .I2(GND_net), .I3(GND_net), .O(n44129));   // verilog/coms.v(104[34:55])
    defparam i29041_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i1_2_lut_4_lut_adj_925 (.I0(n47), .I1(n2_adj_3220), .I2(n6_adj_3221), 
            .I3(\FRAME_MATCHER.state [16]), .O(n39436));
    defparam i1_2_lut_4_lut_adj_925.LUT_INIT = 16'hfe00;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_3_i6_4_lut (.I0(\data_out_frame[5] [3]), 
            .I1(n44129), .I2(byte_transmit_counter_c[2]), .I3(byte_transmit_counter[0]), 
            .O(n6_adj_3229));   // verilog/coms.v(104[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_3_i6_4_lut.LUT_INIT = 16'haf0c;
    SB_LUT4 i1_2_lut_4_lut_adj_926 (.I0(n47), .I1(n2_adj_3220), .I2(n6_adj_3221), 
            .I3(\FRAME_MATCHER.state [17]), .O(n39522));
    defparam i1_2_lut_4_lut_adj_926.LUT_INIT = 16'hfe00;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_3_i5_3_lut (.I0(\data_out_frame[6] [3]), 
            .I1(\data_out_frame[7] [3]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n5_adj_3230));   // verilog/coms.v(104[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_3_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i26696_3_lut (.I0(n5_adj_3230), .I1(n6_adj_3229), .I2(n43966), 
            .I3(GND_net), .O(n42215));
    defparam i26696_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i26698_4_lut (.I0(n42215), .I1(n47024), .I2(byte_transmit_counter_c[4]), 
            .I3(byte_transmit_counter_c[3]), .O(n42217));
    defparam i26698_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i26697_3_lut (.I0(n46958), .I1(n46952), .I2(byte_transmit_counter_c[2]), 
            .I3(GND_net), .O(n42216));
    defparam i26697_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_4_lut_adj_927 (.I0(n47), .I1(n2_adj_3220), .I2(n6_adj_3221), 
            .I3(\FRAME_MATCHER.state [18]), .O(n39512));
    defparam i1_2_lut_4_lut_adj_927.LUT_INIT = 16'hfe00;
    SB_LUT4 i1_2_lut_4_lut_adj_928 (.I0(n47), .I1(n2_adj_3220), .I2(n6_adj_3221), 
            .I3(\FRAME_MATCHER.state [19]), .O(n39556));
    defparam i1_2_lut_4_lut_adj_928.LUT_INIT = 16'hfe00;
    SB_LUT4 i1_2_lut_4_lut_adj_929 (.I0(n47), .I1(n2_adj_3220), .I2(n6_adj_3221), 
            .I3(\FRAME_MATCHER.state [21]), .O(n39554));
    defparam i1_2_lut_4_lut_adj_929.LUT_INIT = 16'hfe00;
    SB_LUT4 i1_2_lut_4_lut_adj_930 (.I0(n47), .I1(n2_adj_3220), .I2(n6_adj_3221), 
            .I3(\FRAME_MATCHER.state [22]), .O(n39552));
    defparam i1_2_lut_4_lut_adj_930.LUT_INIT = 16'hfe00;
    SB_LUT4 i29309_2_lut (.I0(\data_out_frame[0][2] ), .I1(byte_transmit_counter[1]), 
            .I2(GND_net), .I3(GND_net), .O(n44126));   // verilog/coms.v(104[34:55])
    defparam i29309_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_2_i19_3_lut (.I0(\data_out_frame[20] [2]), 
            .I1(\data_out_frame[21] [2]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n19_adj_3231));   // verilog/coms.v(104[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_2_i19_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_2_i6_4_lut (.I0(\data_out_frame[5][2] ), 
            .I1(n44126), .I2(byte_transmit_counter_c[2]), .I3(byte_transmit_counter[0]), 
            .O(n6_adj_3232));   // verilog/coms.v(104[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_2_i6_4_lut.LUT_INIT = 16'ha00c;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_2_i5_3_lut (.I0(\data_out_frame[6] [2]), 
            .I1(\data_out_frame[7] [2]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n5_adj_3233));   // verilog/coms.v(104[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_2_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_4_lut_adj_931 (.I0(n47), .I1(n2_adj_3220), .I2(n6_adj_3221), 
            .I3(\FRAME_MATCHER.state [23]), .O(n39494));
    defparam i1_2_lut_4_lut_adj_931.LUT_INIT = 16'hfe00;
    SB_LUT4 i26721_4_lut (.I0(n19_adj_3231), .I1(\data_out_frame[22] [2]), 
            .I2(byte_transmit_counter[1]), .I3(byte_transmit_counter[0]), 
            .O(n42240));
    defparam i26721_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i26722_3_lut (.I0(n46946), .I1(n42240), .I2(byte_transmit_counter_c[2]), 
            .I3(GND_net), .O(n42241));
    defparam i26722_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i26693_3_lut (.I0(n5_adj_3233), .I1(n6_adj_3232), .I2(n43966), 
            .I3(GND_net), .O(n42212));
    defparam i26693_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i26695_4_lut (.I0(n42212), .I1(n42241), .I2(byte_transmit_counter_c[4]), 
            .I3(byte_transmit_counter_c[3]), .O(n42214));
    defparam i26695_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i26694_3_lut (.I0(n46970), .I1(n46964), .I2(byte_transmit_counter_c[2]), 
            .I3(GND_net), .O(n42213));
    defparam i26694_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_4_lut_adj_932 (.I0(n47), .I1(n2_adj_3220), .I2(n6_adj_3221), 
            .I3(\FRAME_MATCHER.state [24]), .O(n39492));
    defparam i1_2_lut_4_lut_adj_932.LUT_INIT = 16'hfe00;
    SB_LUT4 i1_2_lut_4_lut_adj_933 (.I0(n47), .I1(n2_adj_3220), .I2(n6_adj_3221), 
            .I3(\FRAME_MATCHER.state [25]), .O(n39496));
    defparam i1_2_lut_4_lut_adj_933.LUT_INIT = 16'hfe00;
    SB_LUT4 i1_2_lut_4_lut_adj_934 (.I0(n47), .I1(n2_adj_3220), .I2(n6_adj_3221), 
            .I3(\FRAME_MATCHER.state [26]), .O(n39516));
    defparam i1_2_lut_4_lut_adj_934.LUT_INIT = 16'hfe00;
    SB_LUT4 i1_2_lut_4_lut_adj_935 (.I0(n47), .I1(n2_adj_3220), .I2(n6_adj_3221), 
            .I3(\FRAME_MATCHER.state [27]), .O(n39550));
    defparam i1_2_lut_4_lut_adj_935.LUT_INIT = 16'hfe00;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_1_i19_3_lut (.I0(\data_out_frame[20] [1]), 
            .I1(\data_out_frame[21] [1]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n19_adj_3234));   // verilog/coms.v(104[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_1_i19_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_4_lut_adj_936 (.I0(n47), .I1(n2_adj_3220), .I2(n6_adj_3221), 
            .I3(\FRAME_MATCHER.state [28]), .O(n39514));
    defparam i1_2_lut_4_lut_adj_936.LUT_INIT = 16'hfe00;
    SB_LUT4 i29036_2_lut (.I0(byte_transmit_counter_c[2]), .I1(\data_out_frame[5] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n44556));   // verilog/coms.v(104[34:55])
    defparam i29036_2_lut.LUT_INIT = 16'hdddd;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_1_i5_3_lut (.I0(\data_out_frame[6] [1]), 
            .I1(\data_out_frame[7] [1]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n5_adj_3235));   // verilog/coms.v(104[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_1_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i26718_4_lut (.I0(n19_adj_3234), .I1(\data_out_frame[22] [1]), 
            .I2(byte_transmit_counter[1]), .I3(byte_transmit_counter[0]), 
            .O(n42237));
    defparam i26718_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i26719_3_lut (.I0(n46940), .I1(n42237), .I2(byte_transmit_counter_c[2]), 
            .I3(GND_net), .O(n42238));
    defparam i26719_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i26690_4_lut (.I0(n5_adj_3235), .I1(n44556), .I2(n43966), 
            .I3(byte_transmit_counter[0]), .O(n42209));
    defparam i26690_4_lut.LUT_INIT = 16'haca0;
    SB_LUT4 i26692_4_lut (.I0(n42209), .I1(n42238), .I2(byte_transmit_counter_c[4]), 
            .I3(byte_transmit_counter_c[3]), .O(n42211));
    defparam i26692_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i1_2_lut_adj_937 (.I0(\FRAME_MATCHER.state [2]), .I1(\FRAME_MATCHER.state [0]), 
            .I2(GND_net), .I3(GND_net), .O(n4_adj_3236));
    defparam i1_2_lut_adj_937.LUT_INIT = 16'h2222;
    SB_LUT4 i1_2_lut_4_lut_adj_938 (.I0(n47), .I1(n2_adj_3220), .I2(n6_adj_3221), 
            .I3(\FRAME_MATCHER.state [29]), .O(n39510));
    defparam i1_2_lut_4_lut_adj_938.LUT_INIT = 16'hfe00;
    SB_LUT4 i1_2_lut_adj_939 (.I0(n36853), .I1(n40828), .I2(GND_net), 
            .I3(GND_net), .O(n40362));
    defparam i1_2_lut_adj_939.LUT_INIT = 16'h6666;
    SB_LUT4 i26691_3_lut (.I0(n46982), .I1(n46976), .I2(byte_transmit_counter_c[2]), 
            .I3(GND_net), .O(n42210));
    defparam i26691_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_4_lut_adj_940 (.I0(n47), .I1(n2_adj_3220), .I2(n6_adj_3221), 
            .I3(\FRAME_MATCHER.state [30]), .O(n39518));
    defparam i1_2_lut_4_lut_adj_940.LUT_INIT = 16'hfe00;
    SB_LUT4 i1_2_lut_4_lut_adj_941 (.I0(n47), .I1(n2_adj_3220), .I2(n6_adj_3221), 
            .I3(\FRAME_MATCHER.state [31]), .O(n39508));
    defparam i1_2_lut_4_lut_adj_941.LUT_INIT = 16'hfe00;
    SB_LUT4 i5_4_lut_adj_942 (.I0(n37239), .I1(n40420), .I2(n37336), .I3(n37237), 
            .O(n12_adj_3237));
    defparam i5_4_lut_adj_942.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_3_lut_adj_943 (.I0(n5_adj_3238), .I1(n43), .I2(\FRAME_MATCHER.state [4]), 
            .I3(GND_net), .O(n39648));
    defparam i1_2_lut_3_lut_adj_943.LUT_INIT = 16'he0e0;
    SB_LUT4 i6_4_lut_adj_944 (.I0(\data_in_frame[17] [7]), .I1(n12_adj_3237), 
            .I2(n40515), .I3(n37248), .O(n41389));
    defparam i6_4_lut_adj_944.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_945 (.I0(\data_in_frame[13] [5]), .I1(n40791), 
            .I2(n40662), .I3(n40339), .O(n37241));
    defparam i3_4_lut_adj_945.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_946 (.I0(\data_in_frame[19] [2]), .I1(\data_in_frame[16] [6]), 
            .I2(n6_adj_3239), .I3(n40752), .O(n40668));
    defparam i1_4_lut_adj_946.LUT_INIT = 16'h9669;
    SB_LUT4 i14298_2_lut_3_lut (.I0(n5_adj_3238), .I1(n43), .I2(\FRAME_MATCHER.state [5]), 
            .I3(GND_net), .O(n27700));
    defparam i14298_2_lut_3_lut.LUT_INIT = 16'he0e0;
    SB_LUT4 i2_2_lut_adj_947 (.I0(n40776), .I1(\data_in_frame[16] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n10_adj_3240));
    defparam i2_2_lut_adj_947.LUT_INIT = 16'h6666;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_3_i31_3_lut_4_lut (.I0(byte_transmit_counter_c[4]), 
            .I1(byte_transmit_counter_c[3]), .I2(n42217), .I3(n42216), 
            .O(tx_data[3]));   // verilog/coms.v(104[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_3_i31_3_lut_4_lut.LUT_INIT = 16'hf4b0;
    SB_LUT4 i6_4_lut_adj_948 (.I0(n40843), .I1(Kp_23__N_516), .I2(n40737), 
            .I3(\data_in_frame[17] [2]), .O(n14_adj_3241));
    defparam i6_4_lut_adj_948.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut_adj_949 (.I0(\data_in_frame[17] [1]), .I1(n14_adj_3241), 
            .I2(n10_adj_3240), .I3(n40653), .O(n37295));
    defparam i7_4_lut_adj_949.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_950 (.I0(n5_adj_3238), .I1(n43), .I2(\FRAME_MATCHER.state [6]), 
            .I3(GND_net), .O(n39584));
    defparam i1_2_lut_3_lut_adj_950.LUT_INIT = 16'he0e0;
    SB_LUT4 i2_3_lut_adj_951 (.I0(n37295), .I1(n40668), .I2(\data_in_frame[19] [3]), 
            .I3(GND_net), .O(n40359));
    defparam i2_3_lut_adj_951.LUT_INIT = 16'h6969;
    SB_LUT4 i1_2_lut_3_lut_adj_952 (.I0(n5_adj_3238), .I1(n43), .I2(\FRAME_MATCHER.state [7]), 
            .I3(GND_net), .O(n39650));
    defparam i1_2_lut_3_lut_adj_952.LUT_INIT = 16'he0e0;
    SB_LUT4 i3_4_lut_adj_953 (.I0(\data_in_frame[18] [1]), .I1(\data_in_frame[16] [1]), 
            .I2(\data_in_frame[18] [2]), .I3(n40487), .O(n40567));   // verilog/coms.v(72[16:43])
    defparam i3_4_lut_adj_953.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_954 (.I0(n5_adj_3238), .I1(n43), .I2(\FRAME_MATCHER.state [8]), 
            .I3(GND_net), .O(n39652));
    defparam i1_2_lut_3_lut_adj_954.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_2_lut_3_lut_adj_955 (.I0(n5_adj_3238), .I1(n43), .I2(\FRAME_MATCHER.state [9]), 
            .I3(GND_net), .O(n39654));
    defparam i1_2_lut_3_lut_adj_955.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_2_lut_adj_956 (.I0(\data_in_frame[9] [5]), .I1(n22641), .I2(GND_net), 
            .I3(GND_net), .O(n6_adj_3242));
    defparam i1_2_lut_adj_956.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_3_lut_adj_957 (.I0(n5_adj_3238), .I1(n43), .I2(\FRAME_MATCHER.state [10]), 
            .I3(GND_net), .O(n39656));
    defparam i1_2_lut_3_lut_adj_957.LUT_INIT = 16'he0e0;
    SB_LUT4 i4_4_lut_adj_958 (.I0(n16), .I1(n40495), .I2(\data_in_frame[12][1] ), 
            .I3(n6_adj_3242), .O(n40864));
    defparam i4_4_lut_adj_958.LUT_INIT = 16'h9669;
    SB_LUT4 i4_4_lut_adj_959 (.I0(n40840), .I1(n40637), .I2(\data_in_frame[7] [7]), 
            .I3(n40864), .O(n10));
    defparam i4_4_lut_adj_959.LUT_INIT = 16'h6996;
    SB_LUT4 i14878_4_lut (.I0(n28279), .I1(\FRAME_MATCHER.state [2]), .I2(\FRAME_MATCHER.state [3]), 
            .I3(n105), .O(n28289));
    defparam i14878_4_lut.LUT_INIT = 16'hfaea;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_0_i31_3_lut_4_lut (.I0(byte_transmit_counter_c[4]), 
            .I1(byte_transmit_counter_c[3]), .I2(n42208), .I3(n42207), 
            .O(tx_data[0]));   // verilog/coms.v(104[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_0_i31_3_lut_4_lut.LUT_INIT = 16'hf4b0;
    SB_LUT4 i11877_4_lut (.I0(n27701), .I1(n28285), .I2(\FRAME_MATCHER.state [1]), 
            .I3(\FRAME_MATCHER.state [0]), .O(n28293));   // verilog/coms.v(110[11:16])
    defparam i11877_4_lut.LUT_INIT = 16'hcfca;
    SB_LUT4 i13_4_lut_adj_960 (.I0(n28279), .I1(n28293), .I2(\FRAME_MATCHER.state [2]), 
            .I3(n40173), .O(n39256));   // verilog/coms.v(147[4] 288[11])
    defparam i13_4_lut_adj_960.LUT_INIT = 16'h3530;
    SB_LUT4 i1_2_lut_adj_961 (.I0(\data_in_frame[14] [7]), .I1(\data_in_frame[15] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n40867));
    defparam i1_2_lut_adj_961.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_3_lut_adj_962 (.I0(n5_adj_3238), .I1(n43), .I2(\FRAME_MATCHER.state [11]), 
            .I3(GND_net), .O(n39658));
    defparam i1_2_lut_3_lut_adj_962.LUT_INIT = 16'he0e0;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_4_i8_3_lut (.I0(\data_out_frame[8] [4]), 
            .I1(\data_out_frame[9] [4]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n8_adj_3205));   // verilog/coms.v(104[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_4_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4_4_lut_adj_963 (.I0(\data_in_frame[14] [6]), .I1(\data_in_frame[12] [6]), 
            .I2(n22816), .I3(n6_adj_3243), .O(n40365));   // verilog/coms.v(69[16:27])
    defparam i4_4_lut_adj_963.LUT_INIT = 16'h6996;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_4_i9_3_lut (.I0(\data_out_frame[10] [4]), 
            .I1(\data_out_frame[11] [4]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n9_adj_3204));   // verilog/coms.v(104[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_4_i9_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_4_i12_3_lut (.I0(\data_out_frame[14] [4]), 
            .I1(\data_out_frame[15] [4]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n12_adj_3203));   // verilog/coms.v(104[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_4_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_4_i11_3_lut (.I0(\data_out_frame[12] [4]), 
            .I1(\data_out_frame[13] [4]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n11));   // verilog/coms.v(104[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_4_i11_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_adj_964 (.I0(\data_in_frame[15] [6]), .I1(\data_in_frame[18] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n40662));
    defparam i1_2_lut_adj_964.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_3_lut_adj_965 (.I0(n5_adj_3238), .I1(n43), .I2(\FRAME_MATCHER.state [12]), 
            .I3(GND_net), .O(n39660));
    defparam i1_2_lut_3_lut_adj_965.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_2_lut_adj_966 (.I0(\data_in_frame[17] [2]), .I1(\data_in_frame[17] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n40671));   // verilog/coms.v(69[16:27])
    defparam i1_2_lut_adj_966.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_3_lut_adj_967 (.I0(n5_adj_3238), .I1(n43), .I2(\FRAME_MATCHER.state [13]), 
            .I3(GND_net), .O(n39662));
    defparam i1_2_lut_3_lut_adj_967.LUT_INIT = 16'he0e0;
    SB_LUT4 i6_4_lut_adj_968 (.I0(n22716), .I1(n40699), .I2(n40450), .I3(n40392), 
            .O(n14_adj_3244));
    defparam i6_4_lut_adj_968.LUT_INIT = 16'h6996;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_1_i31_3_lut_4_lut (.I0(byte_transmit_counter_c[4]), 
            .I1(byte_transmit_counter_c[3]), .I2(n42211), .I3(n42210), 
            .O(tx_data[1]));   // verilog/coms.v(104[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_1_i31_3_lut_4_lut.LUT_INIT = 16'hf4b0;
    SB_LUT4 i7_4_lut_adj_969 (.I0(n40460), .I1(n14_adj_3244), .I2(n10_adj_3245), 
            .I3(n23120), .O(Kp_23__N_908));
    defparam i7_4_lut_adj_969.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_970 (.I0(n22873), .I1(\data_in_frame[8] [1]), .I2(\data_in_frame[10] [1]), 
            .I3(\data_in_frame[12] [3]), .O(n40637));
    defparam i3_4_lut_adj_970.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_971 (.I0(\data_in_frame[14] [5]), .I1(n40637), 
            .I2(\data_in_frame[9] [7]), .I3(\data_in_frame[7] [5]), .O(n40776));
    defparam i3_4_lut_adj_971.LUT_INIT = 16'h6996;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_2_i31_3_lut_4_lut (.I0(byte_transmit_counter_c[4]), 
            .I1(byte_transmit_counter_c[3]), .I2(n42214), .I3(n42213), 
            .O(tx_data[2]));   // verilog/coms.v(104[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_2_i31_3_lut_4_lut.LUT_INIT = 16'hf4b0;
    SB_LUT4 i3_4_lut_adj_972 (.I0(\data_in_frame[16] [6]), .I1(\data_in_frame[16] [1]), 
            .I2(\data_in_frame[16] [3]), .I3(n22794), .O(n40693));
    defparam i3_4_lut_adj_972.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_973 (.I0(n5_adj_3238), .I1(n43), .I2(\FRAME_MATCHER.state [14]), 
            .I3(GND_net), .O(n39664));
    defparam i1_2_lut_3_lut_adj_973.LUT_INIT = 16'he0e0;
    SB_LUT4 i4_4_lut_adj_974 (.I0(n40776), .I1(n40466), .I2(n22648), .I3(n6), 
            .O(n36853));
    defparam i4_4_lut_adj_974.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_975 (.I0(\data_in_frame[10] [2]), .I1(\data_in_frame[14] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n40843));
    defparam i1_2_lut_adj_975.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_976 (.I0(\data_in_frame[8] [6]), .I1(\data_in_frame[8] [7]), 
            .I2(n40285), .I3(GND_net), .O(n41155));   // verilog/coms.v(69[16:27])
    defparam i2_3_lut_adj_976.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_977 (.I0(\FRAME_MATCHER.state [0]), .I1(n11_adj_3246), 
            .I2(\FRAME_MATCHER.state [1]), .I3(GND_net), .O(\FRAME_MATCHER.i_31__N_1821 ));   // verilog/coms.v(126[12] 289[6])
    defparam i1_2_lut_3_lut_adj_977.LUT_INIT = 16'h0202;
    SB_LUT4 i22_4_lut (.I0(\data_in_frame[6][0] ), .I1(\data_in_frame[11] [4]), 
            .I2(\data_in_frame[9] [2]), .I3(\data_in_frame[13] [0]), .O(n52));
    defparam i22_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i20_4_lut (.I0(n40867), .I1(n40788), .I2(n40840), .I3(n40755), 
            .O(n50));
    defparam i20_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_978 (.I0(n5_adj_3238), .I1(n43), .I2(\FRAME_MATCHER.state [15]), 
            .I3(GND_net), .O(n39666));
    defparam i1_2_lut_3_lut_adj_978.LUT_INIT = 16'he0e0;
    SB_LUT4 i21_4_lut (.I0(n40731), .I1(n40584), .I2(n40647), .I3(n40450), 
            .O(n51));
    defparam i21_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i19_4_lut (.I0(n41155), .I1(Kp_23__N_839), .I2(\data_in_frame[13] [1]), 
            .I3(\data_in_frame[15] [5]), .O(n49));
    defparam i19_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i16_4_lut (.I0(n40876), .I1(n40734), .I2(n40417), .I3(n22873), 
            .O(n46));
    defparam i16_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i18_4_lut (.I0(n40843), .I1(n40650), .I2(n40782), .I3(n40460), 
            .O(n48));
    defparam i18_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i17_4_lut (.I0(n40800), .I1(n22873), .I2(n40595), .I3(\data_in_frame[15] [1]), 
            .O(n47_adj_3247));
    defparam i17_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i28_4_lut (.I0(n49), .I1(n51), .I2(n50), .I3(n52), .O(n58));
    defparam i28_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_979 (.I0(\FRAME_MATCHER.state [0]), .I1(n11_adj_3246), 
            .I2(\FRAME_MATCHER.state [1]), .I3(GND_net), .O(\FRAME_MATCHER.i_31__N_1827 ));   // verilog/coms.v(126[12] 289[6])
    defparam i1_2_lut_3_lut_adj_979.LUT_INIT = 16'h2020;
    SB_LUT4 i23_3_lut (.I0(\data_in_frame[15] [4]), .I1(n46), .I2(\data_in_frame[15] [3]), 
            .I3(GND_net), .O(n53));
    defparam i23_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 i29_4_lut (.I0(n53), .I1(n58), .I2(n47_adj_3247), .I3(n48), 
            .O(n37228));
    defparam i29_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_980 (.I0(n63), .I1(\FRAME_MATCHER.state [2]), .I2(n63_adj_3248), 
            .I3(n63_adj_3249), .O(n40193));
    defparam i1_4_lut_adj_980.LUT_INIT = 16'h8a0a;
    SB_LUT4 i1_2_lut_adj_981 (.I0(\FRAME_MATCHER.i_31__N_1821 ), .I1(n740), 
            .I2(GND_net), .I3(GND_net), .O(n5_adj_3250));
    defparam i1_2_lut_adj_981.LUT_INIT = 16'h2222;
    SB_LUT4 i1_2_lut_adj_982 (.I0(\data_in_frame[16] [7]), .I1(n37228), 
            .I2(GND_net), .I3(GND_net), .O(n40598));
    defparam i1_2_lut_adj_982.LUT_INIT = 16'h6666;
    SB_LUT4 data_in_frame_18__7__I_0_3252_2_lut (.I0(\data_in_frame[18] [7]), 
            .I1(\data_in_frame[18] [6]), .I2(GND_net), .I3(GND_net), .O(Kp_23__N_786));   // verilog/coms.v(76[16:27])
    defparam data_in_frame_18__7__I_0_3252_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_983 (.I0(\data_in_frame[17] [1]), .I1(\data_in_frame[17] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n40797));
    defparam i1_2_lut_adj_983.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_984 (.I0(n41003), .I1(n15_adj_3251), .I2(\FRAME_MATCHER.i_31__N_1825 ), 
            .I3(n5_adj_3250), .O(n41586));
    defparam i3_4_lut_adj_984.LUT_INIT = 16'hfffd;
    SB_LUT4 i2_3_lut_adj_985 (.I0(n36853), .I1(\data_in_frame[15] [5]), 
            .I2(\data_in_frame[17] [5]), .I3(GND_net), .O(n37304));
    defparam i2_3_lut_adj_985.LUT_INIT = 16'h9696;
    SB_LUT4 i2_4_lut_adj_986 (.I0(\FRAME_MATCHER.i_31__N_1823 ), .I1(\FRAME_MATCHER.i_31__N_1827 ), 
            .I2(n40193), .I3(n3761), .O(n6_adj_3252));
    defparam i2_4_lut_adj_986.LUT_INIT = 16'heeea;
    SB_LUT4 i2_3_lut_adj_987 (.I0(n22250), .I1(\FRAME_MATCHER.i [31]), .I2(\FRAME_MATCHER.i_31__N_1825 ), 
            .I3(GND_net), .O(n41620));
    defparam i2_3_lut_adj_987.LUT_INIT = 16'h2020;
    SB_LUT4 i3_4_lut_adj_988 (.I0(n41620), .I1(n6_adj_3252), .I2(n41586), 
            .I3(n40193), .O(n47027));
    defparam i3_4_lut_adj_988.LUT_INIT = 16'hfeee;
    SB_LUT4 i5_4_lut_adj_989 (.I0(n40570), .I1(n40671), .I2(Kp_23__N_908), 
            .I3(n47038), .O(n12_adj_3253));
    defparam i5_4_lut_adj_989.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_990 (.I0(n37304), .I1(n12_adj_3253), .I2(n40797), 
            .I3(\data_in_frame[17] [4]), .O(n41987));
    defparam i6_4_lut_adj_990.LUT_INIT = 16'h6996;
    SB_LUT4 i2_2_lut_3_lut (.I0(\FRAME_MATCHER.state [0]), .I1(n11_adj_3246), 
            .I2(\FRAME_MATCHER.i_31__N_1825 ), .I3(GND_net), .O(n1498));   // verilog/coms.v(126[12] 289[6])
    defparam i2_2_lut_3_lut.LUT_INIT = 16'hf2f2;
    SB_LUT4 i5_4_lut_adj_991 (.I0(n40398), .I1(n40567), .I2(n41987), .I3(n40377), 
            .O(n12_adj_3254));
    defparam i5_4_lut_adj_991.LUT_INIT = 16'h9669;
    SB_LUT4 i6_4_lut_adj_992 (.I0(Kp_23__N_786), .I1(n12_adj_3254), .I2(n40598), 
            .I3(n40258), .O(n37310));
    defparam i6_4_lut_adj_992.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_993 (.I0(\data_in_frame[19] [4]), .I1(n23257), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_3255));   // verilog/coms.v(69[16:27])
    defparam i1_2_lut_adj_993.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_994 (.I0(n40365), .I1(n22648), .I2(n40671), .I3(n6_adj_3255), 
            .O(n40573));   // verilog/coms.v(69[16:27])
    defparam i4_4_lut_adj_994.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_995 (.I0(n5_adj_3238), .I1(n43), .I2(\FRAME_MATCHER.state [16]), 
            .I3(GND_net), .O(n39668));
    defparam i1_2_lut_3_lut_adj_995.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_2_lut_3_lut_adj_996 (.I0(n5_adj_3238), .I1(n43), .I2(\FRAME_MATCHER.state [17]), 
            .I3(GND_net), .O(n39670));
    defparam i1_2_lut_3_lut_adj_996.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_2_lut_3_lut_adj_997 (.I0(n5_adj_3238), .I1(n43), .I2(\FRAME_MATCHER.state [18]), 
            .I3(GND_net), .O(n39672));
    defparam i1_2_lut_3_lut_adj_997.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_2_lut_3_lut_adj_998 (.I0(n5_adj_3238), .I1(n43), .I2(\FRAME_MATCHER.state [19]), 
            .I3(GND_net), .O(n39674));
    defparam i1_2_lut_3_lut_adj_998.LUT_INIT = 16'he0e0;
    SB_LUT4 i6_4_lut_adj_999 (.I0(\data_in_frame[11] [0]), .I1(n37304), 
            .I2(n40662), .I3(n40540), .O(n16_adj_3256));
    defparam i6_4_lut_adj_999.LUT_INIT = 16'h9669;
    SB_LUT4 i3_4_lut_adj_1000 (.I0(\data_in_frame[20] [5]), .I1(n40377), 
            .I2(\data_in_frame[16] [1]), .I3(n21050), .O(n41706));
    defparam i3_4_lut_adj_1000.LUT_INIT = 16'h6996;
    SB_LUT4 i5_2_lut (.I0(\data_in_frame[13] [1]), .I1(n37310), .I2(GND_net), 
            .I3(GND_net), .O(n15_adj_3257));
    defparam i5_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i1_2_lut_3_lut_adj_1001 (.I0(n5_adj_3238), .I1(n43), .I2(\FRAME_MATCHER.state [20]), 
            .I3(GND_net), .O(n39676));
    defparam i1_2_lut_3_lut_adj_1001.LUT_INIT = 16'he0e0;
    SB_LUT4 i7_4_lut_adj_1002 (.I0(n36562), .I1(n40619), .I2(n40794), 
            .I3(n23094), .O(n17_adj_3258));
    defparam i7_4_lut_adj_1002.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1003 (.I0(\data_in_frame[19] [7]), .I1(n17_adj_3258), 
            .I2(n15_adj_3257), .I3(n16_adj_3256), .O(n40828));
    defparam i1_4_lut_adj_1003.LUT_INIT = 16'h9669;
    SB_LUT4 i7_4_lut_adj_1004 (.I0(\data_in_frame[17] [0]), .I1(n37336), 
            .I2(n40693), .I3(\data_in_frame[18] [7]), .O(n18_adj_3259));   // verilog/coms.v(83[17:28])
    defparam i7_4_lut_adj_1004.LUT_INIT = 16'h9669;
    SB_LUT4 i9_4_lut_adj_1005 (.I0(n40653), .I1(n18_adj_3259), .I2(\data_in_frame[19] [1]), 
            .I3(n40332), .O(n20_adj_3260));   // verilog/coms.v(83[17:28])
    defparam i9_4_lut_adj_1005.LUT_INIT = 16'h6996;
    SB_LUT4 i10_4_lut_adj_1006 (.I0(n15), .I1(n20_adj_3260), .I2(n37228), 
            .I3(\data_in_frame[14] [6]), .O(n40352));   // verilog/coms.v(83[17:28])
    defparam i10_4_lut_adj_1006.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_3_lut_adj_1007 (.I0(n5_adj_3238), .I1(n43), .I2(\FRAME_MATCHER.state [21]), 
            .I3(GND_net), .O(n39684));
    defparam i1_2_lut_3_lut_adj_1007.LUT_INIT = 16'he0e0;
    SB_LUT4 i2_4_lut_adj_1008 (.I0(n40352), .I1(n40828), .I2(n40573), 
            .I3(n40746), .O(n41807));
    defparam i2_4_lut_adj_1008.LUT_INIT = 16'h6996;
    SB_LUT4 i2_4_lut_adj_1009 (.I0(n22997), .I1(n40359), .I2(n40554), 
            .I3(n41807), .O(n37284));
    defparam i2_4_lut_adj_1009.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1010 (.I0(\FRAME_MATCHER.state [2]), .I1(n1_c), 
            .I2(\FRAME_MATCHER.state [3]), .I3(GND_net), .O(n11_adj_3246));
    defparam i1_2_lut_3_lut_adj_1010.LUT_INIT = 16'hfefe;
    SB_LUT4 i1_2_lut_adj_1011 (.I0(\data_in_frame[16] [4]), .I1(\data_in_frame[16] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n22794));   // verilog/coms.v(83[17:63])
    defparam i1_2_lut_adj_1011.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_1012 (.I0(\data_in_frame[18] [5]), .I1(n22794), 
            .I2(n36591), .I3(n37239), .O(n40398));
    defparam i3_4_lut_adj_1012.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1013 (.I0(\data_in_frame[15] [4]), .I1(n22721), 
            .I2(GND_net), .I3(GND_net), .O(n40794));
    defparam i1_2_lut_adj_1013.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1014 (.I0(\data_in_frame[10] [7]), .I1(\data_in_frame[13] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n40728));   // verilog/coms.v(72[16:43])
    defparam i1_2_lut_adj_1014.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1015 (.I0(\data_in_frame[10] [6]), .I1(\data_in_frame[13] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n40849));   // verilog/coms.v(70[16:41])
    defparam i1_2_lut_adj_1015.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1016 (.I0(n23101), .I1(\data_in_frame[11] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n40855));   // verilog/coms.v(69[16:27])
    defparam i1_2_lut_adj_1016.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_1017 (.I0(\data_in_frame[5] [5]), .I1(n40308), 
            .I2(\data_in_frame[3] [3]), .I3(\data_in_frame[3] [4]), .O(n22641));   // verilog/coms.v(71[16:34])
    defparam i3_4_lut_adj_1017.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1018 (.I0(\data_in_frame[10] [4]), .I1(\data_in_frame[12] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n40876));
    defparam i1_2_lut_adj_1018.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_3_lut_adj_1019 (.I0(n5_adj_3238), .I1(n43), .I2(\FRAME_MATCHER.state [22]), 
            .I3(GND_net), .O(n39686));
    defparam i1_2_lut_3_lut_adj_1019.LUT_INIT = 16'he0e0;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_31387 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[18] [5]), .I2(\data_out_frame[19] [5]), 
            .I3(byte_transmit_counter[1]), .O(n46901));
    defparam byte_transmit_counter_0__bdd_4_lut_31387.LUT_INIT = 16'he4aa;
    SB_LUT4 i4_4_lut_adj_1020 (.I0(n22641), .I1(\data_in_frame[10] [3]), 
            .I2(\data_in_frame[7] [7]), .I3(n6_adj_3261), .O(n40332));   // verilog/coms.v(69[16:27])
    defparam i4_4_lut_adj_1020.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_1021 (.I0(\data_in_frame[14] [7]), .I1(\data_in_frame[15] [1]), 
            .I2(\data_in_frame[10] [5]), .I3(n6_adj_3262), .O(n40737));   // verilog/coms.v(69[16:27])
    defparam i4_4_lut_adj_1021.LUT_INIT = 16'h6996;
    SB_LUT4 n46901_bdd_4_lut (.I0(n46901), .I1(\data_out_frame[17] [5]), 
            .I2(\data_out_frame[16] [5]), .I3(byte_transmit_counter[1]), 
            .O(n46904));
    defparam n46901_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_2_lut_3_lut_adj_1022 (.I0(n5_adj_3238), .I1(n43), .I2(\FRAME_MATCHER.state [23]), 
            .I3(GND_net), .O(n39744));
    defparam i1_2_lut_3_lut_adj_1022.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_2_lut_adj_1023 (.I0(\data_in_frame[11] [0]), .I1(\data_in_frame[6] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n40677));   // verilog/coms.v(72[16:43])
    defparam i1_2_lut_adj_1023.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1024 (.I0(n10_adj_3263), .I1(\data_in_frame[6] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n23224));   // verilog/coms.v(70[16:41])
    defparam i1_2_lut_adj_1024.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_4_lut_adj_1025 (.I0(n102), .I1(\FRAME_MATCHER.state [0]), 
            .I2(n1_c), .I3(\FRAME_MATCHER.state [1]), .O(\FRAME_MATCHER.i_31__N_1825 ));   // verilog/coms.v(126[12] 289[6])
    defparam i1_2_lut_4_lut_adj_1025.LUT_INIT = 16'h0008;
    SB_LUT4 i1_2_lut_adj_1026 (.I0(n10_adj_3263), .I1(n22716), .I2(GND_net), 
            .I3(GND_net), .O(n23098));   // verilog/coms.v(72[16:43])
    defparam i1_2_lut_adj_1026.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1027 (.I0(Kp_23__N_459), .I1(\data_in_frame[10] [4]), 
            .I2(n40322), .I3(\data_in_frame[5] [6]), .O(n10_adj_3264));   // verilog/coms.v(70[16:41])
    defparam i4_4_lut_adj_1027.LUT_INIT = 16'h6996;
    SB_LUT4 i5_3_lut_adj_1028 (.I0(\data_in_frame[5] [7]), .I1(n10_adj_3264), 
            .I2(n40481), .I3(GND_net), .O(n22816));   // verilog/coms.v(70[16:41])
    defparam i5_3_lut_adj_1028.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1029 (.I0(n22721), .I1(\data_in_frame[6] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n40392));
    defparam i1_2_lut_adj_1029.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1030 (.I0(\data_in_frame[8] [4]), .I1(n23275), 
            .I2(GND_net), .I3(GND_net), .O(n40616));   // verilog/coms.v(70[16:41])
    defparam i1_2_lut_adj_1030.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1031 (.I0(\data_in_frame[1] [5]), .I1(\data_in_frame[1] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_3265));   // verilog/coms.v(230[9:81])
    defparam i1_2_lut_adj_1031.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1032 (.I0(\data_in_frame[3] [7]), .I1(\data_in_frame[4] [1]), 
            .I2(\data_in_frame[2] [0]), .I3(n6_adj_3265), .O(n10_adj_3263));   // verilog/coms.v(230[9:81])
    defparam i4_4_lut_adj_1032.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1033 (.I0(\data_in_frame[10] [5]), .I1(\data_in_frame[8] [3]), 
            .I2(n10_adj_3263), .I3(\data_in_frame[8] [4]), .O(n40595));   // verilog/coms.v(70[16:41])
    defparam i3_4_lut_adj_1033.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1034 (.I0(n5_adj_3238), .I1(n43), .I2(\FRAME_MATCHER.state [24]), 
            .I3(GND_net), .O(n39632));
    defparam i1_2_lut_3_lut_adj_1034.LUT_INIT = 16'he0e0;
    SB_LUT4 i4_4_lut_adj_1035 (.I0(\data_in_frame[6] [3]), .I1(\data_in_frame[6][1] ), 
            .I2(n23094), .I3(n40595), .O(n10_adj_3266));   // verilog/coms.v(70[16:41])
    defparam i4_4_lut_adj_1035.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1036 (.I0(n5_adj_3238), .I1(n43), .I2(\FRAME_MATCHER.state [25]), 
            .I3(GND_net), .O(n39634));
    defparam i1_2_lut_3_lut_adj_1036.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_2_lut_3_lut_adj_1037 (.I0(n5_adj_3238), .I1(n43), .I2(\FRAME_MATCHER.state [26]), 
            .I3(GND_net), .O(n39636));
    defparam i1_2_lut_3_lut_adj_1037.LUT_INIT = 16'he0e0;
    SB_LUT4 i2_3_lut_adj_1038 (.I0(n22670), .I1(n40531), .I2(\data_in_frame[10] [7]), 
            .I3(GND_net), .O(n23350));   // verilog/coms.v(69[16:27])
    defparam i2_3_lut_adj_1038.LUT_INIT = 16'h9696;
    SB_LUT4 i3_4_lut_adj_1039 (.I0(n40677), .I1(\data_in_frame[12] [7]), 
            .I2(\data_in_frame[15] [2]), .I3(\data_in_frame[12] [6]), .O(n40800));   // verilog/coms.v(69[16:27])
    defparam i3_4_lut_adj_1039.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_1040 (.I0(n40800), .I1(n23350), .I2(n40326), 
            .I3(n22), .O(n14_adj_3268));   // verilog/coms.v(72[16:43])
    defparam i6_4_lut_adj_1040.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1041 (.I0(n5_adj_3238), .I1(n43), .I2(\FRAME_MATCHER.state [27]), 
            .I3(GND_net), .O(n39638));
    defparam i1_2_lut_3_lut_adj_1041.LUT_INIT = 16'he0e0;
    SB_LUT4 i7_4_lut_adj_1042 (.I0(n22816), .I1(n14_adj_3268), .I2(n10_adj_3269), 
            .I3(n23098), .O(n23257));   // verilog/coms.v(72[16:43])
    defparam i7_4_lut_adj_1042.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1043 (.I0(\data_in_frame[19] [6]), .I1(\data_in_frame[17] [4]), 
            .I2(n23257), .I3(\data_in_frame[17] [5]), .O(n40554));
    defparam i3_4_lut_adj_1043.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1044 (.I0(\data_in_frame[17] [4]), .I1(n40540), 
            .I2(GND_net), .I3(GND_net), .O(n14_adj_3270));   // verilog/coms.v(69[16:27])
    defparam i1_2_lut_adj_1044.LUT_INIT = 16'h6666;
    SB_LUT4 i9_4_lut_adj_1045 (.I0(n40737), .I1(\data_in_frame[8] [7]), 
            .I2(\data_in_frame[6][0] ), .I3(n40326), .O(n22_adj_3271));   // verilog/coms.v(69[16:27])
    defparam i9_4_lut_adj_1045.LUT_INIT = 16'h6996;
    SB_LUT4 i14281_2_lut_3_lut (.I0(n5_adj_3238), .I1(n43), .I2(\FRAME_MATCHER.state [28]), 
            .I3(GND_net), .O(n27682));
    defparam i14281_2_lut_3_lut.LUT_INIT = 16'he0e0;
    SB_LUT4 i8_4_lut_adj_1046 (.I0(n8_adj_3128), .I1(\data_in_frame[17] [3]), 
            .I2(n40819), .I3(n40332), .O(n21_adj_3272));   // verilog/coms.v(69[16:27])
    defparam i8_4_lut_adj_1046.LUT_INIT = 16'h6996;
    SB_LUT4 i10_4_lut_adj_1047 (.I0(n40855), .I1(n23224), .I2(n40650), 
            .I3(n14_adj_3270), .O(n23));   // verilog/coms.v(69[16:27])
    defparam i10_4_lut_adj_1047.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1048 (.I0(\data_in_frame[19] [5]), .I1(n23), .I2(n21_adj_3272), 
            .I3(n22_adj_3271), .O(n40746));
    defparam i1_4_lut_adj_1048.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_adj_1049 (.I0(n102), .I1(\FRAME_MATCHER.state [0]), 
            .I2(n1_c), .I3(\FRAME_MATCHER.state [1]), .O(\FRAME_MATCHER.i_31__N_1824 ));   // verilog/coms.v(126[12] 289[6])
    defparam i1_2_lut_4_lut_adj_1049.LUT_INIT = 16'h0800;
    SB_LUT4 i5_4_lut_adj_1050 (.I0(n40728), .I1(n40794), .I2(\data_in_frame[6] [3]), 
            .I3(n40677), .O(n12_adj_3273));   // verilog/coms.v(70[16:41])
    defparam i5_4_lut_adj_1050.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1051 (.I0(n5_adj_3238), .I1(n43), .I2(\FRAME_MATCHER.state [29]), 
            .I3(GND_net), .O(n39640));
    defparam i1_2_lut_3_lut_adj_1051.LUT_INIT = 16'he0e0;
    SB_LUT4 i6_4_lut_adj_1052 (.I0(n40285), .I1(n12_adj_3273), .I2(n40849), 
            .I3(n40616), .O(n22997));   // verilog/coms.v(70[16:41])
    defparam i6_4_lut_adj_1052.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1053 (.I0(\data_in_frame[7] [3]), .I1(n36582), 
            .I2(GND_net), .I3(GND_net), .O(n40495));
    defparam i1_2_lut_adj_1053.LUT_INIT = 16'h6666;
    SB_LUT4 i10168_3_lut_4_lut (.I0(n8_adj_3123), .I1(n40212), .I2(rx_data[0]), 
            .I3(\data_in_frame[0] [0]), .O(n23586));
    defparam i10168_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 data_in_frame_13__7__I_0_2_lut (.I0(\data_in_frame[13] [7]), .I1(\data_in_frame[13] [6]), 
            .I2(GND_net), .I3(GND_net), .O(Kp_23__N_839));   // verilog/coms.v(68[16:27])
    defparam data_in_frame_13__7__I_0_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_1054 (.I0(\data_in_frame[4] [3]), .I1(n40261), 
            .I2(\data_in_frame[1] [7]), .I3(\data_in_frame[2] [1]), .O(n22716));   // verilog/coms.v(230[9:81])
    defparam i3_4_lut_adj_1054.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1055 (.I0(\data_in_frame[11] [3]), .I1(n22716), 
            .I2(\data_in_frame[7] [1]), .I3(GND_net), .O(n40731));
    defparam i2_3_lut_adj_1055.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1056 (.I0(n5_adj_3238), .I1(n43), .I2(\FRAME_MATCHER.state [30]), 
            .I3(GND_net), .O(n39642));
    defparam i1_2_lut_3_lut_adj_1056.LUT_INIT = 16'he0e0;
    SB_LUT4 i5_4_lut_adj_1057 (.I0(\data_in_frame[4] [7]), .I1(n40528), 
            .I2(\data_in_frame[8] [7]), .I3(\data_in_frame[6] [5]), .O(n12_adj_3274));
    defparam i5_4_lut_adj_1057.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_1058 (.I0(Kp_23__N_329), .I1(n12_adj_3274), .I2(n40731), 
            .I3(\data_in_frame[9] [1]), .O(n23120));
    defparam i6_4_lut_adj_1058.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1059 (.I0(\data_in_frame[14] [0]), .I1(\data_in_frame[11] [6]), 
            .I2(\data_in_frame[11] [5]), .I3(\data_in_frame[15] [7]), .O(n40755));
    defparam i3_4_lut_adj_1059.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1060 (.I0(n40674), .I1(\data_in_frame[5] [1]), 
            .I2(n40371), .I3(GND_net), .O(n36582));
    defparam i2_3_lut_adj_1060.LUT_INIT = 16'h9696;
    SB_LUT4 i3_4_lut_adj_1061 (.I0(\data_in_frame[0] [0]), .I1(\data_in_frame[4] [4]), 
            .I2(n4_adj_3275), .I3(n40261), .O(n22721));   // verilog/coms.v(166[9:87])
    defparam i3_4_lut_adj_1061.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1062 (.I0(\data_in_frame[9] [3]), .I1(\data_in_frame[7] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n40734));
    defparam i1_2_lut_adj_1062.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_1063 (.I0(n23290), .I1(\data_in_frame[6] [7]), 
            .I2(\data_in_frame[9] [2]), .I3(\data_in_frame[6] [6]), .O(n40528));
    defparam i3_4_lut_adj_1063.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_1064 (.I0(\data_in_frame[11] [4]), .I1(n40734), 
            .I2(n22721), .I3(n36582), .O(n10_adj_3276));
    defparam i4_4_lut_adj_1064.LUT_INIT = 16'h6996;
    SB_LUT4 i5_3_lut_adj_1065 (.I0(n40528), .I1(n10_adj_3276), .I2(\data_in_frame[7] [0]), 
            .I3(GND_net), .O(n40339));
    defparam i5_3_lut_adj_1065.LUT_INIT = 16'h9696;
    SB_LUT4 i1_3_lut (.I0(\data_in_frame[13] [5]), .I1(n23120), .I2(n40339), 
            .I3(GND_net), .O(n36562));
    defparam i1_3_lut.LUT_INIT = 16'h6969;
    SB_LUT4 i2_4_lut_adj_1066 (.I0(n40339), .I1(\data_in_frame[14] [0]), 
            .I2(n40659), .I3(n37268), .O(n36591));
    defparam i2_4_lut_adj_1066.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1067 (.I0(n40755), .I1(n40858), .I2(GND_net), 
            .I3(GND_net), .O(n6_adj_3277));
    defparam i1_2_lut_adj_1067.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1068 (.I0(n36562), .I1(Kp_23__N_326), .I2(n40831), 
            .I3(n6_adj_3277), .O(n21050));
    defparam i4_4_lut_adj_1068.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1069 (.I0(n5_adj_3238), .I1(n43), .I2(\FRAME_MATCHER.state [31]), 
            .I3(GND_net), .O(n39646));
    defparam i1_2_lut_3_lut_adj_1069.LUT_INIT = 16'he0e0;
    SB_LUT4 i10513_3_lut_4_lut (.I0(n8_adj_3123), .I1(n40212), .I2(rx_data[7]), 
            .I3(\data_in_frame[0] [7]), .O(n23931));
    defparam i10513_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_1070 (.I0(\data_in_frame[15] [6]), .I1(\data_in_frame[13] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n40788));   // verilog/coms.v(72[16:43])
    defparam i1_2_lut_adj_1070.LUT_INIT = 16'h6666;
    SB_LUT4 i16_4_lut_adj_1071 (.I0(n27), .I1(n42187), .I2(n28), .I3(n30), 
            .O(\FRAME_MATCHER.state_31__N_1925 [3]));
    defparam i16_4_lut_adj_1071.LUT_INIT = 16'h2000;
    SB_LUT4 i4_4_lut_adj_1072 (.I0(\data_in_frame[21] [4]), .I1(\data_in_frame[21] [6]), 
            .I2(n40359), .I3(n47033), .O(n13_adj_3278));
    defparam i4_4_lut_adj_1072.LUT_INIT = 16'h1248;
    SB_LUT4 i2_4_lut_adj_1073 (.I0(\FRAME_MATCHER.state [2]), .I1(n41005), 
            .I2(\FRAME_MATCHER.state [1]), .I3(\FRAME_MATCHER.state [3]), 
            .O(n5021));
    defparam i2_4_lut_adj_1073.LUT_INIT = 16'h0032;
    SB_LUT4 i6_4_lut_adj_1074 (.I0(n11_adj_3216), .I1(\data_in_frame[21] [1]), 
            .I2(n41676), .I3(n37284), .O(n15_adj_3279));
    defparam i6_4_lut_adj_1074.LUT_INIT = 16'h0802;
    SB_LUT4 i1_2_lut_adj_1075 (.I0(n5021), .I1(\FRAME_MATCHER.state_31__N_1925 [3]), 
            .I2(GND_net), .I3(GND_net), .O(n22338));
    defparam i1_2_lut_adj_1075.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_3_lut_adj_1076 (.I0(n63_adj_3249), .I1(n63_adj_3248), 
            .I2(n63), .I3(GND_net), .O(n20075));
    defparam i1_2_lut_3_lut_adj_1076.LUT_INIT = 16'h8080;
    SB_LUT4 i14600_2_lut_3_lut (.I0(n63_adj_3249), .I1(n63_adj_3248), .I2(\FRAME_MATCHER.state [1]), 
            .I3(GND_net), .O(n7[1]));
    defparam i14600_2_lut_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 i30692_2_lut_3_lut (.I0(r_SM_Main_2__N_2756[0]), .I1(tx_active), 
            .I2(n28275), .I3(GND_net), .O(tx_transmit_N_2648));
    defparam i30692_2_lut_3_lut.LUT_INIT = 16'h0101;
    SB_LUT4 i3_4_lut_adj_1077 (.I0(\data_in_frame[1] [6]), .I1(\data_in_frame[2] [1]), 
            .I2(\data_in_frame[0] [0]), .I3(\data_in_frame[2] [0]), .O(n40383));   // verilog/coms.v(68[16:27])
    defparam i3_4_lut_adj_1077.LUT_INIT = 16'h6996;
    SB_LUT4 i8_4_lut_adj_1078 (.I0(n15_adj_3279), .I1(n13_adj_3278), .I2(n41706), 
            .I3(n10_adj_3218), .O(Kp_23__N_152));
    defparam i8_4_lut_adj_1078.LUT_INIT = 16'h0800;
    SB_LUT4 i1_2_lut_adj_1079 (.I0(\data_in_frame[6] [6]), .I1(\data_in_frame[9] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n40699));   // verilog/coms.v(69[16:27])
    defparam i1_2_lut_adj_1079.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_3_lut_adj_1080 (.I0(r_SM_Main_2__N_2756[0]), .I1(tx_active), 
            .I2(n28275), .I3(GND_net), .O(n736));
    defparam i1_2_lut_3_lut_adj_1080.LUT_INIT = 16'hefef;
    SB_LUT4 i1_2_lut_adj_1081 (.I0(\data_in_frame[4] [2]), .I1(n40383), 
            .I2(GND_net), .I3(GND_net), .O(n23094));   // verilog/coms.v(68[16:27])
    defparam i1_2_lut_adj_1081.LUT_INIT = 16'h6666;
    SB_LUT4 i10514_3_lut_4_lut (.I0(n8_adj_3123), .I1(n40212), .I2(rx_data[6]), 
            .I3(\data_in_frame[0] [6]), .O(n23932));
    defparam i10514_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_4_lut_adj_1082 (.I0(\FRAME_MATCHER.i [4]), .I1(n22347), 
            .I2(n22400), .I3(\FRAME_MATCHER.i [2]), .O(n4_adj_3280));   // verilog/coms.v(154[7:23])
    defparam i1_2_lut_4_lut_adj_1082.LUT_INIT = 16'hfffe;
    SB_LUT4 i5_4_lut_adj_1083 (.I0(n40819), .I1(\data_in_frame[11] [2]), 
            .I2(\data_in_frame[6] [7]), .I3(Kp_23__N_326), .O(n12_adj_3281));   // verilog/coms.v(72[16:43])
    defparam i5_4_lut_adj_1083.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_1084 (.I0(\data_in_frame[7] [0]), .I1(n12_adj_3281), 
            .I2(\data_in_frame[9] [1]), .I3(\data_in_frame[4] [6]), .O(n40285));   // verilog/coms.v(72[16:43])
    defparam i6_4_lut_adj_1084.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_adj_1085 (.I0(\FRAME_MATCHER.i [4]), .I1(n22347), 
            .I2(n22400), .I3(n27743), .O(n22250));   // verilog/coms.v(154[7:23])
    defparam i1_2_lut_4_lut_adj_1085.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1086 (.I0(n7[1]), .I1(n63), .I2(n41992), 
            .I3(n15_adj_3251), .O(n39504));
    defparam i1_2_lut_3_lut_4_lut_adj_1086.LUT_INIT = 16'hbb0b;
    SB_LUT4 i2_3_lut_adj_1087 (.I0(n40619), .I1(\data_in_frame[13] [4]), 
            .I2(n40285), .I3(GND_net), .O(n40791));   // verilog/coms.v(76[16:50])
    defparam i2_3_lut_adj_1087.LUT_INIT = 16'h9696;
    SB_LUT4 i10369_3_lut_4_lut (.I0(n8_adj_3124), .I1(n40205), .I2(rx_data[7]), 
            .I3(\data_in_frame[18] [7]), .O(n23787));
    defparam i10369_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i3_4_lut_adj_1088 (.I0(Kp_23__N_839), .I1(n40495), .I2(n40758), 
            .I3(n40591), .O(n40659));
    defparam i3_4_lut_adj_1088.LUT_INIT = 16'h9669;
    SB_LUT4 i10370_3_lut_4_lut (.I0(n8_adj_3124), .I1(n40205), .I2(rx_data[6]), 
            .I3(\data_in_frame[18] [6]), .O(n23788));
    defparam i10370_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10515_3_lut_4_lut (.I0(n8_adj_3123), .I1(n40212), .I2(rx_data[5]), 
            .I3(\data_in_frame[0] [5]), .O(n23933));
    defparam i10515_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10371_3_lut_4_lut (.I0(n8_adj_3124), .I1(n40205), .I2(rx_data[5]), 
            .I3(\data_in_frame[18] [5]), .O(n23789));
    defparam i10371_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_1089 (.I0(n40659), .I1(n40791), .I2(GND_net), 
            .I3(GND_net), .O(n6_adj_3282));   // verilog/coms.v(72[16:43])
    defparam i1_2_lut_adj_1089.LUT_INIT = 16'h6666;
    SB_LUT4 i4048_2_lut (.I0(\FRAME_MATCHER.state [0]), .I1(\FRAME_MATCHER.state [1]), 
            .I2(GND_net), .I3(GND_net), .O(n19614));
    defparam i4048_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i29331_4_lut (.I0(n27693), .I1(n102), .I2(n28279), .I3(\FRAME_MATCHER.state [0]), 
            .O(n44105));   // verilog/coms.v(110[11:16])
    defparam i29331_4_lut.LUT_INIT = 16'h0c04;
    SB_LUT4 i10372_3_lut_4_lut (.I0(n8_adj_3124), .I1(n40205), .I2(rx_data[4]), 
            .I3(\data_in_frame[18] [4]), .O(n23790));
    defparam i10372_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i4_4_lut_adj_1090 (.I0(\data_in_frame[16] [0]), .I1(\data_in_frame[14] [0]), 
            .I2(n40788), .I3(n6_adj_3282), .O(n40487));   // verilog/coms.v(72[16:43])
    defparam i4_4_lut_adj_1090.LUT_INIT = 16'h6996;
    SB_LUT4 i11817_4_lut (.I0(n8_adj_3283), .I1(n44105), .I2(\FRAME_MATCHER.state [1]), 
            .I3(n41005), .O(n23400));   // verilog/coms.v(110[11:16])
    defparam i11817_4_lut.LUT_INIT = 16'hc0ca;
    SB_LUT4 i10373_3_lut_4_lut (.I0(n8_adj_3124), .I1(n40205), .I2(rx_data[3]), 
            .I3(\data_in_frame[18] [3]), .O(n23791));
    defparam i10373_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_1091 (.I0(n21050), .I1(n36591), .I2(GND_net), 
            .I3(GND_net), .O(n40420));
    defparam i1_2_lut_adj_1091.LUT_INIT = 16'h6666;
    SB_LUT4 i10374_3_lut_4_lut (.I0(n8_adj_3124), .I1(n40205), .I2(rx_data[2]), 
            .I3(\data_in_frame[18] [2]), .O(n23792));
    defparam i10374_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_3_lut_adj_1092 (.I0(\data_in_frame[0] [2]), .I1(\data_in_frame[2] [3]), 
            .I2(\data_in_frame[0] [1]), .I3(GND_net), .O(n4_adj_3275));   // verilog/coms.v(166[9:87])
    defparam i2_3_lut_adj_1092.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_adj_1093 (.I0(\data_in_frame[4] [5]), .I1(n5_adj_3135), 
            .I2(n4_adj_3275), .I3(GND_net), .O(n23101));   // verilog/coms.v(230[9:81])
    defparam i2_3_lut_adj_1093.LUT_INIT = 16'h9696;
    SB_LUT4 i3_4_lut_adj_1094 (.I0(n41662), .I1(\data_in_frame[0] [5]), 
            .I2(\data_in_frame[0] [7]), .I3(\data_in_frame[1] [0]), .O(n40371));   // verilog/coms.v(68[16:69])
    defparam i3_4_lut_adj_1094.LUT_INIT = 16'h6996;
    SB_LUT4 i10375_3_lut_4_lut (.I0(n8_adj_3124), .I1(n40205), .I2(rx_data[1]), 
            .I3(\data_in_frame[18] [1]), .O(n23793));
    defparam i10375_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10376_3_lut_4_lut (.I0(n8_adj_3124), .I1(n40205), .I2(rx_data[0]), 
            .I3(\data_in_frame[18] [0]), .O(n23794));
    defparam i10376_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i5_4_lut_adj_1095 (.I0(\data_out_frame[20][7] ), .I1(n40279), 
            .I2(n40612), .I3(n40761), .O(n12_adj_3284));
    defparam i5_4_lut_adj_1095.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_1096 (.I0(\data_out_frame[7] [0]), .I1(\data_out_frame[7] [1]), 
            .I2(\data_out_frame[7] [3]), .I3(\data_out_frame[7] [2]), .O(n40628));
    defparam i2_3_lut_4_lut_adj_1096.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_1097 (.I0(\data_out_frame[7] [0]), .I1(\data_out_frame[7] [1]), 
            .I2(n40292), .I3(n23166), .O(n41642));
    defparam i2_3_lut_4_lut_adj_1097.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_adj_1098 (.I0(n40401), .I1(n10_adj_3285), .I2(n40282), 
            .I3(n40380), .O(n37253));   // verilog/coms.v(71[16:27])
    defparam i1_2_lut_4_lut_adj_1098.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_1099 (.I0(\data_out_frame[20] [6]), .I1(n12_adj_3284), 
            .I2(n40822), .I3(\data_out_frame[14] [0]), .O(n41847));
    defparam i6_4_lut_adj_1099.LUT_INIT = 16'h6996;
    SB_LUT4 i10516_3_lut_4_lut (.I0(n8_adj_3123), .I1(n40212), .I2(rx_data[4]), 
            .I3(\data_in_frame[0] [4]), .O(n23934));
    defparam i10516_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i3_4_lut_adj_1100 (.I0(n41673), .I1(n41806), .I2(\data_out_frame[20][7] ), 
            .I3(n36572), .O(n8_adj_3286));
    defparam i3_4_lut_adj_1100.LUT_INIT = 16'h9669;
    SB_LUT4 i4_3_lut (.I0(n36494), .I1(n8_adj_3286), .I2(n22729), .I3(GND_net), 
            .O(n41498));
    defparam i4_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 i4_4_lut_adj_1101 (.I0(n40690), .I1(\data_out_frame[18] [6]), 
            .I2(n40415), .I3(n40810), .O(n10_adj_3287));
    defparam i4_4_lut_adj_1101.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_adj_1102 (.I0(n36991), .I1(n40490), .I2(GND_net), 
            .I3(GND_net), .O(n36572));
    defparam i1_2_lut_adj_1102.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_1103 (.I0(\data_out_frame[17] [1]), .I1(n40329), 
            .I2(n23285), .I3(n36572), .O(n41672));   // verilog/coms.v(76[16:27])
    defparam i3_4_lut_adj_1103.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_adj_1104 (.I0(n40401), .I1(n10_adj_3285), .I2(n40282), 
            .I3(\data_out_frame[13] [6]), .O(n36529));   // verilog/coms.v(71[16:27])
    defparam i1_2_lut_4_lut_adj_1104.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1105 (.I0(\data_out_frame[17] [1]), .I1(n40535), 
            .I2(n40490), .I3(\data_out_frame[19] [2]), .O(n41339));
    defparam i3_4_lut_adj_1105.LUT_INIT = 16'h9669;
    SB_LUT4 i2_2_lut_adj_1106 (.I0(n36532), .I1(\data_out_frame[16] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n10_adj_3288));
    defparam i2_2_lut_adj_1106.LUT_INIT = 16'h6666;
    SB_LUT4 i6_4_lut_adj_1107 (.I0(n40356), .I1(n22729), .I2(\data_out_frame[15] [1]), 
            .I3(n22132), .O(n14_adj_3289));
    defparam i6_4_lut_adj_1107.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut_adj_1108 (.I0(n40551), .I1(n14_adj_3289), .I2(n10_adj_3288), 
            .I3(n1695), .O(n41673));
    defparam i7_4_lut_adj_1108.LUT_INIT = 16'h6996;
    SB_LUT4 i1_3_lut_adj_1109 (.I0(n23285), .I1(n41673), .I2(\data_out_frame[19][3] ), 
            .I3(GND_net), .O(n40535));   // verilog/coms.v(71[16:42])
    defparam i1_3_lut_adj_1109.LUT_INIT = 16'h9696;
    SB_LUT4 i10517_3_lut_4_lut (.I0(n8_adj_3123), .I1(n40212), .I2(rx_data[3]), 
            .I3(\data_in_frame[0] [3]), .O(n23935));
    defparam i10517_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_3_lut_adj_1110 (.I0(n40561), .I1(n40641), .I2(n40535), 
            .I3(GND_net), .O(n41129));   // verilog/coms.v(71[16:42])
    defparam i2_3_lut_adj_1110.LUT_INIT = 16'h9696;
    SB_LUT4 i3_4_lut_adj_1111 (.I0(\data_out_frame[12] [6]), .I1(n40785), 
            .I2(n40656), .I3(n1695), .O(n23285));
    defparam i3_4_lut_adj_1111.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1112 (.I0(\data_out_frame[19] [4]), .I1(\data_out_frame[17] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n40641));   // verilog/coms.v(71[16:42])
    defparam i1_2_lut_adj_1112.LUT_INIT = 16'h6666;
    SB_LUT4 i5_4_lut_adj_1113 (.I0(n23316), .I1(n40311), .I2(n36597), 
            .I3(\data_out_frame[17] [4]), .O(n12_adj_3290));   // verilog/coms.v(71[16:42])
    defparam i5_4_lut_adj_1113.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_1114 (.I0(\data_out_frame[19] [5]), .I1(n12_adj_3290), 
            .I2(n40641), .I3(n23285), .O(n41124));   // verilog/coms.v(71[16:42])
    defparam i6_4_lut_adj_1114.LUT_INIT = 16'h6996;
    SB_LUT4 i5_4_lut_adj_1115 (.I0(n40767), .I1(n40837), .I2(\data_out_frame[8] [5]), 
            .I3(n40631), .O(n12_adj_3291));
    defparam i5_4_lut_adj_1115.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_adj_1116 (.I0(n40401), .I1(n10_adj_3285), .I2(n40282), 
            .I3(\data_out_frame[16] [2]), .O(n40822));   // verilog/coms.v(71[16:27])
    defparam i1_2_lut_4_lut_adj_1116.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_1117 (.I0(\data_out_frame[6] [3]), .I1(n12_adj_3291), 
            .I2(n40861), .I3(n22132), .O(n36532));
    defparam i6_4_lut_adj_1117.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1118 (.I0(\data_out_frame[14] [7]), .I1(n36532), 
            .I2(\data_out_frame[15] [1]), .I3(GND_net), .O(n36597));
    defparam i2_3_lut_adj_1118.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1119 (.I0(\data_out_frame[5] [5]), .I1(\data_out_frame[7] [7]), 
            .I2(\data_out_frame[9] [7]), .I3(GND_net), .O(n40723));   // verilog/coms.v(73[16:27])
    defparam i1_2_lut_3_lut_adj_1119.LUT_INIT = 16'h9696;
    SB_LUT4 i2_2_lut_3_lut_4_lut (.I0(\data_out_frame[5] [5]), .I1(\data_out_frame[7] [7]), 
            .I2(n40665), .I3(n40349), .O(n22047));   // verilog/coms.v(73[16:27])
    defparam i2_2_lut_3_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1120 (.I0(\data_out_frame[17] [3]), .I1(n23316), 
            .I2(GND_net), .I3(GND_net), .O(n40561));
    defparam i1_2_lut_adj_1120.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1121 (.I0(n40561), .I1(\data_out_frame[19] [5]), 
            .I2(n36494), .I3(n36629), .O(n10_adj_3292));
    defparam i4_4_lut_adj_1121.LUT_INIT = 16'h6996;
    SB_LUT4 i5_3_lut_adj_1122 (.I0(\data_out_frame[19] [6]), .I1(n10_adj_3292), 
            .I2(n41402), .I3(GND_net), .O(n41732));
    defparam i5_3_lut_adj_1122.LUT_INIT = 16'h6969;
    SB_LUT4 i1_2_lut_adj_1123 (.I0(n36837), .I1(\data_out_frame[18] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n40761));
    defparam i1_2_lut_adj_1123.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1124 (.I0(\data_out_frame[5] [5]), .I1(\data_out_frame[7] [7]), 
            .I2(n40506), .I3(n40349), .O(n40474));   // verilog/coms.v(73[16:27])
    defparam i1_2_lut_3_lut_4_lut_adj_1124.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1125 (.I0(\data_out_frame[19] [2]), .I1(\data_out_frame[19] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n40329));   // verilog/coms.v(76[16:27])
    defparam i1_2_lut_adj_1125.LUT_INIT = 16'h6666;
    SB_LUT4 i13_4_lut_adj_1126 (.I0(\data_out_frame[17] [6]), .I1(\data_out_frame[18] [7]), 
            .I2(n37234), .I3(n18_adj_3293), .O(n30_adj_3294));
    defparam i13_4_lut_adj_1126.LUT_INIT = 16'h6996;
    SB_LUT4 i11_4_lut_adj_1127 (.I0(\data_out_frame[17] [5]), .I1(n40714), 
            .I2(\data_out_frame[18][3] ), .I3(\data_out_frame[17] [7]), 
            .O(n28_adj_3295));
    defparam i11_4_lut_adj_1127.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1128 (.I0(\data_out_frame[5] [4]), .I1(\data_out_frame[8] [0]), 
            .I2(\data_out_frame[5] [6]), .I3(GND_net), .O(n22635));
    defparam i1_2_lut_3_lut_adj_1128.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_4_lut_adj_1129 (.I0(\data_out_frame[5] [4]), .I1(\data_out_frame[8] [0]), 
            .I2(n40764), .I3(\data_out_frame[8] [1]), .O(n40609));
    defparam i2_3_lut_4_lut_adj_1129.LUT_INIT = 16'h6996;
    SB_LUT4 i12_4_lut (.I0(n23383), .I1(n40588), .I2(n40761), .I3(\data_out_frame[16] [5]), 
            .O(n29));
    defparam i12_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_1130 (.I0(\data_out_frame[9] [2]), .I1(\data_out_frame[9] [0]), 
            .I2(\data_out_frame[7] [4]), .I3(\data_out_frame[11] [6]), .O(n40622));
    defparam i2_3_lut_4_lut_adj_1130.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_1131 (.I0(\data_out_frame[9] [2]), .I1(\data_out_frame[9] [0]), 
            .I2(\data_out_frame[5] [0]), .I3(n40870), .O(n40292));
    defparam i2_3_lut_4_lut_adj_1131.LUT_INIT = 16'h6996;
    SB_LUT4 i10_4_lut_adj_1132 (.I0(\data_out_frame[19][3] ), .I1(\data_out_frame[19] [4]), 
            .I2(n40581), .I3(n40368), .O(n27_adj_3296));
    defparam i10_4_lut_adj_1132.LUT_INIT = 16'h6996;
    SB_LUT4 i16_4_lut_adj_1133 (.I0(n27_adj_3296), .I1(n29), .I2(n28_adj_3295), 
            .I3(n30_adj_3294), .O(n41806));
    defparam i16_4_lut_adj_1133.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1134 (.I0(\data_out_frame[20] [2]), .I1(n37246), 
            .I2(n36588), .I3(GND_net), .O(n40448));
    defparam i1_2_lut_3_lut_adj_1134.LUT_INIT = 16'h9696;
    SB_LUT4 i10518_3_lut_4_lut (.I0(n8_adj_3123), .I1(n40212), .I2(rx_data[2]), 
            .I3(\data_in_frame[0] [2]), .O(n23936));
    defparam i10518_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_1135 (.I0(\data_out_frame[12] [5]), .I1(\data_out_frame[14] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n40356));
    defparam i1_2_lut_adj_1135.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1136 (.I0(\data_out_frame[17] [5]), .I1(n1787), 
            .I2(GND_net), .I3(GND_net), .O(n40558));
    defparam i1_2_lut_adj_1136.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1137 (.I0(\data_out_frame[18] [7]), .I1(\data_out_frame[16] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n40690));
    defparam i1_2_lut_adj_1137.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1138 (.I0(\data_out_frame[20] [2]), .I1(n37246), 
            .I2(n41416), .I3(\data_out_frame[20] [1]), .O(n40449));
    defparam i1_2_lut_3_lut_4_lut_adj_1138.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1139 (.I0(n22840), .I1(n40813), .I2(n40690), 
            .I3(n40576), .O(n42020));
    defparam i3_4_lut_adj_1139.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1140 (.I0(n40825), .I1(\data_out_frame[16] [3]), 
            .I2(n42020), .I3(n40577), .O(n36991));
    defparam i3_4_lut_adj_1140.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_3_lut_adj_1141 (.I0(\data_out_frame[11] [0]), .I1(n40861), 
            .I2(\data_out_frame[12] [6]), .I3(GND_net), .O(n40770));   // verilog/coms.v(72[16:27])
    defparam i1_2_lut_3_lut_adj_1141.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1142 (.I0(\data_out_frame[11] [0]), .I1(n40861), 
            .I2(\data_out_frame[6] [6]), .I3(GND_net), .O(n6_adj_3297));   // verilog/coms.v(72[16:27])
    defparam i1_2_lut_3_lut_adj_1142.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1143 (.I0(n36991), .I1(\data_out_frame[19] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n40810));
    defparam i1_2_lut_adj_1143.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_1144 (.I0(\data_out_frame[15] [0]), .I1(n40474), 
            .I2(n40298), .I3(n22666), .O(n40785));
    defparam i3_4_lut_adj_1144.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1145 (.I0(\data_out_frame[16] [4]), .I1(\data_out_frame[16] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n40612));
    defparam i1_2_lut_adj_1145.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1146 (.I0(n40453), .I1(\data_out_frame[20][7] ), 
            .I2(n37308), .I3(n40703), .O(n10_adj_3298));
    defparam i4_4_lut_adj_1146.LUT_INIT = 16'h6996;
    SB_LUT4 i5_3_lut_adj_1147 (.I0(\data_out_frame[20] [2]), .I1(n10_adj_3298), 
            .I2(\data_out_frame[20] [1]), .I3(GND_net), .O(n41192));
    defparam i5_3_lut_adj_1147.LUT_INIT = 16'h9696;
    SB_LUT4 i3_4_lut_adj_1148 (.I0(n37246), .I1(n41416), .I2(n41192), 
            .I3(n22071), .O(n36629));
    defparam i3_4_lut_adj_1148.LUT_INIT = 16'h6996;
    SB_LUT4 i10_4_lut_adj_1149 (.I0(n40813), .I1(n22047), .I2(n36837), 
            .I3(\data_out_frame[18] [7]), .O(n28_adj_3299));
    defparam i10_4_lut_adj_1149.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1150 (.I0(\data_out_frame[20] [1]), .I1(n41416), 
            .I2(n41402), .I3(GND_net), .O(n40375));
    defparam i1_2_lut_3_lut_adj_1150.LUT_INIT = 16'h6969;
    SB_LUT4 i12_4_lut_adj_1151 (.I0(n22134), .I1(\data_out_frame[15] [0]), 
            .I2(n40429), .I3(n40558), .O(n30_adj_3300));
    defparam i12_4_lut_adj_1151.LUT_INIT = 16'h6996;
    SB_LUT4 i13_4_lut_adj_1152 (.I0(\data_out_frame[17] [0]), .I1(n40785), 
            .I2(n40408), .I3(n40810), .O(n31));
    defparam i13_4_lut_adj_1152.LUT_INIT = 16'h6996;
    SB_LUT4 i11_4_lut_adj_1153 (.I0(n40356), .I1(n41806), .I2(\data_out_frame[18] [5]), 
            .I3(n23169), .O(n29_adj_3301));
    defparam i11_4_lut_adj_1153.LUT_INIT = 16'h9669;
    SB_LUT4 i17_4_lut_adj_1154 (.I0(n29_adj_3301), .I1(n31), .I2(n30_adj_3300), 
            .I3(n32), .O(n37255));
    defparam i17_4_lut_adj_1154.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1155 (.I0(n37255), .I1(n36629), .I2(GND_net), 
            .I3(GND_net), .O(n40513));
    defparam i1_2_lut_adj_1155.LUT_INIT = 16'h6666;
    SB_LUT4 i5_3_lut_4_lut (.I0(\data_out_frame[17] [3]), .I1(n22729), .I2(n37234), 
            .I3(n10_adj_3302), .O(n41416));
    defparam i5_3_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_1156 (.I0(\data_out_frame[5] [7]), .I1(n40343), 
            .I2(n22666), .I3(\data_out_frame[10] [5]), .O(n40429));
    defparam i2_3_lut_4_lut_adj_1156.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1157 (.I0(\data_out_frame[6] [4]), .I1(\data_out_frame[13] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n40837));
    defparam i1_2_lut_adj_1157.LUT_INIT = 16'h6666;
    SB_LUT4 i1_4_lut_adj_1158 (.I0(n40110), .I1(n31577), .I2(n40247), 
            .I3(n40106), .O(n1_c));
    defparam i1_4_lut_adj_1158.LUT_INIT = 16'hfffe;
    SB_LUT4 i3_4_lut_adj_1159 (.I0(n22515), .I1(n40423), .I2(n1595), .I3(\data_out_frame[13] [1]), 
            .O(n1787));   // verilog/coms.v(71[16:42])
    defparam i3_4_lut_adj_1159.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_1160 (.I0(\data_out_frame[8] [6]), .I1(n40770), 
            .I2(n40665), .I3(n6_adj_3303), .O(n41850));   // verilog/coms.v(73[16:27])
    defparam i4_4_lut_adj_1160.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_1161 (.I0(\data_out_frame[13] [1]), .I1(n41850), 
            .I2(n40837), .I3(\data_out_frame[15] [2]), .O(n23316));   // verilog/coms.v(73[16:27])
    defparam i6_4_lut_adj_1161.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1162 (.I0(\data_out_frame[19] [6]), .I1(\data_out_frame[19] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n40581));
    defparam i1_2_lut_adj_1162.LUT_INIT = 16'h6666;
    SB_LUT4 i5_4_lut_adj_1163 (.I0(n23107), .I1(n40581), .I2(\data_out_frame[20] [0]), 
            .I3(n40577), .O(n12_adj_3304));
    defparam i5_4_lut_adj_1163.LUT_INIT = 16'h9669;
    SB_LUT4 i6_4_lut_adj_1164 (.I0(n23316), .I1(n12_adj_3304), .I2(n40749), 
            .I3(n1787), .O(n41402));
    defparam i6_4_lut_adj_1164.LUT_INIT = 16'h6996;
    SB_LUT4 mux_923_i1_3_lut_4_lut (.I0(\FRAME_MATCHER.state [1]), .I1(n27693), 
            .I2(\data_in_frame[3] [0]), .I3(\data_in_frame[16] [0]), .O(n3792));
    defparam mux_923_i1_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i939_2_lut (.I0(\data_out_frame[14] [7]), .I1(\data_out_frame[14] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n1695));   // verilog/coms.v(69[16:27])
    defparam i939_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1165 (.I0(\data_out_frame[15] [3]), .I1(\data_out_frame[15] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n40423));   // verilog/coms.v(71[16:42])
    defparam i1_2_lut_adj_1165.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_1166 (.I0(\data_out_frame[10] [2]), .I1(n40496), 
            .I2(\data_out_frame[14] [4]), .I3(GND_net), .O(n36837));
    defparam i2_3_lut_adj_1166.LUT_INIT = 16'h9696;
    SB_LUT4 i14299_2_lut (.I0(Kp_23__N_152), .I1(n27691), .I2(GND_net), 
            .I3(GND_net), .O(n27701));
    defparam i14299_2_lut.LUT_INIT = 16'hdddd;
    SB_LUT4 i1_2_lut_adj_1167 (.I0(\data_out_frame[10] [2]), .I1(n22095), 
            .I2(GND_net), .I3(GND_net), .O(n40408));   // verilog/coms.v(73[16:27])
    defparam i1_2_lut_adj_1167.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1168 (.I0(\data_out_frame[12] [3]), .I1(n40723), 
            .I2(n40408), .I3(\data_out_frame[10] [1]), .O(n10_adj_3305));   // verilog/coms.v(73[16:27])
    defparam i4_4_lut_adj_1168.LUT_INIT = 16'h6996;
    SB_LUT4 i10519_3_lut_4_lut (.I0(n8_adj_3123), .I1(n40212), .I2(rx_data[1]), 
            .I3(\data_in_frame[0] [1]), .O(n23937));
    defparam i10519_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1816_3_lut (.I0(Kp_23__N_152), .I1(n31_adj_3306), .I2(\FRAME_MATCHER.state [1]), 
            .I3(GND_net), .O(n19864));
    defparam i1816_3_lut.LUT_INIT = 16'hc5c5;
    SB_LUT4 i1_2_lut_adj_1169 (.I0(\data_out_frame[14] [5]), .I1(n22134), 
            .I2(GND_net), .I3(GND_net), .O(n40414));
    defparam i1_2_lut_adj_1169.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_1170 (.I0(Kp_23__N_326), .I1(n22641), .I2(\data_in_frame[4] [6]), 
            .I3(GND_net), .O(n6_adj_3307));   // verilog/coms.v(230[9:81])
    defparam i2_3_lut_adj_1170.LUT_INIT = 16'h7b7b;
    SB_LUT4 i1_2_lut_adj_1171 (.I0(\data_out_frame[10] [3]), .I1(n40474), 
            .I2(GND_net), .I3(GND_net), .O(n22132));
    defparam i1_2_lut_adj_1171.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_1172 (.I0(Kp_23__N_459), .I1(n6_adj_3307), .I2(n22842), 
            .I3(\data_in_frame[5] [6]), .O(n41802));   // verilog/coms.v(230[9:81])
    defparam i3_4_lut_adj_1172.LUT_INIT = 16'hdfef;
    SB_LUT4 i1_2_lut_adj_1173 (.I0(\data_out_frame[5] [6]), .I1(\data_out_frame[5] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n23038));   // verilog/coms.v(71[16:34])
    defparam i1_2_lut_adj_1173.LUT_INIT = 16'h6666;
    SB_LUT4 i9_4_lut_adj_1174 (.I0(n23290), .I1(n22716), .I2(n16), .I3(n22721), 
            .O(n22_adj_3308));   // verilog/coms.v(230[9:81])
    defparam i9_4_lut_adj_1174.LUT_INIT = 16'hfffe;
    SB_LUT4 i3_4_lut_adj_1175 (.I0(\data_out_frame[12] [2]), .I1(n22095), 
            .I2(\data_out_frame[12] [3]), .I3(n23000), .O(n40496));
    defparam i3_4_lut_adj_1175.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1176 (.I0(\data_out_frame[12] [4]), .I1(\data_out_frame[10] [3]), 
            .I2(\data_out_frame[10] [2]), .I3(GND_net), .O(n40335));
    defparam i2_3_lut_adj_1176.LUT_INIT = 16'h9696;
    SB_LUT4 i7_3_lut (.I0(n36582), .I1(n10_adj_3263), .I2(n23157), .I3(GND_net), 
            .O(n20_adj_3309));   // verilog/coms.v(230[9:81])
    defparam i7_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i1_2_lut_adj_1177 (.I0(\data_out_frame[6] [3]), .I1(\data_out_frame[6] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n22666));   // verilog/coms.v(72[16:27])
    defparam i1_2_lut_adj_1177.LUT_INIT = 16'h6666;
    SB_LUT4 i11_4_lut_adj_1178 (.I0(n23094), .I1(n22_adj_3308), .I2(n16_adj_3310), 
            .I3(n41802), .O(n24));   // verilog/coms.v(230[9:81])
    defparam i11_4_lut_adj_1178.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_adj_1179 (.I0(\data_out_frame[6] [2]), .I1(\data_out_frame[6] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n23248));   // verilog/coms.v(69[16:62])
    defparam i1_2_lut_adj_1179.LUT_INIT = 16'h6666;
    SB_LUT4 i12_4_lut_adj_1180 (.I0(n22873), .I1(n24), .I2(n20_adj_3309), 
            .I3(n23275), .O(n31_adj_3306));   // verilog/coms.v(230[9:81])
    defparam i12_4_lut_adj_1180.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_adj_1181 (.I0(\data_out_frame[6] [1]), .I1(\data_out_frame[8] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n40349));   // verilog/coms.v(71[16:34])
    defparam i1_2_lut_adj_1181.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1182 (.I0(\data_out_frame[12] [5]), .I1(\data_out_frame[12] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n40631));
    defparam i1_2_lut_adj_1182.LUT_INIT = 16'h6666;
    SB_LUT4 i17_4_lut_adj_1183 (.I0(n40631), .I1(n40770), .I2(n40349), 
            .I3(n40518), .O(n48_adj_3311));
    defparam i17_4_lut_adj_1183.LUT_INIT = 16'h6996;
    SB_LUT4 i14292_2_lut (.I0(n31_adj_3306), .I1(n27691), .I2(GND_net), 
            .I3(GND_net), .O(n27693));
    defparam i14292_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i23_4_lut (.I0(n23248), .I1(\data_out_frame[6] [4]), .I2(n40604), 
            .I3(\data_out_frame[6] [5]), .O(n54));
    defparam i23_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 mux_923_i2_3_lut_4_lut (.I0(\FRAME_MATCHER.state [1]), .I1(n27693), 
            .I2(\data_in_frame[3] [1]), .I3(\data_in_frame[16] [1]), .O(n3793));
    defparam mux_923_i2_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i21_4_lut_adj_1184 (.I0(n40609), .I1(n40628), .I2(n23004), 
            .I3(n40401), .O(n52_adj_3312));
    defparam i21_4_lut_adj_1184.LUT_INIT = 16'h6996;
    SB_LUT4 i22_4_lut_adj_1185 (.I0(\data_out_frame[7] [7]), .I1(n22630), 
            .I2(n22666), .I3(n40282), .O(n53_adj_3313));
    defparam i22_4_lut_adj_1185.LUT_INIT = 16'h6996;
    SB_LUT4 i20_4_lut_adj_1186 (.I0(\data_out_frame[5] [0]), .I1(n40335), 
            .I2(\data_out_frame[11] [4]), .I3(n40343), .O(n51_adj_3314));
    defparam i20_4_lut_adj_1186.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1187 (.I0(n27691), .I1(n28279), .I2(n93), .I3(n19864), 
            .O(n23430));
    defparam i3_4_lut_adj_1187.LUT_INIT = 16'h0010;
    SB_LUT4 i19_4_lut_adj_1188 (.I0(n40622), .I1(n40496), .I2(n40506), 
            .I3(n40386), .O(n50_adj_3315));
    defparam i19_4_lut_adj_1188.LUT_INIT = 16'h6996;
    SB_LUT4 i25_4_lut (.I0(n40429), .I1(n50_adj_3315), .I2(n36), .I3(\data_out_frame[8] [2]), 
            .O(n56));
    defparam i25_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i29_4_lut_adj_1189 (.I0(n51_adj_3314), .I1(n53_adj_3313), .I2(n52_adj_3312), 
            .I3(n54), .O(n60));
    defparam i29_4_lut_adj_1189.LUT_INIT = 16'h6996;
    SB_LUT4 i24_4_lut (.I0(n23038), .I1(n48_adj_3311), .I2(\data_out_frame[11] [3]), 
            .I3(n40499), .O(n55));
    defparam i24_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1190 (.I0(n55), .I1(\data_out_frame[13] [0]), .I2(n60), 
            .I3(n56), .O(n37341));
    defparam i1_4_lut_adj_1190.LUT_INIT = 16'h6996;
    SB_LUT4 mux_923_i3_3_lut_4_lut (.I0(\FRAME_MATCHER.state [1]), .I1(n27693), 
            .I2(\data_in_frame[3] [2]), .I3(\data_in_frame[16] [2]), .O(n3794));
    defparam mux_923_i3_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 mux_923_i4_3_lut_4_lut (.I0(\FRAME_MATCHER.state [1]), .I1(n27693), 
            .I2(\data_in_frame[3] [3]), .I3(\data_in_frame[16] [3]), .O(n3795));
    defparam mux_923_i4_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i6_4_lut_adj_1191 (.I0(n1664), .I1(n37341), .I2(n40852), .I3(n40720), 
            .O(n16_adj_3316));
    defparam i6_4_lut_adj_1191.LUT_INIT = 16'h9669;
    SB_LUT4 i7_4_lut_adj_1192 (.I0(\data_out_frame[13] [3]), .I1(n40806), 
            .I2(n40873), .I3(n40499), .O(n17_adj_3317));
    defparam i7_4_lut_adj_1192.LUT_INIT = 16'h6996;
    SB_LUT4 i11_4_lut_adj_1193 (.I0(n1515), .I1(n40414), .I2(\data_out_frame[15] [2]), 
            .I3(\data_out_frame[15] [1]), .O(n30_adj_3318));
    defparam i11_4_lut_adj_1193.LUT_INIT = 16'h6996;
    SB_LUT4 i9_4_lut_adj_1194 (.I0(n17_adj_3317), .I1(n22511), .I2(n16_adj_3316), 
            .I3(\data_out_frame[13] [5]), .O(n41479));
    defparam i9_4_lut_adj_1194.LUT_INIT = 16'h6996;
    SB_LUT4 mux_923_i5_3_lut_4_lut (.I0(\FRAME_MATCHER.state [1]), .I1(n27693), 
            .I2(\data_in_frame[3] [4]), .I3(\data_in_frame[16] [4]), .O(n3796));
    defparam mux_923_i5_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i15_4_lut (.I0(n41479), .I1(n30_adj_3318), .I2(n40443), .I3(\data_out_frame[15] [7]), 
            .O(n34));
    defparam i15_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_1195 (.I0(n1498), .I1(n164), .I2(\FRAME_MATCHER.i [4]), 
            .I3(n22347), .O(n40205));
    defparam i2_3_lut_4_lut_adj_1195.LUT_INIT = 16'hff7f;
    SB_LUT4 i2_3_lut_4_lut_adj_1196 (.I0(n1498), .I1(n164), .I2(\FRAME_MATCHER.i [3]), 
            .I3(n9), .O(n40221));
    defparam i2_3_lut_4_lut_adj_1196.LUT_INIT = 16'hff7f;
    SB_LUT4 mux_923_i6_3_lut_4_lut (.I0(\FRAME_MATCHER.state [1]), .I1(n27693), 
            .I2(\data_in_frame[3] [5]), .I3(\data_in_frame[16] [5]), .O(n3797));
    defparam mux_923_i6_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i13_4_lut_adj_1197 (.I0(\data_out_frame[13] [5]), .I1(n40415), 
            .I2(n1695), .I3(n40471), .O(n32_adj_3319));
    defparam i13_4_lut_adj_1197.LUT_INIT = 16'h9669;
    SB_LUT4 i14_4_lut (.I0(n22051), .I1(n1716), .I2(n40711), .I3(n22840), 
            .O(n33));
    defparam i14_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 mux_923_i7_3_lut_4_lut (.I0(\FRAME_MATCHER.state [1]), .I1(n27693), 
            .I2(\data_in_frame[3] [6]), .I3(\data_in_frame[16] [6]), .O(n3798));
    defparam mux_923_i7_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i12_4_lut_adj_1198 (.I0(\data_out_frame[15] [5]), .I1(\data_out_frame[15] [6]), 
            .I2(n40423), .I3(\data_out_frame[15] [0]), .O(n31_adj_3320));
    defparam i12_4_lut_adj_1198.LUT_INIT = 16'h6996;
    SB_LUT4 i18_4_lut_adj_1199 (.I0(n31_adj_3320), .I1(n33), .I2(n32_adj_3319), 
            .I3(n34), .O(n40825));
    defparam i18_4_lut_adj_1199.LUT_INIT = 16'h6996;
    SB_LUT4 mux_923_i8_3_lut_4_lut (.I0(\FRAME_MATCHER.state [1]), .I1(n27693), 
            .I2(\data_in_frame[3] [7]), .I3(\data_in_frame[16] [7]), .O(n3799));
    defparam mux_923_i8_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i2_3_lut_adj_1200 (.I0(n40415), .I1(\data_out_frame[17] [0]), 
            .I2(\data_out_frame[16] [6]), .I3(GND_net), .O(n40490));
    defparam i2_3_lut_adj_1200.LUT_INIT = 16'h6969;
    SB_LUT4 mux_923_i9_3_lut_4_lut (.I0(\FRAME_MATCHER.state [1]), .I1(n27693), 
            .I2(\data_in_frame[2] [0]), .I3(\data_in_frame[15] [0]), .O(n3800));
    defparam mux_923_i9_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1_2_lut_adj_1201 (.I0(\data_out_frame[16] [3]), .I1(\data_out_frame[16] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n40717));
    defparam i1_2_lut_adj_1201.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1202 (.I0(n40490), .I1(n40825), .I2(GND_net), 
            .I3(GND_net), .O(n6_adj_3321));
    defparam i1_2_lut_adj_1202.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1203 (.I0(n40717), .I1(\data_out_frame[16] [4]), 
            .I2(n23383), .I3(n6_adj_3321), .O(n37264));
    defparam i4_4_lut_adj_1203.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1204 (.I0(\data_out_frame[17] [1]), .I1(\data_out_frame[17] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n22729));   // verilog/coms.v(76[16:27])
    defparam i1_2_lut_adj_1204.LUT_INIT = 16'h6666;
    SB_LUT4 mux_923_i10_3_lut_4_lut (.I0(\FRAME_MATCHER.state [1]), .I1(n27693), 
            .I2(\data_in_frame[2] [1]), .I3(\data_in_frame[15] [1]), .O(n3801));
    defparam mux_923_i10_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1_2_lut_adj_1205 (.I0(\data_out_frame[8] [3]), .I1(\data_out_frame[8] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n40343));
    defparam i1_2_lut_adj_1205.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_4_lut_adj_1206 (.I0(n1498), .I1(n164), .I2(\FRAME_MATCHER.i [3]), 
            .I3(n9), .O(n40212));
    defparam i2_3_lut_4_lut_adj_1206.LUT_INIT = 16'hfff7;
    SB_LUT4 i1_2_lut_adj_1207 (.I0(\data_out_frame[6] [1]), .I1(n40298), 
            .I2(GND_net), .I3(GND_net), .O(n40767));
    defparam i1_2_lut_adj_1207.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1208 (.I0(\data_out_frame[13] [1]), .I1(\data_out_frame[13] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n22511));   // verilog/coms.v(71[16:42])
    defparam i1_2_lut_adj_1208.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_1209 (.I0(\data_out_frame[12] [7]), .I1(n40634), 
            .I2(n40249), .I3(\data_out_frame[11] [0]), .O(n1595));   // verilog/coms.v(72[16:27])
    defparam i3_4_lut_adj_1209.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1210 (.I0(\data_out_frame[15] [3]), .I1(n1506), 
            .I2(n1595), .I3(n22511), .O(n40311));   // verilog/coms.v(71[16:42])
    defparam i3_4_lut_adj_1210.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1211 (.I0(n37264), .I1(n40576), .I2(GND_net), 
            .I3(GND_net), .O(n40577));
    defparam i1_2_lut_adj_1211.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1212 (.I0(n37222), .I1(n37264), .I2(GND_net), 
            .I3(GND_net), .O(n40749));
    defparam i1_2_lut_adj_1212.LUT_INIT = 16'h9999;
    SB_LUT4 i4_4_lut_adj_1213 (.I0(n40684), .I1(\data_out_frame[17] [4]), 
            .I2(\data_out_frame[19] [7]), .I3(n40749), .O(n10_adj_3302));
    defparam i4_4_lut_adj_1213.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1214 (.I0(\data_out_frame[8] [4]), .I1(\data_out_frame[10] [6]), 
            .I2(\data_out_frame[6] [2]), .I3(GND_net), .O(n40861));   // verilog/coms.v(72[16:27])
    defparam i2_3_lut_adj_1214.LUT_INIT = 16'h9696;
    SB_LUT4 i4_4_lut_adj_1215 (.I0(n23004), .I1(\data_out_frame[11] [1]), 
            .I2(\data_out_frame[9] [0]), .I3(n6_adj_3297), .O(n1506));   // verilog/coms.v(72[16:27])
    defparam i4_4_lut_adj_1215.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1216 (.I0(\data_out_frame[17] [7]), .I1(\data_out_frame[17] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n23218));
    defparam i1_2_lut_adj_1216.LUT_INIT = 16'h6666;
    SB_LUT4 i7_4_lut_adj_1217 (.I0(n40548), .I1(n40292), .I2(\data_out_frame[15] [4]), 
            .I3(\data_out_frame[13] [5]), .O(n18_adj_3322));   // verilog/coms.v(72[16:27])
    defparam i7_4_lut_adj_1217.LUT_INIT = 16'h6996;
    SB_LUT4 mux_923_i11_3_lut_4_lut (.I0(\FRAME_MATCHER.state [1]), .I1(n27693), 
            .I2(\data_in_frame[2] [2]), .I3(\data_in_frame[15] [2]), .O(n3802));
    defparam mux_923_i11_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i5_2_lut_adj_1218 (.I0(\data_out_frame[5] [1]), .I1(n1506), 
            .I2(GND_net), .I3(GND_net), .O(n16_adj_3323));   // verilog/coms.v(72[16:27])
    defparam i5_2_lut_adj_1218.LUT_INIT = 16'h6666;
    SB_LUT4 i9_4_lut_adj_1219 (.I0(n23218), .I1(n18_adj_3322), .I2(\data_out_frame[18] [0]), 
            .I3(\data_out_frame[13] [2]), .O(n20_adj_3324));   // verilog/coms.v(72[16:27])
    defparam i9_4_lut_adj_1219.LUT_INIT = 16'h6996;
    SB_LUT4 equal_59_i8_2_lut_3_lut (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(\FRAME_MATCHER.i [0]), .I3(GND_net), .O(n8_adj_3123));   // verilog/coms.v(154[7:23])
    defparam equal_59_i8_2_lut_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i10_4_lut_adj_1220 (.I0(n40740), .I1(n20_adj_3324), .I2(n16_adj_3323), 
            .I3(n40521), .O(n40684));   // verilog/coms.v(72[16:27])
    defparam i10_4_lut_adj_1220.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1221 (.I0(n22051), .I1(n40684), .I2(GND_net), 
            .I3(GND_net), .O(n40588));
    defparam i1_2_lut_adj_1221.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1222 (.I0(\data_out_frame[18] [1]), .I1(n37222), 
            .I2(n37253), .I3(n6_adj_3325), .O(n37246));
    defparam i4_4_lut_adj_1222.LUT_INIT = 16'h9669;
    SB_LUT4 mux_923_i12_3_lut_4_lut (.I0(\FRAME_MATCHER.state [1]), .I1(n27693), 
            .I2(\data_in_frame[2] [3]), .I3(\data_in_frame[15] [3]), .O(n3803));
    defparam mux_923_i12_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1_2_lut_adj_1223 (.I0(\data_out_frame[18] [1]), .I1(n40816), 
            .I2(GND_net), .I3(GND_net), .O(n40368));
    defparam i1_2_lut_adj_1223.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1224 (.I0(\data_out_frame[8] [6]), .I1(\data_out_frame[8] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n40249));   // verilog/coms.v(72[16:27])
    defparam i1_2_lut_adj_1224.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1225 (.I0(\data_out_frame[10] [7]), .I1(\data_out_frame[11] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n4_adj_3326));
    defparam i1_2_lut_adj_1225.LUT_INIT = 16'h6666;
    SB_LUT4 i2_4_lut_adj_1226 (.I0(\data_out_frame[9] [1]), .I1(\data_out_frame[6] [3]), 
            .I2(\data_out_frame[11] [1]), .I3(n4_adj_3326), .O(n40386));   // verilog/coms.v(73[16:27])
    defparam i2_4_lut_adj_1226.LUT_INIT = 16'h6996;
    SB_LUT4 mux_923_i13_3_lut_4_lut (.I0(\FRAME_MATCHER.state [1]), .I1(n27693), 
            .I2(\data_in_frame[2] [4]), .I3(\data_in_frame[15] [4]), .O(n3804));
    defparam mux_923_i13_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i3_4_lut_adj_1227 (.I0(\data_out_frame[13] [3]), .I1(n40386), 
            .I2(n23323), .I3(n23004), .O(n22515));   // verilog/coms.v(73[16:27])
    defparam i3_4_lut_adj_1227.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1228 (.I0(\data_out_frame[13] [4]), .I1(n22515), 
            .I2(GND_net), .I3(GND_net), .O(n40548));
    defparam i1_2_lut_adj_1228.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_1229 (.I0(\data_out_frame[17] [7]), .I1(\data_out_frame[15] [5]), 
            .I2(n40548), .I3(n41642), .O(n37222));
    defparam i3_4_lut_adj_1229.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1230 (.I0(\data_out_frame[20] [3]), .I1(n37222), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_3327));
    defparam i1_2_lut_adj_1230.LUT_INIT = 16'h6666;
    SB_LUT4 mux_923_i14_3_lut_4_lut (.I0(\FRAME_MATCHER.state [1]), .I1(n27693), 
            .I2(\data_in_frame[2] [5]), .I3(\data_in_frame[15] [5]), .O(n3805));
    defparam mux_923_i14_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4_4_lut_adj_1231 (.I0(\data_out_frame[16] [1]), .I1(n40381), 
            .I2(n40368), .I3(n6_adj_3327), .O(n36588));
    defparam i4_4_lut_adj_1231.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_adj_1232 (.I0(n36588), .I1(n40456), .I2(GND_net), 
            .I3(GND_net), .O(n40703));
    defparam i1_2_lut_adj_1232.LUT_INIT = 16'h6666;
    SB_LUT4 mux_923_i15_3_lut_4_lut (.I0(\FRAME_MATCHER.state [1]), .I1(n27693), 
            .I2(\data_in_frame[2] [6]), .I3(\data_in_frame[15] [6]), .O(n3806));
    defparam mux_923_i15_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1_2_lut_adj_1233 (.I0(\data_out_frame[7] [3]), .I1(\data_out_frame[13] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n40852));   // verilog/coms.v(71[16:27])
    defparam i1_2_lut_adj_1233.LUT_INIT = 16'h6666;
    SB_LUT4 mux_923_i16_3_lut_4_lut (.I0(\FRAME_MATCHER.state [1]), .I1(n27693), 
            .I2(\data_in_frame[2] [7]), .I3(\data_in_frame[15] [7]), .O(n3807));
    defparam mux_923_i16_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1_2_lut_adj_1234 (.I0(\data_out_frame[7] [2]), .I1(\data_out_frame[15] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n40740));   // verilog/coms.v(72[16:27])
    defparam i1_2_lut_adj_1234.LUT_INIT = 16'h6666;
    SB_LUT4 mux_923_i17_3_lut_4_lut (.I0(\FRAME_MATCHER.state [1]), .I1(n27693), 
            .I2(\data_in_frame[1] [0]), .I3(\data_in_frame[14] [0]), .O(n3808));
    defparam mux_923_i17_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i2_3_lut_adj_1235 (.I0(\data_out_frame[11] [2]), .I1(\data_out_frame[8] [6]), 
            .I2(\data_out_frame[6] [4]), .I3(GND_net), .O(n40870));   // verilog/coms.v(71[16:27])
    defparam i2_3_lut_adj_1235.LUT_INIT = 16'h9696;
    SB_LUT4 i7_4_lut_adj_1236 (.I0(\data_out_frame[15] [7]), .I1(n40870), 
            .I2(n40803), .I3(n40622), .O(n18_adj_3328));   // verilog/coms.v(71[16:27])
    defparam i7_4_lut_adj_1236.LUT_INIT = 16'h6996;
    SB_LUT4 i9_4_lut_adj_1237 (.I0(n36529), .I1(n18_adj_3328), .I2(n37253), 
            .I3(\data_out_frame[18] [2]), .O(n20_adj_3329));   // verilog/coms.v(71[16:27])
    defparam i9_4_lut_adj_1237.LUT_INIT = 16'h6996;
    SB_LUT4 mux_923_i18_3_lut_4_lut (.I0(\FRAME_MATCHER.state [1]), .I1(n27693), 
            .I2(\data_in_frame[1] [1]), .I3(\data_in_frame[14] [1]), .O(n3809));
    defparam mux_923_i18_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i10_4_lut_adj_1238 (.I0(n23166), .I1(n20_adj_3329), .I2(n16_adj_3330), 
            .I3(n40852), .O(n40816));   // verilog/coms.v(71[16:27])
    defparam i10_4_lut_adj_1238.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1239 (.I0(\data_out_frame[16] [1]), .I1(\data_out_frame[16] [2]), 
            .I2(\data_out_frame[16] [0]), .I3(GND_net), .O(n40443));
    defparam i2_3_lut_adj_1239.LUT_INIT = 16'h9696;
    SB_LUT4 mux_923_i19_3_lut_4_lut (.I0(\FRAME_MATCHER.state [1]), .I1(n27693), 
            .I2(\data_in_frame[1] [2]), .I3(\data_in_frame[14] [2]), .O(n3810));
    defparam mux_923_i19_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1_2_lut_adj_1240 (.I0(\data_out_frame[20] [4]), .I1(n22051), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_3331));
    defparam i1_2_lut_adj_1240.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1241 (.I0(n40696), .I1(n40443), .I2(n40816), 
            .I3(n6_adj_3331), .O(n40456));
    defparam i4_4_lut_adj_1241.LUT_INIT = 16'h6996;
    SB_LUT4 mux_923_i20_3_lut_4_lut (.I0(\FRAME_MATCHER.state [1]), .I1(n27693), 
            .I2(\data_in_frame[1] [3]), .I3(\data_in_frame[14] [3]), .O(n3811));
    defparam mux_923_i20_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i2_3_lut_adj_1242 (.I0(n37308), .I1(n40456), .I2(\data_out_frame[20] [5]), 
            .I3(GND_net), .O(n41743));
    defparam i2_3_lut_adj_1242.LUT_INIT = 16'h9696;
    SB_LUT4 mux_923_i21_3_lut_4_lut (.I0(\FRAME_MATCHER.state [1]), .I1(n27693), 
            .I2(\data_in_frame[1] [4]), .I3(\data_in_frame[14] [4]), .O(n3812));
    defparam mux_923_i21_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 mux_923_i22_3_lut_4_lut (.I0(\FRAME_MATCHER.state [1]), .I1(n27693), 
            .I2(\data_in_frame[1] [5]), .I3(\data_in_frame[14] [5]), .O(n3813));
    defparam mux_923_i22_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 mux_923_i24_3_lut_4_lut (.I0(\FRAME_MATCHER.state [1]), .I1(n27693), 
            .I2(\data_in_frame[1] [7]), .I3(\data_in_frame[14] [7]), .O(n3815));
    defparam mux_923_i24_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1_2_lut_adj_1243 (.I0(\data_out_frame[12] [1]), .I1(\data_out_frame[12] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n23029));
    defparam i1_2_lut_adj_1243.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_1244 (.I0(\data_out_frame[7] [3]), .I1(\data_out_frame[9] [5]), 
            .I2(\data_out_frame[10] [1]), .I3(\data_out_frame[11] [7]), 
            .O(n40518));   // verilog/coms.v(71[16:27])
    defparam i3_4_lut_adj_1244.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1245 (.I0(\data_out_frame[5] [4]), .I1(\data_out_frame[5][2] ), 
            .I2(GND_net), .I3(GND_net), .O(n22630));   // verilog/coms.v(72[16:27])
    defparam i1_2_lut_adj_1245.LUT_INIT = 16'h6666;
    SB_LUT4 mux_923_i23_3_lut_4_lut (.I0(\FRAME_MATCHER.state [1]), .I1(n27693), 
            .I2(\data_in_frame[1] [6]), .I3(\data_in_frame[14] [6]), .O(n3814));
    defparam mux_923_i23_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1246 (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(n40205), .I3(\FRAME_MATCHER.i [0]), .O(n40209));   // verilog/coms.v(154[7:23])
    defparam i1_2_lut_3_lut_4_lut_adj_1246.LUT_INIT = 16'hfeff;
    SB_LUT4 i5_3_lut_adj_1247 (.I0(\data_out_frame[12] [2]), .I1(\data_out_frame[12] [1]), 
            .I2(n22635), .I3(GND_net), .O(n14_adj_3332));   // verilog/coms.v(71[16:27])
    defparam i5_3_lut_adj_1247.LUT_INIT = 16'h9696;
    SB_LUT4 i6_4_lut_adj_1248 (.I0(n40723), .I1(\data_out_frame[14] [3]), 
            .I2(n22630), .I3(n40518), .O(n15_adj_3333));   // verilog/coms.v(71[16:27])
    defparam i6_4_lut_adj_1248.LUT_INIT = 16'h6996;
    SB_LUT4 i8_4_lut_adj_1249 (.I0(n15_adj_3333), .I1(\data_out_frame[5] [1]), 
            .I2(n14_adj_3332), .I3(\data_out_frame[9] [6]), .O(n23383));   // verilog/coms.v(71[16:27])
    defparam i8_4_lut_adj_1249.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1250 (.I0(n23383), .I1(n40440), .I2(GND_net), 
            .I3(GND_net), .O(n1716));
    defparam i1_2_lut_adj_1250.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1251 (.I0(\data_out_frame[14] [0]), .I1(n23169), 
            .I2(GND_net), .I3(GND_net), .O(n40471));
    defparam i1_2_lut_adj_1251.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1252 (.I0(\data_out_frame[18] [5]), .I1(\data_out_frame[18] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n40714));
    defparam i1_2_lut_adj_1252.LUT_INIT = 16'h6666;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_31382 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[18] [4]), .I2(\data_out_frame[19] [4]), 
            .I3(byte_transmit_counter[1]), .O(n46895));
    defparam byte_transmit_counter_0__bdd_4_lut_31382.LUT_INIT = 16'he4aa;
    SB_LUT4 i1_2_lut_adj_1253 (.I0(\data_out_frame[6] [7]), .I1(\data_out_frame[6] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n40282));   // verilog/coms.v(71[16:27])
    defparam i1_2_lut_adj_1253.LUT_INIT = 16'h6666;
    SB_LUT4 i908_2_lut (.I0(\data_out_frame[13] [7]), .I1(\data_out_frame[13] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n1664));   // verilog/coms.v(83[17:28])
    defparam i908_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1254 (.I0(\data_out_frame[11] [6]), .I1(\data_out_frame[9] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n40681));   // verilog/coms.v(71[16:27])
    defparam i1_2_lut_adj_1254.LUT_INIT = 16'h6666;
    SB_LUT4 i5_3_lut_4_lut_adj_1255 (.I0(\data_out_frame[7] [5]), .I1(n22635), 
            .I2(\data_out_frame[5] [3]), .I3(n10_adj_3305), .O(n40551));   // verilog/coms.v(73[16:27])
    defparam i5_3_lut_4_lut_adj_1255.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_1256 (.I0(n40681), .I1(n40295), .I2(\data_out_frame[9] [3]), 
            .I3(n40803), .O(n10_adj_3285));   // verilog/coms.v(71[16:27])
    defparam i4_4_lut_adj_1256.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1257 (.I0(\data_out_frame[11] [3]), .I1(\data_out_frame[8] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n23166));
    defparam i1_2_lut_adj_1257.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_1258 (.I0(\data_out_frame[11] [4]), .I1(\data_out_frame[9] [3]), 
            .I2(\data_out_frame[9] [1]), .I3(\data_out_frame[6] [5]), .O(n40521));   // verilog/coms.v(69[16:27])
    defparam i3_4_lut_adj_1258.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1259 (.I0(\data_out_frame[5] [1]), .I1(\data_out_frame[7] [1]), 
            .I2(\data_out_frame[6] [7]), .I3(GND_net), .O(n40499));
    defparam i2_3_lut_adj_1259.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1260 (.I0(\data_out_frame[7] [0]), .I1(\data_out_frame[6] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n23323));   // verilog/coms.v(69[16:27])
    defparam i1_2_lut_adj_1260.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1261 (.I0(n23323), .I1(n40499), .I2(n40521), 
            .I3(n6_adj_3334), .O(n1515));
    defparam i4_4_lut_adj_1261.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1262 (.I0(n36529), .I1(\data_out_frame[13] [5]), 
            .I2(n1515), .I3(GND_net), .O(n40711));
    defparam i2_3_lut_adj_1262.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1263 (.I0(\data_out_frame[14] [0]), .I1(n40380), 
            .I2(GND_net), .I3(GND_net), .O(n40381));
    defparam i1_2_lut_adj_1263.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1264 (.I0(\data_out_frame[7] [4]), .I1(\data_out_frame[5] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n40401));   // verilog/coms.v(72[16:27])
    defparam i1_2_lut_adj_1264.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1265 (.I0(\data_out_frame[5] [5]), .I1(\data_out_frame[7] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n40764));   // verilog/coms.v(72[16:27])
    defparam i1_2_lut_adj_1265.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1266 (.I0(n40625), .I1(\data_out_frame[5][2] ), 
            .I2(\data_out_frame[10] [0]), .I3(n40764), .O(n10_adj_3335));   // verilog/coms.v(72[16:27])
    defparam i4_4_lut_adj_1266.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1267 (.I0(\data_out_frame[5] [1]), .I1(\data_out_frame[5] [0]), 
            .I2(\data_out_frame[5] [3]), .I3(GND_net), .O(n40604));   // verilog/coms.v(71[16:27])
    defparam i2_3_lut_adj_1267.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1268 (.I0(\data_out_frame[5][2] ), .I1(\data_out_frame[9] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n40806));
    defparam i1_2_lut_adj_1268.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_1269 (.I0(\data_out_frame[11] [5]), .I1(\data_out_frame[9] [3]), 
            .I2(\data_out_frame[5] [0]), .I3(GND_net), .O(n40720));
    defparam i2_3_lut_adj_1269.LUT_INIT = 16'h9696;
    SB_LUT4 i3_4_lut_adj_1270 (.I0(\data_out_frame[6] [7]), .I1(n40720), 
            .I2(\data_out_frame[5] [3]), .I3(\data_out_frame[9] [5]), .O(n40289));   // verilog/coms.v(71[16:27])
    defparam i3_4_lut_adj_1270.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1271 (.I0(\data_out_frame[5] [4]), .I1(\data_out_frame[9] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n40625));   // verilog/coms.v(71[16:27])
    defparam i1_2_lut_adj_1271.LUT_INIT = 16'h6666;
    SB_LUT4 i5_3_lut_adj_1272 (.I0(\data_out_frame[13] [7]), .I1(\data_out_frame[9] [4]), 
            .I2(\data_out_frame[7] [1]), .I3(GND_net), .O(n14_adj_3336));   // verilog/coms.v(71[16:27])
    defparam i5_3_lut_adj_1272.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1273 (.I0(n22047), .I1(n40656), .I2(n40551), 
            .I3(GND_net), .O(n22134));
    defparam i1_2_lut_3_lut_adj_1273.LUT_INIT = 16'h9696;
    SB_LUT4 i6_4_lut_adj_1274 (.I0(n40625), .I1(\data_out_frame[14] [1]), 
            .I2(\data_out_frame[11] [7]), .I3(n40289), .O(n15_adj_3337));   // verilog/coms.v(71[16:27])
    defparam i6_4_lut_adj_1274.LUT_INIT = 16'h6996;
    SB_LUT4 i8_4_lut_adj_1275 (.I0(n15_adj_3337), .I1(\data_out_frame[7] [5]), 
            .I2(n14_adj_3336), .I3(\data_out_frame[12] [0]), .O(n23169));   // verilog/coms.v(71[16:27])
    defparam i8_4_lut_adj_1275.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1276 (.I0(\data_out_frame[11] [5]), .I1(n40628), 
            .I2(n40295), .I3(\data_out_frame[6] [6]), .O(n22051));
    defparam i3_4_lut_adj_1276.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1277 (.I0(\data_out_frame[16] [3]), .I1(\data_out_frame[18] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n40279));
    defparam i1_2_lut_adj_1277.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_3_lut_adj_1278 (.I0(n22047), .I1(n40656), .I2(n40873), 
            .I3(GND_net), .O(n22840));
    defparam i1_2_lut_3_lut_adj_1278.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1279 (.I0(n22051), .I1(n23169), .I2(GND_net), 
            .I3(GND_net), .O(n4_adj_3338));
    defparam i1_2_lut_adj_1279.LUT_INIT = 16'h6666;
    SB_LUT4 i2_4_lut_adj_1280 (.I0(\data_out_frame[16] [1]), .I1(n40381), 
            .I2(n4_adj_3338), .I3(\data_out_frame[18][3] ), .O(n40696));
    defparam i2_4_lut_adj_1280.LUT_INIT = 16'h9669;
    SB_LUT4 select_267_Select_0_i3_2_lut_3_lut (.I0(n1498), .I1(n19_adj_3206), 
            .I2(\FRAME_MATCHER.i [0]), .I3(GND_net), .O(n3_adj_3217));
    defparam select_267_Select_0_i3_2_lut_3_lut.LUT_INIT = 16'h4040;
    SB_LUT4 i4_4_lut_adj_1281 (.I0(n40604), .I1(n40806), .I2(n23000), 
            .I3(\data_out_frame[7] [4]), .O(n10_adj_3339));
    defparam i4_4_lut_adj_1281.LUT_INIT = 16'h6996;
    SB_LUT4 select_267_Select_1_i3_2_lut_3_lut (.I0(n1498), .I1(n19_adj_3206), 
            .I2(\FRAME_MATCHER.i [1]), .I3(GND_net), .O(n3_adj_3200));
    defparam select_267_Select_1_i3_2_lut_3_lut.LUT_INIT = 16'h4040;
    SB_LUT4 select_267_Select_2_i3_2_lut_3_lut (.I0(n1498), .I1(n19_adj_3206), 
            .I2(\FRAME_MATCHER.i [2]), .I3(GND_net), .O(n3_adj_3199));
    defparam select_267_Select_2_i3_2_lut_3_lut.LUT_INIT = 16'h4040;
    SB_LUT4 i2_4_lut_adj_1282 (.I0(\data_out_frame[14] [2]), .I1(n23029), 
            .I2(n9_adj_3340), .I3(n10_adj_3339), .O(n40440));
    defparam i2_4_lut_adj_1282.LUT_INIT = 16'h6996;
    SB_LUT4 select_267_Select_3_i3_2_lut_3_lut (.I0(n1498), .I1(n19_adj_3206), 
            .I2(\FRAME_MATCHER.i [3]), .I3(GND_net), .O(n3_adj_3198));
    defparam select_267_Select_3_i3_2_lut_3_lut.LUT_INIT = 16'h4040;
    SB_LUT4 i3_4_lut_adj_1283 (.I0(n40411), .I1(n40822), .I2(n40714), 
            .I3(n40471), .O(n22071));
    defparam i3_4_lut_adj_1283.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1284 (.I0(\data_out_frame[20] [6]), .I1(\data_out_frame[20] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n40453));
    defparam i1_2_lut_adj_1284.LUT_INIT = 16'h6666;
    SB_LUT4 select_267_Select_4_i3_2_lut_3_lut (.I0(n1498), .I1(n19_adj_3206), 
            .I2(\FRAME_MATCHER.i [4]), .I3(GND_net), .O(n3_adj_3197));
    defparam select_267_Select_4_i3_2_lut_3_lut.LUT_INIT = 16'h4040;
    SB_LUT4 select_267_Select_5_i3_2_lut_3_lut (.I0(n1498), .I1(n19_adj_3206), 
            .I2(\FRAME_MATCHER.i [5]), .I3(GND_net), .O(n3_adj_3196));
    defparam select_267_Select_5_i3_2_lut_3_lut.LUT_INIT = 16'h4040;
    SB_LUT4 select_267_Select_6_i3_2_lut_3_lut (.I0(n1498), .I1(n19_adj_3206), 
            .I2(\FRAME_MATCHER.i [6]), .I3(GND_net), .O(n3_adj_3195));
    defparam select_267_Select_6_i3_2_lut_3_lut.LUT_INIT = 16'h4040;
    SB_LUT4 i30694_2_lut (.I0(n5021), .I1(n5019), .I2(GND_net), .I3(GND_net), 
            .O(n23452));
    defparam i30694_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 select_267_Select_7_i3_2_lut_3_lut (.I0(n1498), .I1(n19_adj_3206), 
            .I2(\FRAME_MATCHER.i [7]), .I3(GND_net), .O(n3_adj_3193));
    defparam select_267_Select_7_i3_2_lut_3_lut.LUT_INIT = 16'h4040;
    SB_LUT4 select_267_Select_8_i3_2_lut_3_lut (.I0(n1498), .I1(n19_adj_3206), 
            .I2(\FRAME_MATCHER.i [8]), .I3(GND_net), .O(n3_adj_3191));
    defparam select_267_Select_8_i3_2_lut_3_lut.LUT_INIT = 16'h4040;
    SB_LUT4 select_267_Select_9_i3_2_lut_3_lut (.I0(n1498), .I1(n19_adj_3206), 
            .I2(\FRAME_MATCHER.i [9]), .I3(GND_net), .O(n3_adj_3189));
    defparam select_267_Select_9_i3_2_lut_3_lut.LUT_INIT = 16'h4040;
    SB_LUT4 select_267_Select_10_i3_2_lut_3_lut (.I0(n1498), .I1(n19_adj_3206), 
            .I2(\FRAME_MATCHER.i [10]), .I3(GND_net), .O(n3_adj_3188));
    defparam select_267_Select_10_i3_2_lut_3_lut.LUT_INIT = 16'h4040;
    SB_LUT4 i1_2_lut_adj_1285 (.I0(\FRAME_MATCHER.i_31__N_1824 ), .I1(n736), 
            .I2(GND_net), .I3(GND_net), .O(n15_adj_3251));
    defparam i1_2_lut_adj_1285.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_1286 (.I0(\FRAME_MATCHER.i_31__N_1827 ), .I1(n3761), 
            .I2(GND_net), .I3(GND_net), .O(n40163));
    defparam i1_2_lut_adj_1286.LUT_INIT = 16'h2222;
    SB_LUT4 select_302_Select_1_i5_4_lut (.I0(n63), .I1(\FRAME_MATCHER.i_31__N_1825 ), 
            .I2(n2857), .I3(n7[1]), .O(n5_adj_3341));
    defparam select_302_Select_1_i5_4_lut.LUT_INIT = 16'hccc4;
    SB_LUT4 select_302_Select_1_i1_4_lut (.I0(n740), .I1(\FRAME_MATCHER.i_31__N_1821 ), 
            .I2(n7[1]), .I3(n63), .O(n1_adj_3342));
    defparam select_302_Select_1_i1_4_lut.LUT_INIT = 16'hc8cc;
    SB_LUT4 select_267_Select_11_i3_2_lut_3_lut (.I0(n1498), .I1(n19_adj_3206), 
            .I2(\FRAME_MATCHER.i [11]), .I3(GND_net), .O(n3_adj_3187));
    defparam select_267_Select_11_i3_2_lut_3_lut.LUT_INIT = 16'h4040;
    SB_LUT4 select_267_Select_12_i3_2_lut_3_lut (.I0(n1498), .I1(n19_adj_3206), 
            .I2(\FRAME_MATCHER.i [12]), .I3(GND_net), .O(n3_adj_3186));
    defparam select_267_Select_12_i3_2_lut_3_lut.LUT_INIT = 16'h4040;
    SB_LUT4 i3_4_lut_adj_1287 (.I0(\FRAME_MATCHER.i_31__N_1823 ), .I1(n36044), 
            .I2(n1_adj_3342), .I3(n5_adj_3341), .O(n47026));
    defparam i3_4_lut_adj_1287.LUT_INIT = 16'hfffe;
    SB_LUT4 select_267_Select_13_i3_2_lut_3_lut (.I0(n1498), .I1(n19_adj_3206), 
            .I2(\FRAME_MATCHER.i [13]), .I3(GND_net), .O(n3_adj_3185));
    defparam select_267_Select_13_i3_2_lut_3_lut.LUT_INIT = 16'h4040;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1288 (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(n40221), .I3(\FRAME_MATCHER.i [0]), .O(n40222));   // verilog/coms.v(154[7:23])
    defparam i1_2_lut_3_lut_4_lut_adj_1288.LUT_INIT = 16'hfeff;
    SB_LUT4 select_267_Select_14_i3_2_lut_3_lut (.I0(n1498), .I1(n19_adj_3206), 
            .I2(\FRAME_MATCHER.i [14]), .I3(GND_net), .O(n3_adj_3184));
    defparam select_267_Select_14_i3_2_lut_3_lut.LUT_INIT = 16'h4040;
    SB_LUT4 select_267_Select_15_i3_2_lut_3_lut (.I0(n1498), .I1(n19_adj_3206), 
            .I2(\FRAME_MATCHER.i [15]), .I3(GND_net), .O(n3_adj_3183));
    defparam select_267_Select_15_i3_2_lut_3_lut.LUT_INIT = 16'h4040;
    SB_LUT4 select_267_Select_16_i3_2_lut_3_lut (.I0(n1498), .I1(n19_adj_3206), 
            .I2(\FRAME_MATCHER.i [16]), .I3(GND_net), .O(n3_adj_3182));
    defparam select_267_Select_16_i3_2_lut_3_lut.LUT_INIT = 16'h4040;
    SB_LUT4 i3_3_lut (.I0(\FRAME_MATCHER.state [0]), .I1(\FRAME_MATCHER.state [1]), 
            .I2(n1_c), .I3(GND_net), .O(n8_adj_3343));
    defparam i3_3_lut.LUT_INIT = 16'h0404;
    SB_LUT4 select_267_Select_17_i3_2_lut_3_lut (.I0(n1498), .I1(n19_adj_3206), 
            .I2(\FRAME_MATCHER.i [17]), .I3(GND_net), .O(n3_adj_3181));
    defparam select_267_Select_17_i3_2_lut_3_lut.LUT_INIT = 16'h4040;
    SB_LUT4 i29304_3_lut (.I0(n43), .I1(n2_adj_3220), .I2(n47), .I3(GND_net), 
            .O(n44171));
    defparam i29304_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 select_267_Select_18_i3_2_lut_3_lut (.I0(n1498), .I1(n19_adj_3206), 
            .I2(\FRAME_MATCHER.i [18]), .I3(GND_net), .O(n3_adj_3180));
    defparam select_267_Select_18_i3_2_lut_3_lut.LUT_INIT = 16'h4040;
    SB_LUT4 i29340_2_lut (.I0(\FRAME_MATCHER.state_31__N_1925 [3]), .I1(\FRAME_MATCHER.state [2]), 
            .I2(GND_net), .I3(GND_net), .O(n44173));
    defparam i29340_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 select_267_Select_19_i3_2_lut_3_lut (.I0(n1498), .I1(n19_adj_3206), 
            .I2(\FRAME_MATCHER.i [19]), .I3(GND_net), .O(n3_adj_3178));
    defparam select_267_Select_19_i3_2_lut_3_lut.LUT_INIT = 16'h4040;
    SB_LUT4 i24_4_lut_adj_1289 (.I0(n44173), .I1(n44171), .I2(\FRAME_MATCHER.state [3]), 
            .I3(n8_adj_3343), .O(n39742));
    defparam i24_4_lut_adj_1289.LUT_INIT = 16'hcac0;
    SB_LUT4 select_267_Select_20_i3_2_lut_3_lut (.I0(n1498), .I1(n19_adj_3206), 
            .I2(\FRAME_MATCHER.i [20]), .I3(GND_net), .O(n3_adj_3176));
    defparam select_267_Select_20_i3_2_lut_3_lut.LUT_INIT = 16'h4040;
    SB_LUT4 i1_3_lut_adj_1290 (.I0(\FRAME_MATCHER.state [3]), .I1(n6_adj_3221), 
            .I2(n5_adj_3238), .I3(GND_net), .O(n39506));
    defparam i1_3_lut_adj_1290.LUT_INIT = 16'ha8a8;
    SB_LUT4 select_267_Select_21_i3_2_lut_3_lut (.I0(n1498), .I1(n19_adj_3206), 
            .I2(\FRAME_MATCHER.i [21]), .I3(GND_net), .O(n3_adj_3174));
    defparam select_267_Select_21_i3_2_lut_3_lut.LUT_INIT = 16'h4040;
    SB_LUT4 i1_2_lut_adj_1291 (.I0(\FRAME_MATCHER.state [4]), .I1(n36224), 
            .I2(GND_net), .I3(GND_net), .O(n39406));
    defparam i1_2_lut_adj_1291.LUT_INIT = 16'h8888;
    SB_LUT4 select_267_Select_22_i3_2_lut_3_lut (.I0(n1498), .I1(n19_adj_3206), 
            .I2(\FRAME_MATCHER.i [22]), .I3(GND_net), .O(n3_adj_3172));
    defparam select_267_Select_22_i3_2_lut_3_lut.LUT_INIT = 16'h4040;
    SB_LUT4 i14752_2_lut (.I0(\FRAME_MATCHER.state [5]), .I1(n36224), .I2(GND_net), 
            .I3(GND_net), .O(n28157));
    defparam i14752_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 select_267_Select_23_i3_2_lut_3_lut (.I0(n1498), .I1(n19_adj_3206), 
            .I2(\FRAME_MATCHER.i [23]), .I3(GND_net), .O(n3_adj_3170));
    defparam select_267_Select_23_i3_2_lut_3_lut.LUT_INIT = 16'h4040;
    SB_LUT4 i14753_2_lut (.I0(\FRAME_MATCHER.state [6]), .I1(n36224), .I2(GND_net), 
            .I3(GND_net), .O(n28159));
    defparam i14753_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 select_267_Select_24_i3_2_lut_3_lut (.I0(n1498), .I1(n19_adj_3206), 
            .I2(\FRAME_MATCHER.i [24]), .I3(GND_net), .O(n3_adj_3168));
    defparam select_267_Select_24_i3_2_lut_3_lut.LUT_INIT = 16'h4040;
    SB_LUT4 i1_2_lut_adj_1292 (.I0(\FRAME_MATCHER.state [8]), .I1(n36224), 
            .I2(GND_net), .I3(GND_net), .O(n39402));
    defparam i1_2_lut_adj_1292.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1293 (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(n40212), .I3(\FRAME_MATCHER.i [0]), .O(n40213));   // verilog/coms.v(154[7:23])
    defparam i1_2_lut_3_lut_4_lut_adj_1293.LUT_INIT = 16'hfeff;
    SB_LUT4 select_267_Select_25_i3_2_lut_3_lut (.I0(n1498), .I1(n19_adj_3206), 
            .I2(\FRAME_MATCHER.i [25]), .I3(GND_net), .O(n3_adj_3166));
    defparam select_267_Select_25_i3_2_lut_3_lut.LUT_INIT = 16'h4040;
    SB_LUT4 i2_3_lut_adj_1294 (.I0(n10_adj_3344), .I1(\FRAME_MATCHER.i_31__N_1823 ), 
            .I2(n1498), .I3(GND_net), .O(n41992));
    defparam i2_3_lut_adj_1294.LUT_INIT = 16'hfefe;
    SB_LUT4 i2_4_lut_adj_1295 (.I0(n47), .I1(n2_adj_3220), .I2(n20075), 
            .I3(n41992), .O(n36224));
    defparam i2_4_lut_adj_1295.LUT_INIT = 16'heefe;
    SB_LUT4 select_267_Select_26_i3_2_lut_3_lut (.I0(n1498), .I1(n19_adj_3206), 
            .I2(\FRAME_MATCHER.i [26]), .I3(GND_net), .O(n3_adj_3164));
    defparam select_267_Select_26_i3_2_lut_3_lut.LUT_INIT = 16'h4040;
    SB_LUT4 i20490_2_lut (.I0(\FRAME_MATCHER.state [20]), .I1(n36224), .I2(GND_net), 
            .I3(GND_net), .O(n35999));
    defparam i20490_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 select_267_Select_27_i3_2_lut_3_lut (.I0(n1498), .I1(n19_adj_3206), 
            .I2(\FRAME_MATCHER.i [27]), .I3(GND_net), .O(n3_adj_3162));
    defparam select_267_Select_27_i3_2_lut_3_lut.LUT_INIT = 16'h4040;
    SB_LUT4 select_267_Select_28_i3_2_lut_3_lut (.I0(n1498), .I1(n19_adj_3206), 
            .I2(\FRAME_MATCHER.i [28]), .I3(GND_net), .O(n3_adj_3160));
    defparam select_267_Select_28_i3_2_lut_3_lut.LUT_INIT = 16'h4040;
    SB_LUT4 select_267_Select_29_i3_2_lut_3_lut (.I0(n1498), .I1(n19_adj_3206), 
            .I2(\FRAME_MATCHER.i [29]), .I3(GND_net), .O(n3_adj_3158));
    defparam select_267_Select_29_i3_2_lut_3_lut.LUT_INIT = 16'h4040;
    SB_LUT4 n46895_bdd_4_lut (.I0(n46895), .I1(\data_out_frame[17] [4]), 
            .I2(\data_out_frame[16] [4]), .I3(byte_transmit_counter[1]), 
            .O(n46898));
    defparam n46895_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_2_lut_adj_1296 (.I0(\FRAME_MATCHER.state [1]), .I1(\FRAME_MATCHER.state [0]), 
            .I2(GND_net), .I3(GND_net), .O(n105));
    defparam i1_2_lut_adj_1296.LUT_INIT = 16'heeee;
    SB_LUT4 i14440_4_lut (.I0(\FRAME_MATCHER.i [0]), .I1(\FRAME_MATCHER.i [31]), 
            .I2(n4_adj_3280), .I3(\FRAME_MATCHER.i [1]), .O(n740));   // verilog/coms.v(157[9:60])
    defparam i14440_4_lut.LUT_INIT = 16'h3230;
    SB_LUT4 i14441_2_lut (.I0(n22250), .I1(\FRAME_MATCHER.i [31]), .I2(GND_net), 
            .I3(GND_net), .O(n2857));   // verilog/coms.v(221[9:54])
    defparam i14441_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i1_3_lut_adj_1297 (.I0(\FRAME_MATCHER.state [1]), .I1(\FRAME_MATCHER.state [2]), 
            .I2(\FRAME_MATCHER.state [0]), .I3(GND_net), .O(n17_adj_3345));   // verilog/coms.v(110[11:16])
    defparam i1_3_lut_adj_1297.LUT_INIT = 16'h8a8a;
    SB_LUT4 i2_4_lut_adj_1298 (.I0(n4_adj_3236), .I1(n1_c), .I2(n17_adj_3345), 
            .I3(\FRAME_MATCHER.state [3]), .O(n10_adj_3344));   // verilog/coms.v(110[11:16])
    defparam i2_4_lut_adj_1298.LUT_INIT = 16'h0032;
    SB_LUT4 select_267_Select_30_i3_2_lut_3_lut (.I0(n1498), .I1(n19_adj_3206), 
            .I2(\FRAME_MATCHER.i [30]), .I3(GND_net), .O(n3_adj_3156));
    defparam select_267_Select_30_i3_2_lut_3_lut.LUT_INIT = 16'h4040;
    SB_LUT4 i25485_2_lut (.I0(n10_adj_3344), .I1(n1498), .I2(GND_net), 
            .I3(GND_net), .O(n41003));
    defparam i25485_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 select_267_Select_31_i3_2_lut_3_lut (.I0(n1498), .I1(n19_adj_3206), 
            .I2(\FRAME_MATCHER.i [31]), .I3(GND_net), .O(n3));
    defparam select_267_Select_31_i3_2_lut_3_lut.LUT_INIT = 16'h4040;
    SB_LUT4 i1_3_lut_adj_1299 (.I0(n20075), .I1(\FRAME_MATCHER.i_31__N_1821 ), 
            .I2(n740), .I3(GND_net), .O(n47));   // verilog/coms.v(113[11:12])
    defparam i1_3_lut_adj_1299.LUT_INIT = 16'h0808;
    SB_LUT4 i2_2_lut_adj_1300 (.I0(\FRAME_MATCHER.i [23]), .I1(\FRAME_MATCHER.i [26]), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_3346));
    defparam i2_2_lut_adj_1300.LUT_INIT = 16'heeee;
    SB_LUT4 i1_4_lut_adj_1301 (.I0(\FRAME_MATCHER.i [7]), .I1(\FRAME_MATCHER.i [20]), 
            .I2(n6_adj_3346), .I3(\FRAME_MATCHER.i [24]), .O(n6_adj_3347));
    defparam i1_4_lut_adj_1301.LUT_INIT = 16'hfffe;
    SB_LUT4 i3_3_lut_adj_1302 (.I0(\FRAME_MATCHER.i [29]), .I1(\FRAME_MATCHER.i [22]), 
            .I2(\FRAME_MATCHER.i [13]), .I3(GND_net), .O(n8_adj_3348));
    defparam i3_3_lut_adj_1302.LUT_INIT = 16'hfefe;
    SB_LUT4 i4_4_lut_adj_1303 (.I0(\FRAME_MATCHER.i [16]), .I1(\FRAME_MATCHER.i [9]), 
            .I2(\FRAME_MATCHER.i [19]), .I3(n6_adj_3347), .O(n42018));
    defparam i4_4_lut_adj_1303.LUT_INIT = 16'hfffe;
    SB_LUT4 i6_4_lut_adj_1304 (.I0(\FRAME_MATCHER.i [27]), .I1(\FRAME_MATCHER.i [10]), 
            .I2(\FRAME_MATCHER.i [21]), .I3(\FRAME_MATCHER.i [6]), .O(n14_adj_3349));
    defparam i6_4_lut_adj_1304.LUT_INIT = 16'hfffe;
    SB_LUT4 i5_4_lut_adj_1305 (.I0(\FRAME_MATCHER.i [8]), .I1(\FRAME_MATCHER.i [28]), 
            .I2(\FRAME_MATCHER.i [25]), .I3(\FRAME_MATCHER.i [11]), .O(n13_adj_3350));
    defparam i5_4_lut_adj_1305.LUT_INIT = 16'hfffe;
    SB_LUT4 i2_4_lut_adj_1306 (.I0(\FRAME_MATCHER.i [12]), .I1(n42018), 
            .I2(n8_adj_3348), .I3(\FRAME_MATCHER.i [30]), .O(n9_adj_3351));
    defparam i2_4_lut_adj_1306.LUT_INIT = 16'hfffe;
    SB_LUT4 i4_4_lut_adj_1307 (.I0(\FRAME_MATCHER.i [14]), .I1(\FRAME_MATCHER.i [18]), 
            .I2(n13_adj_3350), .I3(n14_adj_3349), .O(n11_adj_3352));
    defparam i4_4_lut_adj_1307.LUT_INIT = 16'hfffe;
    SB_LUT4 i6_4_lut_adj_1308 (.I0(n11_adj_3352), .I1(n9_adj_3351), .I2(\FRAME_MATCHER.i [15]), 
            .I3(\FRAME_MATCHER.i [17]), .O(n22400));
    defparam i6_4_lut_adj_1308.LUT_INIT = 16'hfffe;
    SB_LUT4 i10497_3_lut_4_lut (.I0(n8_adj_3124), .I1(n40212), .I2(rx_data[7]), 
            .I3(\data_in_frame[2] [7]), .O(n23915));
    defparam i10497_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i14442_4_lut (.I0(n10_adj_3353), .I1(\FRAME_MATCHER.i [31]), 
            .I2(\FRAME_MATCHER.i [5]), .I3(n22400), .O(n3761));   // verilog/coms.v(249[9:58])
    defparam i14442_4_lut.LUT_INIT = 16'h3332;
    SB_LUT4 i10498_3_lut_4_lut (.I0(n8_adj_3124), .I1(n40212), .I2(rx_data[6]), 
            .I3(\data_in_frame[2] [6]), .O(n23916));
    defparam i10498_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i27200_2_lut (.I0(byte_transmit_counter_c[2]), .I1(byte_transmit_counter[1]), 
            .I2(GND_net), .I3(GND_net), .O(n43966));
    defparam i27200_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i5_3_lut_adj_1309 (.I0(\data_in[0] [3]), .I1(\data_in[1] [4]), 
            .I2(\data_in[1] [5]), .I3(GND_net), .O(n14_adj_3354));
    defparam i5_3_lut_adj_1309.LUT_INIT = 16'hdfdf;
    SB_LUT4 i6_4_lut_adj_1310 (.I0(\data_in[0] [6]), .I1(n22476), .I2(\data_in[2] [4]), 
            .I3(\data_in[1] [0]), .O(n15_adj_3355));
    defparam i6_4_lut_adj_1310.LUT_INIT = 16'hfeff;
    SB_LUT4 i8_4_lut_adj_1311 (.I0(n15_adj_3355), .I1(\data_in[3] [0]), 
            .I2(n14_adj_3354), .I3(\data_in[2] [2]), .O(n22256));
    defparam i8_4_lut_adj_1311.LUT_INIT = 16'hfbff;
    SB_LUT4 i6_4_lut_adj_1312 (.I0(\data_in[1] [3]), .I1(\data_in[0] [1]), 
            .I2(\data_in[3] [2]), .I3(\data_in[0] [5]), .O(n16_adj_3356));
    defparam i6_4_lut_adj_1312.LUT_INIT = 16'hfffe;
    SB_LUT4 i7_4_lut_adj_1313 (.I0(\data_in[2] [6]), .I1(\data_in[2] [5]), 
            .I2(\data_in[2] [0]), .I3(\data_in[1] [2]), .O(n17_adj_3357));
    defparam i7_4_lut_adj_1313.LUT_INIT = 16'hfffd;
    SB_LUT4 i9_4_lut_adj_1314 (.I0(n17_adj_3357), .I1(\data_in[1] [6]), 
            .I2(n16_adj_3356), .I3(\data_in[3] [7]), .O(n22341));
    defparam i9_4_lut_adj_1314.LUT_INIT = 16'hfbff;
    SB_LUT4 i4_4_lut_adj_1315 (.I0(\data_in[1] [7]), .I1(\data_in[0] [0]), 
            .I2(\data_in[1] [1]), .I3(\data_in[0] [4]), .O(n10_adj_3358));
    defparam i4_4_lut_adj_1315.LUT_INIT = 16'hfdff;
    SB_LUT4 i5_3_lut_adj_1316 (.I0(\data_in[3] [4]), .I1(n10_adj_3358), 
            .I2(\data_in[2] [7]), .I3(GND_net), .O(n22476));
    defparam i5_3_lut_adj_1316.LUT_INIT = 16'hdfdf;
    SB_LUT4 i4_2_lut (.I0(\data_in[3] [1]), .I1(\data_in[0] [7]), .I2(GND_net), 
            .I3(GND_net), .O(n12_adj_3359));
    defparam i4_2_lut.LUT_INIT = 16'hbbbb;
    SB_LUT4 i5_4_lut_adj_1317 (.I0(\data_in[3] [5]), .I1(\data_in[2] [1]), 
            .I2(\data_in[2] [3]), .I3(\data_in[3] [3]), .O(n13_adj_3360));
    defparam i5_4_lut_adj_1317.LUT_INIT = 16'hfffe;
    SB_LUT4 i7_4_lut_adj_1318 (.I0(n13_adj_3360), .I1(\data_in[3] [6]), 
            .I2(n12_adj_3359), .I3(\data_in[0] [2]), .O(n22374));
    defparam i7_4_lut_adj_1318.LUT_INIT = 16'hfffb;
    SB_LUT4 i7_4_lut_adj_1319 (.I0(\data_in[2] [4]), .I1(n22374), .I2(\data_in[1] [5]), 
            .I3(n22476), .O(n18_adj_3361));
    defparam i7_4_lut_adj_1319.LUT_INIT = 16'hfffd;
    SB_LUT4 i9_4_lut_adj_1320 (.I0(\data_in[0] [6]), .I1(n18_adj_3361), 
            .I2(\data_in[3] [0]), .I3(n22341), .O(n20_adj_3362));
    defparam i9_4_lut_adj_1320.LUT_INIT = 16'hfffd;
    SB_LUT4 i4_2_lut_adj_1321 (.I0(\data_in[1] [0]), .I1(\data_in[0] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n15_adj_3363));
    defparam i4_2_lut_adj_1321.LUT_INIT = 16'heeee;
    SB_LUT4 i10_4_lut_adj_1322 (.I0(n15_adj_3363), .I1(n20_adj_3362), .I2(\data_in[2] [2]), 
            .I3(\data_in[1] [4]), .O(n63_adj_3248));
    defparam i10_4_lut_adj_1322.LUT_INIT = 16'hfeff;
    SB_LUT4 i6_4_lut_adj_1323 (.I0(\data_in[3] [6]), .I1(\data_in[0] [7]), 
            .I2(\data_in[2] [1]), .I3(n22256), .O(n16_adj_3364));
    defparam i6_4_lut_adj_1323.LUT_INIT = 16'hffef;
    SB_LUT4 i7_4_lut_adj_1324 (.I0(n22341), .I1(\data_in[2] [3]), .I2(\data_in[0] [2]), 
            .I3(\data_in[3] [1]), .O(n17_adj_3365));
    defparam i7_4_lut_adj_1324.LUT_INIT = 16'hbfff;
    SB_LUT4 i9_4_lut_adj_1325 (.I0(n17_adj_3365), .I1(\data_in[3] [5]), 
            .I2(n16_adj_3364), .I3(\data_in[3] [3]), .O(n63_adj_3249));
    defparam i9_4_lut_adj_1325.LUT_INIT = 16'hfbff;
    SB_LUT4 i8_4_lut_adj_1326 (.I0(n22374), .I1(\data_in[1] [3]), .I2(n22256), 
            .I3(\data_in[2] [0]), .O(n20_adj_3366));
    defparam i8_4_lut_adj_1326.LUT_INIT = 16'hfbff;
    SB_LUT4 i7_4_lut_adj_1327 (.I0(\data_in[2] [6]), .I1(\data_in[1] [6]), 
            .I2(\data_in[3] [7]), .I3(\data_in[0] [1]), .O(n19_adj_3367));
    defparam i7_4_lut_adj_1327.LUT_INIT = 16'hfeff;
    SB_LUT4 i26660_4_lut (.I0(\data_in[1] [2]), .I1(\data_in[3] [2]), .I2(\data_in[2] [5]), 
            .I3(\data_in[0] [5]), .O(n42179));
    defparam i26660_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i11_3_lut_adj_1328 (.I0(n42179), .I1(n19_adj_3367), .I2(n20_adj_3366), 
            .I3(GND_net), .O(n63));
    defparam i11_3_lut_adj_1328.LUT_INIT = 16'hfdfd;
    SB_LUT4 i1_3_lut_adj_1329 (.I0(n736), .I1(\FRAME_MATCHER.i_31__N_1824 ), 
            .I2(n20075), .I3(GND_net), .O(n43));
    defparam i1_3_lut_adj_1329.LUT_INIT = 16'h8080;
    SB_LUT4 i1_3_lut_adj_1330 (.I0(n3761), .I1(\FRAME_MATCHER.i_31__N_1827 ), 
            .I2(n20075), .I3(GND_net), .O(n5_adj_3238));
    defparam i1_3_lut_adj_1330.LUT_INIT = 16'h4040;
    SB_LUT4 i10499_3_lut_4_lut (.I0(n8_adj_3124), .I1(n40212), .I2(rx_data[5]), 
            .I3(\data_in_frame[2] [5]), .O(n23917));
    defparam i10499_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10622_3_lut_4_lut (.I0(\FRAME_MATCHER.state [2]), .I1(n22338), 
            .I2(encoder0_position[1]), .I3(\data_out_frame[8] [1]), .O(n24040));
    defparam i10622_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i10623_3_lut_4_lut (.I0(\FRAME_MATCHER.state [2]), .I1(n22338), 
            .I2(encoder0_position[0]), .I3(\data_out_frame[8] [0]), .O(n24041));
    defparam i10623_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i10626_3_lut_4_lut (.I0(\FRAME_MATCHER.state [2]), .I1(n22338), 
            .I2(encoder0_position[13]), .I3(\data_out_frame[7] [5]), .O(n24044));
    defparam i10626_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i10522_3_lut_4_lut (.I0(\FRAME_MATCHER.state [2]), .I1(n22338), 
            .I2(displacement[5]), .I3(\data_out_frame[20] [5]), .O(n23940));
    defparam i10522_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 equal_61_i8_2_lut_3_lut (.I0(\FRAME_MATCHER.i [0]), .I1(\FRAME_MATCHER.i [1]), 
            .I2(\FRAME_MATCHER.i [2]), .I3(GND_net), .O(n8_adj_3122));   // verilog/coms.v(154[7:23])
    defparam equal_61_i8_2_lut_3_lut.LUT_INIT = 16'hbfbf;
    SB_LUT4 i14345_2_lut_3_lut (.I0(\FRAME_MATCHER.i [0]), .I1(\FRAME_MATCHER.i [1]), 
            .I2(\FRAME_MATCHER.i [2]), .I3(GND_net), .O(n27747));
    defparam i14345_2_lut_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 i10590_3_lut_4_lut (.I0(\FRAME_MATCHER.state [2]), .I1(n22338), 
            .I2(setpoint[17]), .I3(\data_out_frame[12] [1]), .O(n24008));
    defparam i10590_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i10595_3_lut_4_lut (.I0(\FRAME_MATCHER.state [2]), .I1(n22338), 
            .I2(encoder1_position[4]), .I3(\data_out_frame[11] [4]), .O(n24013));
    defparam i10595_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i10591_3_lut_4_lut (.I0(\FRAME_MATCHER.state [2]), .I1(n22338), 
            .I2(setpoint[16]), .I3(\data_out_frame[12] [0]), .O(n24009));
    defparam i10591_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i10592_3_lut_4_lut (.I0(\FRAME_MATCHER.state [2]), .I1(n22338), 
            .I2(encoder1_position[7]), .I3(\data_out_frame[11] [7]), .O(n24010));
    defparam i10592_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i10593_3_lut_4_lut (.I0(\FRAME_MATCHER.state [2]), .I1(n22338), 
            .I2(encoder1_position[6]), .I3(\data_out_frame[11] [6]), .O(n24011));
    defparam i10593_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i10596_3_lut_4_lut (.I0(\FRAME_MATCHER.state [2]), .I1(n22338), 
            .I2(encoder1_position[3]), .I3(\data_out_frame[11] [3]), .O(n24014));
    defparam i10596_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i10597_3_lut_4_lut (.I0(\FRAME_MATCHER.state [2]), .I1(n22338), 
            .I2(encoder1_position[2]), .I3(\data_out_frame[11] [2]), .O(n24015));
    defparam i10597_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i10598_3_lut_4_lut (.I0(\FRAME_MATCHER.state [2]), .I1(n22338), 
            .I2(encoder1_position[1]), .I3(\data_out_frame[11] [1]), .O(n24016));
    defparam i10598_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i1_2_lut_adj_1331 (.I0(\FRAME_MATCHER.i [3]), .I1(\FRAME_MATCHER.i [5]), 
            .I2(GND_net), .I3(GND_net), .O(n22347));   // verilog/coms.v(154[7:23])
    defparam i1_2_lut_adj_1331.LUT_INIT = 16'heeee;
    SB_LUT4 i3_4_lut_adj_1332 (.I0(\FRAME_MATCHER.state [1]), .I1(n27701), 
            .I2(n93), .I3(n1_c), .O(n23399));
    defparam i3_4_lut_adj_1332.LUT_INIT = 16'h0010;
    SB_LUT4 i30697_2_lut_3_lut_4_lut (.I0(n20075), .I1(n11_adj_3246), .I2(\FRAME_MATCHER.state [1]), 
            .I3(\FRAME_MATCHER.state [0]), .O(n40886));
    defparam i30697_2_lut_3_lut_4_lut.LUT_INIT = 16'h5557;
    SB_LUT4 i10631_3_lut_4_lut (.I0(\FRAME_MATCHER.state [2]), .I1(n22338), 
            .I2(encoder0_position[8]), .I3(\data_out_frame[7] [0]), .O(n24049));
    defparam i10631_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i10500_3_lut_4_lut (.I0(n8_adj_3124), .I1(n40212), .I2(rx_data[4]), 
            .I3(\data_in_frame[2] [4]), .O(n23918));
    defparam i10500_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10501_3_lut_4_lut (.I0(n8_adj_3124), .I1(n40212), .I2(rx_data[3]), 
            .I3(\data_in_frame[2] [3]), .O(n23919));
    defparam i10501_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10632_3_lut_4_lut (.I0(\FRAME_MATCHER.state [2]), .I1(n22338), 
            .I2(encoder0_position[23]), .I3(\data_out_frame[6] [7]), .O(n24050));
    defparam i10632_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i10633_3_lut_4_lut (.I0(\FRAME_MATCHER.state [2]), .I1(n22338), 
            .I2(encoder0_position[22]), .I3(\data_out_frame[6] [6]), .O(n24051));
    defparam i10633_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i10634_3_lut_4_lut (.I0(\FRAME_MATCHER.state [2]), .I1(n22338), 
            .I2(encoder0_position[21]), .I3(\data_out_frame[6] [5]), .O(n24052));
    defparam i10634_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i10635_3_lut_4_lut (.I0(\FRAME_MATCHER.state [2]), .I1(n22338), 
            .I2(encoder0_position[20]), .I3(\data_out_frame[6] [4]), .O(n24053));
    defparam i10635_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i10636_3_lut_4_lut (.I0(\FRAME_MATCHER.state [2]), .I1(n22338), 
            .I2(encoder0_position[19]), .I3(\data_out_frame[6] [3]), .O(n24054));
    defparam i10636_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i26756_3_lut (.I0(\data_out_frame[8] [7]), .I1(\data_out_frame[9] [7]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n42275));
    defparam i26756_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10534_3_lut_4_lut (.I0(\FRAME_MATCHER.state [2]), .I1(n22338), 
            .I2(displacement[9]), .I3(\data_out_frame[19] [1]), .O(n23952));
    defparam i10534_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i26757_3_lut (.I0(\data_out_frame[10] [7]), .I1(\data_out_frame[11] [7]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n42276));
    defparam i26757_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i26760_3_lut (.I0(\data_out_frame[14] [7]), .I1(\data_out_frame[15] [7]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n42279));
    defparam i26760_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i26759_3_lut (.I0(\data_out_frame[12] [7]), .I1(\data_out_frame[13] [7]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n42278));
    defparam i26759_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10638_3_lut_4_lut (.I0(\FRAME_MATCHER.state [2]), .I1(n22338), 
            .I2(encoder0_position[17]), .I3(\data_out_frame[6] [1]), .O(n24056));
    defparam i10638_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i10640_3_lut_4_lut (.I0(\FRAME_MATCHER.state [2]), .I1(n22338), 
            .I2(control_mode[7]), .I3(\data_out_frame[5] [7]), .O(n24058));
    defparam i10640_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i10502_3_lut_4_lut (.I0(n8_adj_3124), .I1(n40212), .I2(rx_data[2]), 
            .I3(\data_in_frame[2] [2]), .O(n23920));
    defparam i10502_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10642_3_lut_4_lut (.I0(\FRAME_MATCHER.state [2]), .I1(n22338), 
            .I2(control_mode[5]), .I3(\data_out_frame[5] [5]), .O(n24060));
    defparam i10642_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i10646_3_lut_4_lut (.I0(\FRAME_MATCHER.state [2]), .I1(n22338), 
            .I2(control_mode[1]), .I3(\data_out_frame[5] [1]), .O(n24064));
    defparam i10646_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i10643_3_lut_4_lut (.I0(\FRAME_MATCHER.state [2]), .I1(n22338), 
            .I2(control_mode[4]), .I3(\data_out_frame[5] [4]), .O(n24061));
    defparam i10643_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i10644_3_lut_4_lut (.I0(\FRAME_MATCHER.state [2]), .I1(n22338), 
            .I2(control_mode[3]), .I3(\data_out_frame[5] [3]), .O(n24062));
    defparam i10644_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i10647_3_lut_4_lut (.I0(\FRAME_MATCHER.state [2]), .I1(n22338), 
            .I2(control_mode[0]), .I3(\data_out_frame[5] [0]), .O(n24065));
    defparam i10647_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i10599_3_lut_4_lut (.I0(\FRAME_MATCHER.state [2]), .I1(n22338), 
            .I2(encoder1_position[0]), .I3(\data_out_frame[11] [0]), .O(n24017));
    defparam i10599_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i10503_3_lut_4_lut (.I0(n8_adj_3124), .I1(n40212), .I2(rx_data[1]), 
            .I3(\data_in_frame[2] [1]), .O(n23921));
    defparam i10503_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10600_3_lut_4_lut (.I0(\FRAME_MATCHER.state [2]), .I1(n22338), 
            .I2(encoder1_position[15]), .I3(\data_out_frame[10] [7]), .O(n24018));
    defparam i10600_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i10601_3_lut_4_lut (.I0(\FRAME_MATCHER.state [2]), .I1(n22338), 
            .I2(encoder1_position[14]), .I3(\data_out_frame[10] [6]), .O(n24019));
    defparam i10601_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i10504_3_lut_4_lut (.I0(n8_adj_3124), .I1(n40212), .I2(rx_data[0]), 
            .I3(\data_in_frame[2] [0]), .O(n23922));
    defparam i10504_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10602_3_lut_4_lut (.I0(\FRAME_MATCHER.state [2]), .I1(n22338), 
            .I2(encoder1_position[13]), .I3(\data_out_frame[10] [5]), .O(n24020));
    defparam i10602_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i10603_3_lut_4_lut (.I0(\FRAME_MATCHER.state [2]), .I1(n22338), 
            .I2(encoder1_position[12]), .I3(\data_out_frame[10] [4]), .O(n24021));
    defparam i10603_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 equal_65_i8_2_lut_3_lut (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(\FRAME_MATCHER.i [0]), .I3(GND_net), .O(n8_adj_3124));   // verilog/coms.v(154[7:23])
    defparam equal_65_i8_2_lut_3_lut.LUT_INIT = 16'hfdfd;
    SB_LUT4 i10604_3_lut_4_lut (.I0(\FRAME_MATCHER.state [2]), .I1(n22338), 
            .I2(encoder1_position[11]), .I3(\data_out_frame[10] [3]), .O(n24022));
    defparam i10604_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i10606_3_lut_4_lut (.I0(\FRAME_MATCHER.state [2]), .I1(n22338), 
            .I2(encoder1_position[9]), .I3(\data_out_frame[10] [1]), .O(n24024));
    defparam i10606_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i10607_3_lut_4_lut (.I0(\FRAME_MATCHER.state [2]), .I1(n22338), 
            .I2(encoder1_position[8]), .I3(\data_out_frame[10] [0]), .O(n24025));
    defparam i10607_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1333 (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(n40212), .I3(\FRAME_MATCHER.i [0]), .O(n40216));   // verilog/coms.v(154[7:23])
    defparam i1_2_lut_3_lut_4_lut_adj_1333.LUT_INIT = 16'hfdff;
    SB_LUT4 i10611_3_lut_4_lut (.I0(\FRAME_MATCHER.state [2]), .I1(n22338), 
            .I2(encoder1_position[20]), .I3(\data_out_frame[9] [4]), .O(n24029));
    defparam i10611_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i10608_3_lut_4_lut (.I0(\FRAME_MATCHER.state [2]), .I1(n22338), 
            .I2(encoder1_position[23]), .I3(\data_out_frame[9] [7]), .O(n24026));
    defparam i10608_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i10609_3_lut_4_lut (.I0(\FRAME_MATCHER.state [2]), .I1(n22338), 
            .I2(encoder1_position[22]), .I3(\data_out_frame[9] [6]), .O(n24027));
    defparam i10609_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i14855_3_lut_4_lut (.I0(byte_transmit_counter_c[2]), .I1(byte_transmit_counter[1]), 
            .I2(byte_transmit_counter_c[4]), .I3(byte_transmit_counter_c[3]), 
            .O(n28265));
    defparam i14855_3_lut_4_lut.LUT_INIT = 16'hf080;
    SB_LUT4 i1814_3_lut_4_lut (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(\FRAME_MATCHER.i [4]), .I3(\FRAME_MATCHER.i [3]), .O(n10_adj_3353));
    defparam i1814_3_lut_4_lut.LUT_INIT = 16'hf080;
    SB_LUT4 i1_3_lut_4_lut (.I0(\FRAME_MATCHER.i_31__N_1825 ), .I1(n22250), 
            .I2(\FRAME_MATCHER.i [31]), .I3(n20075), .O(n2_adj_3220));   // verilog/coms.v(126[12] 289[6])
    defparam i1_3_lut_4_lut.LUT_INIT = 16'ha200;
    SB_LUT4 i2_3_lut_4_lut_adj_1334 (.I0(\FRAME_MATCHER.i_31__N_1823 ), .I1(n10_adj_3344), 
            .I2(n1498), .I3(n20075), .O(n6_adj_3221));
    defparam i2_3_lut_4_lut_adj_1334.LUT_INIT = 16'h0100;
    SB_LUT4 i1_2_lut_3_lut_adj_1335 (.I0(\FRAME_MATCHER.state [3]), .I1(\FRAME_MATCHER.state [1]), 
            .I2(\FRAME_MATCHER.state [0]), .I3(GND_net), .O(n40173));   // verilog/coms.v(126[12] 289[6])
    defparam i1_2_lut_3_lut_adj_1335.LUT_INIT = 16'h0202;
    SB_LUT4 i1_3_lut_4_lut_adj_1336 (.I0(n7[1]), .I1(\FRAME_MATCHER.i_31__N_1827 ), 
            .I2(n3761), .I3(n63), .O(n36044));
    defparam i1_3_lut_4_lut_adj_1336.LUT_INIT = 16'h080c;
    SB_LUT4 i2_3_lut_4_lut_adj_1337 (.I0(n37308), .I1(\data_out_frame[20] [6]), 
            .I2(\data_out_frame[20] [5]), .I3(n22071), .O(n41574));
    defparam i2_3_lut_4_lut_adj_1337.LUT_INIT = 16'h9669;
    SB_LUT4 i2_3_lut_4_lut_adj_1338 (.I0(n40440), .I1(n40696), .I2(\data_out_frame[16] [3]), 
            .I3(\data_out_frame[18] [4]), .O(n37308));
    defparam i2_3_lut_4_lut_adj_1338.LUT_INIT = 16'h6996;
    SB_LUT4 i3_2_lut_3_lut (.I0(\data_out_frame[11] [6]), .I1(\data_out_frame[9] [5]), 
            .I2(\data_out_frame[7] [2]), .I3(GND_net), .O(n9_adj_3340));
    defparam i3_2_lut_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_4_lut_adj_1339 (.I0(\data_out_frame[9] [2]), .I1(\data_out_frame[5][2] ), 
            .I2(\data_out_frame[9] [4]), .I3(\data_out_frame[11] [4]), .O(n40295));
    defparam i2_3_lut_4_lut_adj_1339.LUT_INIT = 16'h6996;
    SB_LUT4 i5_3_lut_4_lut_adj_1340 (.I0(\data_out_frame[7] [4]), .I1(\data_out_frame[5] [3]), 
            .I2(n10_adj_3335), .I3(\data_out_frame[9] [7]), .O(n23000));   // verilog/coms.v(72[16:27])
    defparam i5_3_lut_4_lut_adj_1340.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_adj_1341 (.I0(\data_out_frame[15] [7]), .I1(n36529), 
            .I2(\data_out_frame[13] [5]), .I3(n1515), .O(n40380));
    defparam i1_2_lut_4_lut_adj_1341.LUT_INIT = 16'h6996;
    SB_LUT4 i5_2_lut_3_lut_4_lut (.I0(\data_out_frame[7] [5]), .I1(n22635), 
            .I2(\data_out_frame[12] [1]), .I3(\data_out_frame[12] [0]), 
            .O(n36));   // verilog/coms.v(73[16:27])
    defparam i5_2_lut_3_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1342 (.I0(\data_out_frame[11] [3]), .I1(\data_out_frame[8] [7]), 
            .I2(\data_out_frame[7] [2]), .I3(GND_net), .O(n6_adj_3334));
    defparam i1_2_lut_3_lut_adj_1342.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1343 (.I0(\data_out_frame[7] [0]), .I1(\data_out_frame[13] [7]), 
            .I2(\data_out_frame[13] [6]), .I3(GND_net), .O(n40803));   // verilog/coms.v(71[16:27])
    defparam i1_2_lut_3_lut_adj_1343.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1344 (.I0(\data_out_frame[16] [4]), .I1(n23383), 
            .I2(n40440), .I3(GND_net), .O(n40411));
    defparam i1_2_lut_3_lut_adj_1344.LUT_INIT = 16'h9696;
    SB_LUT4 i5_2_lut_3_lut (.I0(\data_out_frame[7] [2]), .I1(\data_out_frame[15] [6]), 
            .I2(n40289), .I3(GND_net), .O(n16_adj_3330));   // verilog/coms.v(71[16:27])
    defparam i5_2_lut_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1345 (.I0(\data_out_frame[8] [7]), .I1(\data_out_frame[8] [6]), 
            .I2(\data_out_frame[8] [5]), .I3(GND_net), .O(n23004));   // verilog/coms.v(72[16:27])
    defparam i1_2_lut_3_lut_adj_1345.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1346 (.I0(\data_out_frame[16] [0]), .I1(n22051), 
            .I2(n40684), .I3(GND_net), .O(n6_adj_3325));
    defparam i1_2_lut_3_lut_adj_1346.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1347 (.I0(n37264), .I1(n40576), .I2(n40311), 
            .I3(GND_net), .O(n37234));
    defparam i1_2_lut_3_lut_adj_1347.LUT_INIT = 16'h6969;
    SB_LUT4 i2_3_lut_4_lut_adj_1348 (.I0(\data_out_frame[10] [7]), .I1(\data_out_frame[6] [1]), 
            .I2(n40298), .I3(\data_out_frame[6] [5]), .O(n40634));   // verilog/coms.v(72[16:27])
    defparam i2_3_lut_4_lut_adj_1348.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_1349 (.I0(\data_out_frame[17] [7]), .I1(\data_out_frame[17] [6]), 
            .I2(n23107), .I3(\data_out_frame[17] [4]), .O(n40576));
    defparam i2_3_lut_4_lut_adj_1349.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_1350 (.I0(\data_out_frame[10] [4]), .I1(\data_out_frame[6] [2]), 
            .I2(\data_out_frame[6] [0]), .I3(\data_out_frame[8] [3]), .O(n40506));   // verilog/coms.v(71[16:34])
    defparam i2_3_lut_4_lut_adj_1350.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_1351 (.I0(\data_out_frame[5] [6]), .I1(\data_out_frame[5] [7]), 
            .I2(n40609), .I3(\data_out_frame[6] [0]), .O(n22095));   // verilog/coms.v(73[16:27])
    defparam i2_3_lut_4_lut_adj_1351.LUT_INIT = 16'h6996;
    SB_LUT4 i3_2_lut_3_lut_adj_1352 (.I0(Kp_23__N_379), .I1(\data_in_frame[5] [7]), 
            .I2(n23101), .I3(GND_net), .O(n16_adj_3310));   // verilog/coms.v(230[9:81])
    defparam i3_2_lut_3_lut_adj_1352.LUT_INIT = 16'hf6f6;
    SB_LUT4 i1_2_lut_3_lut_adj_1353 (.I0(\data_out_frame[12] [5]), .I1(\data_out_frame[10] [3]), 
            .I2(n40474), .I3(GND_net), .O(n40873));
    defparam i1_2_lut_3_lut_adj_1353.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_4_lut_adj_1354 (.I0(\data_out_frame[12] [4]), .I1(\data_out_frame[10] [3]), 
            .I2(\data_out_frame[10] [2]), .I3(n22095), .O(n40656));
    defparam i1_2_lut_4_lut_adj_1354.LUT_INIT = 16'h6996;
    SB_LUT4 i10610_3_lut_4_lut (.I0(\FRAME_MATCHER.state [2]), .I1(n22338), 
            .I2(encoder1_position[21]), .I3(\data_out_frame[9] [5]), .O(n24028));
    defparam i10610_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i1_2_lut_3_lut_adj_1355 (.I0(\data_out_frame[8] [2]), .I1(\data_out_frame[5] [6]), 
            .I2(\data_out_frame[5] [7]), .I3(GND_net), .O(n40665));   // verilog/coms.v(71[16:34])
    defparam i1_2_lut_3_lut_adj_1355.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1356 (.I0(n36837), .I1(\data_out_frame[14] [5]), 
            .I2(n22134), .I3(GND_net), .O(n40415));
    defparam i1_2_lut_3_lut_adj_1356.LUT_INIT = 16'h9696;
    SB_LUT4 i2_2_lut_3_lut_adj_1357 (.I0(\FRAME_MATCHER.state [3]), .I1(\FRAME_MATCHER.state [2]), 
            .I2(\FRAME_MATCHER.state [0]), .I3(GND_net), .O(n93));
    defparam i2_2_lut_3_lut_adj_1357.LUT_INIT = 16'h0404;
    SB_LUT4 i10612_3_lut_4_lut (.I0(\FRAME_MATCHER.state [2]), .I1(n22338), 
            .I2(encoder1_position[19]), .I3(\data_out_frame[9] [3]), .O(n24030));
    defparam i10612_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i10613_3_lut_4_lut (.I0(\FRAME_MATCHER.state [2]), .I1(n22338), 
            .I2(encoder1_position[18]), .I3(\data_out_frame[9] [2]), .O(n24031));
    defparam i10613_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i10614_3_lut_4_lut (.I0(\FRAME_MATCHER.state [2]), .I1(n22338), 
            .I2(encoder1_position[17]), .I3(\data_out_frame[9] [1]), .O(n24032));
    defparam i10614_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i10615_3_lut_4_lut (.I0(\FRAME_MATCHER.state [2]), .I1(n22338), 
            .I2(encoder1_position[16]), .I3(\data_out_frame[9] [0]), .O(n24033));
    defparam i10615_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i10616_3_lut_4_lut (.I0(\FRAME_MATCHER.state [2]), .I1(n22338), 
            .I2(encoder0_position[7]), .I3(\data_out_frame[8] [7]), .O(n24034));
    defparam i10616_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1358 (.I0(\data_out_frame[5] [7]), .I1(\data_out_frame[8] [3]), 
            .I2(\data_out_frame[8] [4]), .I3(\data_out_frame[10] [5]), .O(n40298));
    defparam i1_2_lut_3_lut_4_lut_adj_1358.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_adj_1359 (.I0(n40506), .I1(\data_out_frame[10] [7]), 
            .I2(n40767), .I3(\data_out_frame[6] [5]), .O(n6_adj_3303));   // verilog/coms.v(73[16:27])
    defparam i1_2_lut_4_lut_adj_1359.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1360 (.I0(\data_out_frame[17] [3]), .I1(\data_out_frame[17] [1]), 
            .I2(\data_out_frame[17] [2]), .I3(\data_out_frame[17] [5]), 
            .O(n23107));
    defparam i1_2_lut_3_lut_4_lut_adj_1360.LUT_INIT = 16'h6996;
    SB_LUT4 i14_3_lut_4_lut (.I0(\data_out_frame[16] [3]), .I1(\data_out_frame[16] [7]), 
            .I2(n28_adj_3299), .I3(\data_out_frame[12] [4]), .O(n32));
    defparam i14_3_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1361 (.I0(\data_out_frame[14] [6]), .I1(\data_out_frame[16] [4]), 
            .I2(\data_out_frame[16] [5]), .I3(GND_net), .O(n40813));
    defparam i1_2_lut_3_lut_adj_1361.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1362 (.I0(\data_out_frame[19] [2]), .I1(\data_out_frame[19] [1]), 
            .I2(\data_out_frame[19] [5]), .I3(GND_net), .O(n18_adj_3293));
    defparam i1_2_lut_3_lut_adj_1362.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1363 (.I0(n41402), .I1(n37255), .I2(n36629), 
            .I3(GND_net), .O(n40514));
    defparam i1_2_lut_3_lut_adj_1363.LUT_INIT = 16'h6969;
    SB_LUT4 i10617_3_lut_4_lut (.I0(\FRAME_MATCHER.state [2]), .I1(n22338), 
            .I2(encoder0_position[6]), .I3(\data_out_frame[8] [6]), .O(n24035));
    defparam i10617_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1364 (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(n40221), .I3(\FRAME_MATCHER.i [0]), .O(n40225));   // verilog/coms.v(154[7:23])
    defparam i1_2_lut_3_lut_4_lut_adj_1364.LUT_INIT = 16'hfdff;
    SB_LUT4 i5_3_lut_4_lut_adj_1365 (.I0(\data_out_frame[16] [4]), .I1(n1716), 
            .I2(n10_adj_3287), .I3(\data_out_frame[19] [1]), .O(n41758));
    defparam i5_3_lut_4_lut_adj_1365.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_1366 (.I0(\data_in_frame[0] [6]), .I1(\data_in_frame[1] [0]), 
            .I2(\data_in_frame[2] [7]), .I3(\data_in_frame[1] [1]), .O(n41662));   // verilog/coms.v(76[16:27])
    defparam i2_3_lut_4_lut_adj_1366.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1367 (.I0(n11_adj_3246), .I1(\FRAME_MATCHER.state [1]), 
            .I2(\FRAME_MATCHER.state [0]), .I3(GND_net), .O(n19_adj_3206));
    defparam i1_2_lut_3_lut_adj_1367.LUT_INIT = 16'hfefe;
    SB_LUT4 i19_3_lut_4_lut (.I0(Kp_23__N_152), .I1(n27691), .I2(\FRAME_MATCHER.state [3]), 
            .I3(\FRAME_MATCHER.state [2]), .O(n8_adj_3283));   // verilog/coms.v(126[12] 289[6])
    defparam i19_3_lut_4_lut.LUT_INIT = 16'h02f0;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1368 (.I0(\FRAME_MATCHER.i_31__N_1824 ), 
            .I1(n736), .I2(n41992), .I3(n5_adj_3250), .O(n5_adj_3219));
    defparam i1_2_lut_3_lut_4_lut_adj_1368.LUT_INIT = 16'hff8f;
    SB_LUT4 i1_2_lut_4_lut_adj_1369 (.I0(\data_in_frame[4] [2]), .I1(n40383), 
            .I2(\data_in_frame[6] [6]), .I3(\data_in_frame[9] [0]), .O(n40819));   // verilog/coms.v(69[16:27])
    defparam i1_2_lut_4_lut_adj_1369.LUT_INIT = 16'h6996;
    SB_LUT4 i10618_3_lut_4_lut (.I0(\FRAME_MATCHER.state [2]), .I1(n22338), 
            .I2(encoder0_position[5]), .I3(\data_out_frame[8] [5]), .O(n24036));
    defparam i10618_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i1_2_lut_4_lut_adj_1370 (.I0(\data_in_frame[15] [3]), .I1(n22670), 
            .I2(n40531), .I3(\data_in_frame[10] [7]), .O(n40540));   // verilog/coms.v(73[16:43])
    defparam i1_2_lut_4_lut_adj_1370.LUT_INIT = 16'h6996;
    SB_LUT4 i2_2_lut_3_lut_adj_1371 (.I0(n22721), .I1(\data_in_frame[6] [5]), 
            .I2(\data_in_frame[8] [6]), .I3(GND_net), .O(n10_adj_3269));   // verilog/coms.v(72[16:43])
    defparam i2_2_lut_3_lut_adj_1371.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_4_lut_adj_1372 (.I0(\data_in_frame[8] [5]), .I1(\data_in_frame[8] [4]), 
            .I2(n23275), .I3(\data_in_frame[13] [1]), .O(n40326));   // verilog/coms.v(69[16:27])
    defparam i2_3_lut_4_lut_adj_1372.LUT_INIT = 16'h6996;
    SB_LUT4 i5_3_lut_4_lut_adj_1373 (.I0(Kp_23__N_379), .I1(\data_in_frame[5] [7]), 
            .I2(n10_adj_3266), .I3(n23275), .O(n22670));   // verilog/coms.v(70[16:41])
    defparam i5_3_lut_4_lut_adj_1373.LUT_INIT = 16'h6996;
    SB_LUT4 i10619_3_lut_4_lut (.I0(\FRAME_MATCHER.state [2]), .I1(n22338), 
            .I2(encoder0_position[4]), .I3(\data_out_frame[8] [4]), .O(n24037));
    defparam i10619_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i2_3_lut_4_lut_adj_1374 (.I0(\data_in_frame[8] [3]), .I1(n10_adj_3263), 
            .I2(\data_in_frame[6] [2]), .I3(\data_in_frame[6][0] ), .O(n40322));   // verilog/coms.v(83[17:28])
    defparam i2_3_lut_4_lut_adj_1374.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1375 (.I0(\data_in_frame[10] [6]), .I1(\data_in_frame[13] [0]), 
            .I2(n40531), .I3(GND_net), .O(n6_adj_3262));   // verilog/coms.v(69[16:27])
    defparam i1_2_lut_3_lut_adj_1375.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1376 (.I0(\data_in_frame[8] [1]), .I1(\data_in_frame[10] [4]), 
            .I2(\data_in_frame[12] [5]), .I3(GND_net), .O(n6_adj_3261));   // verilog/coms.v(69[16:27])
    defparam i1_2_lut_3_lut_adj_1376.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1377 (.I0(\FRAME_MATCHER.state [2]), 
            .I1(n1_c), .I2(\FRAME_MATCHER.state [3]), .I3(n105), .O(\FRAME_MATCHER.i_31__N_1823 ));
    defparam i1_2_lut_3_lut_4_lut_adj_1377.LUT_INIT = 16'h0010;
    SB_LUT4 i2_3_lut_4_lut_adj_1378 (.I0(\data_in_frame[16] [7]), .I1(n37228), 
            .I2(n40693), .I3(\data_in_frame[16] [5]), .O(n37237));
    defparam i2_3_lut_4_lut_adj_1378.LUT_INIT = 16'h6996;
    SB_LUT4 i2_2_lut_4_lut (.I0(\data_in_frame[8] [7]), .I1(n10_adj_3263), 
            .I2(n22716), .I3(\data_in_frame[6] [4]), .O(n10_adj_3245));
    defparam i2_2_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1379 (.I0(n10_adj_3263), .I1(n22716), .I2(\data_in_frame[6] [4]), 
            .I3(GND_net), .O(n40705));   // verilog/coms.v(72[16:43])
    defparam i1_2_lut_3_lut_adj_1379.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1380 (.I0(n22721), .I1(n23101), .I2(\data_in_frame[11] [1]), 
            .I3(GND_net), .O(n40450));   // verilog/coms.v(69[16:27])
    defparam i1_2_lut_3_lut_adj_1380.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_4_lut_adj_1381 (.I0(n8_adj_3128), .I1(n10_adj_3266), 
            .I2(n23275), .I3(n40867), .O(n6_adj_3243));   // verilog/coms.v(69[16:27])
    defparam i1_2_lut_4_lut_adj_1381.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_adj_1382 (.I0(\data_in_frame[6][1] ), .I1(\data_in_frame[8] [3]), 
            .I2(n23224), .I3(\data_in_frame[6][0] ), .O(n40653));   // verilog/coms.v(83[17:28])
    defparam i1_2_lut_4_lut_adj_1382.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_1383 (.I0(\data_in_frame[18] [3]), .I1(\data_in_frame[16] [3]), 
            .I2(n40515), .I3(\data_in_frame[18] [4]), .O(n40377));
    defparam i2_3_lut_4_lut_adj_1383.LUT_INIT = 16'h6996;
    SB_LUT4 i2_2_lut_3_lut_adj_1384 (.I0(\data_in_frame[17] [1]), .I1(\data_in_frame[17] [0]), 
            .I2(n40365), .I3(GND_net), .O(n6_adj_3239));
    defparam i2_2_lut_3_lut_adj_1384.LUT_INIT = 16'h9696;
    SB_LUT4 i10620_3_lut_4_lut (.I0(\FRAME_MATCHER.state [2]), .I1(n22338), 
            .I2(encoder0_position[3]), .I3(\data_out_frame[8] [3]), .O(n24038));
    defparam i10620_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i10621_3_lut_4_lut (.I0(\FRAME_MATCHER.state [2]), .I1(n22338), 
            .I2(encoder0_position[2]), .I3(\data_out_frame[8] [2]), .O(n24039));
    defparam i10621_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i10624_3_lut_4_lut (.I0(\FRAME_MATCHER.state [2]), .I1(n22338), 
            .I2(encoder0_position[15]), .I3(\data_out_frame[7] [7]), .O(n24042));
    defparam i10624_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i10627_3_lut_4_lut (.I0(\FRAME_MATCHER.state [2]), .I1(n22338), 
            .I2(encoder0_position[12]), .I3(\data_out_frame[7] [4]), .O(n24045));
    defparam i10627_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1385 (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(n40205), .I3(\FRAME_MATCHER.i [0]), .O(n40211));   // verilog/coms.v(154[7:23])
    defparam i1_2_lut_3_lut_4_lut_adj_1385.LUT_INIT = 16'hfdff;
    SB_LUT4 i1_2_lut_3_lut_adj_1386 (.I0(\data_in_frame[18] [7]), .I1(\data_in_frame[18] [6]), 
            .I2(n23301), .I3(GND_net), .O(n40564));
    defparam i1_2_lut_3_lut_adj_1386.LUT_INIT = 16'h9696;
    SB_LUT4 i10520_3_lut_4_lut (.I0(\FRAME_MATCHER.state [2]), .I1(n22338), 
            .I2(displacement[7]), .I3(\data_out_frame[20][7] ), .O(n23938));
    defparam i10520_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i10521_3_lut_4_lut (.I0(\FRAME_MATCHER.state [2]), .I1(n22338), 
            .I2(displacement[6]), .I3(\data_out_frame[20] [6]), .O(n23939));
    defparam i10521_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i10523_3_lut_4_lut (.I0(\FRAME_MATCHER.state [2]), .I1(n22338), 
            .I2(displacement[4]), .I3(\data_out_frame[20] [4]), .O(n23941));
    defparam i10523_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i10524_3_lut_4_lut (.I0(\FRAME_MATCHER.state [2]), .I1(n22338), 
            .I2(displacement[3]), .I3(\data_out_frame[20] [3]), .O(n23942));
    defparam i10524_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i10529_3_lut_4_lut (.I0(\FRAME_MATCHER.state [2]), .I1(n22338), 
            .I2(displacement[14]), .I3(\data_out_frame[19] [6]), .O(n23947));
    defparam i10529_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i1_3_lut_4_lut_adj_1387 (.I0(n23290), .I1(n22842), .I2(Kp_23__N_326), 
            .I3(n40318), .O(n40758));
    defparam i1_3_lut_4_lut_adj_1387.LUT_INIT = 16'h9669;
    SB_LUT4 i10526_3_lut_4_lut (.I0(\FRAME_MATCHER.state [2]), .I1(n22338), 
            .I2(displacement[1]), .I3(\data_out_frame[20] [1]), .O(n23944));
    defparam i10526_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i10527_3_lut_4_lut (.I0(\FRAME_MATCHER.state [2]), .I1(n22338), 
            .I2(displacement[0]), .I3(\data_out_frame[20] [0]), .O(n23945));
    defparam i10527_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i10528_3_lut_4_lut (.I0(\FRAME_MATCHER.state [2]), .I1(n22338), 
            .I2(displacement[15]), .I3(\data_out_frame[19] [7]), .O(n23946));
    defparam i10528_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i10530_3_lut_4_lut (.I0(\FRAME_MATCHER.state [2]), .I1(n22338), 
            .I2(displacement[13]), .I3(\data_out_frame[19] [5]), .O(n23948));
    defparam i10530_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i10531_3_lut_4_lut (.I0(\FRAME_MATCHER.state [2]), .I1(n22338), 
            .I2(displacement[12]), .I3(\data_out_frame[19] [4]), .O(n23949));
    defparam i10531_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i10532_3_lut_4_lut (.I0(\FRAME_MATCHER.state [2]), .I1(n22338), 
            .I2(displacement[11]), .I3(\data_out_frame[19][3] ), .O(n23950));
    defparam i10532_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i10533_3_lut_4_lut (.I0(\FRAME_MATCHER.state [2]), .I1(n22338), 
            .I2(displacement[10]), .I3(\data_out_frame[19] [2]), .O(n23951));
    defparam i10533_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i10535_3_lut_4_lut (.I0(\FRAME_MATCHER.state [2]), .I1(n22338), 
            .I2(displacement[8]), .I3(\data_out_frame[19] [0]), .O(n23953));
    defparam i10535_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i2_3_lut_4_lut_adj_1388 (.I0(n23290), .I1(n22842), .I2(\data_in_frame[9] [4]), 
            .I3(\data_in_frame[14] [1]), .O(n40782));
    defparam i2_3_lut_4_lut_adj_1388.LUT_INIT = 16'h6996;
    SB_LUT4 i10536_3_lut_4_lut (.I0(\FRAME_MATCHER.state [2]), .I1(n22338), 
            .I2(displacement[23]), .I3(\data_out_frame[18] [7]), .O(n23954));
    defparam i10536_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i10537_3_lut_4_lut (.I0(\FRAME_MATCHER.state [2]), .I1(n22338), 
            .I2(displacement[22]), .I3(\data_out_frame[18] [6]), .O(n23955));
    defparam i10537_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i10538_3_lut_4_lut (.I0(\FRAME_MATCHER.state [2]), .I1(n22338), 
            .I2(displacement[21]), .I3(\data_out_frame[18] [5]), .O(n23956));
    defparam i10538_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i10539_3_lut_4_lut (.I0(\FRAME_MATCHER.state [2]), .I1(n22338), 
            .I2(displacement[20]), .I3(\data_out_frame[18] [4]), .O(n23957));
    defparam i10539_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_31377 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[14] [5]), .I2(\data_out_frame[15] [5]), 
            .I3(byte_transmit_counter[1]), .O(n46889));
    defparam byte_transmit_counter_0__bdd_4_lut_31377.LUT_INIT = 16'he4aa;
    SB_LUT4 i10540_3_lut_4_lut (.I0(\FRAME_MATCHER.state [2]), .I1(n22338), 
            .I2(displacement[19]), .I3(\data_out_frame[18][3] ), .O(n23958));
    defparam i10540_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i10541_3_lut_4_lut (.I0(\FRAME_MATCHER.state [2]), .I1(n22338), 
            .I2(displacement[18]), .I3(\data_out_frame[18] [2]), .O(n23959));
    defparam i10541_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i10542_3_lut_4_lut (.I0(\FRAME_MATCHER.state [2]), .I1(n22338), 
            .I2(displacement[17]), .I3(\data_out_frame[18] [1]), .O(n23960));
    defparam i10542_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i10543_3_lut_4_lut (.I0(\FRAME_MATCHER.state [2]), .I1(n22338), 
            .I2(displacement[16]), .I3(\data_out_frame[18] [0]), .O(n23961));
    defparam i10543_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i2_2_lut_3_lut_4_lut_adj_1389 (.I0(\data_in_frame[3] [0]), .I1(\data_in_frame[0] [7]), 
            .I2(\data_in_frame[0] [6]), .I3(\data_in_frame[1] [0]), .O(n6_adj_3130));   // verilog/coms.v(69[16:69])
    defparam i2_2_lut_3_lut_4_lut_adj_1389.LUT_INIT = 16'h6996;
    SB_LUT4 i26750_3_lut (.I0(\data_out_frame[8] [6]), .I1(\data_out_frame[9] [6]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n42269));
    defparam i26750_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i26751_3_lut (.I0(\data_out_frame[10] [6]), .I1(\data_out_frame[11] [6]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n42270));
    defparam i26751_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i26754_3_lut (.I0(\data_out_frame[14] [6]), .I1(\data_out_frame[15] [6]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n42273));
    defparam i26754_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10544_3_lut_4_lut (.I0(\FRAME_MATCHER.state [2]), .I1(n22338), 
            .I2(pwm[7]), .I3(\data_out_frame[17] [7]), .O(n23962));
    defparam i10544_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i26753_3_lut (.I0(\data_out_frame[12] [6]), .I1(\data_out_frame[13] [6]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n42272));
    defparam i26753_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10546_3_lut_4_lut (.I0(\FRAME_MATCHER.state [2]), .I1(n22338), 
            .I2(pwm[5]), .I3(\data_out_frame[17] [5]), .O(n23964));
    defparam i10546_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_4_i5_3_lut (.I0(\data_out_frame[6] [4]), 
            .I1(\data_out_frame[7] [4]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n5_adj_3142));   // verilog/coms.v(104[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_4_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i29056_2_lut (.I0(\data_out_frame[5] [4]), .I1(byte_transmit_counter[0]), 
            .I2(GND_net), .I3(GND_net), .O(n44143));
    defparam i29056_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_3_i16_3_lut (.I0(\data_out_frame[16] [3]), 
            .I1(\data_out_frame[17] [3]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n16_adj_3140));   // verilog/coms.v(104[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_3_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i29339_2_lut (.I0(\data_out_frame[22] [3]), .I1(byte_transmit_counter[0]), 
            .I2(GND_net), .I3(GND_net), .O(n44182));
    defparam i29339_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_3_i19_3_lut (.I0(\data_out_frame[20] [3]), 
            .I1(\data_out_frame[21] [3]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n19_adj_3139));   // verilog/coms.v(104[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_3_i19_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10547_3_lut_4_lut (.I0(\FRAME_MATCHER.state [2]), .I1(n22338), 
            .I2(pwm[4]), .I3(\data_out_frame[17] [4]), .O(n23965));
    defparam i10547_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i10549_3_lut_4_lut (.I0(\FRAME_MATCHER.state [2]), .I1(n22338), 
            .I2(pwm[2]), .I3(\data_out_frame[17] [2]), .O(n23967));
    defparam i10549_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 n46889_bdd_4_lut (.I0(n46889), .I1(\data_out_frame[13] [5]), 
            .I2(\data_out_frame[12] [5]), .I3(byte_transmit_counter[1]), 
            .O(n46892));
    defparam n46889_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i10550_3_lut_4_lut (.I0(\FRAME_MATCHER.state [2]), .I1(n22338), 
            .I2(pwm[1]), .I3(\data_out_frame[17] [1]), .O(n23968));
    defparam i10550_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i12051_3_lut_4_lut (.I0(\FRAME_MATCHER.state [2]), .I1(n22338), 
            .I2(pwm[0]), .I3(\data_out_frame[17] [0]), .O(n23969));
    defparam i12051_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i10552_3_lut_4_lut (.I0(\FRAME_MATCHER.state [2]), .I1(n22338), 
            .I2(pwm[15]), .I3(\data_out_frame[16] [7]), .O(n23970));
    defparam i10552_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i3_4_lut_adj_1390 (.I0(n37268), .I1(n41875), .I2(n40758), 
            .I3(n40834), .O(n40515));
    defparam i3_4_lut_adj_1390.LUT_INIT = 16'h6996;
    SB_LUT4 i10554_3_lut_4_lut (.I0(\FRAME_MATCHER.state [2]), .I1(n22338), 
            .I2(pwm[13]), .I3(\data_out_frame[16] [5]), .O(n23972));
    defparam i10554_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i10559_3_lut_4_lut (.I0(\FRAME_MATCHER.state [2]), .I1(n22338), 
            .I2(pwm[8]), .I3(\data_out_frame[16] [0]), .O(n23977));
    defparam i10559_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i10555_3_lut_4_lut (.I0(\FRAME_MATCHER.state [2]), .I1(n22338), 
            .I2(pwm[12]), .I3(\data_out_frame[16] [4]), .O(n23973));
    defparam i10555_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i10556_3_lut_4_lut (.I0(\FRAME_MATCHER.state [2]), .I1(n22338), 
            .I2(pwm[11]), .I3(\data_out_frame[16] [3]), .O(n23974));
    defparam i10556_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i10557_3_lut_4_lut (.I0(\FRAME_MATCHER.state [2]), .I1(n22338), 
            .I2(pwm[10]), .I3(\data_out_frame[16] [2]), .O(n23975));
    defparam i10557_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i10558_3_lut_4_lut (.I0(\FRAME_MATCHER.state [2]), .I1(n22338), 
            .I2(pwm[9]), .I3(\data_out_frame[16] [1]), .O(n23976));
    defparam i10558_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i10560_3_lut_4_lut (.I0(\FRAME_MATCHER.state [2]), .I1(n22338), 
            .I2(pwm[23]), .I3(\data_out_frame[15] [7]), .O(n23978));
    defparam i10560_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i10561_3_lut_4_lut (.I0(\FRAME_MATCHER.state [2]), .I1(n22338), 
            .I2(pwm[22]), .I3(\data_out_frame[15] [6]), .O(n23979));
    defparam i10561_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i10563_3_lut_4_lut (.I0(\FRAME_MATCHER.state [2]), .I1(n22338), 
            .I2(pwm[20]), .I3(\data_out_frame[15] [4]), .O(n23981));
    defparam i10563_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i10564_3_lut_4_lut (.I0(\FRAME_MATCHER.state [2]), .I1(n22338), 
            .I2(pwm[19]), .I3(\data_out_frame[15] [3]), .O(n23982));
    defparam i10564_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i10565_3_lut_4_lut (.I0(\FRAME_MATCHER.state [2]), .I1(n22338), 
            .I2(pwm[18]), .I3(\data_out_frame[15] [2]), .O(n23983));
    defparam i10565_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i14741_2_lut_4_lut (.I0(n27691), .I1(Kp_23__N_152), .I2(n31_adj_3306), 
            .I3(\FRAME_MATCHER.state [1]), .O(n28145));
    defparam i14741_2_lut_4_lut.LUT_INIT = 16'hfabb;
    SB_LUT4 i10566_3_lut_4_lut (.I0(\FRAME_MATCHER.state [2]), .I1(n22338), 
            .I2(pwm[17]), .I3(\data_out_frame[15] [1]), .O(n23984));
    defparam i10566_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i10567_3_lut_4_lut (.I0(\FRAME_MATCHER.state [2]), .I1(n22338), 
            .I2(pwm[16]), .I3(\data_out_frame[15] [0]), .O(n23985));
    defparam i10567_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i10568_3_lut_4_lut (.I0(\FRAME_MATCHER.state [2]), .I1(n22338), 
            .I2(setpoint[7]), .I3(\data_out_frame[14] [7]), .O(n23986));
    defparam i10568_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i10481_3_lut_4_lut (.I0(n8), .I1(n40212), .I2(rx_data[7]), 
            .I3(\data_in_frame[4] [7]), .O(n23899));
    defparam i10481_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10569_3_lut_4_lut (.I0(\FRAME_MATCHER.state [2]), .I1(n22338), 
            .I2(setpoint[6]), .I3(\data_out_frame[14] [6]), .O(n23987));
    defparam i10569_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i10570_3_lut_4_lut (.I0(\FRAME_MATCHER.state [2]), .I1(n22338), 
            .I2(setpoint[5]), .I3(\data_out_frame[14] [5]), .O(n23988));
    defparam i10570_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i10571_3_lut_4_lut (.I0(\FRAME_MATCHER.state [2]), .I1(n22338), 
            .I2(setpoint[4]), .I3(\data_out_frame[14] [4]), .O(n23989));
    defparam i10571_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i10572_3_lut_4_lut (.I0(\FRAME_MATCHER.state [2]), .I1(n22338), 
            .I2(setpoint[3]), .I3(\data_out_frame[14] [3]), .O(n23990));
    defparam i10572_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i10482_3_lut_4_lut (.I0(n8), .I1(n40212), .I2(rx_data[6]), 
            .I3(\data_in_frame[4] [6]), .O(n23900));
    defparam i10482_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10573_3_lut_4_lut (.I0(\FRAME_MATCHER.state [2]), .I1(n22338), 
            .I2(setpoint[2]), .I3(\data_out_frame[14] [2]), .O(n23991));
    defparam i10573_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i10574_3_lut_4_lut (.I0(\FRAME_MATCHER.state [2]), .I1(n22338), 
            .I2(setpoint[1]), .I3(\data_out_frame[14] [1]), .O(n23992));
    defparam i10574_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i10575_3_lut_4_lut (.I0(\FRAME_MATCHER.state [2]), .I1(n22338), 
            .I2(setpoint[0]), .I3(\data_out_frame[14] [0]), .O(n23993));
    defparam i10575_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i10576_3_lut_4_lut (.I0(\FRAME_MATCHER.state [2]), .I1(n22338), 
            .I2(setpoint[15]), .I3(\data_out_frame[13] [7]), .O(n23994));
    defparam i10576_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i10483_3_lut_4_lut (.I0(n8), .I1(n40212), .I2(rx_data[5]), 
            .I3(\data_in_frame[4] [5]), .O(n23901));
    defparam i10483_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10628_3_lut_4_lut (.I0(\FRAME_MATCHER.state [2]), .I1(n22338), 
            .I2(encoder0_position[11]), .I3(\data_out_frame[7] [3]), .O(n24046));
    defparam i10628_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i10577_3_lut_4_lut (.I0(\FRAME_MATCHER.state [2]), .I1(n22338), 
            .I2(setpoint[14]), .I3(\data_out_frame[13] [6]), .O(n23995));
    defparam i10577_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i10578_3_lut_4_lut (.I0(\FRAME_MATCHER.state [2]), .I1(n22338), 
            .I2(setpoint[13]), .I3(\data_out_frame[13] [5]), .O(n23996));
    defparam i10578_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i2_3_lut_4_lut_adj_1391 (.I0(\data_in_frame[21] [0]), .I1(Kp_23__N_786), 
            .I2(n23301), .I3(n37284), .O(n41462));
    defparam i2_3_lut_4_lut_adj_1391.LUT_INIT = 16'h6996;
    SB_LUT4 i10579_3_lut_4_lut (.I0(\FRAME_MATCHER.state [2]), .I1(n22338), 
            .I2(setpoint[12]), .I3(\data_out_frame[13] [4]), .O(n23997));
    defparam i10579_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i10580_3_lut_4_lut (.I0(\FRAME_MATCHER.state [2]), .I1(n22338), 
            .I2(setpoint[11]), .I3(\data_out_frame[13] [3]), .O(n23998));
    defparam i10580_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i10581_3_lut_4_lut (.I0(\FRAME_MATCHER.state [2]), .I1(n22338), 
            .I2(setpoint[10]), .I3(\data_out_frame[13] [2]), .O(n23999));
    defparam i10581_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i10582_3_lut_4_lut (.I0(\FRAME_MATCHER.state [2]), .I1(n22338), 
            .I2(setpoint[9]), .I3(\data_out_frame[13] [1]), .O(n24000));
    defparam i10582_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i10484_3_lut_4_lut (.I0(n8), .I1(n40212), .I2(rx_data[4]), 
            .I3(\data_in_frame[4] [4]), .O(n23902));
    defparam i10484_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10583_3_lut_4_lut (.I0(\FRAME_MATCHER.state [2]), .I1(n22338), 
            .I2(setpoint[8]), .I3(\data_out_frame[13] [0]), .O(n24001));
    defparam i10583_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i10584_3_lut_4_lut (.I0(\FRAME_MATCHER.state [2]), .I1(n22338), 
            .I2(setpoint[23]), .I3(\data_out_frame[12] [7]), .O(n24002));
    defparam i10584_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i10485_3_lut_4_lut (.I0(n8), .I1(n40212), .I2(rx_data[3]), 
            .I3(\data_in_frame[4] [3]), .O(n23903));
    defparam i10485_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10585_3_lut_4_lut (.I0(\FRAME_MATCHER.state [2]), .I1(n22338), 
            .I2(setpoint[22]), .I3(\data_out_frame[12] [6]), .O(n24003));
    defparam i10585_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i10486_3_lut_4_lut (.I0(n8), .I1(n40212), .I2(rx_data[2]), 
            .I3(\data_in_frame[4] [2]), .O(n23904));
    defparam i10486_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10586_3_lut_4_lut (.I0(\FRAME_MATCHER.state [2]), .I1(n22338), 
            .I2(setpoint[21]), .I3(\data_out_frame[12] [5]), .O(n24004));
    defparam i10586_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i10587_3_lut_4_lut (.I0(\FRAME_MATCHER.state [2]), .I1(n22338), 
            .I2(setpoint[20]), .I3(\data_out_frame[12] [4]), .O(n24005));
    defparam i10587_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i10487_3_lut_4_lut (.I0(n8), .I1(n40212), .I2(rx_data[1]), 
            .I3(\data_in_frame[4] [1]), .O(n23905));
    defparam i10487_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10588_3_lut_4_lut (.I0(\FRAME_MATCHER.state [2]), .I1(n22338), 
            .I2(setpoint[19]), .I3(\data_out_frame[12] [3]), .O(n24006));
    defparam i10588_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i10488_3_lut_4_lut (.I0(n8), .I1(n40212), .I2(rx_data[0]), 
            .I3(\data_in_frame[4] [0]), .O(n23906));
    defparam i10488_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10605_3_lut_4_lut (.I0(\FRAME_MATCHER.state [2]), .I1(n22338), 
            .I2(encoder1_position[10]), .I3(\data_out_frame[10] [2]), .O(n24023));
    defparam i10605_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i10641_3_lut_4_lut (.I0(\FRAME_MATCHER.state [2]), .I1(n22338), 
            .I2(control_mode[6]), .I3(\data_out_frame[5] [6]), .O(n24059));
    defparam i10641_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i6_3_lut_4_lut (.I0(\data_in_frame[0] [5]), .I1(\data_in_frame[0] [7]), 
            .I2(\data_in_frame[0] [4]), .I3(\data_in_frame[0] [6]), .O(n14_adj_3144));   // verilog/coms.v(232[13:35])
    defparam i6_3_lut_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_3_lut_adj_1392 (.I0(\data_in_frame[16] [6]), .I1(n22648), 
            .I2(n40752), .I3(GND_net), .O(n40258));
    defparam i1_2_lut_3_lut_adj_1392.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1393 (.I0(\data_in_frame[0] [4]), .I1(\data_in_frame[0] [5]), 
            .I2(\data_in_frame[2] [6]), .I3(GND_net), .O(n4_c));   // verilog/coms.v(74[16:27])
    defparam i1_2_lut_3_lut_adj_1393.LUT_INIT = 16'h9696;
    SB_LUT4 i3_2_lut_4_lut (.I0(\data_in_frame[3] [2]), .I1(\data_in_frame[3] [3]), 
            .I2(\data_in_frame[0] [7]), .I3(\data_in_frame[3] [1]), .O(n9_adj_3134));   // verilog/coms.v(71[16:34])
    defparam i3_2_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_adj_1394 (.I0(\data_in_frame[1] [2]), .I1(\data_in_frame[1] [4]), 
            .I2(\data_in_frame[3] [5]), .I3(\data_in_frame[3] [4]), .O(Kp_23__N_459));   // verilog/coms.v(74[16:43])
    defparam i1_2_lut_4_lut_adj_1394.LUT_INIT = 16'h6996;
    SB_LUT4 i2_2_lut_4_lut_adj_1395 (.I0(\data_in_frame[7] [6]), .I1(\data_in_frame[7] [7]), 
            .I2(n40773), .I3(\data_in_frame[6][1] ), .O(n10_adj_3129));
    defparam i2_2_lut_4_lut_adj_1395.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_adj_1396 (.I0(\data_in_frame[14] [4]), .I1(\data_in_frame[9] [6]), 
            .I2(\data_in_frame[12] [2]), .I3(Kp_23__N_459), .O(n40584));
    defparam i1_2_lut_4_lut_adj_1396.LUT_INIT = 16'h6996;
    SB_LUT4 i10639_3_lut_4_lut (.I0(\FRAME_MATCHER.state [2]), .I1(n22338), 
            .I2(encoder0_position[16]), .I3(\data_out_frame[6] [0]), .O(n24057));
    defparam i10639_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i1_2_lut_3_lut_adj_1397 (.I0(\data_in_frame[7] [6]), .I1(\data_in_frame[7] [7]), 
            .I2(n40773), .I3(GND_net), .O(n40466));
    defparam i1_2_lut_3_lut_adj_1397.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_4_lut_adj_1398 (.I0(Kp_23__N_379), .I1(\data_in_frame[5] [7]), 
            .I2(\data_in_frame[10] [2]), .I3(\data_in_frame[6][0] ), .O(n40773));
    defparam i2_3_lut_4_lut_adj_1398.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1399 (.I0(\data_in_frame[5] [6]), .I1(\data_in_frame[7] [6]), 
            .I2(\data_in_frame[7] [7]), .I3(GND_net), .O(n40417));   // verilog/coms.v(83[17:28])
    defparam i1_2_lut_3_lut_adj_1399.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_4_lut_adj_1400 (.I0(n37255), .I1(\data_out_frame[17] [5]), 
            .I2(n1787), .I3(n36597), .O(n36494));
    defparam i2_3_lut_4_lut_adj_1400.LUT_INIT = 16'h6996;
    SB_LUT4 i10637_3_lut_4_lut (.I0(\FRAME_MATCHER.state [2]), .I1(n22338), 
            .I2(encoder0_position[18]), .I3(\data_out_frame[6] [2]), .O(n24055));
    defparam i10637_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i14341_2_lut (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(GND_net), .I3(GND_net), .O(n27743));
    defparam i14341_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1401 (.I0(\data_in_frame[6] [5]), .I1(\data_in_frame[6] [4]), 
            .I2(\data_in_frame[10] [6]), .I3(\data_in_frame[13] [2]), .O(n40650));   // verilog/coms.v(72[16:43])
    defparam i1_2_lut_3_lut_4_lut_adj_1401.LUT_INIT = 16'h6996;
    SB_LUT4 i10553_3_lut_4_lut (.I0(\FRAME_MATCHER.state [2]), .I1(n22338), 
            .I2(pwm[14]), .I3(\data_out_frame[16] [6]), .O(n23971));
    defparam i10553_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i10548_3_lut_4_lut (.I0(\FRAME_MATCHER.state [2]), .I1(n22338), 
            .I2(pwm[3]), .I3(\data_out_frame[17] [3]), .O(n23966));
    defparam i10548_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i10630_3_lut_4_lut (.I0(\FRAME_MATCHER.state [2]), .I1(n22338), 
            .I2(encoder0_position[9]), .I3(\data_out_frame[7] [1]), .O(n24048));
    defparam i10630_3_lut_4_lut.LUT_INIT = 16'hfb40;
    uart_tx tx (.n313(n313), .r_Clock_Count({\r_Clock_Count[8] , \r_Clock_Count[7] , 
            \r_Clock_Count[6] , \r_Clock_Count[5] , \r_Clock_Count[4] , 
            \r_Clock_Count[3] , \r_Clock_Count[2] , \r_Clock_Count[1] , 
            Open_6}), .GND_net(GND_net), .n314(n314), .n23624(n23624), 
            .clk32MHz(clk32MHz), .n23627(n23627), .n23630(n23630), .n23633(n23633), 
            .n23636(n23636), .n23639(n23639), .n23642(n23642), .n23645(n23645), 
            .n23649(n23649), .r_Bit_Index({r_Bit_Index}), .n23652(n23652), 
            .n23695(n23695), .tx_data({tx_data}), .n315(n315), .n316(n316), 
            .n317(n317), .n318(n318), .n319(n319), .n320(n320), .VCC_net(VCC_net), 
            .n23644(n23644), .\r_SM_Main[2] (\r_SM_Main[2] ), .tx_active(tx_active), 
            .tx_o(tx_o), .byte_transmit_counter({byte_transmit_counter_c[7:2], 
            byte_transmit_counter[1:0]}), .n44012(n44012), .n23400(n23400), 
            .n24177(n24177), .\r_SM_Main_2__N_2756[0] (r_SM_Main_2__N_2756[0]), 
            .tx_enable(tx_enable), .n23477(n23477), .n23562(n23562), .n4034(n4034), 
            .n19614(n19614), .n2238(n2236[6]), .n24178(n24178), .n2239(n2236[5]), 
            .n23680(n23680), .n2240(n2236[4]), .n23677(n23677), .n28265(n28265), 
            .n28275(n28275), .n2241(n2236[3]), .n23674(n23674), .n2242(n2236[2]), 
            .n23671(n23671), .n2243(n2236[1]), .n23668(n23668), .n2244(n2236[0]), 
            .n24234(n24234), .n31(n31_adj_3306), .n27691(n27691), .tx_transmit_N_2648(tx_transmit_N_2648), 
            .\FRAME_MATCHER.state[0] (\FRAME_MATCHER.state [0]), .n28285(n28285)) /* synthesis lattice_noprune=1, syn_preserve=0, syn_module_defined=1, syn_noprune=0 */ ;   // verilog/coms.v(105[10:70])
    uart_rx rx (.GND_net(GND_net), .r_Rx_Data(r_Rx_Data), .\r_SM_Main[2] (\r_SM_Main[2]_adj_3 ), 
            .\r_SM_Main[1] (\r_SM_Main[1] ), .clk32MHz(clk32MHz), .n23655(n23655), 
            .r_Bit_Index({r_Bit_Index_adj_9}), .n23658(n23658), .n28263(n28263), 
            .n23698(n23698), .n24171(n24171), .rx_data({rx_data}), .PIN_13_N_26(PIN_13_N_26), 
            .VCC_net(VCC_net), .rx_data_ready(rx_data_ready), .n23665(n23665), 
            .n23664(n23664), .n23663(n23663), .n23662(n23662), .n23661(n23661), 
            .n23660(n23660), .n23659(n23659), .n23594(n23594), .n22466(n22466), 
            .n4(n4), .n28231(n28231), .n1(n1), .n27725(n27725), .n4_adj_1(n4_adj_7), 
            .n4_adj_2(n4_adj_8), .n22471(n22471), .n44134(n44134), .n44133(n44133), 
            .n23471(n23471), .n23560(n23560), .n4012(n4012)) /* synthesis lattice_noprune=1, syn_preserve=0, syn_module_defined=1, syn_noprune=0 */ ;   // verilog/coms.v(91[10:44])
    
endmodule
//
// Verilog Description of module uart_tx
//

module uart_tx (n313, r_Clock_Count, GND_net, n314, n23624, clk32MHz, 
            n23627, n23630, n23633, n23636, n23639, n23642, n23645, 
            n23649, r_Bit_Index, n23652, n23695, tx_data, n315, 
            n316, n317, n318, n319, n320, VCC_net, n23644, \r_SM_Main[2] , 
            tx_active, tx_o, byte_transmit_counter, n44012, n23400, 
            n24177, \r_SM_Main_2__N_2756[0] , tx_enable, n23477, n23562, 
            n4034, n19614, n2238, n24178, n2239, n23680, n2240, 
            n23677, n28265, n28275, n2241, n23674, n2242, n23671, 
            n2243, n23668, n2244, n24234, n31, n27691, tx_transmit_N_2648, 
            \FRAME_MATCHER.state[0] , n28285) /* synthesis lattice_noprune=1, syn_preserve=0, syn_module_defined=1, syn_noprune=0 */ ;
    output n313;
    output [8:0]r_Clock_Count;
    input GND_net;
    output n314;
    input n23624;
    input clk32MHz;
    input n23627;
    input n23630;
    input n23633;
    input n23636;
    input n23639;
    input n23642;
    input n23645;
    input n23649;
    output [2:0]r_Bit_Index;
    input n23652;
    input n23695;
    input [7:0]tx_data;
    output n315;
    output n316;
    output n317;
    output n318;
    output n319;
    output n320;
    input VCC_net;
    output n23644;
    output \r_SM_Main[2] ;
    output tx_active;
    output tx_o;
    input [7:0]byte_transmit_counter;
    input n44012;
    input n23400;
    output n24177;
    input \r_SM_Main_2__N_2756[0] ;
    output tx_enable;
    output n23477;
    output n23562;
    output n4034;
    input n19614;
    input n2238;
    output n24178;
    input n2239;
    output n23680;
    input n2240;
    output n23677;
    input n28265;
    output n28275;
    input n2241;
    output n23674;
    input n2242;
    output n23671;
    input n2243;
    output n23668;
    input n2244;
    output n24234;
    input n31;
    input n27691;
    input tx_transmit_N_2648;
    input \FRAME_MATCHER.state[0] ;
    output n28285;
    
    wire clk32MHz /* synthesis SET_AS_NETWORK=clk32MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(34[8:16])
    
    wire n34076, n34075, n39986;
    wire [2:0]r_SM_Main;   // verilog/uart_tx.v(31[16:25])
    
    wire n39902;
    wire [8:0]r_Clock_Count_c;   // verilog/uart_tx.v(32[16:29])
    
    wire n19942;
    wire [7:0]r_Tx_Data;   // verilog/uart_tx.v(34[16:25])
    
    wire n34074, n34073, n34072, n34071, n34070, n34069, n44181, 
        n42287, n42288, n46925, n42219, n42218, o_Tx_Serial_N_2784, 
        n41171, n23598, n23597, n10, n12, n16856, n108, n23425, 
        n27837;
    wire [2:0]r_SM_Main_2__N_2753;
    
    wire n49, n115, n10_adj_3117, n53, n10_adj_3118, n9;
    
    SB_LUT4 add_59_10_lut (.I0(GND_net), .I1(r_Clock_Count[8]), .I2(GND_net), 
            .I3(n34076), .O(n313)) /* synthesis syn_instantiated=1 */ ;
    defparam add_59_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_59_9_lut (.I0(GND_net), .I1(r_Clock_Count[7]), .I2(GND_net), 
            .I3(n34075), .O(n314)) /* synthesis syn_instantiated=1 */ ;
    defparam add_59_9_lut.LUT_INIT = 16'hC33C;
    SB_DFF r_Clock_Count__i8 (.Q(r_Clock_Count[8]), .C(clk32MHz), .D(n23624));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFF r_Clock_Count__i7 (.Q(r_Clock_Count[7]), .C(clk32MHz), .D(n23627));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFF r_Clock_Count__i6 (.Q(r_Clock_Count[6]), .C(clk32MHz), .D(n23630));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFF r_Clock_Count__i5 (.Q(r_Clock_Count[5]), .C(clk32MHz), .D(n23633));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFF r_Clock_Count__i4 (.Q(r_Clock_Count[4]), .C(clk32MHz), .D(n23636));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFF r_Clock_Count__i3 (.Q(r_Clock_Count[3]), .C(clk32MHz), .D(n23639));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFF r_Clock_Count__i2 (.Q(r_Clock_Count[2]), .C(clk32MHz), .D(n23642));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFF r_Clock_Count__i1 (.Q(r_Clock_Count[1]), .C(clk32MHz), .D(n23645));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFF r_Bit_Index_i2 (.Q(r_Bit_Index[2]), .C(clk32MHz), .D(n23649));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFF r_Bit_Index_i1 (.Q(r_Bit_Index[1]), .C(clk32MHz), .D(n23652));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFF r_SM_Main_i1 (.Q(r_SM_Main[1]), .C(clk32MHz), .D(n39986));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFF r_Clock_Count__i0 (.Q(r_Clock_Count_c[0]), .C(clk32MHz), .D(n39902));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFF r_Bit_Index_i0 (.Q(r_Bit_Index[0]), .C(clk32MHz), .D(n23695));   // verilog/uart_tx.v(40[10] 143[8])
    SB_CARRY add_59_9 (.CI(n34075), .I0(r_Clock_Count[7]), .I1(GND_net), 
            .CO(n34076));
    SB_DFFE r_Tx_Data_i0 (.Q(r_Tx_Data[0]), .C(clk32MHz), .E(n19942), 
            .D(tx_data[0]));   // verilog/uart_tx.v(40[10] 143[8])
    SB_LUT4 add_59_8_lut (.I0(GND_net), .I1(r_Clock_Count[6]), .I2(GND_net), 
            .I3(n34074), .O(n315)) /* synthesis syn_instantiated=1 */ ;
    defparam add_59_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_59_8 (.CI(n34074), .I0(r_Clock_Count[6]), .I1(GND_net), 
            .CO(n34075));
    SB_LUT4 add_59_7_lut (.I0(GND_net), .I1(r_Clock_Count[5]), .I2(GND_net), 
            .I3(n34073), .O(n316)) /* synthesis syn_instantiated=1 */ ;
    defparam add_59_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_59_7 (.CI(n34073), .I0(r_Clock_Count[5]), .I1(GND_net), 
            .CO(n34074));
    SB_LUT4 add_59_6_lut (.I0(GND_net), .I1(r_Clock_Count[4]), .I2(GND_net), 
            .I3(n34072), .O(n317)) /* synthesis syn_instantiated=1 */ ;
    defparam add_59_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_59_6 (.CI(n34072), .I0(r_Clock_Count[4]), .I1(GND_net), 
            .CO(n34073));
    SB_LUT4 add_59_5_lut (.I0(GND_net), .I1(r_Clock_Count[3]), .I2(GND_net), 
            .I3(n34071), .O(n318)) /* synthesis syn_instantiated=1 */ ;
    defparam add_59_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_59_5 (.CI(n34071), .I0(r_Clock_Count[3]), .I1(GND_net), 
            .CO(n34072));
    SB_LUT4 add_59_4_lut (.I0(GND_net), .I1(r_Clock_Count[2]), .I2(GND_net), 
            .I3(n34070), .O(n319)) /* synthesis syn_instantiated=1 */ ;
    defparam add_59_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_59_4 (.CI(n34070), .I0(r_Clock_Count[2]), .I1(GND_net), 
            .CO(n34071));
    SB_LUT4 add_59_3_lut (.I0(GND_net), .I1(r_Clock_Count[1]), .I2(GND_net), 
            .I3(n34069), .O(n320)) /* synthesis syn_instantiated=1 */ ;
    defparam add_59_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_59_3 (.CI(n34069), .I0(r_Clock_Count[1]), .I1(GND_net), 
            .CO(n34070));
    SB_LUT4 add_59_2_lut (.I0(n23644), .I1(r_Clock_Count_c[0]), .I2(GND_net), 
            .I3(VCC_net), .O(n44181)) /* synthesis syn_instantiated=1 */ ;
    defparam add_59_2_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_59_2 (.CI(VCC_net), .I0(r_Clock_Count_c[0]), .I1(GND_net), 
            .CO(n34069));
    SB_LUT4 r_Bit_Index_1__bdd_4_lut (.I0(r_Bit_Index[1]), .I1(n42287), 
            .I2(n42288), .I3(r_Bit_Index[2]), .O(n46925));
    defparam r_Bit_Index_1__bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_LUT4 n46925_bdd_4_lut (.I0(n46925), .I1(n42219), .I2(n42218), .I3(r_Bit_Index[2]), 
            .O(o_Tx_Serial_N_2784));
    defparam n46925_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFFE r_Tx_Data_i1 (.Q(r_Tx_Data[1]), .C(clk32MHz), .E(n19942), 
            .D(tx_data[1]));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFE r_Tx_Data_i2 (.Q(r_Tx_Data[2]), .C(clk32MHz), .E(n19942), 
            .D(tx_data[2]));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFE r_Tx_Data_i3 (.Q(r_Tx_Data[3]), .C(clk32MHz), .E(n19942), 
            .D(tx_data[3]));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFE r_Tx_Data_i4 (.Q(r_Tx_Data[4]), .C(clk32MHz), .E(n19942), 
            .D(tx_data[4]));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFE r_Tx_Data_i5 (.Q(r_Tx_Data[5]), .C(clk32MHz), .E(n19942), 
            .D(tx_data[5]));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFE r_Tx_Data_i6 (.Q(r_Tx_Data[6]), .C(clk32MHz), .E(n19942), 
            .D(tx_data[6]));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFE r_Tx_Data_i7 (.Q(r_Tx_Data[7]), .C(clk32MHz), .E(n19942), 
            .D(tx_data[7]));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFF r_SM_Main_i2 (.Q(\r_SM_Main[2] ), .C(clk32MHz), .D(n41171));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFF r_SM_Main_i0 (.Q(r_SM_Main[0]), .C(clk32MHz), .D(n23598));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFF r_Tx_Active_47 (.Q(tx_active), .C(clk32MHz), .D(n23597));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFF o_Tx_Serial_45 (.Q(tx_o), .C(clk32MHz), .D(n10));   // verilog/uart_tx.v(40[10] 143[8])
    SB_LUT4 i25_3_lut (.I0(r_Clock_Count_c[0]), .I1(n44181), .I2(\r_SM_Main[2] ), 
            .I3(GND_net), .O(n39902));
    defparam i25_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i11706_3_lut (.I0(byte_transmit_counter[7]), .I1(n44012), .I2(n23400), 
            .I3(GND_net), .O(n24177));
    defparam i11706_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i26_3_lut (.I0(r_SM_Main[0]), .I1(o_Tx_Serial_N_2784), .I2(r_SM_Main[1]), 
            .I3(GND_net), .O(n12));
    defparam i26_3_lut.LUT_INIT = 16'h1a1a;
    SB_LUT4 i25_3_lut_adj_829 (.I0(n12), .I1(tx_o), .I2(\r_SM_Main[2] ), 
            .I3(GND_net), .O(n10));
    defparam i25_3_lut_adj_829.LUT_INIT = 16'hc5c5;
    SB_LUT4 i1_2_lut (.I0(r_SM_Main[0]), .I1(\r_SM_Main_2__N_2756[0] ), 
            .I2(GND_net), .I3(GND_net), .O(n16856));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i1_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i2_4_lut (.I0(n16856), .I1(\r_SM_Main[2] ), .I2(r_SM_Main[1]), 
            .I3(n108), .O(n23425));
    defparam i2_4_lut.LUT_INIT = 16'h3202;
    SB_LUT4 i12286_3_lut (.I0(n23425), .I1(r_SM_Main[1]), .I2(tx_active), 
            .I3(GND_net), .O(n23597));   // verilog/uart_tx.v(31[16:25])
    defparam i12286_3_lut.LUT_INIT = 16'h7272;
    SB_LUT4 i47_4_lut (.I0(\r_SM_Main_2__N_2756[0] ), .I1(n27837), .I2(r_SM_Main[1]), 
            .I3(r_SM_Main_2__N_2753[1]), .O(n49));   // verilog/uart_tx.v(31[16:25])
    defparam i47_4_lut.LUT_INIT = 16'hca0a;
    SB_LUT4 i1_4_lut (.I0(\r_SM_Main[2] ), .I1(n49), .I2(r_SM_Main_2__N_2753[1]), 
            .I3(r_SM_Main[0]), .O(n23598));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i1_4_lut.LUT_INIT = 16'h0544;
    SB_LUT4 i26699_3_lut (.I0(r_Tx_Data[0]), .I1(r_Tx_Data[1]), .I2(r_Bit_Index[0]), 
            .I3(GND_net), .O(n42218));
    defparam i26699_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i26700_3_lut (.I0(r_Tx_Data[2]), .I1(r_Tx_Data[3]), .I2(r_Bit_Index[0]), 
            .I3(GND_net), .O(n42219));
    defparam i26700_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i26769_3_lut (.I0(r_Tx_Data[6]), .I1(r_Tx_Data[7]), .I2(r_Bit_Index[0]), 
            .I3(GND_net), .O(n42288));
    defparam i26769_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i26768_3_lut (.I0(r_Tx_Data[4]), .I1(r_Tx_Data[5]), .I2(r_Bit_Index[0]), 
            .I3(GND_net), .O(n42287));
    defparam i26768_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 o_Tx_Serial_I_0_1_lut (.I0(tx_o), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(tx_enable));   // verilog/uart_tx.v(38[24:36])
    defparam o_Tx_Serial_I_0_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1_2_lut_adj_830 (.I0(r_SM_Main[0]), .I1(r_SM_Main_2__N_2753[1]), 
            .I2(GND_net), .I3(GND_net), .O(n108));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i1_2_lut_adj_830.LUT_INIT = 16'h8888;
    SB_LUT4 i2_3_lut (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[2]), .I2(r_Bit_Index[0]), 
            .I3(GND_net), .O(n27837));
    defparam i2_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 i4_4_lut (.I0(n115), .I1(r_Clock_Count[4]), .I2(r_Clock_Count[8]), 
            .I3(r_Clock_Count[5]), .O(n10_adj_3117));   // verilog/uart_tx.v(32[16:29])
    defparam i4_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i5_3_lut (.I0(r_Clock_Count[7]), .I1(n10_adj_3117), .I2(r_Clock_Count[6]), 
            .I3(GND_net), .O(r_SM_Main_2__N_2753[1]));   // verilog/uart_tx.v(32[16:29])
    defparam i5_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i2_4_lut_adj_831 (.I0(r_SM_Main[0]), .I1(\r_SM_Main[2] ), .I2(r_SM_Main[1]), 
            .I3(r_SM_Main_2__N_2753[1]), .O(n23477));
    defparam i2_4_lut_adj_831.LUT_INIT = 16'h1101;
    SB_LUT4 i10144_3_lut (.I0(n23477), .I1(r_SM_Main[1]), .I2(n27837), 
            .I3(GND_net), .O(n23562));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i10144_3_lut.LUT_INIT = 16'ha2a2;
    SB_LUT4 i1094_2_lut (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[0]), .I2(GND_net), 
            .I3(GND_net), .O(n4034));   // verilog/uart_tx.v(98[36:51])
    defparam i1094_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_832 (.I0(r_SM_Main[1]), .I1(r_SM_Main[0]), .I2(GND_net), 
            .I3(GND_net), .O(n53));   // verilog/uart_tx.v(31[16:25])
    defparam i1_2_lut_adj_832.LUT_INIT = 16'heeee;
    SB_LUT4 i3_4_lut (.I0(r_Clock_Count[2]), .I1(r_Clock_Count_c[0]), .I2(r_Clock_Count[3]), 
            .I3(r_Clock_Count[1]), .O(n115));   // verilog/uart_tx.v(32[16:29])
    defparam i3_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i4_4_lut_adj_833 (.I0(r_Clock_Count[5]), .I1(r_Clock_Count[7]), 
            .I2(n115), .I3(r_Clock_Count[8]), .O(n10_adj_3118));
    defparam i4_4_lut_adj_833.LUT_INIT = 16'hfffe;
    SB_LUT4 i3_2_lut (.I0(r_Clock_Count[4]), .I1(r_Clock_Count[6]), .I2(GND_net), 
            .I3(GND_net), .O(n9));
    defparam i3_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i1_4_lut_adj_834 (.I0(\r_SM_Main[2] ), .I1(n9), .I2(n53), 
            .I3(n10_adj_3118), .O(n23644));   // verilog/uart_tx.v(31[16:25])
    defparam i1_4_lut_adj_834.LUT_INIT = 16'haaba;
    SB_LUT4 i1_4_lut_4_lut (.I0(n23400), .I1(n19614), .I2(n2238), .I3(byte_transmit_counter[6]), 
            .O(n24178));
    defparam i1_4_lut_4_lut.LUT_INIT = 16'hd580;
    SB_LUT4 i10262_4_lut_4_lut (.I0(n23400), .I1(n19614), .I2(n2239), 
            .I3(byte_transmit_counter[5]), .O(n23680));
    defparam i10262_4_lut_4_lut.LUT_INIT = 16'hd580;
    SB_LUT4 i1_4_lut_4_lut_adj_835 (.I0(n23400), .I1(n19614), .I2(n2240), 
            .I3(byte_transmit_counter[4]), .O(n23677));
    defparam i1_4_lut_4_lut_adj_835.LUT_INIT = 16'hd580;
    SB_LUT4 i3_4_lut_adj_836 (.I0(byte_transmit_counter[6]), .I1(n28265), 
            .I2(byte_transmit_counter[5]), .I3(byte_transmit_counter[7]), 
            .O(n28275));
    defparam i3_4_lut_adj_836.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_4_lut_adj_837 (.I0(n23400), .I1(n19614), .I2(n2241), 
            .I3(byte_transmit_counter[3]), .O(n23674));
    defparam i1_4_lut_4_lut_adj_837.LUT_INIT = 16'hd580;
    SB_LUT4 i1_4_lut_4_lut_adj_838 (.I0(n23400), .I1(n19614), .I2(n2242), 
            .I3(byte_transmit_counter[2]), .O(n23671));
    defparam i1_4_lut_4_lut_adj_838.LUT_INIT = 16'hd580;
    SB_LUT4 i10250_4_lut_4_lut (.I0(n23400), .I1(n19614), .I2(n2243), 
            .I3(byte_transmit_counter[1]), .O(n23668));
    defparam i10250_4_lut_4_lut.LUT_INIT = 16'hd580;
    SB_LUT4 i10816_4_lut_4_lut (.I0(n23400), .I1(n19614), .I2(n2244), 
            .I3(byte_transmit_counter[0]), .O(n24234));
    defparam i10816_4_lut_4_lut.LUT_INIT = 16'hd580;
    SB_LUT4 i1_3_lut_4_lut (.I0(\r_SM_Main[2] ), .I1(r_SM_Main[0]), .I2(r_SM_Main_2__N_2753[1]), 
            .I3(r_SM_Main[1]), .O(n39986));   // verilog/uart_tx.v(31[16:25])
    defparam i1_3_lut_4_lut.LUT_INIT = 16'h1540;
    SB_LUT4 i11695_3_lut_4_lut (.I0(n31), .I1(n27691), .I2(tx_transmit_N_2648), 
            .I3(\FRAME_MATCHER.state[0] ), .O(n28285));   // verilog/coms.v(110[11:16])
    defparam i11695_3_lut_4_lut.LUT_INIT = 16'h0fee;
    SB_LUT4 i2_3_lut_4_lut (.I0(r_SM_Main[0]), .I1(r_SM_Main_2__N_2753[1]), 
            .I2(r_SM_Main[1]), .I3(\r_SM_Main[2] ), .O(n41171));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i2_3_lut_4_lut.LUT_INIT = 16'h0080;
    SB_LUT4 i2_3_lut_4_lut_adj_839 (.I0(r_SM_Main[1]), .I1(r_SM_Main[0]), 
            .I2(\r_SM_Main[2] ), .I3(\r_SM_Main_2__N_2756[0] ), .O(n19942));
    defparam i2_3_lut_4_lut_adj_839.LUT_INIT = 16'h0100;
    
endmodule
//
// Verilog Description of module uart_rx
//

module uart_rx (GND_net, r_Rx_Data, \r_SM_Main[2] , \r_SM_Main[1] , 
            clk32MHz, n23655, r_Bit_Index, n23658, n28263, n23698, 
            n24171, rx_data, PIN_13_N_26, VCC_net, rx_data_ready, 
            n23665, n23664, n23663, n23662, n23661, n23660, n23659, 
            n23594, n22466, n4, n28231, n1, n27725, n4_adj_1, 
            n4_adj_2, n22471, n44134, n44133, n23471, n23560, n4012) /* synthesis lattice_noprune=1, syn_preserve=0, syn_module_defined=1, syn_noprune=0 */ ;
    input GND_net;
    output r_Rx_Data;
    output \r_SM_Main[2] ;
    output \r_SM_Main[1] ;
    input clk32MHz;
    input n23655;
    output [2:0]r_Bit_Index;
    input n23658;
    input n28263;
    input n23698;
    input n24171;
    output [7:0]rx_data;
    input PIN_13_N_26;
    input VCC_net;
    output rx_data_ready;
    input n23665;
    input n23664;
    input n23663;
    input n23662;
    input n23661;
    input n23660;
    input n23659;
    input n23594;
    output n22466;
    output n4;
    output n28231;
    output n1;
    output n27725;
    output n4_adj_1;
    output n4_adj_2;
    output n22471;
    output n44134;
    output n44133;
    output n23471;
    output n23560;
    output n4012;
    
    wire clk32MHz /* synthesis SET_AS_NETWORK=clk32MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(34[8:16])
    wire [7:0]r_Clock_Count;   // verilog/uart_rx.v(32[17:30])
    
    wire n44103, n23505, n23621, n44169, n39586, n44010, n23615, 
        n44011, n23612, n44013, n23609, n44102, n23606, n40167, 
        n8;
    wire [2:0]r_SM_Main;   // verilog/uart_rx.v(36[17:26])
    
    wire n151, n44175, n44176, n28, n28152;
    wire [2:0]r_SM_Main_2__N_2688;
    
    wire n41980, n44108, n23603, n23689, r_Rx_Data_R, n39692;
    wire [2:0]r_SM_Main_2__N_2682;
    
    wire n40171, n34068, n131, n34067, n34066, n34065, n34064, 
        n34063, n34062, n44009, n22219, n28196, n23412;
    
    SB_LUT4 i15985_3_lut (.I0(r_Clock_Count[1]), .I1(n44103), .I2(n23505), 
            .I3(GND_net), .O(n23621));
    defparam i15985_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11_3_lut (.I0(r_Clock_Count[2]), .I1(n44169), .I2(n23505), 
            .I3(GND_net), .O(n39586));
    defparam i11_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16005_3_lut (.I0(r_Clock_Count[3]), .I1(n44010), .I2(n23505), 
            .I3(GND_net), .O(n23615));
    defparam i16005_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16011_3_lut (.I0(r_Clock_Count[4]), .I1(n44011), .I2(n23505), 
            .I3(GND_net), .O(n23612));
    defparam i16011_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16017_3_lut (.I0(r_Clock_Count[5]), .I1(n44013), .I2(n23505), 
            .I3(GND_net), .O(n23609));
    defparam i16017_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15979_3_lut (.I0(r_Clock_Count[6]), .I1(n44102), .I2(n23505), 
            .I3(GND_net), .O(n23606));
    defparam i15979_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2_3_lut (.I0(r_Clock_Count[2]), .I1(r_Clock_Count[0]), .I2(r_Clock_Count[1]), 
            .I3(GND_net), .O(n40167));
    defparam i2_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 i3_3_lut (.I0(r_Clock_Count[3]), .I1(n40167), .I2(r_Clock_Count[7]), 
            .I3(GND_net), .O(n8));
    defparam i3_3_lut.LUT_INIT = 16'h0404;
    SB_LUT4 i29335_4_lut (.I0(r_Rx_Data), .I1(r_SM_Main[0]), .I2(n8), 
            .I3(n151), .O(n44175));
    defparam i29335_4_lut.LUT_INIT = 16'h3373;
    SB_LUT4 i1_4_lut (.I0(\r_SM_Main[2] ), .I1(n44175), .I2(n44176), .I3(\r_SM_Main[1] ), 
            .O(n28));
    defparam i1_4_lut.LUT_INIT = 16'h5044;
    SB_LUT4 i1_3_lut (.I0(r_Clock_Count[5]), .I1(r_Clock_Count[6]), .I2(r_Clock_Count[4]), 
            .I3(GND_net), .O(n151));
    defparam i1_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i2_3_lut_adj_824 (.I0(r_Clock_Count[0]), .I1(r_Clock_Count[1]), 
            .I2(r_Clock_Count[2]), .I3(GND_net), .O(n28152));
    defparam i2_3_lut_adj_824.LUT_INIT = 16'h8080;
    SB_LUT4 i3_4_lut (.I0(\r_SM_Main[1] ), .I1(r_SM_Main_2__N_2688[0]), 
            .I2(r_Rx_Data), .I3(r_SM_Main[0]), .O(n41980));
    defparam i3_4_lut.LUT_INIT = 16'h1000;
    SB_LUT4 i1_3_lut_adj_825 (.I0(\r_SM_Main[2] ), .I1(n28), .I2(n41980), 
            .I3(GND_net), .O(n23505));
    defparam i1_3_lut_adj_825.LUT_INIT = 16'hcdcd;
    SB_LUT4 i15993_3_lut (.I0(r_Clock_Count[7]), .I1(n44108), .I2(n23505), 
            .I3(GND_net), .O(n23603));
    defparam i15993_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF r_Clock_Count__i7 (.Q(r_Clock_Count[7]), .C(clk32MHz), .D(n23603));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Clock_Count__i6 (.Q(r_Clock_Count[6]), .C(clk32MHz), .D(n23606));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Clock_Count__i5 (.Q(r_Clock_Count[5]), .C(clk32MHz), .D(n23609));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Clock_Count__i4 (.Q(r_Clock_Count[4]), .C(clk32MHz), .D(n23612));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Clock_Count__i3 (.Q(r_Clock_Count[3]), .C(clk32MHz), .D(n23615));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Clock_Count__i2 (.Q(r_Clock_Count[2]), .C(clk32MHz), .D(n39586));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Clock_Count__i1 (.Q(r_Clock_Count[1]), .C(clk32MHz), .D(n23621));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Bit_Index_i2 (.Q(r_Bit_Index[2]), .C(clk32MHz), .D(n23655));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Bit_Index_i1 (.Q(r_Bit_Index[1]), .C(clk32MHz), .D(n23658));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_SM_Main_i1 (.Q(\r_SM_Main[1] ), .C(clk32MHz), .D(n28263));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Clock_Count__i0 (.Q(r_Clock_Count[0]), .C(clk32MHz), .D(n23689));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Bit_Index_i0 (.Q(r_Bit_Index[0]), .C(clk32MHz), .D(n23698));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_Byte_i0 (.Q(rx_data[0]), .C(clk32MHz), .D(n24171));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_Data_50 (.Q(r_Rx_Data), .C(clk32MHz), .D(r_Rx_Data_R));   // verilog/uart_rx.v(41[10] 45[8])
    SB_DFF r_Rx_Data_R_49 (.Q(r_Rx_Data_R), .C(clk32MHz), .D(PIN_13_N_26));   // verilog/uart_rx.v(41[10] 45[8])
    SB_DFFE r_Rx_DV_52 (.Q(rx_data_ready), .C(clk32MHz), .E(VCC_net), 
            .D(n39692));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFFSR r_SM_Main_i2 (.Q(\r_SM_Main[2] ), .C(clk32MHz), .D(r_SM_Main_2__N_2682[2]), 
            .R(n40171));   // verilog/uart_rx.v(49[10] 144[8])
    SB_LUT4 add_62_9_lut (.I0(n131), .I1(r_Clock_Count[7]), .I2(GND_net), 
            .I3(n34068), .O(n44108)) /* synthesis syn_instantiated=1 */ ;
    defparam add_62_9_lut.LUT_INIT = 16'h8228;
    SB_LUT4 add_62_8_lut (.I0(n131), .I1(r_Clock_Count[6]), .I2(GND_net), 
            .I3(n34067), .O(n44102)) /* synthesis syn_instantiated=1 */ ;
    defparam add_62_8_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_62_8 (.CI(n34067), .I0(r_Clock_Count[6]), .I1(GND_net), 
            .CO(n34068));
    SB_LUT4 add_62_7_lut (.I0(n131), .I1(r_Clock_Count[5]), .I2(GND_net), 
            .I3(n34066), .O(n44013)) /* synthesis syn_instantiated=1 */ ;
    defparam add_62_7_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_62_7 (.CI(n34066), .I0(r_Clock_Count[5]), .I1(GND_net), 
            .CO(n34067));
    SB_LUT4 add_62_6_lut (.I0(n131), .I1(r_Clock_Count[4]), .I2(GND_net), 
            .I3(n34065), .O(n44011)) /* synthesis syn_instantiated=1 */ ;
    defparam add_62_6_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_62_6 (.CI(n34065), .I0(r_Clock_Count[4]), .I1(GND_net), 
            .CO(n34066));
    SB_LUT4 add_62_5_lut (.I0(n131), .I1(r_Clock_Count[3]), .I2(GND_net), 
            .I3(n34064), .O(n44010)) /* synthesis syn_instantiated=1 */ ;
    defparam add_62_5_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_62_5 (.CI(n34064), .I0(r_Clock_Count[3]), .I1(GND_net), 
            .CO(n34065));
    SB_LUT4 add_62_4_lut (.I0(n131), .I1(r_Clock_Count[2]), .I2(GND_net), 
            .I3(n34063), .O(n44169)) /* synthesis syn_instantiated=1 */ ;
    defparam add_62_4_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_62_4 (.CI(n34063), .I0(r_Clock_Count[2]), .I1(GND_net), 
            .CO(n34064));
    SB_LUT4 add_62_3_lut (.I0(n131), .I1(r_Clock_Count[1]), .I2(GND_net), 
            .I3(n34062), .O(n44103)) /* synthesis syn_instantiated=1 */ ;
    defparam add_62_3_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_62_3 (.CI(n34062), .I0(r_Clock_Count[1]), .I1(GND_net), 
            .CO(n34063));
    SB_LUT4 add_62_2_lut (.I0(n131), .I1(r_Clock_Count[0]), .I2(GND_net), 
            .I3(VCC_net), .O(n44009)) /* synthesis syn_instantiated=1 */ ;
    defparam add_62_2_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_62_2 (.CI(VCC_net), .I0(r_Clock_Count[0]), .I1(GND_net), 
            .CO(n34062));
    SB_DFF r_Rx_Byte_i1 (.Q(rx_data[1]), .C(clk32MHz), .D(n23665));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_Byte_i2 (.Q(rx_data[2]), .C(clk32MHz), .D(n23664));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_Byte_i3 (.Q(rx_data[3]), .C(clk32MHz), .D(n23663));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_Byte_i4 (.Q(rx_data[4]), .C(clk32MHz), .D(n23662));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_Byte_i5 (.Q(rx_data[5]), .C(clk32MHz), .D(n23661));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_Byte_i6 (.Q(rx_data[6]), .C(clk32MHz), .D(n23660));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_Byte_i7 (.Q(rx_data[7]), .C(clk32MHz), .D(n23659));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_SM_Main_i0 (.Q(r_SM_Main[0]), .C(clk32MHz), .D(n23594));   // verilog/uart_rx.v(49[10] 144[8])
    SB_LUT4 i3_4_lut_adj_826 (.I0(\r_SM_Main[1] ), .I1(r_SM_Main[0]), .I2(\r_SM_Main[2] ), 
            .I3(r_SM_Main_2__N_2682[2]), .O(n22219));   // verilog/uart_rx.v(52[7] 143[14])
    defparam i3_4_lut_adj_826.LUT_INIT = 16'hfdff;
    SB_LUT4 i1_2_lut (.I0(r_Bit_Index[0]), .I1(n22219), .I2(GND_net), 
            .I3(GND_net), .O(n22466));   // verilog/uart_rx.v(52[7] 143[14])
    defparam i1_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 equal_75_i4_2_lut (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[2]), 
            .I2(GND_net), .I3(GND_net), .O(n4));   // verilog/uart_rx.v(97[17:39])
    defparam equal_75_i4_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i15999_3_lut (.I0(r_Clock_Count[0]), .I1(n44009), .I2(n23505), 
            .I3(GND_net), .O(n23689));
    defparam i15999_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 r_SM_Main_2__I_0_56_Mux_0_i2_3_lut (.I0(n28196), .I1(r_SM_Main_2__N_2682[2]), 
            .I2(r_SM_Main[0]), .I3(GND_net), .O(n28231));   // verilog/uart_rx.v(52[7] 143[14])
    defparam r_SM_Main_2__I_0_56_Mux_0_i2_3_lut.LUT_INIT = 16'hc7c7;
    SB_LUT4 r_SM_Main_2__I_0_56_Mux_0_i1_3_lut (.I0(r_Rx_Data), .I1(r_SM_Main_2__N_2688[0]), 
            .I2(r_SM_Main[0]), .I3(GND_net), .O(n1));   // verilog/uart_rx.v(52[7] 143[14])
    defparam r_SM_Main_2__I_0_56_Mux_0_i1_3_lut.LUT_INIT = 16'hc5c5;
    SB_LUT4 i14323_2_lut (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[2]), .I2(GND_net), 
            .I3(GND_net), .O(n27725));
    defparam i14323_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 equal_71_i4_2_lut (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[2]), 
            .I2(GND_net), .I3(GND_net), .O(n4_adj_1));   // verilog/uart_rx.v(97[17:39])
    defparam equal_71_i4_2_lut.LUT_INIT = 16'hbbbb;
    SB_LUT4 equal_73_i4_2_lut (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[2]), 
            .I2(GND_net), .I3(GND_net), .O(n4_adj_2));   // verilog/uart_rx.v(97[17:39])
    defparam equal_73_i4_2_lut.LUT_INIT = 16'hdddd;
    SB_LUT4 i1_2_lut_adj_827 (.I0(n22219), .I1(r_Bit_Index[0]), .I2(GND_net), 
            .I3(GND_net), .O(n22471));   // verilog/uart_rx.v(52[7] 143[14])
    defparam i1_2_lut_adj_827.LUT_INIT = 16'hbbbb;
    SB_LUT4 i14433_3_lut_4_lut (.I0(n151), .I1(r_Clock_Count[7]), .I2(n40167), 
            .I3(r_Clock_Count[3]), .O(r_SM_Main_2__N_2682[2]));
    defparam i14433_3_lut_4_lut.LUT_INIT = 16'hfeee;
    SB_LUT4 i29325_2_lut (.I0(r_SM_Main_2__N_2682[2]), .I1(r_SM_Main[0]), 
            .I2(GND_net), .I3(GND_net), .O(n44134));   // verilog/uart_rx.v(52[7] 143[14])
    defparam i29325_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i29065_3_lut (.I0(r_SM_Main[0]), .I1(r_SM_Main_2__N_2688[0]), 
            .I2(r_Rx_Data), .I3(GND_net), .O(n44133));   // verilog/uart_rx.v(52[7] 143[14])
    defparam i29065_3_lut.LUT_INIT = 16'hfdfd;
    SB_LUT4 i2_3_lut_adj_828 (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[2]), 
            .I2(r_Bit_Index[0]), .I3(GND_net), .O(n28196));
    defparam i2_3_lut_adj_828.LUT_INIT = 16'h8080;
    SB_LUT4 i2_4_lut (.I0(\r_SM_Main[2] ), .I1(r_SM_Main_2__N_2682[2]), 
            .I2(r_SM_Main[0]), .I3(\r_SM_Main[1] ), .O(n23471));
    defparam i2_4_lut.LUT_INIT = 16'h0405;
    SB_LUT4 i10142_3_lut (.I0(n23471), .I1(n28196), .I2(\r_SM_Main[1] ), 
            .I3(GND_net), .O(n23560));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i10142_3_lut.LUT_INIT = 16'h8a8a;
    SB_LUT4 i1072_2_lut (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[0]), .I2(GND_net), 
            .I3(GND_net), .O(n4012));   // verilog/uart_rx.v(102[36:51])
    defparam i1072_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i29337_3_lut_4_lut (.I0(n151), .I1(r_Clock_Count[7]), .I2(r_Clock_Count[3]), 
            .I3(n28152), .O(n44176));
    defparam i29337_3_lut_4_lut.LUT_INIT = 16'hfeee;
    SB_LUT4 i29_1_lut_4_lut (.I0(\r_SM_Main[2] ), .I1(n44175), .I2(n44176), 
            .I3(\r_SM_Main[1] ), .O(n131));
    defparam i29_1_lut_4_lut.LUT_INIT = 16'hafbb;
    SB_LUT4 i1_3_lut_4_lut (.I0(n151), .I1(r_Clock_Count[7]), .I2(n28152), 
            .I3(r_Clock_Count[3]), .O(r_SM_Main_2__N_2688[0]));
    defparam i1_3_lut_4_lut.LUT_INIT = 16'hffef;
    SB_LUT4 i31362_2_lut_3_lut (.I0(\r_SM_Main[1] ), .I1(\r_SM_Main[2] ), 
            .I2(r_SM_Main[0]), .I3(GND_net), .O(n40171));   // verilog/uart_rx.v(52[7] 143[14])
    defparam i31362_2_lut_3_lut.LUT_INIT = 16'hdfdf;
    SB_LUT4 i13_4_lut_4_lut (.I0(\r_SM_Main[1] ), .I1(\r_SM_Main[2] ), .I2(r_SM_Main_2__N_2682[2]), 
            .I3(r_SM_Main[0]), .O(n23412));   // verilog/uart_rx.v(52[7] 143[14])
    defparam i13_4_lut_4_lut.LUT_INIT = 16'h2055;
    SB_LUT4 i12_3_lut_4_lut (.I0(\r_SM_Main[1] ), .I1(\r_SM_Main[2] ), .I2(n23412), 
            .I3(rx_data_ready), .O(n39692));   // verilog/uart_rx.v(52[7] 143[14])
    defparam i12_3_lut_4_lut.LUT_INIT = 16'h2f20;
    
endmodule
//
// Verilog Description of module \quad(DEBOUNCE_TICKS=100)_U1 
//

module \quad(DEBOUNCE_TICKS=100)_U1  (n2276, encoder0_position, GND_net, 
            data_o, clk32MHz, n23721, n23720, n23719, n23718, n23717, 
            n23716, n23715, n23714, n23713, n23712, n23711, n23710, 
            n23709, n23708, n23707, n23706, n23705, n23704, n23703, 
            n23702, n23701, n23700, n23699, n23591, count_enable, 
            n24229, reg_B, PIN_23_c_1, PIN_24_c_0, n23593, n41998) /* synthesis lattice_noprune=1, syn_preserve=0, syn_module_defined=1, syn_noprune=0 */ ;
    output [23:0]n2276;
    output [23:0]encoder0_position;
    input GND_net;
    output [1:0]data_o;
    input clk32MHz;
    input n23721;
    input n23720;
    input n23719;
    input n23718;
    input n23717;
    input n23716;
    input n23715;
    input n23714;
    input n23713;
    input n23712;
    input n23711;
    input n23710;
    input n23709;
    input n23708;
    input n23707;
    input n23706;
    input n23705;
    input n23704;
    input n23703;
    input n23702;
    input n23701;
    input n23700;
    input n23699;
    input n23591;
    output count_enable;
    input n24229;
    output [1:0]reg_B;
    input PIN_23_c_1;
    input PIN_24_c_0;
    input n23593;
    output n41998;
    
    wire clk32MHz /* synthesis SET_AS_NETWORK=clk32MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(34[8:16])
    
    wire n2272, n34081, n34082, n34080, n34079, n34078, count_direction, 
        n34077, B_delayed, A_delayed, n34100, n34099, n34098, n34097, 
        n34096, n34095, n34094, n34093, n34092, n34091, n34090, 
        n34089, n34088, n34087, n34086, n34085, n34083, n34084;
    
    SB_LUT4 add_533_6_lut (.I0(GND_net), .I1(encoder0_position[4]), .I2(n2272), 
            .I3(n34081), .O(n2276[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_533_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_533_6 (.CI(n34081), .I0(encoder0_position[4]), .I1(n2272), 
            .CO(n34082));
    SB_LUT4 add_533_5_lut (.I0(GND_net), .I1(encoder0_position[3]), .I2(n2272), 
            .I3(n34080), .O(n2276[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_533_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_533_5 (.CI(n34080), .I0(encoder0_position[3]), .I1(n2272), 
            .CO(n34081));
    SB_LUT4 add_533_4_lut (.I0(GND_net), .I1(encoder0_position[2]), .I2(n2272), 
            .I3(n34079), .O(n2276[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_533_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_533_4 (.CI(n34079), .I0(encoder0_position[2]), .I1(n2272), 
            .CO(n34080));
    SB_LUT4 add_533_3_lut (.I0(GND_net), .I1(encoder0_position[1]), .I2(n2272), 
            .I3(n34078), .O(n2276[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_533_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_533_3 (.CI(n34078), .I0(encoder0_position[1]), .I1(n2272), 
            .CO(n34079));
    SB_LUT4 add_533_2_lut (.I0(GND_net), .I1(encoder0_position[0]), .I2(count_direction), 
            .I3(n34077), .O(n2276[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_533_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_533_2 (.CI(n34077), .I0(encoder0_position[0]), .I1(count_direction), 
            .CO(n34078));
    SB_CARRY add_533_1 (.CI(GND_net), .I0(n2272), .I1(n2272), .CO(n34077));
    SB_DFF B_delayed_16 (.Q(B_delayed), .C(clk32MHz), .D(data_o[0]));   // quad.v(23[10:54])
    SB_DFF A_delayed_15 (.Q(A_delayed), .C(clk32MHz), .D(data_o[1]));   // quad.v(22[10:54])
    SB_LUT4 add_533_25_lut (.I0(GND_net), .I1(encoder0_position[23]), .I2(n2272), 
            .I3(n34100), .O(n2276[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_533_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_533_24_lut (.I0(GND_net), .I1(encoder0_position[22]), .I2(n2272), 
            .I3(n34099), .O(n2276[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_533_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_533_24 (.CI(n34099), .I0(encoder0_position[22]), .I1(n2272), 
            .CO(n34100));
    SB_LUT4 add_533_23_lut (.I0(GND_net), .I1(encoder0_position[21]), .I2(n2272), 
            .I3(n34098), .O(n2276[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_533_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_533_23 (.CI(n34098), .I0(encoder0_position[21]), .I1(n2272), 
            .CO(n34099));
    SB_LUT4 add_533_22_lut (.I0(GND_net), .I1(encoder0_position[20]), .I2(n2272), 
            .I3(n34097), .O(n2276[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_533_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_533_22 (.CI(n34097), .I0(encoder0_position[20]), .I1(n2272), 
            .CO(n34098));
    SB_LUT4 add_533_21_lut (.I0(GND_net), .I1(encoder0_position[19]), .I2(n2272), 
            .I3(n34096), .O(n2276[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_533_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_533_21 (.CI(n34096), .I0(encoder0_position[19]), .I1(n2272), 
            .CO(n34097));
    SB_LUT4 add_533_20_lut (.I0(GND_net), .I1(encoder0_position[18]), .I2(n2272), 
            .I3(n34095), .O(n2276[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_533_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_533_20 (.CI(n34095), .I0(encoder0_position[18]), .I1(n2272), 
            .CO(n34096));
    SB_LUT4 add_533_19_lut (.I0(GND_net), .I1(encoder0_position[17]), .I2(n2272), 
            .I3(n34094), .O(n2276[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_533_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_533_19 (.CI(n34094), .I0(encoder0_position[17]), .I1(n2272), 
            .CO(n34095));
    SB_LUT4 add_533_18_lut (.I0(GND_net), .I1(encoder0_position[16]), .I2(n2272), 
            .I3(n34093), .O(n2276[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_533_18_lut.LUT_INIT = 16'hC33C;
    SB_DFF count_i0_i1 (.Q(encoder0_position[1]), .C(clk32MHz), .D(n23721));   // quad.v(35[10] 41[6])
    SB_CARRY add_533_18 (.CI(n34093), .I0(encoder0_position[16]), .I1(n2272), 
            .CO(n34094));
    SB_DFF count_i0_i2 (.Q(encoder0_position[2]), .C(clk32MHz), .D(n23720));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i3 (.Q(encoder0_position[3]), .C(clk32MHz), .D(n23719));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i4 (.Q(encoder0_position[4]), .C(clk32MHz), .D(n23718));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i5 (.Q(encoder0_position[5]), .C(clk32MHz), .D(n23717));   // quad.v(35[10] 41[6])
    SB_LUT4 add_533_17_lut (.I0(GND_net), .I1(encoder0_position[15]), .I2(n2272), 
            .I3(n34092), .O(n2276[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_533_17_lut.LUT_INIT = 16'hC33C;
    SB_DFF count_i0_i6 (.Q(encoder0_position[6]), .C(clk32MHz), .D(n23716));   // quad.v(35[10] 41[6])
    SB_CARRY add_533_17 (.CI(n34092), .I0(encoder0_position[15]), .I1(n2272), 
            .CO(n34093));
    SB_DFF count_i0_i7 (.Q(encoder0_position[7]), .C(clk32MHz), .D(n23715));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i8 (.Q(encoder0_position[8]), .C(clk32MHz), .D(n23714));   // quad.v(35[10] 41[6])
    SB_LUT4 add_533_16_lut (.I0(GND_net), .I1(encoder0_position[14]), .I2(n2272), 
            .I3(n34091), .O(n2276[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_533_16_lut.LUT_INIT = 16'hC33C;
    SB_DFF count_i0_i9 (.Q(encoder0_position[9]), .C(clk32MHz), .D(n23713));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i10 (.Q(encoder0_position[10]), .C(clk32MHz), .D(n23712));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i11 (.Q(encoder0_position[11]), .C(clk32MHz), .D(n23711));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i12 (.Q(encoder0_position[12]), .C(clk32MHz), .D(n23710));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i13 (.Q(encoder0_position[13]), .C(clk32MHz), .D(n23709));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i14 (.Q(encoder0_position[14]), .C(clk32MHz), .D(n23708));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i15 (.Q(encoder0_position[15]), .C(clk32MHz), .D(n23707));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i16 (.Q(encoder0_position[16]), .C(clk32MHz), .D(n23706));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i17 (.Q(encoder0_position[17]), .C(clk32MHz), .D(n23705));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i18 (.Q(encoder0_position[18]), .C(clk32MHz), .D(n23704));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i19 (.Q(encoder0_position[19]), .C(clk32MHz), .D(n23703));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i20 (.Q(encoder0_position[20]), .C(clk32MHz), .D(n23702));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i21 (.Q(encoder0_position[21]), .C(clk32MHz), .D(n23701));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i22 (.Q(encoder0_position[22]), .C(clk32MHz), .D(n23700));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i23 (.Q(encoder0_position[23]), .C(clk32MHz), .D(n23699));   // quad.v(35[10] 41[6])
    SB_CARRY add_533_16 (.CI(n34091), .I0(encoder0_position[14]), .I1(n2272), 
            .CO(n34092));
    SB_LUT4 add_533_15_lut (.I0(GND_net), .I1(encoder0_position[13]), .I2(n2272), 
            .I3(n34090), .O(n2276[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_533_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_533_15 (.CI(n34090), .I0(encoder0_position[13]), .I1(n2272), 
            .CO(n34091));
    SB_LUT4 add_533_14_lut (.I0(GND_net), .I1(encoder0_position[12]), .I2(n2272), 
            .I3(n34089), .O(n2276[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_533_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_533_14 (.CI(n34089), .I0(encoder0_position[12]), .I1(n2272), 
            .CO(n34090));
    SB_LUT4 add_533_13_lut (.I0(GND_net), .I1(encoder0_position[11]), .I2(n2272), 
            .I3(n34088), .O(n2276[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_533_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_533_13 (.CI(n34088), .I0(encoder0_position[11]), .I1(n2272), 
            .CO(n34089));
    SB_LUT4 add_533_12_lut (.I0(GND_net), .I1(encoder0_position[10]), .I2(n2272), 
            .I3(n34087), .O(n2276[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_533_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_533_12 (.CI(n34087), .I0(encoder0_position[10]), .I1(n2272), 
            .CO(n34088));
    SB_LUT4 add_533_11_lut (.I0(GND_net), .I1(encoder0_position[9]), .I2(n2272), 
            .I3(n34086), .O(n2276[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_533_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_533_11 (.CI(n34086), .I0(encoder0_position[9]), .I1(n2272), 
            .CO(n34087));
    SB_LUT4 add_533_10_lut (.I0(GND_net), .I1(encoder0_position[8]), .I2(n2272), 
            .I3(n34085), .O(n2276[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_533_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_533_10 (.CI(n34085), .I0(encoder0_position[8]), .I1(n2272), 
            .CO(n34086));
    SB_LUT4 add_533_7_lut (.I0(GND_net), .I1(encoder0_position[5]), .I2(n2272), 
            .I3(n34082), .O(n2276[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_533_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_533_8 (.CI(n34083), .I0(encoder0_position[6]), .I1(n2272), 
            .CO(n34084));
    SB_LUT4 add_533_8_lut (.I0(GND_net), .I1(encoder0_position[6]), .I2(n2272), 
            .I3(n34083), .O(n2276[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_533_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_533_9 (.CI(n34084), .I0(encoder0_position[7]), .I1(n2272), 
            .CO(n34085));
    SB_LUT4 add_533_9_lut (.I0(GND_net), .I1(encoder0_position[7]), .I2(n2272), 
            .I3(n34084), .O(n2276[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_533_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_533_7 (.CI(n34082), .I0(encoder0_position[5]), .I1(n2272), 
            .CO(n34083));
    SB_DFF count_i0_i0 (.Q(encoder0_position[0]), .C(clk32MHz), .D(n23591));   // quad.v(35[10] 41[6])
    SB_LUT4 quadA_debounced_I_0_2_lut (.I0(data_o[1]), .I1(B_delayed), .I2(GND_net), 
            .I3(GND_net), .O(count_direction));   // quad.v(26[26:53])
    defparam quadA_debounced_I_0_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut (.I0(data_o[1]), .I1(data_o[0]), .I2(B_delayed), 
            .I3(A_delayed), .O(count_enable));   // quad.v(25[23:80])
    defparam i3_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i757_1_lut_2_lut (.I0(data_o[1]), .I1(B_delayed), .I2(GND_net), 
            .I3(GND_net), .O(n2272));   // quad.v(37[5] 40[8])
    defparam i757_1_lut_2_lut.LUT_INIT = 16'h9999;
    \grp_debouncer(2,5)_U0  debounce (.n24229(n24229), .data_o({data_o}), 
            .clk32MHz(clk32MHz), .reg_B({reg_B}), .PIN_23_c_1(PIN_23_c_1), 
            .PIN_24_c_0(PIN_24_c_0), .n23593(n23593), .GND_net(GND_net), 
            .n41998(n41998)) /* synthesis lattice_noprune=1, syn_preserve=0, syn_noprune=0 */ ;   // quad.v(15[24] 19[4])
    
endmodule
//
// Verilog Description of module \grp_debouncer(2,5)_U0 
//

module \grp_debouncer(2,5)_U0  (n24229, data_o, clk32MHz, reg_B, PIN_23_c_1, 
            PIN_24_c_0, n23593, GND_net, n41998) /* synthesis lattice_noprune=1, syn_preserve=0, syn_noprune=0 */ ;
    input n24229;
    output [1:0]data_o;
    input clk32MHz;
    output [1:0]reg_B;
    input PIN_23_c_1;
    input PIN_24_c_0;
    input n23593;
    input GND_net;
    output n41998;
    
    wire clk32MHz /* synthesis SET_AS_NETWORK=clk32MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(34[8:16])
    wire [1:0]reg_A;   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(142[12:17])
    wire [2:0]n17;
    wire [2:0]cnt_reg;   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(149[12:19])
    
    wire cnt_next_2__N_3113, n2;
    
    SB_DFF reg_out_i0_i1 (.Q(data_o[1]), .C(clk32MHz), .D(n24229));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(186[9] 190[16])
    SB_DFF reg_B_i0 (.Q(reg_B[0]), .C(clk32MHz), .D(reg_A[0]));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(178[9] 184[16])
    SB_DFF reg_A_i1 (.Q(reg_A[1]), .C(clk32MHz), .D(PIN_23_c_1));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(178[9] 184[16])
    SB_DFFSR cnt_reg_1018__i0 (.Q(cnt_reg[0]), .C(clk32MHz), .D(n17[0]), 
            .R(cnt_next_2__N_3113));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[78:85])
    SB_DFF reg_B_i1 (.Q(reg_B[1]), .C(clk32MHz), .D(reg_A[1]));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(178[9] 184[16])
    SB_DFF reg_A_i0 (.Q(reg_A[0]), .C(clk32MHz), .D(PIN_24_c_0));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(178[9] 184[16])
    SB_DFF reg_out_i0_i0 (.Q(data_o[0]), .C(clk32MHz), .D(n23593));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(186[9] 190[16])
    SB_DFFSR cnt_reg_1018__i1 (.Q(cnt_reg[1]), .C(clk32MHz), .D(n17[1]), 
            .R(cnt_next_2__N_3113));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[78:85])
    SB_DFFSR cnt_reg_1018__i2 (.Q(cnt_reg[2]), .C(clk32MHz), .D(n17[2]), 
            .R(cnt_next_2__N_3113));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[78:85])
    SB_LUT4 i20426_3_lut (.I0(cnt_reg[2]), .I1(cnt_reg[1]), .I2(cnt_reg[0]), 
            .I3(GND_net), .O(n17[2]));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[78:85])
    defparam i20426_3_lut.LUT_INIT = 16'h6a6a;
    SB_LUT4 i20419_2_lut (.I0(cnt_reg[1]), .I1(cnt_reg[0]), .I2(GND_net), 
            .I3(GND_net), .O(n17[1]));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[78:85])
    defparam i20419_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut (.I0(cnt_reg[0]), .I1(cnt_reg[2]), .I2(cnt_reg[1]), 
            .I3(GND_net), .O(n41998));
    defparam i2_3_lut.LUT_INIT = 16'hf7f7;
    SB_LUT4 reg_B_1__I_0_i2_2_lut (.I0(reg_B[1]), .I1(reg_A[1]), .I2(GND_net), 
            .I3(GND_net), .O(n2));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(193[46:60])
    defparam reg_B_1__I_0_i2_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i2_4_lut (.I0(reg_B[0]), .I1(n41998), .I2(reg_A[0]), .I3(n2), 
            .O(cnt_next_2__N_3113));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[40:72])
    defparam i2_4_lut.LUT_INIT = 16'hff7b;
    SB_LUT4 i20417_1_lut (.I0(cnt_reg[0]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n17[0]));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[78:85])
    defparam i20417_1_lut.LUT_INIT = 16'h5555;
    
endmodule
//
// Verilog Description of module \quad(DEBOUNCE_TICKS=100) 
//

module \quad(DEBOUNCE_TICKS=100)  (n24204, encoder1_position, clk32MHz, 
            n24203, n24202, n24201, n24200, n24199, n24198, n24197, 
            n24196, n24195, n24194, n24193, n24192, n24191, n24190, 
            n24189, n24188, n24187, n24186, n24185, n24184, n24183, 
            n24170, data_o, n2226, GND_net, n23592, count_enable, 
            n24231, reg_B, PIN_18_c_1, PIN_19_c_0, n23595, n41767) /* synthesis lattice_noprune=1, syn_preserve=0, syn_module_defined=1, syn_noprune=0 */ ;
    input n24204;
    output [23:0]encoder1_position;
    input clk32MHz;
    input n24203;
    input n24202;
    input n24201;
    input n24200;
    input n24199;
    input n24198;
    input n24197;
    input n24196;
    input n24195;
    input n24194;
    input n24193;
    input n24192;
    input n24191;
    input n24190;
    input n24189;
    input n24188;
    input n24187;
    input n24186;
    input n24185;
    input n24184;
    input n24183;
    input n24170;
    output [1:0]data_o;
    output [23:0]n2226;
    input GND_net;
    input n23592;
    output count_enable;
    input n24231;
    output [1:0]reg_B;
    input PIN_18_c_1;
    input PIN_19_c_0;
    input n23595;
    output n41767;
    
    wire clk32MHz /* synthesis SET_AS_NETWORK=clk32MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(34[8:16])
    
    wire B_delayed, A_delayed, n2216, n34190, n34189, n34188, n34187, 
        n34186, n34185, n34184, n34183, n34182, n34181, n34180, 
        n34179, n34178, n34177, n34176, n34175, n34174, n34173, 
        n34172, n34171, n34170, n34169, n34168, count_direction, 
        n34167;
    
    SB_DFF count_i0_i23 (.Q(encoder1_position[23]), .C(clk32MHz), .D(n24204));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i22 (.Q(encoder1_position[22]), .C(clk32MHz), .D(n24203));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i21 (.Q(encoder1_position[21]), .C(clk32MHz), .D(n24202));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i20 (.Q(encoder1_position[20]), .C(clk32MHz), .D(n24201));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i19 (.Q(encoder1_position[19]), .C(clk32MHz), .D(n24200));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i18 (.Q(encoder1_position[18]), .C(clk32MHz), .D(n24199));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i17 (.Q(encoder1_position[17]), .C(clk32MHz), .D(n24198));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i16 (.Q(encoder1_position[16]), .C(clk32MHz), .D(n24197));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i15 (.Q(encoder1_position[15]), .C(clk32MHz), .D(n24196));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i14 (.Q(encoder1_position[14]), .C(clk32MHz), .D(n24195));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i13 (.Q(encoder1_position[13]), .C(clk32MHz), .D(n24194));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i12 (.Q(encoder1_position[12]), .C(clk32MHz), .D(n24193));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i11 (.Q(encoder1_position[11]), .C(clk32MHz), .D(n24192));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i10 (.Q(encoder1_position[10]), .C(clk32MHz), .D(n24191));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i9 (.Q(encoder1_position[9]), .C(clk32MHz), .D(n24190));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i8 (.Q(encoder1_position[8]), .C(clk32MHz), .D(n24189));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i7 (.Q(encoder1_position[7]), .C(clk32MHz), .D(n24188));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i6 (.Q(encoder1_position[6]), .C(clk32MHz), .D(n24187));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i5 (.Q(encoder1_position[5]), .C(clk32MHz), .D(n24186));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i4 (.Q(encoder1_position[4]), .C(clk32MHz), .D(n24185));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i3 (.Q(encoder1_position[3]), .C(clk32MHz), .D(n24184));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i2 (.Q(encoder1_position[2]), .C(clk32MHz), .D(n24183));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i1 (.Q(encoder1_position[1]), .C(clk32MHz), .D(n24170));   // quad.v(35[10] 41[6])
    SB_DFF B_delayed_16 (.Q(B_delayed), .C(clk32MHz), .D(data_o[0]));   // quad.v(23[10:54])
    SB_DFF A_delayed_15 (.Q(A_delayed), .C(clk32MHz), .D(data_o[1]));   // quad.v(22[10:54])
    SB_LUT4 add_507_25_lut (.I0(GND_net), .I1(encoder1_position[23]), .I2(n2216), 
            .I3(n34190), .O(n2226[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_507_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_507_24_lut (.I0(GND_net), .I1(encoder1_position[22]), .I2(n2216), 
            .I3(n34189), .O(n2226[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_507_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_507_24 (.CI(n34189), .I0(encoder1_position[22]), .I1(n2216), 
            .CO(n34190));
    SB_LUT4 add_507_23_lut (.I0(GND_net), .I1(encoder1_position[21]), .I2(n2216), 
            .I3(n34188), .O(n2226[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_507_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_507_23 (.CI(n34188), .I0(encoder1_position[21]), .I1(n2216), 
            .CO(n34189));
    SB_LUT4 add_507_22_lut (.I0(GND_net), .I1(encoder1_position[20]), .I2(n2216), 
            .I3(n34187), .O(n2226[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_507_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_507_22 (.CI(n34187), .I0(encoder1_position[20]), .I1(n2216), 
            .CO(n34188));
    SB_LUT4 add_507_21_lut (.I0(GND_net), .I1(encoder1_position[19]), .I2(n2216), 
            .I3(n34186), .O(n2226[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_507_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_507_21 (.CI(n34186), .I0(encoder1_position[19]), .I1(n2216), 
            .CO(n34187));
    SB_LUT4 add_507_20_lut (.I0(GND_net), .I1(encoder1_position[18]), .I2(n2216), 
            .I3(n34185), .O(n2226[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_507_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_507_20 (.CI(n34185), .I0(encoder1_position[18]), .I1(n2216), 
            .CO(n34186));
    SB_LUT4 add_507_19_lut (.I0(GND_net), .I1(encoder1_position[17]), .I2(n2216), 
            .I3(n34184), .O(n2226[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_507_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_507_19 (.CI(n34184), .I0(encoder1_position[17]), .I1(n2216), 
            .CO(n34185));
    SB_LUT4 add_507_18_lut (.I0(GND_net), .I1(encoder1_position[16]), .I2(n2216), 
            .I3(n34183), .O(n2226[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_507_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_507_18 (.CI(n34183), .I0(encoder1_position[16]), .I1(n2216), 
            .CO(n34184));
    SB_LUT4 add_507_17_lut (.I0(GND_net), .I1(encoder1_position[15]), .I2(n2216), 
            .I3(n34182), .O(n2226[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_507_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_507_17 (.CI(n34182), .I0(encoder1_position[15]), .I1(n2216), 
            .CO(n34183));
    SB_LUT4 add_507_16_lut (.I0(GND_net), .I1(encoder1_position[14]), .I2(n2216), 
            .I3(n34181), .O(n2226[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_507_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_507_16 (.CI(n34181), .I0(encoder1_position[14]), .I1(n2216), 
            .CO(n34182));
    SB_LUT4 add_507_15_lut (.I0(GND_net), .I1(encoder1_position[13]), .I2(n2216), 
            .I3(n34180), .O(n2226[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_507_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_507_15 (.CI(n34180), .I0(encoder1_position[13]), .I1(n2216), 
            .CO(n34181));
    SB_LUT4 add_507_14_lut (.I0(GND_net), .I1(encoder1_position[12]), .I2(n2216), 
            .I3(n34179), .O(n2226[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_507_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_507_14 (.CI(n34179), .I0(encoder1_position[12]), .I1(n2216), 
            .CO(n34180));
    SB_LUT4 add_507_13_lut (.I0(GND_net), .I1(encoder1_position[11]), .I2(n2216), 
            .I3(n34178), .O(n2226[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_507_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_507_13 (.CI(n34178), .I0(encoder1_position[11]), .I1(n2216), 
            .CO(n34179));
    SB_LUT4 add_507_12_lut (.I0(GND_net), .I1(encoder1_position[10]), .I2(n2216), 
            .I3(n34177), .O(n2226[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_507_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_507_12 (.CI(n34177), .I0(encoder1_position[10]), .I1(n2216), 
            .CO(n34178));
    SB_LUT4 add_507_11_lut (.I0(GND_net), .I1(encoder1_position[9]), .I2(n2216), 
            .I3(n34176), .O(n2226[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_507_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_507_11 (.CI(n34176), .I0(encoder1_position[9]), .I1(n2216), 
            .CO(n34177));
    SB_LUT4 add_507_10_lut (.I0(GND_net), .I1(encoder1_position[8]), .I2(n2216), 
            .I3(n34175), .O(n2226[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_507_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_507_10 (.CI(n34175), .I0(encoder1_position[8]), .I1(n2216), 
            .CO(n34176));
    SB_LUT4 add_507_9_lut (.I0(GND_net), .I1(encoder1_position[7]), .I2(n2216), 
            .I3(n34174), .O(n2226[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_507_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_507_9 (.CI(n34174), .I0(encoder1_position[7]), .I1(n2216), 
            .CO(n34175));
    SB_LUT4 add_507_8_lut (.I0(GND_net), .I1(encoder1_position[6]), .I2(n2216), 
            .I3(n34173), .O(n2226[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_507_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_507_8 (.CI(n34173), .I0(encoder1_position[6]), .I1(n2216), 
            .CO(n34174));
    SB_LUT4 add_507_7_lut (.I0(GND_net), .I1(encoder1_position[5]), .I2(n2216), 
            .I3(n34172), .O(n2226[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_507_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_507_7 (.CI(n34172), .I0(encoder1_position[5]), .I1(n2216), 
            .CO(n34173));
    SB_LUT4 add_507_6_lut (.I0(GND_net), .I1(encoder1_position[4]), .I2(n2216), 
            .I3(n34171), .O(n2226[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_507_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_507_6 (.CI(n34171), .I0(encoder1_position[4]), .I1(n2216), 
            .CO(n34172));
    SB_LUT4 add_507_5_lut (.I0(GND_net), .I1(encoder1_position[3]), .I2(n2216), 
            .I3(n34170), .O(n2226[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_507_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_507_5 (.CI(n34170), .I0(encoder1_position[3]), .I1(n2216), 
            .CO(n34171));
    SB_LUT4 add_507_4_lut (.I0(GND_net), .I1(encoder1_position[2]), .I2(n2216), 
            .I3(n34169), .O(n2226[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_507_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_507_4 (.CI(n34169), .I0(encoder1_position[2]), .I1(n2216), 
            .CO(n34170));
    SB_LUT4 add_507_3_lut (.I0(GND_net), .I1(encoder1_position[1]), .I2(n2216), 
            .I3(n34168), .O(n2226[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_507_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_507_3 (.CI(n34168), .I0(encoder1_position[1]), .I1(n2216), 
            .CO(n34169));
    SB_LUT4 add_507_2_lut (.I0(GND_net), .I1(encoder1_position[0]), .I2(count_direction), 
            .I3(n34167), .O(n2226[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_507_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_507_2 (.CI(n34167), .I0(encoder1_position[0]), .I1(count_direction), 
            .CO(n34168));
    SB_CARRY add_507_1 (.CI(GND_net), .I0(n2216), .I1(n2216), .CO(n34167));
    SB_DFF count_i0_i0 (.Q(encoder1_position[0]), .C(clk32MHz), .D(n23592));   // quad.v(35[10] 41[6])
    SB_LUT4 i3_4_lut (.I0(data_o[1]), .I1(A_delayed), .I2(B_delayed), 
            .I3(data_o[0]), .O(count_enable));   // quad.v(25[23:80])
    defparam i3_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i775_1_lut_2_lut (.I0(data_o[1]), .I1(B_delayed), .I2(GND_net), 
            .I3(GND_net), .O(n2216));   // quad.v(37[5] 40[8])
    defparam i775_1_lut_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 quadA_debounced_I_0_2_lut (.I0(data_o[1]), .I1(B_delayed), .I2(GND_net), 
            .I3(GND_net), .O(count_direction));   // quad.v(26[26:53])
    defparam quadA_debounced_I_0_2_lut.LUT_INIT = 16'h6666;
    \grp_debouncer(2,5)  debounce (.n24231(n24231), .data_o({data_o}), .clk32MHz(clk32MHz), 
            .reg_B({reg_B}), .PIN_18_c_1(PIN_18_c_1), .PIN_19_c_0(PIN_19_c_0), 
            .n23595(n23595), .GND_net(GND_net), .n41767(n41767)) /* synthesis lattice_noprune=1, syn_preserve=0, syn_noprune=0 */ ;   // quad.v(15[24] 19[4])
    
endmodule
//
// Verilog Description of module \grp_debouncer(2,5) 
//

module \grp_debouncer(2,5)  (n24231, data_o, clk32MHz, reg_B, PIN_18_c_1, 
            PIN_19_c_0, n23595, GND_net, n41767) /* synthesis lattice_noprune=1, syn_preserve=0, syn_noprune=0 */ ;
    input n24231;
    output [1:0]data_o;
    input clk32MHz;
    output [1:0]reg_B;
    input PIN_18_c_1;
    input PIN_19_c_0;
    input n23595;
    input GND_net;
    output n41767;
    
    wire clk32MHz /* synthesis SET_AS_NETWORK=clk32MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(34[8:16])
    wire [1:0]reg_A;   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(142[12:17])
    wire [2:0]n17;
    wire [2:0]cnt_reg;   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(149[12:19])
    
    wire cnt_next_2__N_3113, n2;
    
    SB_DFF reg_out_i0_i1 (.Q(data_o[1]), .C(clk32MHz), .D(n24231));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(186[9] 190[16])
    SB_DFF reg_B_i0 (.Q(reg_B[0]), .C(clk32MHz), .D(reg_A[0]));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(178[9] 184[16])
    SB_DFFSR cnt_reg_1019__i0 (.Q(cnt_reg[0]), .C(clk32MHz), .D(n17[0]), 
            .R(cnt_next_2__N_3113));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[78:85])
    SB_DFF reg_A_i1 (.Q(reg_A[1]), .C(clk32MHz), .D(PIN_18_c_1));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(178[9] 184[16])
    SB_DFF reg_B_i1 (.Q(reg_B[1]), .C(clk32MHz), .D(reg_A[1]));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(178[9] 184[16])
    SB_DFF reg_A_i0 (.Q(reg_A[0]), .C(clk32MHz), .D(PIN_19_c_0));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(178[9] 184[16])
    SB_DFF reg_out_i0_i0 (.Q(data_o[0]), .C(clk32MHz), .D(n23595));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(186[9] 190[16])
    SB_DFFSR cnt_reg_1019__i1 (.Q(cnt_reg[1]), .C(clk32MHz), .D(n17[1]), 
            .R(cnt_next_2__N_3113));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[78:85])
    SB_DFFSR cnt_reg_1019__i2 (.Q(cnt_reg[2]), .C(clk32MHz), .D(n17[2]), 
            .R(cnt_next_2__N_3113));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[78:85])
    SB_LUT4 i20448_3_lut (.I0(cnt_reg[2]), .I1(cnt_reg[1]), .I2(cnt_reg[0]), 
            .I3(GND_net), .O(n17[2]));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[78:85])
    defparam i20448_3_lut.LUT_INIT = 16'h6a6a;
    SB_LUT4 i20441_2_lut (.I0(cnt_reg[1]), .I1(cnt_reg[0]), .I2(GND_net), 
            .I3(GND_net), .O(n17[1]));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[78:85])
    defparam i20441_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut (.I0(cnt_reg[0]), .I1(cnt_reg[2]), .I2(cnt_reg[1]), 
            .I3(GND_net), .O(n41767));
    defparam i2_3_lut.LUT_INIT = 16'hf7f7;
    SB_LUT4 reg_B_1__I_0_i2_2_lut (.I0(reg_B[1]), .I1(reg_A[1]), .I2(GND_net), 
            .I3(GND_net), .O(n2));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(193[46:60])
    defparam reg_B_1__I_0_i2_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i2_4_lut (.I0(reg_B[0]), .I1(n41767), .I2(reg_A[0]), .I3(n2), 
            .O(cnt_next_2__N_3113));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[40:72])
    defparam i2_4_lut.LUT_INIT = 16'hff7b;
    SB_LUT4 i20439_1_lut (.I0(cnt_reg[0]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n17[0]));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[78:85])
    defparam i20439_1_lut.LUT_INIT = 16'h5555;
    
endmodule
