// Verilog netlist produced by program LSE :  version Diamond Version 0.0.0
// Netlist written on Mon Jan 17 19:50:21 2022
//
// Verilog Description of module TinyFPGA_B
//

module TinyFPGA_B (CLK, USBPU, ENCODER0_A, ENCODER0_B, ENCODER1_A, 
            ENCODER1_B, HALL1, HALL2, HALL3, FAULT_N, DE, TX, 
            RX, CS_CLK, CS, CS_MISO, SCL, SDA, INLC, INHC, INLB, 
            INHB, INLA, INHA) /* synthesis syn_module_defined=1 */ ;   // verilog/TinyFPGA_B.v(2[8:18])
    input CLK;   // verilog/TinyFPGA_B.v(3[9:12])
    output USBPU;   // verilog/TinyFPGA_B.v(4[10:15])
    input ENCODER0_A;   // verilog/TinyFPGA_B.v(5[9:19])
    input ENCODER0_B;   // verilog/TinyFPGA_B.v(6[9:19])
    input ENCODER1_A;   // verilog/TinyFPGA_B.v(7[9:19])
    input ENCODER1_B;   // verilog/TinyFPGA_B.v(8[9:19])
    input HALL1 /* synthesis black_box_pad_pin=1 */ ;   // verilog/TinyFPGA_B.v(9[9:14])
    input HALL2 /* synthesis black_box_pad_pin=1 */ ;   // verilog/TinyFPGA_B.v(10[9:14])
    input HALL3 /* synthesis black_box_pad_pin=1 */ ;   // verilog/TinyFPGA_B.v(11[9:14])
    input FAULT_N;   // verilog/TinyFPGA_B.v(12[9:16])
    output DE;   // verilog/TinyFPGA_B.v(13[10:12])
    output TX /* synthesis black_box_pad_pin=1 */ ;   // verilog/TinyFPGA_B.v(14[10:12])
    input RX;   // verilog/TinyFPGA_B.v(15[9:11])
    output CS_CLK;   // verilog/TinyFPGA_B.v(16[10:16])
    output CS;   // verilog/TinyFPGA_B.v(17[10:12])
    input CS_MISO;   // verilog/TinyFPGA_B.v(18[9:16])
    inout SCL /* synthesis black_box_pad_pin=1 */ ;   // verilog/TinyFPGA_B.v(19[9:12])
    inout SDA /* synthesis black_box_pad_pin=1 */ ;   // verilog/TinyFPGA_B.v(20[9:12])
    output INLC;   // verilog/TinyFPGA_B.v(21[10:14])
    output INHC;   // verilog/TinyFPGA_B.v(22[10:14])
    output INLB;   // verilog/TinyFPGA_B.v(23[10:14])
    output INHB;   // verilog/TinyFPGA_B.v(24[10:14])
    output INLA;   // verilog/TinyFPGA_B.v(25[10:14])
    output INHA;   // verilog/TinyFPGA_B.v(26[10:14])
    
    wire clk16MHz /* synthesis SET_AS_NETWORK=clk16MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(31[6:14])
    wire clk32MHz /* synthesis SET_AS_NETWORK=clk32MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(31[16:24])
    
    wire GND_net, VCC_net, ENCODER0_A_N, ENCODER0_B_N, ENCODER1_A_N, 
        ENCODER1_B_N, DE_c, RX_c, CS_CLK_c, CS_c, CS_MISO_c, INLC_c_0, 
        INHC_c_0, INLB_c_0, INHB_c_0, INLA_c_0, INHA_c_0;
    wire [7:0]ID;   // verilog/TinyFPGA_B.v(44[12:14])
    
    wire reset, hall1, hall2, hall3, pwm_out, dir, GHA, GHB, 
        GHC;
    wire [23:0]pwm_setpoint;   // verilog/TinyFPGA_B.v(83[20:32])
    wire [23:0]duty;   // verilog/TinyFPGA_B.v(84[21:25])
    wire [7:0]commutation_state;   // verilog/TinyFPGA_B.v(119[12:29])
    wire [7:0]commutation_state_prev;   // verilog/TinyFPGA_B.v(120[12:34])
    
    wire dti;
    wire [7:0]dti_counter;   // verilog/TinyFPGA_B.v(129[12:23])
    
    wire tx_o, tx_enable, n26535, n52782, n52823;
    wire [23:0]setpoint;   // verilog/TinyFPGA_B.v(230[22:30])
    wire [23:0]Kp;   // verilog/TinyFPGA_B.v(231[22:24])
    wire [23:0]Ki;   // verilog/TinyFPGA_B.v(232[22:24])
    wire [7:0]control_mode;   // verilog/TinyFPGA_B.v(234[14:26])
    wire [23:0]PWMLimit;   // verilog/TinyFPGA_B.v(235[22:30])
    wire [23:0]IntegralLimit;   // verilog/TinyFPGA_B.v(236[22:35])
    wire [23:0]deadband;   // verilog/TinyFPGA_B.v(237[22:30])
    wire [15:0]current;   // verilog/TinyFPGA_B.v(238[22:29])
    wire [15:0]current_limit;   // verilog/TinyFPGA_B.v(239[22:35])
    wire [31:0]baudrate;   // verilog/TinyFPGA_B.v(241[15:23])
    wire [23:0]motor_state;   // verilog/TinyFPGA_B.v(268[22:33])
    
    wire data_ready, sda_out, sda_enable, scl, scl_enable;
    wire [31:0]delay_counter;   // verilog/TinyFPGA_B.v(338[11:24])
    
    wire read;
    wire [2:0]\ID_READOUT_FSM.state ;   // verilog/TinyFPGA_B.v(346[15:20])
    
    wire pwm_setpoint_23__N_159, n15, n259, n22431, n293, n297, 
        n298, n299, n300, n301, n302, n303, n304, n305, n306, 
        n307, n308, n63587, n9482, n26534, n26533;
    wire [23:0]pwm_setpoint_23__N_1;
    
    wire n19639;
    wire [7:0]commutation_state_7__N_160;
    
    wire commutation_state_7__N_168, n26532, n26531;
    wire [31:0]encoder0_position;   // verilog/TinyFPGA_B.v(225[11:28])
    
    wire GHA_N_307, GLA_N_324, GHB_N_329, GLB_N_338, GHC_N_343, GLC_N_352, 
        dti_N_356, n26530, RX_N_42, n1507, n60533, n63581, n60513, 
        n60509, n60505, n60499, n1048, n1049, n1050, n1051, n1052, 
        n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, 
        n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, 
        n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, 
        n1077, n1078, n1079, read_N_361, n52313, n35339, n1159, 
        n61749, n4551, n1, n19, n17, n16, n15_adj_5463, n13, 
        n12, n11, n10, n9, n8, n7, n6, n5, n4, n1548;
    wire [31:0]encoder1_position;   // verilog/TinyFPGA_B.v(227[11:28])
    
    wire n2, n14, n15_adj_5464, n16_adj_5465, n17_adj_5466, n18, 
        n19_adj_5467, n20, n21, n22, n23, n24, n25, rx_data_ready;
    wire [7:0]rx_data;   // verilog/coms.v(92[13:20])
    wire [7:0]\data_in_frame[21] ;   // verilog/coms.v(97[12:25])
    wire [7:0]\data_in_frame[20] ;   // verilog/coms.v(97[12:25])
    wire [7:0]\data_in_frame[18] ;   // verilog/coms.v(97[12:25])
    wire [7:0]\data_in_frame[11] ;   // verilog/coms.v(97[12:25])
    wire [7:0]\data_in_frame[4] ;   // verilog/coms.v(97[12:25])
    wire [7:0]\data_in_frame[3] ;   // verilog/coms.v(97[12:25])
    wire [7:0]\data_in_frame[1] ;   // verilog/coms.v(97[12:25])
    wire [7:0]\data_out_frame[27] ;   // verilog/coms.v(98[12:26])
    wire [7:0]\data_out_frame[26] ;   // verilog/coms.v(98[12:26])
    wire [7:0]\data_out_frame[22] ;   // verilog/coms.v(98[12:26])
    wire [7:0]\data_out_frame[21] ;   // verilog/coms.v(98[12:26])
    wire [7:0]\data_out_frame[17] ;   // verilog/coms.v(98[12:26])
    wire [7:0]\data_out_frame[16] ;   // verilog/coms.v(98[12:26])
    wire [7:0]\data_out_frame[15] ;   // verilog/coms.v(98[12:26])
    wire [7:0]\data_out_frame[14] ;   // verilog/coms.v(98[12:26])
    wire [7:0]\data_out_frame[13] ;   // verilog/coms.v(98[12:26])
    wire [7:0]\data_out_frame[12] ;   // verilog/coms.v(98[12:26])
    wire [7:0]\data_out_frame[11] ;   // verilog/coms.v(98[12:26])
    wire [7:0]\data_out_frame[10] ;   // verilog/coms.v(98[12:26])
    wire [7:0]\data_out_frame[9] ;   // verilog/coms.v(98[12:26])
    wire [7:0]\data_out_frame[8] ;   // verilog/coms.v(98[12:26])
    wire [7:0]\data_out_frame[7] ;   // verilog/coms.v(98[12:26])
    wire [7:0]\data_out_frame[6] ;   // verilog/coms.v(98[12:26])
    wire [7:0]\data_out_frame[5] ;   // verilog/coms.v(98[12:26])
    wire [7:0]\data_out_frame[4] ;   // verilog/coms.v(98[12:26])
    wire [7:0]\data_out_frame[3] ;   // verilog/coms.v(98[12:26])
    wire [7:0]\data_out_frame[1] ;   // verilog/coms.v(98[12:26])
    wire [7:0]\data_out_frame[0] ;   // verilog/coms.v(98[12:26])
    wire [7:0]byte_transmit_counter;   // verilog/coms.v(103[12:33])
    wire [31:0]\FRAME_MATCHER.state ;   // verilog/coms.v(113[11:16])
    
    wire n4550, n4549, \FRAME_MATCHER.rx_data_ready_prev , n4529, n4528, 
        n4530, n4531, n4532, n4533, n4534, n4535, n4536, n4537, 
        n4538, n4539, n4540, n4541, n4542, n4543, n4544, n4545, 
        n4546, n4547, n4548, n4834, n61479, n2568, n63575, n46118, 
        n61715, n46043, n46102, n32007, n35347, n46117, n46116, 
        n46115, n2533, n46114, n46042, n46113, n52710, n52712, 
        n52713, n52714, n52715, n52790, n52716, n52717, n52718, 
        n52719, n52720, n52721, n52722, n52723, n52724, n52725, 
        n52726, n52727, n52728, n52729, n52730, n52731, n52732, 
        n52733, n52681, n52734, n52735, n52736, n52737, n52738, 
        n52739, n52740, n52741, n25663, n52742, n52743, n52744, 
        n52745, n52746, n52747, n52748, n52749, n52750, n52751, 
        n52752, n52753, n52754, n52755, n52756, n52757, n52758, 
        n25620, n52759, n52760, n52761, n52762, n52763, n52764, 
        n52765, n52766, n52777, n52767, n52770, n52771, n52772, 
        n52773, n52774, n52775, n52778, n52779, n52780, n52781, 
        n52783, n52776, n52796, n52784, n46112, n26516, n52680, 
        n63569, n46111, n35411, n61681, n46110, n35713, n35402, 
        n61675, n46109, n14_adj_5468, n10_adj_5469, n61659, n46108, 
        n46107, n46106, n46105, n46104, n46101, n46100, n63563, 
        n46041, n46099, n46098, n46103, n46026, n46040, n46097, 
        n46096, n46025, n4_adj_5470, n4_adj_5471, n35211, n55221, 
        n15_adj_5472, n14_adj_5473, n46254, n46253, n46252, n46251, 
        n46250, n46249, n46248, n46247, n46246, n46245, n46244, 
        n46243, n4_adj_5474, n46242, n9484, n9522, n9520, n9518, 
        n61855, n62, \FRAME_MATCHER.i_31__N_2320 , n15_adj_5475, n18203, 
        n8_adj_5476, n26445, n26443, n63545, n26439, n26437, n26435, 
        n26433, n26430, n26428, n26427, n26424, n26422, n26420, 
        n26418, n26416, n26414, n26294, n26291, n26274, n26271, 
        n26268, n26265, n26262, n26253, n26250, n26245, n26244, 
        n26243, n26242, n26238, n26211, n26205, n26202, n26199, 
        n26196, n26193, n26190, n26186, n62647, n19_adj_5477, n17_adj_5478, 
        n16_adj_5479, n15_adj_5480, n13_adj_5481, n11_adj_5482, n9_adj_5483, 
        n8_adj_5484, n7_adj_5485, n6_adj_5486, n5_adj_5487, n4_adj_5488, 
        n30, n62374, n23_adj_5489, n21_adj_5490, n19_adj_5491, n17_adj_5492, 
        n16_adj_5493, n15_adj_5494, n13_adj_5495, n11_adj_5496, n10_adj_5497, 
        n9_adj_5498, n8_adj_5499, n7_adj_5500, n6_adj_5501, n4_adj_5502, 
        n7_adj_5503, n47, n36763, n46039, n4_adj_5504, n4_adj_5505, 
        n6_adj_5506, n27051, n27035, control_update;
    wire [23:0]\PID_CONTROLLER.integral ;   // verilog/motorControl.v(36[23:31])
    
    wire n46038, n240, n258, n284, n292, n336, n337, n338, n339, 
        n340, n341, n343, n344, n345, n346, n347, n348, n349, 
        n350, n351, n352, n353, n354, n355, n356, n357, n358, 
        n359, n46037, n26142, n26970, n6_adj_5507;
    wire [1:0]a_new;   // vhdl/quadrature_decoder.vhd(39[9:14])
    wire [1:0]b_new;   // vhdl/quadrature_decoder.vhd(40[9:14])
    
    wire a_prev, b_prev, debounce_cnt_N_3606, position_31__N_3609, n63539, 
        n5_adj_5508, n26139;
    wire [1:0]a_new_adj_5613;   // vhdl/quadrature_decoder.vhd(39[9:14])
    wire [1:0]b_new_adj_5614;   // vhdl/quadrature_decoder.vhd(40[9:14])
    
    wire a_prev_adj_5511, b_prev_adj_5512, debounce_cnt_N_3606_adj_5513, 
        n26911, n26910, n26909, n26908, n26907, n26906, position_31__N_3609_adj_5514, 
        n26905, n26904, n26903, n26902, n26901, n26900, n26899, 
        n26898, n26897, n26896, n26895, n26894;
    wire [7:0]data_adj_5627;   // verilog/eeprom.v(23[12:16])
    
    wire rw;
    wire [7:0]state_adj_5628;   // verilog/eeprom.v(27[11:16])
    
    wire n46036, n26136, n26133, n26130, n26127, n24_adj_5515, n19770, 
        n26870, n26869, n26868, n11_adj_5516, n26867, n9_adj_5517, 
        n26866, n26865, n26864, n26863, n26862, n26861, n26860, 
        n26859, n26858, n26857, n26856, n26855, n46024, n26854;
    wire [15:0]data_adj_5634;   // verilog/tli4970.v(27[14:18])
    
    wire n26853, n26852, n26851, n26850, n26849, n56512, n26840, 
        n26837, n22357, n26836, n26832, n26829, n26826, n6504, 
        state_7__N_4092, n62259, r_Rx_Data;
    wire [7:0]r_Clock_Count;   // verilog/uart_rx.v(33[17:30])
    wire [2:0]r_Bit_Index;   // verilog/uart_rx.v(34[17:28])
    wire [2:0]r_SM_Main;   // verilog/uart_rx.v(37[17:26])
    
    wire n22269, n4837, n26780, n9486, n9488, n9490, n31535, n6_adj_5526;
    wire [24:0]o_Rx_DV_N_3261;
    
    wire n9492, n9494, n9496, n9498, n9500, n9502, n9504, n9506;
    wire [2:0]r_SM_Main_2__N_3219;
    
    wire n62258, n26767;
    wire [8:0]r_Clock_Count_adj_5650;   // verilog/uart_tx.v(33[16:29])
    wire [2:0]r_Bit_Index_adj_5651;   // verilog/uart_tx.v(34[16:27])
    
    wire n46035, n9508, n9510, n9512, n9514, n9516;
    wire [7:0]state_adj_5663;   // verilog/i2c_controller.v(33[12:17])
    wire [7:0]saved_addr;   // verilog/i2c_controller.v(34[12:22])
    
    wire enable_slow_N_3986;
    wire [7:0]state_7__N_3883;
    
    wire n22369, n6319;
    wire [7:0]state_7__N_3899;
    
    wire n61221, n26710, n26709, n62264, n35374, n5617, n6_adj_5537, 
        n26111, n26702, n9470, n26699, n24669, n26696, n26693, 
        n15_adj_5538, n19_adj_5539, n35, n63521, n62278, n26690, 
        n24621, n52711, n46034, n63515, n57010, n24612, n46033, 
        n46023, n46022, n55498, n6_adj_5540, n46032, n46021, n26687, 
        n46031, n46030, n35277, n22404, n62373, n61973, n61081, 
        n46029, n61079, n1_adj_5541, n12_adj_5542, n9480, n61069, 
        n60201, n4_adj_5543, n6_adj_5544, n8_adj_5545, n9_adj_5546, 
        n25915, n46520, n52769, n46519, n4_adj_5547, n6_adj_5548, 
        n8_adj_5549, n9_adj_5550, n11_adj_5551, n13_adj_5552, n15_adj_5553, 
        n46518, n24535, n6_adj_5554, n46517, n46516, n52819, n24517, 
        n52787, n46515, n46514, n1_adj_5555, n417, n38, n39, n40, 
        n41, n42, n43, n44, n45, n26092, n52818, n24502, n24501, 
        n22377, n22361, n22380, n26091, n4_adj_5556, n3, n4_adj_5557, 
        n52817, n52816, n35435, n24487, n52815, n9409, n9407, 
        n52814, n24463, n52813, n52812, n52811, n52810, n52809, 
        n52808, n52807, n52806, n52797, n52798, n52799, n52800, 
        n52801, n52802, n52803, n52804, n52805, n52683, n52682, 
        n52684, n52685, n52686, n52687, n52688, n52689, n52694, 
        n52693, n52692, n52691, n52690, n52701, n52702, n52794, 
        n52793, n52785, n52786, n52788, n52789, n52795, n52791, 
        n52792, n52695, n52696, n52697, n52698, n25161, n25157, 
        n25141, n25127, n25123, n25559, n25556, n53097, n344_adj_5558, 
        n62817, n46028, n271, n198, n26655, n26649, n26646, n26643, 
        n26640, n26634, n52699, n26090, n26089, n48858, n53, n125, 
        n54542, n60184, n60162, n26085, n61972, n22373, n26083, 
        n26080, n26079, n26078, n26077, n26076, n26587, n48959, 
        n35258, n46020, n46027, n46049, n26567, n26566, n26565, 
        n26564, n26563, n26562, n26561, n26560, n26075, n26074, 
        n52768, n26540, n26539, n26538, n26537, n26536, n52700, 
        n63975, n22256, n46048, n55461, n52703, n46047, n52704, 
        n46019, n10_adj_5559, n55183, n46046, n52705, n52706, n46045, 
        n24840, n52707, n46044, n56726, n26062, n54628, n22253, 
        n52708, n52709, n490, n63009, n47777, n33792, n62372, 
        n6_adj_5560, n60765, n60734, n62218, n60551, n59928, n59927, 
        n59914, n63671, n6_adj_5561, n63006, n51215, n24_adj_5562, 
        n17_adj_5563, n25_adj_5564, n4_adj_5565, n59891, n59888, n5_adj_5566, 
        n51303, n62739, n59865, n63665, n52908, n54590, n62114, 
        n53789, n52872, n63659, n56008, n56002, n62959, n55996, 
        n62948, n55082, n53474, n54544, n55992, n62947, n55986, 
        n62926, n62925, n55980, n55976, n55970, n62479, n55964, 
        n55960, n55954, n55948, n55944, n55938, n53662, n55932, 
        n55928, n55922, n55916, n55912, n55906, n55900, n55896, 
        n55890, n55884, n63647, n62719, n63641, n62124, n57016, 
        n57014, n63635, n62128, n57013, n52055, n55814, n55808, 
        n55525, n34, n33, n18_adj_5567, n17_adj_5568, n16_adj_5569, 
        n14_adj_5570, n12_adj_5571, n62588, n62587, n63629, n8_adj_5572, 
        n62574, n59720, n14_adj_5573, n13_adj_5574, n62540, n63623, 
        n62657, n7_adj_5575, n63617, n29, n27, n23_adj_5576, n55718, 
        n55370, n55666, n62279, n63599, n52431, n63593, n6_adj_5577;
    
    VCC i2 (.Y(VCC_net));
    SB_IO hall2_input (.PACKAGE_PIN(HALL2), .LATCH_INPUT_VALUE(GND_net), 
          .INPUT_CLK(GND_net), .OUTPUT_CLK(GND_net), .OUTPUT_ENABLE(GND_net), 
          .D_OUT_1(GND_net), .D_OUT_0(GND_net), .D_IN_0(hall2)) /* synthesis syn_instantiated=1 */ ;   // /home/administrator/lscc/iCEcube2.2020.12/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam hall2_input.PIN_TYPE = 6'b000001;
    defparam hall2_input.PULLUP = 1'b1;
    defparam hall2_input.NEG_TRIGGER = 1'b0;
    defparam hall2_input.IO_STANDARD = "SB_LVCMOS";
    SB_IO hall3_input (.PACKAGE_PIN(HALL3), .LATCH_INPUT_VALUE(GND_net), 
          .INPUT_CLK(GND_net), .OUTPUT_CLK(GND_net), .OUTPUT_ENABLE(GND_net), 
          .D_OUT_1(GND_net), .D_OUT_0(GND_net), .D_IN_0(hall3)) /* synthesis syn_instantiated=1 */ ;   // /home/administrator/lscc/iCEcube2.2020.12/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam hall3_input.PIN_TYPE = 6'b000001;
    defparam hall3_input.PULLUP = 1'b1;
    defparam hall3_input.NEG_TRIGGER = 1'b0;
    defparam hall3_input.IO_STANDARD = "SB_LVCMOS";
    SB_IO tx_output (.PACKAGE_PIN(TX), .LATCH_INPUT_VALUE(GND_net), .INPUT_CLK(GND_net), 
          .OUTPUT_CLK(GND_net), .OUTPUT_ENABLE(tx_enable), .D_OUT_1(GND_net), 
          .D_OUT_0(tx_o)) /* synthesis syn_instantiated=1 */ ;   // /home/administrator/lscc/iCEcube2.2020.12/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam tx_output.PIN_TYPE = 6'b101001;
    defparam tx_output.PULLUP = 1'b1;
    defparam tx_output.NEG_TRIGGER = 1'b0;
    defparam tx_output.IO_STANDARD = "SB_LVCMOS";
    SB_DFF dir_178 (.Q(dir), .C(clk16MHz), .D(pwm_setpoint_23__N_159));   // verilog/TinyFPGA_B.v(92[9] 117[5])
    SB_DFFE dti_180 (.Q(dti), .C(clk16MHz), .E(n24463), .D(dti_N_356));   // verilog/TinyFPGA_B.v(131[9] 210[5])
    SB_LUT4 i47545_3_lut (.I0(n4_adj_5547), .I1(o_Rx_DV_N_3261[5]), .I2(n11_adj_5551), 
            .I3(GND_net), .O(n62258));   // verilog/uart_tx.v(117[17:57])
    defparam i47545_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF pwm_setpoint_i0 (.Q(pwm_setpoint[0]), .C(clk16MHz), .D(pwm_setpoint_23__N_1[0]));   // verilog/TinyFPGA_B.v(92[9] 117[5])
    SB_IO sda_output (.PACKAGE_PIN(SDA), .LATCH_INPUT_VALUE(GND_net), .INPUT_CLK(GND_net), 
          .OUTPUT_CLK(GND_net), .OUTPUT_ENABLE(sda_enable), .D_OUT_1(GND_net), 
          .D_OUT_0(sda_out), .D_IN_0(state_7__N_3899[3])) /* synthesis syn_instantiated=1 */ ;   // /home/administrator/lscc/iCEcube2.2020.12/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam sda_output.PIN_TYPE = 6'b101001;
    defparam sda_output.PULLUP = 1'b1;
    defparam sda_output.NEG_TRIGGER = 1'b0;
    defparam sda_output.IO_STANDARD = "SB_LVCMOS";
    SB_IO scl_output (.PACKAGE_PIN(SCL), .LATCH_INPUT_VALUE(GND_net), .INPUT_CLK(GND_net), 
          .OUTPUT_CLK(GND_net), .OUTPUT_ENABLE(scl_enable), .D_OUT_1(GND_net), 
          .D_OUT_0(scl)) /* synthesis syn_instantiated=1 */ ;   // /home/administrator/lscc/iCEcube2.2020.12/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam scl_output.PIN_TYPE = 6'b101001;
    defparam scl_output.PULLUP = 1'b1;
    defparam scl_output.NEG_TRIGGER = 1'b0;
    defparam scl_output.IO_STANDARD = "SB_LVCMOS";
    SB_IO hall1_input (.PACKAGE_PIN(HALL1), .LATCH_INPUT_VALUE(GND_net), 
          .INPUT_CLK(GND_net), .OUTPUT_CLK(GND_net), .OUTPUT_ENABLE(GND_net), 
          .D_OUT_1(GND_net), .D_OUT_0(GND_net), .D_IN_0(hall1)) /* synthesis syn_instantiated=1 */ ;   // /home/administrator/lscc/iCEcube2.2020.12/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam hall1_input.PIN_TYPE = 6'b000001;
    defparam hall1_input.PULLUP = 1'b1;
    defparam hall1_input.NEG_TRIGGER = 1'b0;
    defparam hall1_input.IO_STANDARD = "SB_LVCMOS";
    EEPROM eeprom (.clk16MHz(clk16MHz), .enable_slow_N_3986(enable_slow_N_3986), 
           .n5616({n5617}), .\state[2] (state_adj_5628[2]), .n52055(n52055), 
           .n26840(n26840), .VCC_net(VCC_net), .\state[0] (state_adj_5628[0]), 
           .\state[1] (state_adj_5628[1]), .GND_net(GND_net), .n3(n3), 
           .n55082(n55082), .n26090(n26090), .rw(rw), .n52313(n52313), 
           .data_ready(data_ready), .ID({ID}), .baudrate({baudrate}), 
           .n26567(n26567), .n26566(n26566), .n26565(n26565), .n26564(n26564), 
           .n26563(n26563), .n26562(n26562), .n26561(n26561), .n26560(n26560), 
           .n35339(n35339), .n55498(n55498), .n4(n4_adj_5474), .\state[0]_adj_21 (state_adj_5663[0]), 
           .n22361(n22361), .read(read), .data({data_adj_5627}), .scl_enable(scl_enable), 
           .\state_7__N_3883[0] (state_7__N_3883[0]), .n26826(n26826), .n8(n8_adj_5572), 
           .n6319(n6319), .sda_enable(sda_enable), .n35402(n35402), .n26091(n26091), 
           .\saved_addr[0] (saved_addr[0]), .n26080(n26080), .n26079(n26079), 
           .n26078(n26078), .n26077(n26077), .n26076(n26076), .n26075(n26075), 
           .n26074(n26074), .n4_adj_22(n4_adj_5504), .n4_adj_23(n4_adj_5505), 
           .n22404(n22404), .n35435(n35435), .n10(n10_adj_5559), .n52872(n52872), 
           .\state_7__N_3899[3] (state_7__N_3899[3]), .scl(scl), .sda_out(sda_out), 
           .n6(n6_adj_5560), .n22380(n22380)) /* synthesis syn_noprune=1, syn_module_defined=1 */ ;   // verilog/TinyFPGA_B.v(377[10] 389[6])
    SB_LUT4 i47546_3_lut (.I0(n62258), .I1(o_Rx_DV_N_3261[6]), .I2(n13_adj_5552), 
            .I3(GND_net), .O(n62259));   // verilog/uart_tx.v(117[17:57])
    defparam i47546_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_1589_i21_3_lut (.I0(duty[23]), .I1(duty[20]), .I2(n259), 
            .I3(GND_net), .O(n9484));   // verilog/TinyFPGA_B.v(105[13] 116[7])
    defparam mux_1589_i21_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 i13036_3_lut (.I0(\data_in_frame[18] [2]), .I1(rx_data[2]), 
            .I2(n25127), .I3(GND_net), .O(n26640));   // verilog/coms.v(128[12] 296[6])
    defparam i13036_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i46766_4_lut (.I0(n13_adj_5552), .I1(n11_adj_5551), .I2(n9_adj_5550), 
            .I3(n60533), .O(n61479));
    defparam i46766_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 LessThan_1094_i8_3_lut (.I0(n6_adj_5548), .I1(o_Rx_DV_N_3261[4]), 
            .I2(n9_adj_5550), .I3(GND_net), .O(n8_adj_5549));   // verilog/uart_tx.v(117[17:57])
    defparam LessThan_1094_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i17860_3_lut (.I0(n25127), .I1(rx_data[1]), .I2(\data_in_frame[18] [1]), 
            .I3(GND_net), .O(n27035));   // verilog/coms.v(92[13:20])
    defparam i17860_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i46508_3_lut (.I0(n62259), .I1(o_Rx_DV_N_3261[7]), .I2(n15_adj_5553), 
            .I3(GND_net), .O(n61221));   // verilog/uart_tx.v(117[17:57])
    defparam i46508_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i47551_4_lut (.I0(n61221), .I1(n8_adj_5549), .I2(n15_adj_5553), 
            .I3(n61479), .O(n62264));   // verilog/uart_tx.v(117[17:57])
    defparam i47551_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i47552_3_lut (.I0(n62264), .I1(o_Rx_DV_N_3261[8]), .I2(r_Clock_Count_adj_5650[8]), 
            .I3(GND_net), .O(n4837));   // verilog/uart_tx.v(117[17:57])
    defparam i47552_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i13030_3_lut (.I0(\data_in_frame[18] [0]), .I1(rx_data[0]), 
            .I2(n25127), .I3(GND_net), .O(n26634));   // verilog/coms.v(128[12] 296[6])
    defparam i13030_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_3_lut (.I0(n23_adj_5576), .I1(o_Rx_DV_N_3261[12]), .I2(n4837), 
            .I3(GND_net), .O(n55666));
    defparam i1_3_lut.LUT_INIT = 16'hfefe;
    SB_CARRY add_146_14 (.CI(n46030), .I0(delay_counter[12]), .I1(GND_net), 
            .CO(n46031));
    SB_LUT4 i1_4_lut (.I0(o_Rx_DV_N_3261[24]), .I1(n27), .I2(n29), .I3(n55666), 
            .O(n36763));
    defparam i1_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 add_146_5_lut (.I0(GND_net), .I1(delay_counter[3]), .I2(GND_net), 
            .I3(n46021), .O(n1076)) /* synthesis syn_instantiated=1 */ ;
    defparam add_146_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_146_13_lut (.I0(GND_net), .I1(delay_counter[11]), .I2(GND_net), 
            .I3(n46029), .O(n1068)) /* synthesis syn_instantiated=1 */ ;
    defparam add_146_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i12658_3_lut (.I0(\data_in_frame[3] [6]), .I1(rx_data[6]), .I2(n25157), 
            .I3(GND_net), .O(n26262));   // verilog/coms.v(128[12] 296[6])
    defparam i12658_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_1668 (.I0(o_Rx_DV_N_3261[12]), .I1(n4834), .I2(o_Rx_DV_N_3261[8]), 
            .I3(n55948), .O(n55954));
    defparam i1_4_lut_adj_1668.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1669 (.I0(o_Rx_DV_N_3261[24]), .I1(n29), .I2(n23_adj_5576), 
            .I3(n55954), .O(n55960));
    defparam i1_4_lut_adj_1669.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut (.I0(n31535), .I1(Ki[1]), .I2(GND_net), .I3(GND_net), 
            .O(n125));
    defparam i1_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i13447_4_lut (.I0(r_Rx_Data), .I1(rx_data[6]), .I2(n55960), 
            .I3(n27), .O(n27051));   // verilog/uart_rx.v(50[10] 145[8])
    defparam i13447_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 mux_1589_i22_3_lut (.I0(duty[23]), .I1(duty[21]), .I2(n259), 
            .I3(GND_net), .O(n9482));   // verilog/TinyFPGA_B.v(105[13] 116[7])
    defparam mux_1589_i22_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 LessThan_11_i23_2_lut (.I0(current[11]), .I1(duty[11]), .I2(GND_net), 
            .I3(GND_net), .O(n23_adj_5489));   // verilog/TinyFPGA_B.v(98[10:22])
    defparam LessThan_11_i23_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_11_i7_2_lut (.I0(current[3]), .I1(duty[3]), .I2(GND_net), 
            .I3(GND_net), .O(n7_adj_5500));   // verilog/TinyFPGA_B.v(98[10:22])
    defparam LessThan_11_i7_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_11_i11_2_lut (.I0(current[5]), .I1(duty[5]), .I2(GND_net), 
            .I3(GND_net), .O(n11_adj_5496));   // verilog/TinyFPGA_B.v(98[10:22])
    defparam LessThan_11_i11_2_lut.LUT_INIT = 16'h6666;
    SB_DFFESR dti_counter_1934__i0 (.Q(dti_counter[0]), .C(clk16MHz), .E(n24669), 
            .D(n45), .R(n25915));   // verilog/TinyFPGA_B.v(162[23:37])
    SB_LUT4 LessThan_11_i13_2_lut (.I0(current[6]), .I1(duty[6]), .I2(GND_net), 
            .I3(GND_net), .O(n13_adj_5495));   // verilog/TinyFPGA_B.v(98[10:22])
    defparam LessThan_11_i13_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_11_i15_2_lut (.I0(current[7]), .I1(duty[7]), .I2(GND_net), 
            .I3(GND_net), .O(n15_adj_5494));   // verilog/TinyFPGA_B.v(98[10:22])
    defparam LessThan_11_i15_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_11_i9_2_lut (.I0(current[4]), .I1(duty[4]), .I2(GND_net), 
            .I3(GND_net), .O(n9_adj_5498));   // verilog/TinyFPGA_B.v(98[10:22])
    defparam LessThan_11_i9_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_11_i17_2_lut (.I0(current[8]), .I1(duty[8]), .I2(GND_net), 
            .I3(GND_net), .O(n17_adj_5492));   // verilog/TinyFPGA_B.v(98[10:22])
    defparam LessThan_11_i17_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_11_i19_2_lut (.I0(current[9]), .I1(duty[9]), .I2(GND_net), 
            .I3(GND_net), .O(n19_adj_5491));   // verilog/TinyFPGA_B.v(98[10:22])
    defparam LessThan_11_i19_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_11_i21_2_lut (.I0(current[10]), .I1(duty[10]), .I2(GND_net), 
            .I3(GND_net), .O(n21_adj_5490));   // verilog/TinyFPGA_B.v(98[10:22])
    defparam LessThan_11_i21_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_17_i15_2_lut (.I0(duty[7]), .I1(n302), .I2(GND_net), 
            .I3(GND_net), .O(n15_adj_5463));   // verilog/TinyFPGA_B.v(109[11:24])
    defparam LessThan_17_i15_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_17_i13_2_lut (.I0(duty[6]), .I1(n303), .I2(GND_net), 
            .I3(GND_net), .O(n13));   // verilog/TinyFPGA_B.v(109[11:24])
    defparam LessThan_17_i13_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_17_i19_2_lut (.I0(duty[9]), .I1(n300), .I2(GND_net), 
            .I3(GND_net), .O(n19));   // verilog/TinyFPGA_B.v(109[11:24])
    defparam LessThan_17_i19_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_17_i17_2_lut (.I0(duty[8]), .I1(n301), .I2(GND_net), 
            .I3(GND_net), .O(n17));   // verilog/TinyFPGA_B.v(109[11:24])
    defparam LessThan_17_i17_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_17_i7_2_lut (.I0(duty[3]), .I1(n306), .I2(GND_net), 
            .I3(GND_net), .O(n7));   // verilog/TinyFPGA_B.v(109[11:24])
    defparam LessThan_17_i7_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_17_i9_2_lut (.I0(duty[4]), .I1(n305), .I2(GND_net), 
            .I3(GND_net), .O(n9));   // verilog/TinyFPGA_B.v(109[11:24])
    defparam LessThan_17_i9_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_17_i11_2_lut (.I0(duty[5]), .I1(n304), .I2(GND_net), 
            .I3(GND_net), .O(n11));   // verilog/TinyFPGA_B.v(109[11:24])
    defparam LessThan_17_i11_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_17_i5_2_lut (.I0(duty[2]), .I1(n307), .I2(GND_net), 
            .I3(GND_net), .O(n5));   // verilog/TinyFPGA_B.v(109[11:24])
    defparam LessThan_17_i5_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i45801_4_lut (.I0(n11), .I1(n9), .I2(n7), .I3(n5), .O(n60513));
    defparam i45801_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 LessThan_17_i8_3_lut (.I0(n305), .I1(n301), .I2(n17), .I3(GND_net), 
            .O(n8));   // verilog/TinyFPGA_B.v(109[11:24])
    defparam LessThan_17_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_17_i6_3_lut (.I0(n307), .I1(n306), .I2(n7), .I3(GND_net), 
            .O(n6));   // verilog/TinyFPGA_B.v(109[11:24])
    defparam LessThan_17_i6_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_17_i16_3_lut (.I0(n8), .I1(n300), .I2(n19), .I3(GND_net), 
            .O(n16));   // verilog/TinyFPGA_B.v(109[11:24])
    defparam LessThan_17_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2_3_lut (.I0(duty[14]), .I1(duty[18]), .I2(n293), .I3(GND_net), 
            .O(n12_adj_5571));   // verilog/TinyFPGA_B.v(109[11:24])
    defparam i2_3_lut.LUT_INIT = 16'h7e7e;
    SB_LUT4 i6_4_lut (.I0(duty[13]), .I1(n12_adj_5571), .I2(duty[19]), 
            .I3(n293), .O(n16_adj_5569));   // verilog/TinyFPGA_B.v(109[11:24])
    defparam i6_4_lut.LUT_INIT = 16'hdffe;
    SB_LUT4 i4_3_lut (.I0(duty[17]), .I1(duty[22]), .I2(n293), .I3(GND_net), 
            .O(n14_adj_5570));   // verilog/TinyFPGA_B.v(109[11:24])
    defparam i4_3_lut.LUT_INIT = 16'h7e7e;
    SB_LUT4 LessThan_17_i10_3_lut (.I0(n304), .I1(n303), .I2(n13), .I3(GND_net), 
            .O(n10));   // verilog/TinyFPGA_B.v(109[11:24])
    defparam LessThan_17_i10_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_17_i4_3_lut (.I0(n59720), .I1(n308), .I2(duty[1]), 
            .I3(GND_net), .O(n4));   // verilog/TinyFPGA_B.v(109[11:24])
    defparam LessThan_17_i4_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 LessThan_17_i12_3_lut (.I0(n10), .I1(n302), .I2(n15_adj_5463), 
            .I3(GND_net), .O(n12));   // verilog/TinyFPGA_B.v(109[11:24])
    defparam LessThan_17_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i45793_4_lut (.I0(n17), .I1(n15_adj_5463), .I2(n13), .I3(n60513), 
            .O(n60505));
    defparam i45793_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i47944_4_lut (.I0(n16), .I1(n6), .I2(n19), .I3(n60499), 
            .O(n62657));   // verilog/TinyFPGA_B.v(109[11:24])
    defparam i47944_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i47142_4_lut (.I0(n12), .I1(n4), .I2(n15_adj_5463), .I3(n60509), 
            .O(n61855));   // verilog/TinyFPGA_B.v(109[11:24])
    defparam i47142_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i48212_4_lut (.I0(n61855), .I1(n62657), .I2(n19), .I3(n60505), 
            .O(n62925));   // verilog/TinyFPGA_B.v(109[11:24])
    defparam i48212_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i48213_3_lut (.I0(n62925), .I1(n299), .I2(duty[10]), .I3(GND_net), 
            .O(n62926));   // verilog/TinyFPGA_B.v(109[11:24])
    defparam i48213_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i48104_3_lut (.I0(n62926), .I1(n298), .I2(duty[11]), .I3(GND_net), 
            .O(n62817));   // verilog/TinyFPGA_B.v(109[11:24])
    defparam i48104_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i8_4_lut (.I0(duty[21]), .I1(n16_adj_5569), .I2(duty[16]), 
            .I3(n293), .O(n18_adj_5567));   // verilog/TinyFPGA_B.v(109[11:24])
    defparam i8_4_lut.LUT_INIT = 16'hdffe;
    SB_LUT4 i7_4_lut (.I0(duty[20]), .I1(n14_adj_5570), .I2(duty[15]), 
            .I3(n293), .O(n17_adj_5568));   // verilog/TinyFPGA_B.v(109[11:24])
    defparam i7_4_lut.LUT_INIT = 16'hdffe;
    SB_LUT4 i47565_3_lut (.I0(n62817), .I1(n297), .I2(duty[12]), .I3(GND_net), 
            .O(n62278));   // verilog/TinyFPGA_B.v(109[11:24])
    defparam i47565_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i47566_4_lut (.I0(n62278), .I1(n293), .I2(n17_adj_5568), .I3(n18_adj_5567), 
            .O(n62279));   // verilog/TinyFPGA_B.v(109[11:24])
    defparam i47566_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i39170_4_lut (.I0(n259), .I1(duty[23]), .I2(n293), .I3(n62279), 
            .O(n9407));
    defparam i39170_4_lut.LUT_INIT = 16'h1151;
    SB_LUT4 i47002_3_lut (.I0(n15_adj_5494), .I1(n13_adj_5495), .I2(n11_adj_5496), 
            .I3(GND_net), .O(n61715));
    defparam i47002_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i46962_4_lut (.I0(current[15]), .I1(duty[13]), .I2(duty[14]), 
            .I3(n61715), .O(n61675));
    defparam i46962_4_lut.LUT_INIT = 16'h7eff;
    SB_LUT4 i46053_4_lut (.I0(n21_adj_5490), .I1(n19_adj_5491), .I2(n17_adj_5492), 
            .I3(n9_adj_5498), .O(n60765));
    defparam i46053_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i47036_4_lut (.I0(n9_adj_5498), .I1(n7_adj_5500), .I2(current[2]), 
            .I3(duty[2]), .O(n61749));
    defparam i47036_4_lut.LUT_INIT = 16'heffe;
    SB_LUT4 i47415_4_lut (.I0(n15_adj_5494), .I1(n13_adj_5495), .I2(n11_adj_5496), 
            .I3(n61749), .O(n62128));
    defparam i47415_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i47411_4_lut (.I0(n21_adj_5490), .I1(n19_adj_5491), .I2(n17_adj_5492), 
            .I3(n62128), .O(n62124));
    defparam i47411_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i48006_4_lut (.I0(current[15]), .I1(n23_adj_5489), .I2(duty[12]), 
            .I3(n62124), .O(n62719));
    defparam i48006_4_lut.LUT_INIT = 16'hffde;
    SB_LUT4 i46968_4_lut (.I0(current[15]), .I1(duty[13]), .I2(duty[14]), 
            .I3(n62719), .O(n61681));
    defparam i46968_4_lut.LUT_INIT = 16'h7eff;
    SB_LUT4 LessThan_11_i4_4_lut (.I0(duty[0]), .I1(duty[1]), .I2(current[1]), 
            .I3(current[0]), .O(n4_adj_5502));   // verilog/TinyFPGA_B.v(98[10:22])
    defparam LessThan_11_i4_4_lut.LUT_INIT = 16'h0c8e;
    SB_LUT4 i47661_3_lut (.I0(n4_adj_5502), .I1(duty[13]), .I2(current[15]), 
            .I3(GND_net), .O(n62374));   // verilog/TinyFPGA_B.v(98[10:22])
    defparam i47661_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i46946_4_lut (.I0(current[15]), .I1(duty[16]), .I2(duty[17]), 
            .I3(n15_adj_5494), .O(n61659));
    defparam i46946_4_lut.LUT_INIT = 16'hff7e;
    SB_LUT4 LessThan_11_i30_4_lut (.I0(duty[7]), .I1(duty[17]), .I2(current[15]), 
            .I3(duty[16]), .O(n30));   // verilog/TinyFPGA_B.v(98[10:22])
    defparam LessThan_11_i30_4_lut.LUT_INIT = 16'h8f0e;
    SB_LUT4 i46022_4_lut (.I0(current[15]), .I1(duty[15]), .I2(duty[16]), 
            .I3(n61675), .O(n60734));
    defparam i46022_4_lut.LUT_INIT = 16'h5adb;
    SB_LUT4 LessThan_11_i35_rep_267_2_lut (.I0(current[15]), .I1(duty[17]), 
            .I2(GND_net), .I3(GND_net), .O(n63975));   // verilog/TinyFPGA_B.v(98[10:22])
    defparam LessThan_11_i35_rep_267_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i48026_3_lut (.I0(n30), .I1(n10_adj_5497), .I2(n61659), .I3(GND_net), 
            .O(n62739));   // verilog/TinyFPGA_B.v(98[10:22])
    defparam i48026_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i46367_4_lut (.I0(n62374), .I1(duty[15]), .I2(current[15]), 
            .I3(duty[14]), .O(n61079));   // verilog/TinyFPGA_B.v(98[10:22])
    defparam i46367_4_lut.LUT_INIT = 16'h8f0e;
    SB_LUT4 i47659_3_lut (.I0(n6_adj_5501), .I1(duty[10]), .I2(n21_adj_5490), 
            .I3(GND_net), .O(n62372));   // verilog/TinyFPGA_B.v(98[10:22])
    defparam i47659_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i47660_3_lut (.I0(n62372), .I1(duty[11]), .I2(n23_adj_5489), 
            .I3(GND_net), .O(n62373));   // verilog/TinyFPGA_B.v(98[10:22])
    defparam i47660_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i47401_4_lut (.I0(current[15]), .I1(n23_adj_5489), .I2(duty[12]), 
            .I3(n60765), .O(n62114));
    defparam i47401_4_lut.LUT_INIT = 16'hffde;
    SB_LUT4 LessThan_11_i16_3_lut (.I0(n8_adj_5499), .I1(duty[9]), .I2(n19_adj_5491), 
            .I3(GND_net), .O(n16_adj_5493));   // verilog/TinyFPGA_B.v(98[10:22])
    defparam LessThan_11_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i46369_3_lut (.I0(n62373), .I1(duty[12]), .I2(current[15]), 
            .I3(GND_net), .O(n61081));   // verilog/TinyFPGA_B.v(98[10:22])
    defparam i46369_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i12926_3_lut (.I0(current[11]), .I1(data_adj_5634[11]), .I2(n24517), 
            .I3(GND_net), .O(n26530));   // verilog/tli4970.v(35[10] 68[6])
    defparam i12926_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i47766_4_lut (.I0(current[15]), .I1(duty[15]), .I2(duty[16]), 
            .I3(n61681), .O(n62479));
    defparam i47766_4_lut.LUT_INIT = 16'hff7e;
    SB_LUT4 i48246_4_lut (.I0(n61079), .I1(n62739), .I2(n63975), .I3(n60734), 
            .O(n62959));   // verilog/TinyFPGA_B.v(98[10:22])
    defparam i48246_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i47505_3_lut (.I0(n61081), .I1(n16_adj_5493), .I2(n62114), 
            .I3(GND_net), .O(n62218));   // verilog/TinyFPGA_B.v(98[10:22])
    defparam i47505_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i48296_4_lut (.I0(n62218), .I1(n62959), .I2(n63975), .I3(n62479), 
            .O(n63009));   // verilog/TinyFPGA_B.v(98[10:22])
    defparam i48296_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i48293_4_lut (.I0(n63009), .I1(duty[19]), .I2(current[15]), 
            .I3(duty[18]), .O(n63006));   // verilog/TinyFPGA_B.v(98[10:22])
    defparam i48293_4_lut.LUT_INIT = 16'h8f0e;
    SB_LUT4 i2_2_lut (.I0(duty[22]), .I1(current[15]), .I2(GND_net), .I3(GND_net), 
            .O(n6_adj_5554));
    defparam i2_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i47827_4_lut (.I0(n63006), .I1(duty[21]), .I2(current[15]), 
            .I3(duty[20]), .O(n62540));   // verilog/TinyFPGA_B.v(98[10:22])
    defparam i47827_4_lut.LUT_INIT = 16'h8f0e;
    SB_LUT4 i7_4_lut_adj_1670 (.I0(n62540), .I1(duty[23]), .I2(n6_adj_5554), 
            .I3(n259), .O(n9409));
    defparam i7_4_lut_adj_1670.LUT_INIT = 16'h3332;
    SB_LUT4 i1_2_lut_adj_1671 (.I0(n31535), .I1(Ki[2]), .I2(GND_net), 
            .I3(GND_net), .O(n198));
    defparam i1_2_lut_adj_1671.LUT_INIT = 16'h8888;
    SB_IO USBPU_pad (.PACKAGE_PIN(USBPU), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(GND_net));   // /home/administrator/lscc/iCEcube2.2020.12/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam USBPU_pad.PIN_TYPE = 6'b011001;
    defparam USBPU_pad.PULLUP = 1'b0;
    defparam USBPU_pad.NEG_TRIGGER = 1'b0;
    defparam USBPU_pad.IO_STANDARD = "SB_LVCMOS";
    SB_GB_IO CLK_pad (.PACKAGE_PIN(CLK), .OUTPUT_ENABLE(VCC_net), .GLOBAL_BUFFER_OUTPUT(clk16MHz));   // verilog/TinyFPGA_B.v(3[9:12])
    defparam CLK_pad.PIN_TYPE = 6'b000001;
    defparam CLK_pad.PULLUP = 1'b0;
    defparam CLK_pad.NEG_TRIGGER = 1'b0;
    defparam CLK_pad.IO_STANDARD = "SB_LVCMOS";
    SB_DFF pwm_setpoint_i3 (.Q(pwm_setpoint[3]), .C(clk16MHz), .D(pwm_setpoint_23__N_1[3]));   // verilog/TinyFPGA_B.v(92[9] 117[5])
    SB_CARRY add_146_13 (.CI(n46029), .I0(delay_counter[11]), .I1(GND_net), 
            .CO(n46030));
    SB_DFF pwm_setpoint_i2 (.Q(pwm_setpoint[2]), .C(clk16MHz), .D(pwm_setpoint_23__N_1[2]));   // verilog/TinyFPGA_B.v(92[9] 117[5])
    SB_DFF pwm_setpoint_i1 (.Q(pwm_setpoint[1]), .C(clk16MHz), .D(pwm_setpoint_23__N_1[1]));   // verilog/TinyFPGA_B.v(92[9] 117[5])
    SB_LUT4 i1_2_lut_adj_1672 (.I0(n31535), .I1(Ki[3]), .I2(GND_net), 
            .I3(GND_net), .O(n271));
    defparam i1_2_lut_adj_1672.LUT_INIT = 16'h8888;
    SB_LUT4 i12649_3_lut (.I0(\data_in_frame[3] [3]), .I1(rx_data[3]), .I2(n25157), 
            .I3(GND_net), .O(n26253));   // verilog/coms.v(128[12] 296[6])
    defparam i12649_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_adj_1673 (.I0(n31535), .I1(Ki[4]), .I2(GND_net), 
            .I3(GND_net), .O(n344_adj_5558));
    defparam i1_2_lut_adj_1673.LUT_INIT = 16'h8888;
    SB_LUT4 add_146_12_lut (.I0(GND_net), .I1(delay_counter[10]), .I2(GND_net), 
            .I3(n46028), .O(n1069)) /* synthesis syn_instantiated=1 */ ;
    defparam add_146_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_146_33_lut (.I0(GND_net), .I1(delay_counter[31]), .I2(GND_net), 
            .I3(n46049), .O(n1048)) /* synthesis syn_instantiated=1 */ ;
    defparam add_146_33_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_146_5 (.CI(n46021), .I0(delay_counter[3]), .I1(GND_net), 
            .CO(n46022));
    SB_CARRY add_146_12 (.CI(n46028), .I0(delay_counter[10]), .I1(GND_net), 
            .CO(n46029));
    SB_LUT4 add_146_32_lut (.I0(GND_net), .I1(delay_counter[30]), .I2(GND_net), 
            .I3(n46048), .O(n1049)) /* synthesis syn_instantiated=1 */ ;
    defparam add_146_32_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_146_32 (.CI(n46048), .I0(delay_counter[30]), .I1(GND_net), 
            .CO(n46049));
    SB_LUT4 add_146_11_lut (.I0(GND_net), .I1(delay_counter[9]), .I2(GND_net), 
            .I3(n46027), .O(n1070)) /* synthesis syn_instantiated=1 */ ;
    defparam add_146_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_146_31_lut (.I0(GND_net), .I1(delay_counter[29]), .I2(GND_net), 
            .I3(n46047), .O(n1050)) /* synthesis syn_instantiated=1 */ ;
    defparam add_146_31_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_146_31 (.CI(n46047), .I0(delay_counter[29]), .I1(GND_net), 
            .CO(n46048));
    SB_DFFESR dti_counter_1934__i7 (.Q(dti_counter[7]), .C(clk16MHz), .E(n24669), 
            .D(n38), .R(n25915));   // verilog/TinyFPGA_B.v(162[23:37])
    SB_LUT4 i12646_3_lut (.I0(\data_in_frame[3] [2]), .I1(rx_data[2]), .I2(n25157), 
            .I3(GND_net), .O(n26250));   // verilog/coms.v(128[12] 296[6])
    defparam i12646_3_lut.LUT_INIT = 16'hacac;
    SB_DFFESR dti_counter_1934__i6 (.Q(dti_counter[6]), .C(clk16MHz), .E(n24669), 
            .D(n39), .R(n25915));   // verilog/TinyFPGA_B.v(162[23:37])
    SB_DFFESR dti_counter_1934__i5 (.Q(dti_counter[5]), .C(clk16MHz), .E(n24669), 
            .D(n40), .R(n25915));   // verilog/TinyFPGA_B.v(162[23:37])
    SB_DFFESR dti_counter_1934__i4 (.Q(dti_counter[4]), .C(clk16MHz), .E(n24669), 
            .D(n41), .R(n25915));   // verilog/TinyFPGA_B.v(162[23:37])
    SB_LUT4 LessThan_14_i13_2_lut (.I0(current[6]), .I1(current_limit[6]), 
            .I2(GND_net), .I3(GND_net), .O(n13_adj_5481));   // verilog/TinyFPGA_B.v(106[9:30])
    defparam LessThan_14_i13_2_lut.LUT_INIT = 16'h6666;
    SB_DFFESR dti_counter_1934__i3 (.Q(dti_counter[3]), .C(clk16MHz), .E(n24669), 
            .D(n42), .R(n25915));   // verilog/TinyFPGA_B.v(162[23:37])
    SB_DFFESR dti_counter_1934__i2 (.Q(dti_counter[2]), .C(clk16MHz), .E(n24669), 
            .D(n43), .R(n25915));   // verilog/TinyFPGA_B.v(162[23:37])
    SB_LUT4 LessThan_14_i15_2_lut (.I0(current[7]), .I1(current_limit[7]), 
            .I2(GND_net), .I3(GND_net), .O(n15_adj_5480));   // verilog/TinyFPGA_B.v(106[9:30])
    defparam LessThan_14_i15_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_14_i19_2_lut (.I0(current[9]), .I1(current_limit[9]), 
            .I2(GND_net), .I3(GND_net), .O(n19_adj_5477));   // verilog/TinyFPGA_B.v(106[9:30])
    defparam LessThan_14_i19_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_14_i17_2_lut (.I0(current[8]), .I1(current_limit[8]), 
            .I2(GND_net), .I3(GND_net), .O(n17_adj_5478));   // verilog/TinyFPGA_B.v(106[9:30])
    defparam LessThan_14_i17_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_14_i7_2_lut (.I0(current[3]), .I1(current_limit[3]), 
            .I2(GND_net), .I3(GND_net), .O(n7_adj_5485));   // verilog/TinyFPGA_B.v(106[9:30])
    defparam LessThan_14_i7_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_14_i9_2_lut (.I0(current[4]), .I1(current_limit[4]), 
            .I2(GND_net), .I3(GND_net), .O(n9_adj_5483));   // verilog/TinyFPGA_B.v(106[9:30])
    defparam LessThan_14_i9_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_14_i11_2_lut (.I0(current[5]), .I1(current_limit[5]), 
            .I2(GND_net), .I3(GND_net), .O(n11_adj_5482));   // verilog/TinyFPGA_B.v(106[9:30])
    defparam LessThan_14_i11_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_146_30_lut (.I0(GND_net), .I1(delay_counter[28]), .I2(GND_net), 
            .I3(n46046), .O(n1051)) /* synthesis syn_instantiated=1 */ ;
    defparam add_146_30_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_14_i5_2_lut (.I0(current[2]), .I1(current_limit[2]), 
            .I2(GND_net), .I3(GND_net), .O(n5_adj_5487));   // verilog/TinyFPGA_B.v(106[9:30])
    defparam LessThan_14_i5_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_146_30 (.CI(n46046), .I0(delay_counter[28]), .I1(GND_net), 
            .CO(n46047));
    SB_LUT4 i45489_4_lut (.I0(n11_adj_5482), .I1(n9_adj_5483), .I2(n7_adj_5485), 
            .I3(n5_adj_5487), .O(n60201));
    defparam i45489_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 LessThan_14_i16_3_lut (.I0(n8_adj_5484), .I1(current_limit[9]), 
            .I2(n19_adj_5477), .I3(GND_net), .O(n16_adj_5479));   // verilog/TinyFPGA_B.v(106[9:30])
    defparam LessThan_14_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_14_i4_4_lut (.I0(current_limit[0]), .I1(current_limit[1]), 
            .I2(current[1]), .I3(current[0]), .O(n4_adj_5488));   // verilog/TinyFPGA_B.v(106[9:30])
    defparam LessThan_14_i4_4_lut.LUT_INIT = 16'h0c8e;
    SB_LUT4 i47259_3_lut (.I0(n4_adj_5488), .I1(current_limit[5]), .I2(n11_adj_5482), 
            .I3(GND_net), .O(n61972));   // verilog/TinyFPGA_B.v(106[9:30])
    defparam i47259_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i47260_3_lut (.I0(n61972), .I1(current_limit[6]), .I2(n13_adj_5481), 
            .I3(GND_net), .O(n61973));   // verilog/TinyFPGA_B.v(106[9:30])
    defparam i47260_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_146_11 (.CI(n46027), .I0(delay_counter[9]), .I1(GND_net), 
            .CO(n46028));
    SB_LUT4 i45472_4_lut (.I0(n17_adj_5478), .I1(n15_adj_5480), .I2(n13_adj_5481), 
            .I3(n60201), .O(n60184));
    defparam i45472_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i47934_4_lut (.I0(n16_adj_5479), .I1(n6_adj_5486), .I2(n19_adj_5477), 
            .I3(n60162), .O(n62647));   // verilog/TinyFPGA_B.v(106[9:30])
    defparam i47934_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i46357_3_lut (.I0(n61973), .I1(current_limit[7]), .I2(n15_adj_5480), 
            .I3(GND_net), .O(n61069));   // verilog/TinyFPGA_B.v(106[9:30])
    defparam i46357_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i48234_4_lut (.I0(n61069), .I1(n62647), .I2(n19_adj_5477), 
            .I3(n60184), .O(n62947));   // verilog/TinyFPGA_B.v(239[22:35])
    defparam i48234_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i48235_3_lut (.I0(n62947), .I1(current_limit[10]), .I2(current[10]), 
            .I3(GND_net), .O(n62948));   // verilog/TinyFPGA_B.v(239[22:35])
    defparam i48235_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i48124_3_lut (.I0(n62948), .I1(current_limit[11]), .I2(current[11]), 
            .I3(GND_net), .O(n1_adj_5555));   // verilog/TinyFPGA_B.v(239[22:35])
    defparam i48124_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i1_4_lut_adj_1674 (.I0(current_limit[13]), .I1(n1_adj_5555), 
            .I2(current_limit[12]), .I3(current_limit[14]), .O(n54542));   // verilog/TinyFPGA_B.v(106[9:30])
    defparam i1_4_lut_adj_1674.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1675 (.I0(current_limit[13]), .I1(n1_adj_5555), 
            .I2(current_limit[12]), .I3(current_limit[14]), .O(n54544));   // verilog/TinyFPGA_B.v(106[9:30])
    defparam i1_4_lut_adj_1675.LUT_INIT = 16'h8000;
    SB_LUT4 i1_4_lut_adj_1676 (.I0(current[15]), .I1(current_limit[15]), 
            .I2(n54544), .I3(n54542), .O(n259));   // verilog/TinyFPGA_B.v(106[9:30])
    defparam i1_4_lut_adj_1676.LUT_INIT = 16'hb3a2;
    SB_LUT4 i1_4_lut_adj_1677 (.I0(hall3), .I1(commutation_state[1]), .I2(hall2), 
            .I3(hall1), .O(n52431));   // verilog/TinyFPGA_B.v(131[9] 210[5])
    defparam i1_4_lut_adj_1677.LUT_INIT = 16'hd054;
    SB_LUT4 i1_2_lut_adj_1678 (.I0(n31535), .I1(Ki[5]), .I2(GND_net), 
            .I3(GND_net), .O(n417));
    defparam i1_2_lut_adj_1678.LUT_INIT = 16'h8888;
    SB_LUT4 i12634_3_lut (.I0(\data_in_frame[3] [1]), .I1(rx_data[1]), .I2(n25157), 
            .I3(GND_net), .O(n26238));   // verilog/coms.v(128[12] 296[6])
    defparam i12634_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_adj_1679 (.I0(n31535), .I1(Ki[6]), .I2(GND_net), 
            .I3(GND_net), .O(n490));
    defparam i1_2_lut_adj_1679.LUT_INIT = 16'h8888;
    SB_LUT4 i9_2_lut (.I0(n292), .I1(n240), .I2(GND_net), .I3(GND_net), 
            .O(n35));
    defparam i9_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_4_lut_adj_1680 (.I0(state_adj_5628[2]), .I1(state_adj_5628[1]), 
            .I2(state_adj_5628[0]), .I3(n35339), .O(n52055));   // verilog/eeprom.v(35[8] 81[4])
    defparam i1_4_lut_adj_1680.LUT_INIT = 16'ha8e8;
    SB_LUT4 mux_1589_i23_3_lut (.I0(duty[23]), .I1(duty[22]), .I2(n259), 
            .I3(GND_net), .O(n9480));   // verilog/TinyFPGA_B.v(105[13] 116[7])
    defparam mux_1589_i23_3_lut.LUT_INIT = 16'h3535;
    SB_DFFESR dti_counter_1934__i1 (.Q(dti_counter[1]), .C(clk16MHz), .E(n24669), 
            .D(n44), .R(n25915));   // verilog/TinyFPGA_B.v(162[23:37])
    SB_DFFE commutation_state_i1 (.Q(commutation_state[1]), .C(clk16MHz), 
            .E(VCC_net), .D(n52431));   // verilog/TinyFPGA_B.v(131[9] 210[5])
    SB_IO CS_MISO_pad (.PACKAGE_PIN(CS_MISO), .OUTPUT_ENABLE(VCC_net), .D_IN_0(CS_MISO_c));   // /home/administrator/lscc/iCEcube2.2020.12/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam CS_MISO_pad.PIN_TYPE = 6'b000001;
    defparam CS_MISO_pad.PULLUP = 1'b0;
    defparam CS_MISO_pad.NEG_TRIGGER = 1'b0;
    defparam CS_MISO_pad.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 add_146_4_lut (.I0(GND_net), .I1(delay_counter[2]), .I2(GND_net), 
            .I3(n46020), .O(n1077)) /* synthesis syn_instantiated=1 */ ;
    defparam add_146_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_146_29_lut (.I0(GND_net), .I1(delay_counter[27]), .I2(GND_net), 
            .I3(n46045), .O(n1052)) /* synthesis syn_instantiated=1 */ ;
    defparam add_146_29_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i12810_4_lut (.I0(CS_MISO_c), .I1(data_adj_5634[1]), .I2(n5_adj_5508), 
            .I3(n4_adj_5565), .O(n26414));   // verilog/tli4970.v(35[10] 68[6])
    defparam i12810_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i12812_4_lut (.I0(CS_MISO_c), .I1(data_adj_5634[2]), .I2(n6_adj_5537), 
            .I3(n22357), .O(n26416));   // verilog/tli4970.v(35[10] 68[6])
    defparam i12812_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 add_146_10_lut (.I0(GND_net), .I1(delay_counter[8]), .I2(GND_net), 
            .I3(n46026), .O(n1071)) /* synthesis syn_instantiated=1 */ ;
    defparam add_146_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i12814_4_lut (.I0(CS_MISO_c), .I1(data_adj_5634[3]), .I2(n6_adj_5537), 
            .I3(n22373), .O(n26418));   // verilog/tli4970.v(35[10] 68[6])
    defparam i12814_4_lut.LUT_INIT = 16'hccca;
    SB_CARRY add_146_29 (.CI(n46045), .I0(delay_counter[27]), .I1(GND_net), 
            .CO(n46046));
    SB_LUT4 i12816_4_lut (.I0(CS_MISO_c), .I1(data_adj_5634[4]), .I2(n9_adj_5517), 
            .I3(n22377), .O(n26420));   // verilog/tli4970.v(35[10] 68[6])
    defparam i12816_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 add_1103_25_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_setpoint_23__N_159), 
            .I3(n46118), .O(n4528)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1103_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_1103_24_lut (.I0(GND_net), .I1(GND_net), .I2(n9480), .I3(n46117), 
            .O(n4529)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1103_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i12818_4_lut (.I0(CS_MISO_c), .I1(data_adj_5634[5]), .I2(n5_adj_5508), 
            .I3(n22377), .O(n26422));   // verilog/tli4970.v(35[10] 68[6])
    defparam i12818_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 n9409_bdd_4_lut (.I0(n9409), .I1(current[15]), .I2(duty[22]), 
            .I3(n9407), .O(n63671));
    defparam n9409_bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_LUT4 i12820_4_lut (.I0(CS_MISO_c), .I1(data_adj_5634[6]), .I2(n6_adj_5507), 
            .I3(n22357), .O(n26424));   // verilog/tli4970.v(35[10] 68[6])
    defparam i12820_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 n63671_bdd_4_lut (.I0(n63671), .I1(duty[19]), .I2(n4532), 
            .I3(n9407), .O(pwm_setpoint_23__N_1[19]));
    defparam n63671_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i12823_4_lut (.I0(CS_MISO_c), .I1(data_adj_5634[7]), .I2(n6_adj_5507), 
            .I3(n22373), .O(n26427));   // verilog/tli4970.v(35[10] 68[6])
    defparam i12823_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i12824_4_lut (.I0(CS_MISO_c), .I1(data_adj_5634[8]), .I2(n9_adj_5517), 
            .I3(n22369), .O(n26428));   // verilog/tli4970.v(35[10] 68[6])
    defparam i12824_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 n9409_bdd_4_lut_48887 (.I0(n9409), .I1(current[15]), .I2(duty[21]), 
            .I3(n9407), .O(n63665));
    defparam n9409_bdd_4_lut_48887.LUT_INIT = 16'he4aa;
    SB_CARRY add_1103_24 (.CI(n46117), .I0(GND_net), .I1(n9480), .CO(n46118));
    SB_LUT4 add_1103_23_lut (.I0(GND_net), .I1(GND_net), .I2(n9482), .I3(n46116), 
            .O(n4530)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1103_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i12826_4_lut (.I0(CS_MISO_c), .I1(data_adj_5634[9]), .I2(n5_adj_5508), 
            .I3(n22369), .O(n26430));   // verilog/tli4970.v(35[10] 68[6])
    defparam i12826_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i12601_3_lut (.I0(\data_in_frame[1] [7]), .I1(rx_data[7]), .I2(n25161), 
            .I3(GND_net), .O(n26205));   // verilog/coms.v(128[12] 296[6])
    defparam i12601_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 n63665_bdd_4_lut (.I0(n63665), .I1(duty[18]), .I2(n4533), 
            .I3(n9407), .O(pwm_setpoint_23__N_1[18]));
    defparam n63665_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i12598_3_lut (.I0(\data_in_frame[1] [6]), .I1(rx_data[6]), .I2(n25161), 
            .I3(GND_net), .O(n26202));   // verilog/coms.v(128[12] 296[6])
    defparam i12598_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12829_4_lut (.I0(CS_MISO_c), .I1(data_adj_5634[10]), .I2(n6_adj_5506), 
            .I3(n22357), .O(n26433));   // verilog/tli4970.v(35[10] 68[6])
    defparam i12829_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i12595_3_lut (.I0(\data_in_frame[1] [5]), .I1(rx_data[5]), .I2(n25161), 
            .I3(GND_net), .O(n26199));   // verilog/coms.v(128[12] 296[6])
    defparam i12595_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12831_4_lut (.I0(CS_MISO_c), .I1(data_adj_5634[11]), .I2(n35347), 
            .I3(n22369), .O(n26435));   // verilog/tli4970.v(35[10] 68[6])
    defparam i12831_4_lut.LUT_INIT = 16'hccac;
    SB_LUT4 i12592_3_lut (.I0(\data_in_frame[1] [4]), .I1(rx_data[4]), .I2(n25161), 
            .I3(GND_net), .O(n26196));   // verilog/coms.v(128[12] 296[6])
    defparam i12592_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 n9409_bdd_4_lut_48882 (.I0(n9409), .I1(current[15]), .I2(duty[20]), 
            .I3(n9407), .O(n63659));
    defparam n9409_bdd_4_lut_48882.LUT_INIT = 16'he4aa;
    SB_LUT4 i12833_4_lut (.I0(CS_MISO_c), .I1(data_adj_5634[12]), .I2(n9_adj_5517), 
            .I3(n4_adj_5470), .O(n26437));   // verilog/tli4970.v(35[10] 68[6])
    defparam i12833_4_lut.LUT_INIT = 16'hccca;
    SB_CARRY add_1103_23 (.CI(n46116), .I0(GND_net), .I1(n9482), .CO(n46117));
    SB_LUT4 add_1103_22_lut (.I0(GND_net), .I1(GND_net), .I2(n9484), .I3(n46115), 
            .O(n4531)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1103_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i12589_3_lut (.I0(\data_in_frame[1] [3]), .I1(rx_data[3]), .I2(n25161), 
            .I3(GND_net), .O(n26193));   // verilog/coms.v(128[12] 296[6])
    defparam i12589_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 n63659_bdd_4_lut (.I0(n63659), .I1(duty[17]), .I2(n4534), 
            .I3(n9407), .O(pwm_setpoint_23__N_1[17]));
    defparam n63659_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i12835_4_lut (.I0(CS_MISO_c), .I1(data_adj_5634[15]), .I2(n35411), 
            .I3(n22373), .O(n26439));   // verilog/tli4970.v(35[10] 68[6])
    defparam i12835_4_lut.LUT_INIT = 16'hccac;
    SB_CARRY add_1103_22 (.CI(n46115), .I0(GND_net), .I1(n9484), .CO(n46116));
    SB_LUT4 add_1103_21_lut (.I0(GND_net), .I1(GND_net), .I2(n9486), .I3(n46114), 
            .O(n4532)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1103_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i12586_3_lut (.I0(\data_in_frame[1] [2]), .I1(rx_data[2]), .I2(n25161), 
            .I3(GND_net), .O(n26190));   // verilog/coms.v(128[12] 296[6])
    defparam i12586_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 add_146_28_lut (.I0(GND_net), .I1(delay_counter[26]), .I2(GND_net), 
            .I3(n46044), .O(n1053)) /* synthesis syn_instantiated=1 */ ;
    defparam add_146_28_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_2_lut_adj_1681 (.I0(r_SM_Main[1]), .I1(r_SM_Main[2]), .I2(GND_net), 
            .I3(GND_net), .O(n52823));   // verilog/uart_rx.v(50[10] 145[8])
    defparam i1_2_lut_adj_1681.LUT_INIT = 16'h2222;
    SB_LUT4 i1_4_lut_adj_1682 (.I0(o_Rx_DV_N_3261[12]), .I1(n4834), .I2(o_Rx_DV_N_3261[8]), 
            .I3(n55932), .O(n55938));
    defparam i1_4_lut_adj_1682.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1683 (.I0(o_Rx_DV_N_3261[24]), .I1(n29), .I2(n23_adj_5576), 
            .I3(n55938), .O(n55944));
    defparam i1_4_lut_adj_1683.LUT_INIT = 16'hfffe;
    SB_LUT4 i12839_4_lut (.I0(r_Rx_Data), .I1(rx_data[1]), .I2(n55944), 
            .I3(n27), .O(n26443));   // verilog/uart_rx.v(50[10] 145[8])
    defparam i12839_4_lut.LUT_INIT = 16'hccca;
    SB_DFF \ID_READOUT_FSM.state__i1  (.Q(\ID_READOUT_FSM.state [1]), .C(clk16MHz), 
           .D(n17_adj_5563));   // verilog/TinyFPGA_B.v(345[10] 375[6])
    SB_DFFE \ID_READOUT_FSM.state__i0  (.Q(\ID_READOUT_FSM.state [0]), .C(clk16MHz), 
            .E(VCC_net), .D(n51215));   // verilog/TinyFPGA_B.v(345[10] 375[6])
    SB_DFF commutation_state_prev_i2 (.Q(commutation_state_prev[2]), .C(clk16MHz), 
           .D(commutation_state[2]));   // verilog/TinyFPGA_B.v(131[9] 210[5])
    SB_CARRY add_1103_21 (.CI(n46114), .I0(GND_net), .I1(n9486), .CO(n46115));
    SB_LUT4 i12690_3_lut (.I0(\data_in_frame[4] [7]), .I1(rx_data[7]), .I2(n7_adj_5575), 
            .I3(GND_net), .O(n26294));   // verilog/coms.v(128[12] 296[6])
    defparam i12690_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 add_1103_20_lut (.I0(GND_net), .I1(GND_net), .I2(n9488), .I3(n46113), 
            .O(n4533)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1103_20_lut.LUT_INIT = 16'hC33C;
    SB_IO RX_pad (.PACKAGE_PIN(RX), .OUTPUT_ENABLE(VCC_net), .D_IN_0(RX_c));   // /home/administrator/lscc/iCEcube2.2020.12/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam RX_pad.PIN_TYPE = 6'b000001;
    defparam RX_pad.PULLUP = 1'b0;
    defparam RX_pad.NEG_TRIGGER = 1'b0;
    defparam RX_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO ENCODER1_B_pad (.PACKAGE_PIN(ENCODER1_B), .OUTPUT_ENABLE(VCC_net), 
          .D_IN_0(ENCODER1_B_N));   // /home/administrator/lscc/iCEcube2.2020.12/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam ENCODER1_B_pad.PIN_TYPE = 6'b000001;
    defparam ENCODER1_B_pad.PULLUP = 1'b0;
    defparam ENCODER1_B_pad.NEG_TRIGGER = 1'b0;
    defparam ENCODER1_B_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO ENCODER1_A_pad (.PACKAGE_PIN(ENCODER1_A), .OUTPUT_ENABLE(VCC_net), 
          .D_IN_0(ENCODER1_A_N));   // /home/administrator/lscc/iCEcube2.2020.12/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam ENCODER1_A_pad.PIN_TYPE = 6'b000001;
    defparam ENCODER1_A_pad.PULLUP = 1'b0;
    defparam ENCODER1_A_pad.NEG_TRIGGER = 1'b0;
    defparam ENCODER1_A_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO ENCODER0_B_pad (.PACKAGE_PIN(ENCODER0_B), .OUTPUT_ENABLE(VCC_net), 
          .D_IN_0(ENCODER0_B_N));   // /home/administrator/lscc/iCEcube2.2020.12/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam ENCODER0_B_pad.PIN_TYPE = 6'b000001;
    defparam ENCODER0_B_pad.PULLUP = 1'b0;
    defparam ENCODER0_B_pad.NEG_TRIGGER = 1'b0;
    defparam ENCODER0_B_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO ENCODER0_A_pad (.PACKAGE_PIN(ENCODER0_A), .OUTPUT_ENABLE(VCC_net), 
          .D_IN_0(ENCODER0_A_N));   // /home/administrator/lscc/iCEcube2.2020.12/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam ENCODER0_A_pad.PIN_TYPE = 6'b000001;
    defparam ENCODER0_A_pad.PULLUP = 1'b0;
    defparam ENCODER0_A_pad.NEG_TRIGGER = 1'b0;
    defparam ENCODER0_A_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO INHA_pad (.PACKAGE_PIN(INHA), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(INHA_c_0));   // /home/administrator/lscc/iCEcube2.2020.12/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam INHA_pad.PIN_TYPE = 6'b011001;
    defparam INHA_pad.PULLUP = 1'b0;
    defparam INHA_pad.NEG_TRIGGER = 1'b0;
    defparam INHA_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO DE_pad (.PACKAGE_PIN(DE), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(DE_c));   // /home/administrator/lscc/iCEcube2.2020.12/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DE_pad.PIN_TYPE = 6'b011001;
    defparam DE_pad.PULLUP = 1'b0;
    defparam DE_pad.NEG_TRIGGER = 1'b0;
    defparam DE_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO INLA_pad (.PACKAGE_PIN(INLA), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(INLA_c_0));   // /home/administrator/lscc/iCEcube2.2020.12/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam INLA_pad.PIN_TYPE = 6'b011001;
    defparam INLA_pad.PULLUP = 1'b0;
    defparam INLA_pad.NEG_TRIGGER = 1'b0;
    defparam INLA_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO INHB_pad (.PACKAGE_PIN(INHB), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(INHB_c_0));   // /home/administrator/lscc/iCEcube2.2020.12/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam INHB_pad.PIN_TYPE = 6'b011001;
    defparam INHB_pad.PULLUP = 1'b0;
    defparam INHB_pad.NEG_TRIGGER = 1'b0;
    defparam INHB_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO INLB_pad (.PACKAGE_PIN(INLB), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(INLB_c_0));   // /home/administrator/lscc/iCEcube2.2020.12/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam INLB_pad.PIN_TYPE = 6'b011001;
    defparam INLB_pad.PULLUP = 1'b0;
    defparam INLB_pad.NEG_TRIGGER = 1'b0;
    defparam INLB_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO INHC_pad (.PACKAGE_PIN(INHC), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(INHC_c_0));   // /home/administrator/lscc/iCEcube2.2020.12/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam INHC_pad.PIN_TYPE = 6'b011001;
    defparam INHC_pad.PULLUP = 1'b0;
    defparam INHC_pad.NEG_TRIGGER = 1'b0;
    defparam INHC_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO INLC_pad (.PACKAGE_PIN(INLC), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(INLC_c_0));   // /home/administrator/lscc/iCEcube2.2020.12/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam INLC_pad.PIN_TYPE = 6'b011001;
    defparam INLC_pad.PULLUP = 1'b0;
    defparam INLC_pad.NEG_TRIGGER = 1'b0;
    defparam INLC_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO CS_pad (.PACKAGE_PIN(CS), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(CS_c));   // /home/administrator/lscc/iCEcube2.2020.12/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam CS_pad.PIN_TYPE = 6'b011001;
    defparam CS_pad.PULLUP = 1'b0;
    defparam CS_pad.NEG_TRIGGER = 1'b0;
    defparam CS_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO CS_CLK_pad (.PACKAGE_PIN(CS_CLK), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(CS_CLK_c));   // /home/administrator/lscc/iCEcube2.2020.12/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam CS_CLK_pad.PIN_TYPE = 6'b011001;
    defparam CS_CLK_pad.PULLUP = 1'b0;
    defparam CS_CLK_pad.NEG_TRIGGER = 1'b0;
    defparam CS_CLK_pad.IO_STANDARD = "SB_LVCMOS";
    SB_CARRY add_1103_20 (.CI(n46113), .I0(GND_net), .I1(n9488), .CO(n46114));
    SB_LUT4 add_1103_19_lut (.I0(GND_net), .I1(GND_net), .I2(n9490), .I3(n46112), 
            .O(n4534)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1103_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_146_28 (.CI(n46044), .I0(delay_counter[26]), .I1(GND_net), 
            .CO(n46045));
    SB_CARRY add_1103_19 (.CI(n46112), .I0(GND_net), .I1(n9490), .CO(n46113));
    SB_LUT4 add_1103_18_lut (.I0(GND_net), .I1(GND_net), .I2(n9492), .I3(n46111), 
            .O(n4535)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1103_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_146_27_lut (.I0(GND_net), .I1(delay_counter[25]), .I2(GND_net), 
            .I3(n46043), .O(n1054)) /* synthesis syn_instantiated=1 */ ;
    defparam add_146_27_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i12687_3_lut (.I0(\data_in_frame[4] [6]), .I1(rx_data[6]), .I2(n7_adj_5575), 
            .I3(GND_net), .O(n26291));   // verilog/coms.v(128[12] 296[6])
    defparam i12687_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY add_1103_18 (.CI(n46111), .I0(GND_net), .I1(n9492), .CO(n46112));
    SB_LUT4 add_1103_17_lut (.I0(GND_net), .I1(GND_net), .I2(n9494), .I3(n46110), 
            .O(n4536)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1103_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1103_17 (.CI(n46110), .I0(GND_net), .I1(n9494), .CO(n46111));
    SB_LUT4 i1_4_lut_adj_1684 (.I0(o_Rx_DV_N_3261[12]), .I1(n4834), .I2(o_Rx_DV_N_3261[8]), 
            .I3(n55900), .O(n55906));
    defparam i1_4_lut_adj_1684.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1685 (.I0(o_Rx_DV_N_3261[24]), .I1(n29), .I2(n23_adj_5576), 
            .I3(n55906), .O(n55912));
    defparam i1_4_lut_adj_1685.LUT_INIT = 16'hfffe;
    SB_LUT4 i12670_3_lut (.I0(\data_in_frame[4] [2]), .I1(rx_data[2]), .I2(n7_adj_5575), 
            .I3(GND_net), .O(n26274));   // verilog/coms.v(128[12] 296[6])
    defparam i12670_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12841_4_lut (.I0(r_Rx_Data), .I1(rx_data[2]), .I2(n55912), 
            .I3(n27), .O(n26445));   // verilog/uart_rx.v(50[10] 145[8])
    defparam i12841_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 add_1103_16_lut (.I0(GND_net), .I1(GND_net), .I2(n9496), .I3(n46109), 
            .O(n4537)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1103_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1103_16 (.CI(n46109), .I0(GND_net), .I1(n9496), .CO(n46110));
    SB_LUT4 i12667_3_lut (.I0(\data_in_frame[4] [1]), .I1(rx_data[1]), .I2(n7_adj_5575), 
            .I3(GND_net), .O(n26271));   // verilog/coms.v(128[12] 296[6])
    defparam i12667_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 add_1103_15_lut (.I0(GND_net), .I1(GND_net), .I2(n9498), .I3(n46108), 
            .O(n4538)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1103_15_lut.LUT_INIT = 16'hC33C;
    SB_DFF commutation_state_prev_i1 (.Q(commutation_state_prev[1]), .C(clk16MHz), 
           .D(commutation_state[1]));   // verilog/TinyFPGA_B.v(131[9] 210[5])
    SB_CARRY add_1103_15 (.CI(n46108), .I0(GND_net), .I1(n9498), .CO(n46109));
    SB_LUT4 add_1103_14_lut (.I0(GND_net), .I1(GND_net), .I2(n9500), .I3(n46107), 
            .O(n4539)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1103_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1103_14 (.CI(n46107), .I0(GND_net), .I1(n9500), .CO(n46108));
    SB_LUT4 i12664_3_lut (.I0(\data_in_frame[4] [0]), .I1(rx_data[0]), .I2(n7_adj_5575), 
            .I3(GND_net), .O(n26268));   // verilog/coms.v(128[12] 296[6])
    defparam i12664_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 add_1103_13_lut (.I0(GND_net), .I1(GND_net), .I2(n9502), .I3(n46106), 
            .O(n4540)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1103_13_lut.LUT_INIT = 16'hC33C;
    SB_DFF pwm_setpoint_i23 (.Q(pwm_setpoint[23]), .C(clk16MHz), .D(pwm_setpoint_23__N_1[23]));   // verilog/TinyFPGA_B.v(92[9] 117[5])
    SB_LUT4 i12661_3_lut (.I0(\data_in_frame[3] [7]), .I1(rx_data[7]), .I2(n25157), 
            .I3(GND_net), .O(n26265));   // verilog/coms.v(128[12] 296[6])
    defparam i12661_3_lut.LUT_INIT = 16'hacac;
    SB_DFF pwm_setpoint_i22 (.Q(pwm_setpoint[22]), .C(clk16MHz), .D(pwm_setpoint_23__N_1[22]));   // verilog/TinyFPGA_B.v(92[9] 117[5])
    SB_DFF pwm_setpoint_i21 (.Q(pwm_setpoint[21]), .C(clk16MHz), .D(pwm_setpoint_23__N_1[21]));   // verilog/TinyFPGA_B.v(92[9] 117[5])
    SB_DFF pwm_setpoint_i20 (.Q(pwm_setpoint[20]), .C(clk16MHz), .D(pwm_setpoint_23__N_1[20]));   // verilog/TinyFPGA_B.v(92[9] 117[5])
    SB_DFF pwm_setpoint_i19 (.Q(pwm_setpoint[19]), .C(clk16MHz), .D(pwm_setpoint_23__N_1[19]));   // verilog/TinyFPGA_B.v(92[9] 117[5])
    SB_DFF pwm_setpoint_i18 (.Q(pwm_setpoint[18]), .C(clk16MHz), .D(pwm_setpoint_23__N_1[18]));   // verilog/TinyFPGA_B.v(92[9] 117[5])
    SB_DFF pwm_setpoint_i17 (.Q(pwm_setpoint[17]), .C(clk16MHz), .D(pwm_setpoint_23__N_1[17]));   // verilog/TinyFPGA_B.v(92[9] 117[5])
    SB_DFF pwm_setpoint_i16 (.Q(pwm_setpoint[16]), .C(clk16MHz), .D(pwm_setpoint_23__N_1[16]));   // verilog/TinyFPGA_B.v(92[9] 117[5])
    SB_DFF pwm_setpoint_i15 (.Q(pwm_setpoint[15]), .C(clk16MHz), .D(pwm_setpoint_23__N_1[15]));   // verilog/TinyFPGA_B.v(92[9] 117[5])
    SB_DFF pwm_setpoint_i14 (.Q(pwm_setpoint[14]), .C(clk16MHz), .D(pwm_setpoint_23__N_1[14]));   // verilog/TinyFPGA_B.v(92[9] 117[5])
    SB_DFF pwm_setpoint_i13 (.Q(pwm_setpoint[13]), .C(clk16MHz), .D(pwm_setpoint_23__N_1[13]));   // verilog/TinyFPGA_B.v(92[9] 117[5])
    SB_DFF pwm_setpoint_i12 (.Q(pwm_setpoint[12]), .C(clk16MHz), .D(pwm_setpoint_23__N_1[12]));   // verilog/TinyFPGA_B.v(92[9] 117[5])
    SB_DFF pwm_setpoint_i11 (.Q(pwm_setpoint[11]), .C(clk16MHz), .D(pwm_setpoint_23__N_1[11]));   // verilog/TinyFPGA_B.v(92[9] 117[5])
    SB_DFF pwm_setpoint_i10 (.Q(pwm_setpoint[10]), .C(clk16MHz), .D(pwm_setpoint_23__N_1[10]));   // verilog/TinyFPGA_B.v(92[9] 117[5])
    SB_CARRY add_1103_13 (.CI(n46106), .I0(GND_net), .I1(n9502), .CO(n46107));
    SB_DFF pwm_setpoint_i9 (.Q(pwm_setpoint[9]), .C(clk16MHz), .D(pwm_setpoint_23__N_1[9]));   // verilog/TinyFPGA_B.v(92[9] 117[5])
    SB_LUT4 n9409_bdd_4_lut_48877 (.I0(n9409), .I1(current[15]), .I2(duty[19]), 
            .I3(n9407), .O(n63647));
    defparam n9409_bdd_4_lut_48877.LUT_INIT = 16'he4aa;
    SB_DFF pwm_setpoint_i8 (.Q(pwm_setpoint[8]), .C(clk16MHz), .D(pwm_setpoint_23__N_1[8]));   // verilog/TinyFPGA_B.v(92[9] 117[5])
    SB_DFF pwm_setpoint_i7 (.Q(pwm_setpoint[7]), .C(clk16MHz), .D(pwm_setpoint_23__N_1[7]));   // verilog/TinyFPGA_B.v(92[9] 117[5])
    SB_DFF pwm_setpoint_i6 (.Q(pwm_setpoint[6]), .C(clk16MHz), .D(pwm_setpoint_23__N_1[6]));   // verilog/TinyFPGA_B.v(92[9] 117[5])
    SB_DFF pwm_setpoint_i5 (.Q(pwm_setpoint[5]), .C(clk16MHz), .D(pwm_setpoint_23__N_1[5]));   // verilog/TinyFPGA_B.v(92[9] 117[5])
    SB_DFF pwm_setpoint_i4 (.Q(pwm_setpoint[4]), .C(clk16MHz), .D(pwm_setpoint_23__N_1[4]));   // verilog/TinyFPGA_B.v(92[9] 117[5])
    SB_LUT4 n63647_bdd_4_lut (.I0(n63647), .I1(duty[16]), .I2(n4535), 
            .I3(n9407), .O(pwm_setpoint_23__N_1[16]));
    defparam n63647_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n9409_bdd_4_lut_48867 (.I0(n9409), .I1(current[15]), .I2(duty[18]), 
            .I3(n9407), .O(n63641));
    defparam n9409_bdd_4_lut_48867.LUT_INIT = 16'he4aa;
    SB_LUT4 n63641_bdd_4_lut (.I0(n63641), .I1(duty[15]), .I2(n4536), 
            .I3(n9407), .O(pwm_setpoint_23__N_1[15]));
    defparam n63641_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n9409_bdd_4_lut_48862 (.I0(n9409), .I1(current[15]), .I2(duty[17]), 
            .I3(n9407), .O(n63635));
    defparam n9409_bdd_4_lut_48862.LUT_INIT = 16'he4aa;
    SB_LUT4 add_1103_12_lut (.I0(GND_net), .I1(GND_net), .I2(n9504), .I3(n46105), 
            .O(n4541)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1103_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1103_12 (.CI(n46105), .I0(GND_net), .I1(n9504), .CO(n46106));
    SB_LUT4 add_1103_11_lut (.I0(GND_net), .I1(GND_net), .I2(n9506), .I3(n46104), 
            .O(n4542)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1103_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1103_11 (.CI(n46104), .I0(GND_net), .I1(n9506), .CO(n46105));
    SB_DFFESR delay_counter__i1 (.Q(delay_counter[1]), .C(clk16MHz), .E(n24501), 
            .D(n1078), .R(n25559));   // verilog/TinyFPGA_B.v(345[10] 375[6])
    SB_DFFESR delay_counter__i2 (.Q(delay_counter[2]), .C(clk16MHz), .E(n24501), 
            .D(n1077), .R(n25559));   // verilog/TinyFPGA_B.v(345[10] 375[6])
    SB_DFFESR delay_counter__i3 (.Q(delay_counter[3]), .C(clk16MHz), .E(n24501), 
            .D(n1076), .R(n25559));   // verilog/TinyFPGA_B.v(345[10] 375[6])
    SB_LUT4 add_1103_10_lut (.I0(GND_net), .I1(GND_net), .I2(n9508), .I3(n46103), 
            .O(n4543)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1103_10_lut.LUT_INIT = 16'hC33C;
    SB_DFFESR delay_counter__i4 (.Q(delay_counter[4]), .C(clk16MHz), .E(n24501), 
            .D(n1075), .R(n25559));   // verilog/TinyFPGA_B.v(345[10] 375[6])
    SB_DFFESR delay_counter__i5 (.Q(delay_counter[5]), .C(clk16MHz), .E(n24501), 
            .D(n1074), .R(n25559));   // verilog/TinyFPGA_B.v(345[10] 375[6])
    SB_DFFESR delay_counter__i6 (.Q(delay_counter[6]), .C(clk16MHz), .E(n24501), 
            .D(n1073), .R(n25559));   // verilog/TinyFPGA_B.v(345[10] 375[6])
    SB_DFFESR delay_counter__i7 (.Q(delay_counter[7]), .C(clk16MHz), .E(n24501), 
            .D(n1072), .R(n25559));   // verilog/TinyFPGA_B.v(345[10] 375[6])
    SB_DFFESR delay_counter__i8 (.Q(delay_counter[8]), .C(clk16MHz), .E(n24501), 
            .D(n1071), .R(n25559));   // verilog/TinyFPGA_B.v(345[10] 375[6])
    SB_DFFESR delay_counter__i9 (.Q(delay_counter[9]), .C(clk16MHz), .E(n24501), 
            .D(n1070), .R(n25559));   // verilog/TinyFPGA_B.v(345[10] 375[6])
    SB_DFFESR delay_counter__i10 (.Q(delay_counter[10]), .C(clk16MHz), .E(n24501), 
            .D(n1069), .R(n25559));   // verilog/TinyFPGA_B.v(345[10] 375[6])
    SB_DFFESR delay_counter__i11 (.Q(delay_counter[11]), .C(clk16MHz), .E(n24501), 
            .D(n1068), .R(n25559));   // verilog/TinyFPGA_B.v(345[10] 375[6])
    SB_DFFESR delay_counter__i12 (.Q(delay_counter[12]), .C(clk16MHz), .E(n24501), 
            .D(n1067), .R(n25559));   // verilog/TinyFPGA_B.v(345[10] 375[6])
    SB_DFFESR delay_counter__i13 (.Q(delay_counter[13]), .C(clk16MHz), .E(n24501), 
            .D(n1066), .R(n25559));   // verilog/TinyFPGA_B.v(345[10] 375[6])
    SB_DFFESR delay_counter__i14 (.Q(delay_counter[14]), .C(clk16MHz), .E(n24501), 
            .D(n1065), .R(n25559));   // verilog/TinyFPGA_B.v(345[10] 375[6])
    SB_DFFESR delay_counter__i15 (.Q(delay_counter[15]), .C(clk16MHz), .E(n24501), 
            .D(n1064), .R(n25559));   // verilog/TinyFPGA_B.v(345[10] 375[6])
    SB_DFFESR delay_counter__i16 (.Q(delay_counter[16]), .C(clk16MHz), .E(n24501), 
            .D(n1063), .R(n25559));   // verilog/TinyFPGA_B.v(345[10] 375[6])
    SB_DFFESR delay_counter__i17 (.Q(delay_counter[17]), .C(clk16MHz), .E(n24501), 
            .D(n1062), .R(n25559));   // verilog/TinyFPGA_B.v(345[10] 375[6])
    SB_DFFESR delay_counter__i18 (.Q(delay_counter[18]), .C(clk16MHz), .E(n24501), 
            .D(n1061), .R(n25559));   // verilog/TinyFPGA_B.v(345[10] 375[6])
    SB_DFFESR delay_counter__i19 (.Q(delay_counter[19]), .C(clk16MHz), .E(n24501), 
            .D(n1060), .R(n25559));   // verilog/TinyFPGA_B.v(345[10] 375[6])
    SB_DFFESR delay_counter__i20 (.Q(delay_counter[20]), .C(clk16MHz), .E(n24501), 
            .D(n1059), .R(n25559));   // verilog/TinyFPGA_B.v(345[10] 375[6])
    SB_DFFESR delay_counter__i21 (.Q(delay_counter[21]), .C(clk16MHz), .E(n24501), 
            .D(n1058), .R(n25559));   // verilog/TinyFPGA_B.v(345[10] 375[6])
    SB_DFFESR delay_counter__i22 (.Q(delay_counter[22]), .C(clk16MHz), .E(n24501), 
            .D(n1057), .R(n25559));   // verilog/TinyFPGA_B.v(345[10] 375[6])
    SB_DFFESR delay_counter__i23 (.Q(delay_counter[23]), .C(clk16MHz), .E(n24501), 
            .D(n1056), .R(n25559));   // verilog/TinyFPGA_B.v(345[10] 375[6])
    SB_DFFESR delay_counter__i24 (.Q(delay_counter[24]), .C(clk16MHz), .E(n24501), 
            .D(n1055), .R(n25559));   // verilog/TinyFPGA_B.v(345[10] 375[6])
    SB_DFFESR delay_counter__i25 (.Q(delay_counter[25]), .C(clk16MHz), .E(n24501), 
            .D(n1054), .R(n25559));   // verilog/TinyFPGA_B.v(345[10] 375[6])
    SB_DFFESR delay_counter__i26 (.Q(delay_counter[26]), .C(clk16MHz), .E(n24501), 
            .D(n1053), .R(n25559));   // verilog/TinyFPGA_B.v(345[10] 375[6])
    SB_DFFESR delay_counter__i27 (.Q(delay_counter[27]), .C(clk16MHz), .E(n24501), 
            .D(n1052), .R(n25559));   // verilog/TinyFPGA_B.v(345[10] 375[6])
    SB_DFFESR delay_counter__i28 (.Q(delay_counter[28]), .C(clk16MHz), .E(n24501), 
            .D(n1051), .R(n25559));   // verilog/TinyFPGA_B.v(345[10] 375[6])
    SB_DFFESR delay_counter__i29 (.Q(delay_counter[29]), .C(clk16MHz), .E(n24501), 
            .D(n1050), .R(n25559));   // verilog/TinyFPGA_B.v(345[10] 375[6])
    SB_DFFESR delay_counter__i30 (.Q(delay_counter[30]), .C(clk16MHz), .E(n24501), 
            .D(n1049), .R(n25559));   // verilog/TinyFPGA_B.v(345[10] 375[6])
    SB_DFFESR delay_counter__i31 (.Q(delay_counter[31]), .C(clk16MHz), .E(n24501), 
            .D(n1048), .R(n25559));   // verilog/TinyFPGA_B.v(345[10] 375[6])
    SB_DFF read_189 (.Q(read), .C(clk16MHz), .D(n55525));   // verilog/TinyFPGA_B.v(345[10] 375[6])
    SB_CARRY add_1103_10 (.CI(n46103), .I0(GND_net), .I1(n9508), .CO(n46104));
    SB_LUT4 add_1103_9_lut (.I0(GND_net), .I1(GND_net), .I2(n9510), .I3(n46102), 
            .O(n4544)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1103_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_146_10 (.CI(n46026), .I0(delay_counter[8]), .I1(GND_net), 
            .CO(n46027));
    SB_LUT4 n63635_bdd_4_lut (.I0(n63635), .I1(duty[14]), .I2(n4537), 
            .I3(n9407), .O(pwm_setpoint_23__N_1[14]));
    defparam n63635_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n9409_bdd_4_lut_48857 (.I0(n9409), .I1(current[15]), .I2(duty[16]), 
            .I3(n9407), .O(n63629));
    defparam n9409_bdd_4_lut_48857.LUT_INIT = 16'he4aa;
    SB_LUT4 n63629_bdd_4_lut (.I0(n63629), .I1(duty[13]), .I2(n4538), 
            .I3(n9407), .O(pwm_setpoint_23__N_1[13]));
    defparam n63629_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n9409_bdd_4_lut_48852 (.I0(n9409), .I1(current[15]), .I2(duty[15]), 
            .I3(n9407), .O(n63623));
    defparam n9409_bdd_4_lut_48852.LUT_INIT = 16'he4aa;
    SB_LUT4 n63623_bdd_4_lut (.I0(n63623), .I1(duty[12]), .I2(n4539), 
            .I3(n9407), .O(pwm_setpoint_23__N_1[12]));
    defparam n63623_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n9409_bdd_4_lut_48847 (.I0(n9409), .I1(current[11]), .I2(duty[14]), 
            .I3(n9407), .O(n63617));
    defparam n9409_bdd_4_lut_48847.LUT_INIT = 16'he4aa;
    SB_LUT4 n63617_bdd_4_lut (.I0(n63617), .I1(duty[11]), .I2(n4540), 
            .I3(n9407), .O(pwm_setpoint_23__N_1[11]));
    defparam n63617_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_CARRY add_1103_9 (.CI(n46102), .I0(GND_net), .I1(n9510), .CO(n46103));
    SB_LUT4 add_1103_8_lut (.I0(GND_net), .I1(GND_net), .I2(n9512), .I3(n46101), 
            .O(n4545)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1103_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 n9409_bdd_4_lut_48842 (.I0(n9409), .I1(current[10]), .I2(duty[13]), 
            .I3(n9407), .O(n63599));
    defparam n9409_bdd_4_lut_48842.LUT_INIT = 16'he4aa;
    SB_CARRY add_146_27 (.CI(n46043), .I0(delay_counter[25]), .I1(GND_net), 
            .CO(n46044));
    SB_CARRY add_1103_8 (.CI(n46101), .I0(GND_net), .I1(n9512), .CO(n46102));
    SB_LUT4 n63599_bdd_4_lut (.I0(n63599), .I1(duty[10]), .I2(n4541), 
            .I3(n9407), .O(pwm_setpoint_23__N_1[10]));
    defparam n63599_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 add_1103_7_lut (.I0(GND_net), .I1(GND_net), .I2(n9514), .I3(n46100), 
            .O(n4546)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1103_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_146_4 (.CI(n46020), .I0(delay_counter[2]), .I1(GND_net), 
            .CO(n46021));
    SB_CARRY add_1103_7 (.CI(n46100), .I0(GND_net), .I1(n9514), .CO(n46101));
    SB_LUT4 add_1103_6_lut (.I0(GND_net), .I1(GND_net), .I2(n9516), .I3(n46099), 
            .O(n4547)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1103_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 n9409_bdd_4_lut_48827 (.I0(n9409), .I1(current[9]), .I2(duty[12]), 
            .I3(n9407), .O(n63593));
    defparam n9409_bdd_4_lut_48827.LUT_INIT = 16'he4aa;
    SB_LUT4 n63593_bdd_4_lut (.I0(n63593), .I1(duty[9]), .I2(n4542), .I3(n9407), 
            .O(pwm_setpoint_23__N_1[9]));
    defparam n63593_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 add_146_9_lut (.I0(GND_net), .I1(delay_counter[7]), .I2(GND_net), 
            .I3(n46025), .O(n1072)) /* synthesis syn_instantiated=1 */ ;
    defparam add_146_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i45821_3_lut_4_lut (.I0(r_Clock_Count_adj_5650[3]), .I1(o_Rx_DV_N_3261[3]), 
            .I2(o_Rx_DV_N_3261[2]), .I3(r_Clock_Count_adj_5650[2]), .O(n60533));   // verilog/uart_tx.v(117[17:57])
    defparam i45821_3_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 LessThan_1094_i6_3_lut_3_lut (.I0(r_Clock_Count_adj_5650[3]), 
            .I1(o_Rx_DV_N_3261[3]), .I2(o_Rx_DV_N_3261[2]), .I3(GND_net), 
            .O(n6_adj_5548));   // verilog/uart_tx.v(117[17:57])
    defparam LessThan_1094_i6_3_lut_3_lut.LUT_INIT = 16'hd4d4;
    SB_LUT4 add_146_26_lut (.I0(GND_net), .I1(delay_counter[24]), .I2(GND_net), 
            .I3(n46042), .O(n1055)) /* synthesis syn_instantiated=1 */ ;
    defparam add_146_26_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i10_3_lut (.I0(n240), .I1(n292), .I2(n284), .I3(GND_net), 
            .O(n6_adj_5526));
    defparam i10_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i6_3_lut (.I0(n6_adj_5526), .I1(IntegralLimit[17]), .I2(n258), 
            .I3(GND_net), .O(n31535));
    defparam i6_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_adj_1686 (.I0(n31535), .I1(Ki[0]), .I2(GND_net), 
            .I3(GND_net), .O(n53));
    defparam i1_2_lut_adj_1686.LUT_INIT = 16'h8888;
    SB_LUT4 n9409_bdd_4_lut_48822 (.I0(n9409), .I1(current[8]), .I2(duty[11]), 
            .I3(n9407), .O(n63587));
    defparam n9409_bdd_4_lut_48822.LUT_INIT = 16'he4aa;
    SB_CARRY add_1103_6 (.CI(n46099), .I0(GND_net), .I1(n9516), .CO(n46100));
    SB_LUT4 add_1103_5_lut (.I0(GND_net), .I1(GND_net), .I2(n9518), .I3(n46098), 
            .O(n4548)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1103_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1103_5 (.CI(n46098), .I0(GND_net), .I1(n9518), .CO(n46099));
    SB_LUT4 n63587_bdd_4_lut (.I0(n63587), .I1(duty[8]), .I2(n4543), .I3(n9407), 
            .O(pwm_setpoint_23__N_1[8]));
    defparam n63587_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFFESR delay_counter__i0 (.Q(delay_counter[0]), .C(clk16MHz), .E(n24501), 
            .D(n1079), .R(n25559));   // verilog/TinyFPGA_B.v(345[10] 375[6])
    SB_DFFESR GHC_187 (.Q(GHC), .C(clk16MHz), .E(n24487), .D(GHC_N_343), 
            .R(n25556));   // verilog/TinyFPGA_B.v(131[9] 210[5])
    SB_DFFESR GHB_185 (.Q(GHB), .C(clk16MHz), .E(n24487), .D(GHB_N_329), 
            .R(n25556));   // verilog/TinyFPGA_B.v(131[9] 210[5])
    SB_DFFESR GHA_183 (.Q(GHA), .C(clk16MHz), .E(n24487), .D(GHA_N_307), 
            .R(n25556));   // verilog/TinyFPGA_B.v(131[9] 210[5])
    SB_DFFESS commutation_state_i0 (.Q(commutation_state[0]), .C(clk16MHz), 
            .E(n6_adj_5577), .D(commutation_state_7__N_160[0]), .S(commutation_state_7__N_168));   // verilog/TinyFPGA_B.v(131[9] 210[5])
    SB_DFFESR GLA_184 (.Q(INLA_c_0), .C(clk16MHz), .E(n24487), .D(GLA_N_324), 
            .R(n25556));   // verilog/TinyFPGA_B.v(131[9] 210[5])
    SB_DFFESR GLB_186 (.Q(INLB_c_0), .C(clk16MHz), .E(n24487), .D(GLB_N_338), 
            .R(n25556));   // verilog/TinyFPGA_B.v(131[9] 210[5])
    SB_DFFESR GLC_188 (.Q(INLC_c_0), .C(clk16MHz), .E(n24487), .D(GLC_N_352), 
            .R(n25556));   // verilog/TinyFPGA_B.v(131[9] 210[5])
    GND i1 (.Y(GND_net));
    SB_CARRY add_146_26 (.CI(n46042), .I0(delay_counter[24]), .I1(GND_net), 
            .CO(n46043));
    SB_CARRY add_146_9 (.CI(n46025), .I0(delay_counter[7]), .I1(GND_net), 
            .CO(n46026));
    SB_LUT4 n9409_bdd_4_lut_48817 (.I0(n9409), .I1(current[7]), .I2(duty[10]), 
            .I3(n9407), .O(n63581));
    defparam n9409_bdd_4_lut_48817.LUT_INIT = 16'he4aa;
    SB_LUT4 n63581_bdd_4_lut (.I0(n63581), .I1(duty[7]), .I2(n4544), .I3(n9407), 
            .O(pwm_setpoint_23__N_1[7]));
    defparam n63581_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 add_1103_4_lut (.I0(GND_net), .I1(GND_net), .I2(n9520), .I3(n46097), 
            .O(n4549)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1103_4_lut.LUT_INIT = 16'hC33C;
    SB_DFF commutation_state_i2 (.Q(commutation_state[2]), .C(clk16MHz), 
           .D(n53662));   // verilog/TinyFPGA_B.v(131[9] 210[5])
    SB_LUT4 add_146_25_lut (.I0(GND_net), .I1(delay_counter[23]), .I2(GND_net), 
            .I3(n46041), .O(n1056)) /* synthesis syn_instantiated=1 */ ;
    defparam add_146_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1103_4 (.CI(n46097), .I0(GND_net), .I1(n9520), .CO(n46098));
    SB_LUT4 add_1103_3_lut (.I0(GND_net), .I1(GND_net), .I2(n9522), .I3(n46096), 
            .O(n4550)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1103_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1103_3 (.CI(n46096), .I0(GND_net), .I1(n9522), .CO(n46097));
    SB_LUT4 add_1103_2_lut (.I0(GND_net), .I1(GND_net), .I2(n9470), .I3(VCC_net), 
            .O(n4551)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1103_2_lut.LUT_INIT = 16'hC33C;
    SB_DFF commutation_state_prev_i0 (.Q(commutation_state_prev[0]), .C(clk16MHz), 
           .D(commutation_state[0]));   // verilog/TinyFPGA_B.v(131[9] 210[5])
    SB_DFF reset_190 (.Q(reset), .C(clk16MHz), .D(n51303));   // verilog/TinyFPGA_B.v(345[10] 375[6])
    SB_CARRY add_146_25 (.CI(n46041), .I0(delay_counter[23]), .I1(GND_net), 
            .CO(n46042));
    SB_LUT4 add_146_24_lut (.I0(GND_net), .I1(delay_counter[22]), .I2(GND_net), 
            .I3(n46040), .O(n1057)) /* synthesis syn_instantiated=1 */ ;
    defparam add_146_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1103_2 (.CI(VCC_net), .I0(GND_net), .I1(n9470), .CO(n46096));
    SB_CARRY add_146_24 (.CI(n46040), .I0(delay_counter[22]), .I1(GND_net), 
            .CO(n46041));
    SB_LUT4 add_146_23_lut (.I0(GND_net), .I1(delay_counter[21]), .I2(GND_net), 
            .I3(n46039), .O(n1058)) /* synthesis syn_instantiated=1 */ ;
    defparam add_146_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_146_3_lut (.I0(GND_net), .I1(delay_counter[1]), .I2(GND_net), 
            .I3(n46019), .O(n1078)) /* synthesis syn_instantiated=1 */ ;
    defparam add_146_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_146_23 (.CI(n46039), .I0(delay_counter[21]), .I1(GND_net), 
            .CO(n46040));
    SB_LUT4 add_146_22_lut (.I0(GND_net), .I1(delay_counter[20]), .I2(GND_net), 
            .I3(n46038), .O(n1059)) /* synthesis syn_instantiated=1 */ ;
    defparam add_146_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_146_22 (.CI(n46038), .I0(delay_counter[20]), .I1(GND_net), 
            .CO(n46039));
    SB_LUT4 add_146_8_lut (.I0(GND_net), .I1(delay_counter[6]), .I2(GND_net), 
            .I3(n46024), .O(n1073)) /* synthesis syn_instantiated=1 */ ;
    defparam add_146_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_16_add_3_15_lut (.I0(GND_net), .I1(GND_net), .I2(n2), 
            .I3(n46254), .O(n293)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_16_add_3_14_lut (.I0(GND_net), .I1(GND_net), .I2(n2), 
            .I3(n46253), .O(n297)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_14 (.CI(n46253), .I0(GND_net), .I1(n2), 
            .CO(n46254));
    SB_LUT4 add_146_21_lut (.I0(GND_net), .I1(delay_counter[19]), .I2(GND_net), 
            .I3(n46037), .O(n1060)) /* synthesis syn_instantiated=1 */ ;
    defparam add_146_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_16_add_3_13_lut (.I0(GND_net), .I1(GND_net), .I2(n14), 
            .I3(n46252), .O(n298)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_13 (.CI(n46252), .I0(GND_net), .I1(n14), 
            .CO(n46253));
    SB_LUT4 unary_minus_16_add_3_12_lut (.I0(GND_net), .I1(GND_net), .I2(n15_adj_5464), 
            .I3(n46251), .O(n299)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_12 (.CI(n46251), .I0(GND_net), .I1(n15_adj_5464), 
            .CO(n46252));
    SB_LUT4 unary_minus_16_add_3_11_lut (.I0(GND_net), .I1(GND_net), .I2(n16_adj_5465), 
            .I3(n46250), .O(n300)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_11 (.CI(n46250), .I0(GND_net), .I1(n16_adj_5465), 
            .CO(n46251));
    SB_LUT4 unary_minus_16_add_3_10_lut (.I0(GND_net), .I1(GND_net), .I2(n17_adj_5466), 
            .I3(n46249), .O(n301)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_10 (.CI(n46249), .I0(GND_net), .I1(n17_adj_5466), 
            .CO(n46250));
    SB_LUT4 unary_minus_16_add_3_9_lut (.I0(GND_net), .I1(GND_net), .I2(n18), 
            .I3(n46248), .O(n302)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_9 (.CI(n46248), .I0(GND_net), .I1(n18), 
            .CO(n46249));
    SB_LUT4 unary_minus_16_add_3_8_lut (.I0(GND_net), .I1(GND_net), .I2(n19_adj_5467), 
            .I3(n46247), .O(n303)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_8 (.CI(n46247), .I0(GND_net), .I1(n19_adj_5467), 
            .CO(n46248));
    SB_LUT4 unary_minus_16_add_3_7_lut (.I0(GND_net), .I1(GND_net), .I2(n20), 
            .I3(n46246), .O(n304)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_7 (.CI(n46246), .I0(GND_net), .I1(n20), 
            .CO(n46247));
    SB_LUT4 unary_minus_16_add_3_6_lut (.I0(GND_net), .I1(GND_net), .I2(n21), 
            .I3(n46245), .O(n305)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_6 (.CI(n46245), .I0(GND_net), .I1(n21), 
            .CO(n46246));
    SB_LUT4 unary_minus_16_add_3_5_lut (.I0(GND_net), .I1(GND_net), .I2(n22), 
            .I3(n46244), .O(n306)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_5 (.CI(n46244), .I0(GND_net), .I1(n22), 
            .CO(n46245));
    SB_LUT4 unary_minus_16_add_3_4_lut (.I0(GND_net), .I1(GND_net), .I2(n23), 
            .I3(n46243), .O(n307)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_4 (.CI(n46243), .I0(GND_net), .I1(n23), 
            .CO(n46244));
    SB_LUT4 dti_counter_1934_add_4_9_lut (.I0(GND_net), .I1(VCC_net), .I2(dti_counter[7]), 
            .I3(n46520), .O(n38)) /* synthesis syn_instantiated=1 */ ;
    defparam dti_counter_1934_add_4_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 dti_counter_1934_add_4_8_lut (.I0(GND_net), .I1(VCC_net), .I2(dti_counter[6]), 
            .I3(n46519), .O(n39)) /* synthesis syn_instantiated=1 */ ;
    defparam dti_counter_1934_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_16_add_3_3_lut (.I0(GND_net), .I1(GND_net), .I2(n24), 
            .I3(n46242), .O(n308)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_3 (.CI(n46242), .I0(GND_net), .I1(n24), 
            .CO(n46243));
    SB_CARRY dti_counter_1934_add_4_8 (.CI(n46519), .I0(VCC_net), .I1(dti_counter[6]), 
            .CO(n46520));
    SB_LUT4 unary_minus_16_add_3_2_lut (.I0(n35713), .I1(GND_net), .I2(n25), 
            .I3(VCC_net), .O(n59720)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_2_lut.LUT_INIT = 16'h8228;
    SB_CARRY unary_minus_16_add_3_2 (.CI(VCC_net), .I0(GND_net), .I1(n25), 
            .CO(n46242));
    SB_LUT4 dti_counter_1934_add_4_7_lut (.I0(GND_net), .I1(VCC_net), .I2(dti_counter[5]), 
            .I3(n46518), .O(n40)) /* synthesis syn_instantiated=1 */ ;
    defparam dti_counter_1934_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY dti_counter_1934_add_4_7 (.CI(n46518), .I0(VCC_net), .I1(dti_counter[5]), 
            .CO(n46519));
    SB_LUT4 dti_counter_1934_add_4_6_lut (.I0(GND_net), .I1(VCC_net), .I2(dti_counter[4]), 
            .I3(n46517), .O(n41)) /* synthesis syn_instantiated=1 */ ;
    defparam dti_counter_1934_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY dti_counter_1934_add_4_6 (.CI(n46517), .I0(VCC_net), .I1(dti_counter[4]), 
            .CO(n46518));
    SB_LUT4 dti_counter_1934_add_4_5_lut (.I0(GND_net), .I1(VCC_net), .I2(dti_counter[3]), 
            .I3(n46516), .O(n42)) /* synthesis syn_instantiated=1 */ ;
    defparam dti_counter_1934_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY dti_counter_1934_add_4_5 (.CI(n46516), .I0(VCC_net), .I1(dti_counter[3]), 
            .CO(n46517));
    SB_LUT4 dti_counter_1934_add_4_4_lut (.I0(GND_net), .I1(VCC_net), .I2(dti_counter[2]), 
            .I3(n46515), .O(n43)) /* synthesis syn_instantiated=1 */ ;
    defparam dti_counter_1934_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY dti_counter_1934_add_4_4 (.CI(n46515), .I0(VCC_net), .I1(dti_counter[2]), 
            .CO(n46516));
    SB_LUT4 dti_counter_1934_add_4_3_lut (.I0(GND_net), .I1(VCC_net), .I2(dti_counter[1]), 
            .I3(n46514), .O(n44)) /* synthesis syn_instantiated=1 */ ;
    defparam dti_counter_1934_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY dti_counter_1934_add_4_3 (.CI(n46514), .I0(VCC_net), .I1(dti_counter[1]), 
            .CO(n46515));
    SB_LUT4 dti_counter_1934_add_4_2_lut (.I0(GND_net), .I1(GND_net), .I2(dti_counter[0]), 
            .I3(VCC_net), .O(n45)) /* synthesis syn_instantiated=1 */ ;
    defparam dti_counter_1934_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY dti_counter_1934_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(dti_counter[0]), 
            .CO(n46514));
    SB_CARRY add_146_3 (.CI(n46019), .I0(delay_counter[1]), .I1(GND_net), 
            .CO(n46020));
    SB_CARRY add_146_8 (.CI(n46024), .I0(delay_counter[6]), .I1(GND_net), 
            .CO(n46025));
    SB_CARRY add_146_21 (.CI(n46037), .I0(delay_counter[19]), .I1(GND_net), 
            .CO(n46038));
    SB_LUT4 add_146_20_lut (.I0(GND_net), .I1(delay_counter[18]), .I2(GND_net), 
            .I3(n46036), .O(n1061)) /* synthesis syn_instantiated=1 */ ;
    defparam add_146_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_146_20 (.CI(n46036), .I0(delay_counter[18]), .I1(GND_net), 
            .CO(n46037));
    SB_LUT4 add_146_19_lut (.I0(GND_net), .I1(delay_counter[17]), .I2(GND_net), 
            .I3(n46035), .O(n1062)) /* synthesis syn_instantiated=1 */ ;
    defparam add_146_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_146_19 (.CI(n46035), .I0(delay_counter[17]), .I1(GND_net), 
            .CO(n46036));
    SB_LUT4 add_146_7_lut (.I0(GND_net), .I1(delay_counter[5]), .I2(GND_net), 
            .I3(n46023), .O(n1074)) /* synthesis syn_instantiated=1 */ ;
    defparam add_146_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_146_18_lut (.I0(GND_net), .I1(delay_counter[16]), .I2(GND_net), 
            .I3(n46034), .O(n1063)) /* synthesis syn_instantiated=1 */ ;
    defparam add_146_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_146_18 (.CI(n46034), .I0(delay_counter[16]), .I1(GND_net), 
            .CO(n46035));
    SB_LUT4 add_146_17_lut (.I0(GND_net), .I1(delay_counter[15]), .I2(GND_net), 
            .I3(n46033), .O(n1064)) /* synthesis syn_instantiated=1 */ ;
    defparam add_146_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_146_7 (.CI(n46023), .I0(delay_counter[5]), .I1(GND_net), 
            .CO(n46024));
    SB_LUT4 add_146_2_lut (.I0(GND_net), .I1(delay_counter[0]), .I2(GND_net), 
            .I3(VCC_net), .O(n1079)) /* synthesis syn_instantiated=1 */ ;
    defparam add_146_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_146_17 (.CI(n46033), .I0(delay_counter[15]), .I1(GND_net), 
            .CO(n46034));
    SB_LUT4 add_146_16_lut (.I0(GND_net), .I1(delay_counter[14]), .I2(GND_net), 
            .I3(n46032), .O(n1065)) /* synthesis syn_instantiated=1 */ ;
    defparam add_146_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_146_6_lut (.I0(GND_net), .I1(delay_counter[4]), .I2(GND_net), 
            .I3(n46022), .O(n1075)) /* synthesis syn_instantiated=1 */ ;
    defparam add_146_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_146_16 (.CI(n46032), .I0(delay_counter[14]), .I1(GND_net), 
            .CO(n46033));
    SB_CARRY add_146_2 (.CI(VCC_net), .I0(delay_counter[0]), .I1(GND_net), 
            .CO(n46019));
    SB_CARRY add_146_6 (.CI(n46022), .I0(delay_counter[4]), .I1(GND_net), 
            .CO(n46023));
    SB_LUT4 add_146_15_lut (.I0(GND_net), .I1(delay_counter[13]), .I2(GND_net), 
            .I3(n46031), .O(n1066)) /* synthesis syn_instantiated=1 */ ;
    defparam add_146_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_146_15 (.CI(n46031), .I0(delay_counter[13]), .I1(GND_net), 
            .CO(n46032));
    SB_LUT4 add_146_14_lut (.I0(GND_net), .I1(delay_counter[12]), .I2(GND_net), 
            .I3(n46030), .O(n1067)) /* synthesis syn_instantiated=1 */ ;
    defparam add_146_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 n9409_bdd_4_lut_48812 (.I0(n9409), .I1(current[6]), .I2(duty[9]), 
            .I3(n9407), .O(n63575));
    defparam n9409_bdd_4_lut_48812.LUT_INIT = 16'he4aa;
    SB_LUT4 i12311_2_lut_4_lut (.I0(commutation_state[0]), .I1(n4_adj_5471), 
            .I2(commutation_state_prev[0]), .I3(n35258), .O(n25915));   // verilog/TinyFPGA_B.v(134[7:48])
    defparam i12311_2_lut_4_lut.LUT_INIT = 16'h00de;
    SB_LUT4 i1_2_lut_4_lut (.I0(commutation_state[0]), .I1(n4_adj_5471), 
            .I2(commutation_state_prev[0]), .I3(n35258), .O(n24669));   // verilog/TinyFPGA_B.v(134[7:48])
    defparam i1_2_lut_4_lut.LUT_INIT = 16'hffde;
    SB_LUT4 i1_2_lut_4_lut_adj_1687 (.I0(commutation_state[0]), .I1(n4_adj_5471), 
            .I2(commutation_state_prev[0]), .I3(dti_N_356), .O(n24463));   // verilog/TinyFPGA_B.v(134[7:48])
    defparam i1_2_lut_4_lut_adj_1687.LUT_INIT = 16'hdeff;
    SB_LUT4 RX_I_0_1_lut (.I0(RX_c), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(RX_N_42));   // verilog/TinyFPGA_B.v(250[11:14])
    defparam RX_I_0_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1_4_lut_adj_1688 (.I0(o_Rx_DV_N_3261[12]), .I1(n4834), .I2(o_Rx_DV_N_3261[8]), 
            .I3(n55461), .O(n55808));
    defparam i1_4_lut_adj_1688.LUT_INIT = 16'hfeff;
    SB_LUT4 i1_4_lut_adj_1689 (.I0(o_Rx_DV_N_3261[24]), .I1(n29), .I2(n23_adj_5576), 
            .I3(n55808), .O(n55814));
    defparam i1_4_lut_adj_1689.LUT_INIT = 16'hfffe;
    SB_LUT4 n63575_bdd_4_lut (.I0(n63575), .I1(duty[6]), .I2(n4545), .I3(n9407), 
            .O(pwm_setpoint_23__N_1[6]));
    defparam n63575_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i46132_4_lut (.I0(\data_out_frame[26] [6]), .I1(n24840), .I2(\data_out_frame[27] [6]), 
            .I3(byte_transmit_counter[0]), .O(n59928));   // verilog/coms.v(103[12:33])
    defparam i46132_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i45905_2_lut (.I0(byte_transmit_counter[0]), .I1(byte_transmit_counter[2]), 
            .I2(GND_net), .I3(GND_net), .O(n59927));   // verilog/coms.v(103[12:33])
    defparam i45905_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 n9409_bdd_4_lut_48807 (.I0(n9409), .I1(current[5]), .I2(duty[8]), 
            .I3(n9407), .O(n63569));
    defparam n9409_bdd_4_lut_48807.LUT_INIT = 16'he4aa;
    SB_LUT4 n63569_bdd_4_lut (.I0(n63569), .I1(duty[5]), .I2(n4546), .I3(n9407), 
            .O(pwm_setpoint_23__N_1[5]));
    defparam n63569_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n9409_bdd_4_lut_48802 (.I0(n9409), .I1(current[4]), .I2(duty[7]), 
            .I3(n9407), .O(n63563));
    defparam n9409_bdd_4_lut_48802.LUT_INIT = 16'he4aa;
    SB_LUT4 n63563_bdd_4_lut (.I0(n63563), .I1(duty[4]), .I2(n4547), .I3(n9407), 
            .O(pwm_setpoint_23__N_1[4]));
    defparam n63563_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 mux_235_i1_4_lut (.I0(encoder0_position[0]), .I1(encoder1_position[0]), 
            .I2(n15), .I3(n15_adj_5475), .O(motor_state[0]));   // verilog/TinyFPGA_B.v(271[5] 274[10])
    defparam mux_235_i1_4_lut.LUT_INIT = 16'hf535;
    SB_LUT4 i21723_4_lut (.I0(encoder0_position[1]), .I1(encoder1_position[1]), 
            .I2(n15), .I3(n15_adj_5475), .O(n1));
    defparam i21723_4_lut.LUT_INIT = 16'hf535;
    SB_LUT4 mux_235_i3_4_lut (.I0(encoder0_position[2]), .I1(encoder1_position[2]), 
            .I2(n15), .I3(n15_adj_5475), .O(motor_state[2]));   // verilog/TinyFPGA_B.v(271[5] 274[10])
    defparam mux_235_i3_4_lut.LUT_INIT = 16'hf535;
    SB_LUT4 mux_235_i4_4_lut (.I0(encoder0_position[3]), .I1(encoder1_position[3]), 
            .I2(n15), .I3(n15_adj_5475), .O(motor_state[3]));   // verilog/TinyFPGA_B.v(271[5] 274[10])
    defparam mux_235_i4_4_lut.LUT_INIT = 16'hf535;
    SB_LUT4 mux_235_i5_4_lut (.I0(encoder0_position[4]), .I1(encoder1_position[4]), 
            .I2(n15), .I3(n15_adj_5475), .O(motor_state[4]));   // verilog/TinyFPGA_B.v(271[5] 274[10])
    defparam mux_235_i5_4_lut.LUT_INIT = 16'hf535;
    SB_LUT4 mux_235_i6_4_lut (.I0(encoder0_position[5]), .I1(encoder1_position[5]), 
            .I2(n15), .I3(n15_adj_5475), .O(motor_state[5]));   // verilog/TinyFPGA_B.v(271[5] 274[10])
    defparam mux_235_i6_4_lut.LUT_INIT = 16'hf535;
    SB_LUT4 mux_235_i8_4_lut (.I0(encoder0_position[7]), .I1(encoder1_position[7]), 
            .I2(n15), .I3(n15_adj_5475), .O(motor_state[7]));   // verilog/TinyFPGA_B.v(271[5] 274[10])
    defparam mux_235_i8_4_lut.LUT_INIT = 16'hf535;
    SB_LUT4 mux_235_i9_4_lut (.I0(encoder0_position[8]), .I1(encoder1_position[8]), 
            .I2(n15), .I3(n15_adj_5475), .O(motor_state[8]));   // verilog/TinyFPGA_B.v(271[5] 274[10])
    defparam mux_235_i9_4_lut.LUT_INIT = 16'hf535;
    SB_LUT4 mux_235_i10_4_lut (.I0(encoder0_position[9]), .I1(encoder1_position[9]), 
            .I2(n15), .I3(n15_adj_5475), .O(motor_state[9]));   // verilog/TinyFPGA_B.v(271[5] 274[10])
    defparam mux_235_i10_4_lut.LUT_INIT = 16'hf535;
    SB_LUT4 mux_235_i11_4_lut (.I0(encoder0_position[10]), .I1(encoder1_position[10]), 
            .I2(n15), .I3(n15_adj_5475), .O(motor_state[10]));   // verilog/TinyFPGA_B.v(271[5] 274[10])
    defparam mux_235_i11_4_lut.LUT_INIT = 16'hf535;
    SB_LUT4 i21698_4_lut (.I0(encoder0_position[11]), .I1(encoder1_position[11]), 
            .I2(n15), .I3(n15_adj_5475), .O(n35211));
    defparam i21698_4_lut.LUT_INIT = 16'hf535;
    SB_LUT4 mux_235_i13_4_lut (.I0(encoder0_position[12]), .I1(encoder1_position[12]), 
            .I2(n15), .I3(n15_adj_5475), .O(motor_state[12]));   // verilog/TinyFPGA_B.v(271[5] 274[10])
    defparam mux_235_i13_4_lut.LUT_INIT = 16'hf535;
    SB_LUT4 mux_235_i14_4_lut (.I0(encoder0_position[13]), .I1(encoder1_position[13]), 
            .I2(n15), .I3(n15_adj_5475), .O(motor_state[13]));   // verilog/TinyFPGA_B.v(271[5] 274[10])
    defparam mux_235_i14_4_lut.LUT_INIT = 16'hf535;
    SB_LUT4 mux_235_i15_4_lut (.I0(encoder0_position[14]), .I1(encoder1_position[14]), 
            .I2(n15), .I3(n15_adj_5475), .O(motor_state[14]));   // verilog/TinyFPGA_B.v(271[5] 274[10])
    defparam mux_235_i15_4_lut.LUT_INIT = 16'hf535;
    SB_LUT4 mux_235_i16_4_lut (.I0(encoder0_position[15]), .I1(encoder1_position[15]), 
            .I2(n15), .I3(n15_adj_5475), .O(motor_state[15]));   // verilog/TinyFPGA_B.v(271[5] 274[10])
    defparam mux_235_i16_4_lut.LUT_INIT = 16'hf535;
    SB_LUT4 mux_235_i17_4_lut (.I0(encoder0_position[16]), .I1(encoder1_position[16]), 
            .I2(n15), .I3(n15_adj_5475), .O(motor_state[16]));   // verilog/TinyFPGA_B.v(271[5] 274[10])
    defparam mux_235_i17_4_lut.LUT_INIT = 16'hf535;
    SB_LUT4 mux_235_i18_4_lut (.I0(encoder0_position[17]), .I1(encoder1_position[17]), 
            .I2(n15), .I3(n15_adj_5475), .O(motor_state[17]));   // verilog/TinyFPGA_B.v(271[5] 274[10])
    defparam mux_235_i18_4_lut.LUT_INIT = 16'hf535;
    SB_LUT4 mux_235_i19_4_lut (.I0(encoder0_position[18]), .I1(encoder1_position[18]), 
            .I2(n15), .I3(n15_adj_5475), .O(motor_state[18]));   // verilog/TinyFPGA_B.v(271[5] 274[10])
    defparam mux_235_i19_4_lut.LUT_INIT = 16'hf535;
    SB_LUT4 mux_235_i20_4_lut (.I0(encoder0_position[19]), .I1(encoder1_position[19]), 
            .I2(n15), .I3(n15_adj_5475), .O(motor_state[19]));   // verilog/TinyFPGA_B.v(271[5] 274[10])
    defparam mux_235_i20_4_lut.LUT_INIT = 16'hf535;
    SB_LUT4 mux_235_i21_4_lut (.I0(encoder0_position[20]), .I1(encoder1_position[20]), 
            .I2(n15), .I3(n15_adj_5475), .O(motor_state[20]));   // verilog/TinyFPGA_B.v(271[5] 274[10])
    defparam mux_235_i21_4_lut.LUT_INIT = 16'hf535;
    SB_LUT4 mux_235_i22_4_lut (.I0(encoder0_position[21]), .I1(encoder1_position[21]), 
            .I2(n15), .I3(n15_adj_5475), .O(motor_state[21]));   // verilog/TinyFPGA_B.v(271[5] 274[10])
    defparam mux_235_i22_4_lut.LUT_INIT = 16'hf535;
    SB_LUT4 mux_235_i23_4_lut (.I0(encoder0_position[22]), .I1(encoder1_position[22]), 
            .I2(n15), .I3(n15_adj_5475), .O(motor_state[22]));   // verilog/TinyFPGA_B.v(271[5] 274[10])
    defparam mux_235_i23_4_lut.LUT_INIT = 16'hf535;
    SB_LUT4 mux_235_i24_4_lut (.I0(encoder0_position[23]), .I1(encoder1_position[23]), 
            .I2(n15), .I3(n15_adj_5475), .O(motor_state[23]));   // verilog/TinyFPGA_B.v(271[5] 274[10])
    defparam mux_235_i24_4_lut.LUT_INIT = 16'hf535;
    SB_LUT4 unary_minus_16_inv_0_i1_1_lut (.I0(current[0]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n25));   // verilog/TinyFPGA_B.v(109[16:24])
    defparam unary_minus_16_inv_0_i1_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_16_inv_0_i2_1_lut (.I0(current[1]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n24));   // verilog/TinyFPGA_B.v(109[16:24])
    defparam unary_minus_16_inv_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_16_inv_0_i3_1_lut (.I0(current[2]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n23));   // verilog/TinyFPGA_B.v(109[16:24])
    defparam unary_minus_16_inv_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_16_inv_0_i4_1_lut (.I0(current[3]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n22));   // verilog/TinyFPGA_B.v(109[16:24])
    defparam unary_minus_16_inv_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i5_2_lut (.I0(PWMLimit[9]), .I1(setpoint[9]), .I2(GND_net), 
            .I3(GND_net), .O(n19_adj_5539));   // verilog/TinyFPGA_B.v(230[22:30])
    defparam i5_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 unary_minus_16_inv_0_i5_1_lut (.I0(current[4]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n21));   // verilog/TinyFPGA_B.v(109[16:24])
    defparam unary_minus_16_inv_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_16_inv_0_i6_1_lut (.I0(current[5]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n20));   // verilog/TinyFPGA_B.v(109[16:24])
    defparam unary_minus_16_inv_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_16_inv_0_i7_1_lut (.I0(current[6]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n19_adj_5467));   // verilog/TinyFPGA_B.v(109[16:24])
    defparam unary_minus_16_inv_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_16_inv_0_i8_1_lut (.I0(current[7]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n18));   // verilog/TinyFPGA_B.v(109[16:24])
    defparam unary_minus_16_inv_0_i8_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_16_inv_0_i9_1_lut (.I0(current[8]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n17_adj_5466));   // verilog/TinyFPGA_B.v(109[16:24])
    defparam unary_minus_16_inv_0_i9_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_16_inv_0_i10_1_lut (.I0(current[9]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n16_adj_5465));   // verilog/TinyFPGA_B.v(109[16:24])
    defparam unary_minus_16_inv_0_i10_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_16_inv_0_i11_1_lut (.I0(current[10]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n15_adj_5464));   // verilog/TinyFPGA_B.v(109[16:24])
    defparam unary_minus_16_inv_0_i11_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_16_inv_0_i12_1_lut (.I0(current[11]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n14));   // verilog/TinyFPGA_B.v(109[16:24])
    defparam unary_minus_16_inv_0_i12_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_16_inv_0_i24_1_lut (.I0(current[15]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n2));   // verilog/TinyFPGA_B.v(109[16:24])
    defparam unary_minus_16_inv_0_i24_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1_4_lut_adj_1690 (.I0(o_Rx_DV_N_3261[12]), .I1(n4834), .I2(o_Rx_DV_N_3261[8]), 
            .I3(n55980), .O(n55986));
    defparam i1_4_lut_adj_1690.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1691 (.I0(o_Rx_DV_N_3261[24]), .I1(n29), .I2(n23_adj_5576), 
            .I3(n55986), .O(n55992));
    defparam i1_4_lut_adj_1691.LUT_INIT = 16'hfffe;
    SB_LUT4 i12458_4_lut (.I0(r_Rx_Data), .I1(rx_data[7]), .I2(n55992), 
            .I3(n27), .O(n26062));   // verilog/uart_rx.v(50[10] 145[8])
    defparam i12458_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 mux_1589_i1_3_lut (.I0(duty[3]), .I1(duty[0]), .I2(n259), 
            .I3(GND_net), .O(n9470));   // verilog/TinyFPGA_B.v(105[13] 116[7])
    defparam mux_1589_i1_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 i12931_3_lut (.I0(current[6]), .I1(data_adj_5634[6]), .I2(n24517), 
            .I3(GND_net), .O(n26535));   // verilog/tli4970.v(35[10] 68[6])
    defparam i12931_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12932_3_lut (.I0(current[5]), .I1(data_adj_5634[5]), .I2(n24517), 
            .I3(GND_net), .O(n26536));   // verilog/tli4970.v(35[10] 68[6])
    defparam i12932_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12933_3_lut (.I0(current[4]), .I1(data_adj_5634[4]), .I2(n24517), 
            .I3(GND_net), .O(n26537));   // verilog/tli4970.v(35[10] 68[6])
    defparam i12933_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12934_3_lut (.I0(current[3]), .I1(data_adj_5634[3]), .I2(n24517), 
            .I3(GND_net), .O(n26538));   // verilog/tli4970.v(35[10] 68[6])
    defparam i12934_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12935_3_lut (.I0(current[2]), .I1(data_adj_5634[2]), .I2(n24517), 
            .I3(GND_net), .O(n26539));   // verilog/tli4970.v(35[10] 68[6])
    defparam i12935_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_1589_i2_3_lut (.I0(duty[4]), .I1(duty[1]), .I2(n259), 
            .I3(GND_net), .O(n9522));   // verilog/TinyFPGA_B.v(105[13] 116[7])
    defparam mux_1589_i2_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 i12936_3_lut (.I0(current[1]), .I1(data_adj_5634[1]), .I2(n24517), 
            .I3(GND_net), .O(n26540));   // verilog/tli4970.v(35[10] 68[6])
    defparam i12936_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12956_3_lut (.I0(baudrate[15]), .I1(data_adj_5627[7]), .I2(n55498), 
            .I3(GND_net), .O(n26560));   // verilog/eeprom.v(35[8] 81[4])
    defparam i12956_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12957_3_lut (.I0(baudrate[14]), .I1(data_adj_5627[6]), .I2(n55498), 
            .I3(GND_net), .O(n26561));   // verilog/eeprom.v(35[8] 81[4])
    defparam i12957_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12958_3_lut (.I0(baudrate[13]), .I1(data_adj_5627[5]), .I2(n55498), 
            .I3(GND_net), .O(n26562));   // verilog/eeprom.v(35[8] 81[4])
    defparam i12958_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12959_3_lut (.I0(baudrate[12]), .I1(data_adj_5627[4]), .I2(n55498), 
            .I3(GND_net), .O(n26563));   // verilog/eeprom.v(35[8] 81[4])
    defparam i12959_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12960_3_lut (.I0(baudrate[11]), .I1(data_adj_5627[3]), .I2(n55498), 
            .I3(GND_net), .O(n26564));   // verilog/eeprom.v(35[8] 81[4])
    defparam i12960_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12961_3_lut (.I0(baudrate[10]), .I1(data_adj_5627[2]), .I2(n55498), 
            .I3(GND_net), .O(n26565));   // verilog/eeprom.v(35[8] 81[4])
    defparam i12961_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12962_3_lut (.I0(baudrate[9]), .I1(data_adj_5627[1]), .I2(n55498), 
            .I3(GND_net), .O(n26566));   // verilog/eeprom.v(35[8] 81[4])
    defparam i12962_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12963_3_lut (.I0(baudrate[8]), .I1(data_adj_5627[0]), .I2(n55498), 
            .I3(GND_net), .O(n26567));   // verilog/eeprom.v(35[8] 81[4])
    defparam i12963_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12470_4_lut (.I0(state_7__N_3899[3]), .I1(data_adj_5627[1]), 
            .I2(n10_adj_5559), .I3(n22404), .O(n26074));   // verilog/i2c_controller.v(91[8] 173[6])
    defparam i12470_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i12471_4_lut (.I0(state_7__N_3899[3]), .I1(data_adj_5627[2]), 
            .I2(n4_adj_5504), .I3(n22380), .O(n26075));   // verilog/i2c_controller.v(91[8] 173[6])
    defparam i12471_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i12472_4_lut (.I0(state_7__N_3899[3]), .I1(data_adj_5627[3]), 
            .I2(n4_adj_5504), .I3(n22404), .O(n26076));   // verilog/i2c_controller.v(91[8] 173[6])
    defparam i12472_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i12473_4_lut (.I0(state_7__N_3899[3]), .I1(data_adj_5627[4]), 
            .I2(n4_adj_5505), .I3(n22380), .O(n26077));   // verilog/i2c_controller.v(91[8] 173[6])
    defparam i12473_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i12474_4_lut (.I0(state_7__N_3899[3]), .I1(data_adj_5627[5]), 
            .I2(n4_adj_5505), .I3(n22404), .O(n26078));   // verilog/i2c_controller.v(91[8] 173[6])
    defparam i12474_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i12475_4_lut (.I0(state_7__N_3899[3]), .I1(data_adj_5627[6]), 
            .I2(n35435), .I3(n22380), .O(n26079));   // verilog/i2c_controller.v(91[8] 173[6])
    defparam i12475_4_lut.LUT_INIT = 16'hccac;
    SB_LUT4 i12476_4_lut (.I0(state_7__N_3899[3]), .I1(data_adj_5627[7]), 
            .I2(n35435), .I3(n22404), .O(n26080));   // verilog/i2c_controller.v(91[8] 173[6])
    defparam i12476_4_lut.LUT_INIT = 16'hccac;
    SB_LUT4 i1_4_lut_adj_1692 (.I0(o_Rx_DV_N_3261[12]), .I1(n4834), .I2(o_Rx_DV_N_3261[8]), 
            .I3(n55996), .O(n56002));
    defparam i1_4_lut_adj_1692.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1693 (.I0(o_Rx_DV_N_3261[24]), .I1(n29), .I2(n23_adj_5576), 
            .I3(n56002), .O(n56008));
    defparam i1_4_lut_adj_1693.LUT_INIT = 16'hfffe;
    SB_LUT4 i12983_4_lut (.I0(r_Rx_Data), .I1(rx_data[4]), .I2(n56008), 
            .I3(n27), .O(n26587));   // verilog/uart_rx.v(50[10] 145[8])
    defparam i12983_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i12479_3_lut (.I0(current_limit[0]), .I1(\data_in_frame[21] [0]), 
            .I2(n19639), .I3(GND_net), .O(n26083));   // verilog/coms.v(128[12] 296[6])
    defparam i12479_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12481_3_lut (.I0(\PID_CONTROLLER.integral [0]), .I1(n359), 
            .I2(n24502), .I3(GND_net), .O(n26085));   // verilog/motorControl.v(42[14] 73[8])
    defparam i12481_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12485_3_lut (.I0(current[0]), .I1(data_adj_5634[0]), .I2(n24517), 
            .I3(GND_net), .O(n26089));   // verilog/tli4970.v(35[10] 68[6])
    defparam i12485_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12486_4_lut (.I0(rw), .I1(state_adj_5628[1]), .I2(state_adj_5628[2]), 
            .I3(n5617), .O(n26090));   // verilog/eeprom.v(35[8] 81[4])
    defparam i12486_4_lut.LUT_INIT = 16'hacaa;
    SB_LUT4 i12487_4_lut (.I0(saved_addr[0]), .I1(rw), .I2(n52872), .I3(state_7__N_3883[0]), 
            .O(n26091));   // verilog/i2c_controller.v(91[8] 173[6])
    defparam i12487_4_lut.LUT_INIT = 16'hacaa;
    SB_LUT4 i12538_3_lut (.I0(\data_in_frame[11] [7]), .I1(rx_data[7]), 
            .I2(n25141), .I3(GND_net), .O(n26142));   // verilog/coms.v(128[12] 296[6])
    defparam i12538_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12535_3_lut (.I0(\data_in_frame[11] [6]), .I1(rx_data[6]), 
            .I2(n25141), .I3(GND_net), .O(n26139));   // verilog/coms.v(128[12] 296[6])
    defparam i12535_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mux_1589_i3_3_lut (.I0(duty[5]), .I1(duty[2]), .I2(n259), 
            .I3(GND_net), .O(n9520));   // verilog/TinyFPGA_B.v(105[13] 116[7])
    defparam mux_1589_i3_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 i14_3_lut (.I0(hall2), .I1(hall3), .I2(hall1), .I3(GND_net), 
            .O(n6_adj_5577));
    defparam i14_3_lut.LUT_INIT = 16'h7e7e;
    SB_LUT4 i1_3_lut_adj_1694 (.I0(hall3), .I1(hall2), .I2(hall1), .I3(GND_net), 
            .O(commutation_state_7__N_160[0]));   // verilog/TinyFPGA_B.v(151[4] 153[7])
    defparam i1_3_lut_adj_1694.LUT_INIT = 16'h1414;
    SB_LUT4 n9409_bdd_4_lut_48797 (.I0(n9409), .I1(current[3]), .I2(duty[6]), 
            .I3(n9407), .O(n63545));
    defparam n9409_bdd_4_lut_48797.LUT_INIT = 16'he4aa;
    SB_LUT4 i11946_2_lut (.I0(n24487), .I1(dti), .I2(GND_net), .I3(GND_net), 
            .O(n25556));   // verilog/TinyFPGA_B.v(131[9] 210[5])
    defparam i11946_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i48300_4_lut (.I0(commutation_state[1]), .I1(n19770), .I2(dti), 
            .I3(commutation_state[2]), .O(n24487));
    defparam i48300_4_lut.LUT_INIT = 16'hc5cf;
    SB_LUT4 n63545_bdd_4_lut (.I0(n63545), .I1(duty[3]), .I2(n4548), .I3(n9407), 
            .O(pwm_setpoint_23__N_1[3]));
    defparam n63545_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1855_4_lut_4_lut (.I0(\ID_READOUT_FSM.state [0]), .I1(\ID_READOUT_FSM.state [1]), 
            .I2(n1159), .I3(n35277), .O(n6504));   // verilog/TinyFPGA_B.v(348[5] 374[12])
    defparam i1855_4_lut_4_lut.LUT_INIT = 16'hcc8c;
    SB_LUT4 i1_2_lut_4_lut_adj_1695 (.I0(delay_counter[18]), .I1(delay_counter[17]), 
            .I2(delay_counter[16]), .I3(delay_counter[15]), .O(n4_adj_5557));
    defparam i1_2_lut_4_lut_adj_1695.LUT_INIT = 16'hfffe;
    SB_LUT4 i2_3_lut_4_lut (.I0(n62), .I1(delay_counter[31]), .I2(data_ready), 
            .I3(\ID_READOUT_FSM.state [0]), .O(n6_adj_5561));   // verilog/TinyFPGA_B.v(345[10] 375[6])
    defparam i2_3_lut_4_lut.LUT_INIT = 16'h2022;
    SB_LUT4 i1_2_lut_4_lut_adj_1696 (.I0(\ID_READOUT_FSM.state [0]), .I1(\ID_READOUT_FSM.state [1]), 
            .I2(n1159), .I3(n35277), .O(n24_adj_5562));   // verilog/TinyFPGA_B.v(345[10] 375[6])
    defparam i1_2_lut_4_lut_adj_1696.LUT_INIT = 16'hffbf;
    SB_LUT4 i1_2_lut_3_lut (.I0(state_adj_5628[2]), .I1(state_adj_5628[0]), 
            .I2(state_adj_5628[1]), .I3(GND_net), .O(n5_adj_5566));   // verilog/eeprom.v(35[8] 81[4])
    defparam i1_2_lut_3_lut.LUT_INIT = 16'h0202;
    SB_LUT4 i12_3_lut_4_lut (.I0(rx_data_ready), .I1(r_SM_Main[1]), .I2(r_SM_Main[2]), 
            .I3(n24535), .O(n48959));   // verilog/uart_rx.v(50[10] 145[8])
    defparam i12_3_lut_4_lut.LUT_INIT = 16'h0caa;
    SB_LUT4 i1_4_lut_4_lut (.I0(\ID_READOUT_FSM.state [0]), .I1(\ID_READOUT_FSM.state [1]), 
            .I2(read_N_361), .I3(n2533), .O(n25_adj_5564));   // verilog/TinyFPGA_B.v(363[7:11])
    defparam i1_4_lut_4_lut.LUT_INIT = 16'h5450;
    SB_LUT4 mux_1589_i4_3_lut (.I0(duty[6]), .I1(duty[3]), .I2(n259), 
            .I3(GND_net), .O(n9518));   // verilog/TinyFPGA_B.v(105[13] 116[7])
    defparam mux_1589_i4_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 i48335_3_lut_3_lut (.I0(\ID_READOUT_FSM.state [0]), .I1(\ID_READOUT_FSM.state [1]), 
            .I2(n35277), .I3(GND_net), .O(n24501));
    defparam i48335_3_lut_3_lut.LUT_INIT = 16'h1515;
    SB_LUT4 i46171_2_lut_3_lut (.I0(n62), .I1(delay_counter[31]), .I2(\ID_READOUT_FSM.state [0]), 
            .I3(GND_net), .O(n59865));
    defparam i46171_2_lut_3_lut.LUT_INIT = 16'hf2f2;
    SB_LUT4 i21864_2_lut_3_lut (.I0(\ID_READOUT_FSM.state [0]), .I1(\ID_READOUT_FSM.state [1]), 
            .I2(n35277), .I3(GND_net), .O(n35374));
    defparam i21864_2_lut_3_lut.LUT_INIT = 16'hfbfb;
    SB_LUT4 i12532_3_lut (.I0(\data_in_frame[11] [5]), .I1(rx_data[5]), 
            .I2(n25141), .I3(GND_net), .O(n26136));   // verilog/coms.v(128[12] 296[6])
    defparam i12532_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12639_3_lut_3_lut (.I0(\FRAME_MATCHER.rx_data_ready_prev ), .I1(rx_data_ready), 
            .I2(reset), .I3(GND_net), .O(n26243));   // verilog/coms.v(128[12] 296[6])
    defparam i12639_3_lut_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12638_3_lut_4_lut (.I0(n1548), .I1(b_prev_adj_5512), .I2(a_new_adj_5613[1]), 
            .I3(position_31__N_3609_adj_5514), .O(n26242));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    defparam i12638_3_lut_4_lut.LUT_INIT = 16'h3caa;
    SB_LUT4 n9409_bdd_4_lut_48782 (.I0(n9409), .I1(current[2]), .I2(duty[5]), 
            .I3(n9407), .O(n63539));
    defparam n9409_bdd_4_lut_48782.LUT_INIT = 16'he4aa;
    SB_LUT4 n63539_bdd_4_lut (.I0(n63539), .I1(duty[2]), .I2(n4549), .I3(n9407), 
            .O(pwm_setpoint_23__N_1[2]));
    defparam n63539_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i4789_3_lut_4_lut_4_lut (.I0(commutation_state[2]), .I1(commutation_state[1]), 
            .I2(dir), .I3(commutation_state[0]), .O(GHA_N_307));   // verilog/TinyFPGA_B.v(167[7] 186[15])
    defparam i4789_3_lut_4_lut_4_lut.LUT_INIT = 16'h12c2;
    SB_LUT4 i4791_3_lut_4_lut_4_lut (.I0(commutation_state[2]), .I1(commutation_state[1]), 
            .I2(dir), .I3(commutation_state[0]), .O(GLA_N_324));   // verilog/TinyFPGA_B.v(167[7] 186[15])
    defparam i4791_3_lut_4_lut_4_lut.LUT_INIT = 16'h212c;
    SB_LUT4 i4793_3_lut_4_lut_4_lut (.I0(commutation_state[2]), .I1(commutation_state[1]), 
            .I2(dir), .I3(commutation_state[0]), .O(GHB_N_329));
    defparam i4793_3_lut_4_lut_4_lut.LUT_INIT = 16'hc121;
    SB_LUT4 i4795_3_lut_4_lut_4_lut (.I0(commutation_state[2]), .I1(commutation_state[1]), 
            .I2(dir), .I3(commutation_state[0]), .O(GLB_N_338));
    defparam i4795_3_lut_4_lut_4_lut.LUT_INIT = 16'h1c12;
    SB_LUT4 i1_2_lut_4_lut_4_lut (.I0(\FRAME_MATCHER.state [3]), .I1(reset), 
            .I2(\FRAME_MATCHER.i_31__N_2320 ), .I3(\data_out_frame[0] [2]), 
            .O(n52768));   // verilog/TinyFPGA_B.v(345[10] 375[6])
    defparam i1_2_lut_4_lut_4_lut.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1697 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2320 ), .I3(\data_out_frame[0] [3]), 
            .O(n52818));   // verilog/TinyFPGA_B.v(345[10] 375[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1697.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1698 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2320 ), .I3(\data_out_frame[0] [4]), 
            .O(n52817));   // verilog/TinyFPGA_B.v(345[10] 375[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1698.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1699 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2320 ), .I3(\data_out_frame[1] [0]), 
            .O(n52816));   // verilog/TinyFPGA_B.v(345[10] 375[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1699.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1700 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2320 ), .I3(\data_out_frame[1] [1]), 
            .O(n52815));   // verilog/TinyFPGA_B.v(345[10] 375[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1700.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1701 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2320 ), .I3(\data_out_frame[1] [3]), 
            .O(n52814));   // verilog/TinyFPGA_B.v(345[10] 375[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1701.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1702 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2320 ), .I3(\data_out_frame[1] [5]), 
            .O(n52819));   // verilog/TinyFPGA_B.v(345[10] 375[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1702.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1703 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2320 ), .I3(\data_out_frame[1] [6]), 
            .O(n52813));   // verilog/TinyFPGA_B.v(345[10] 375[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1703.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1704 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2320 ), .I3(\data_out_frame[1] [7]), 
            .O(n52812));   // verilog/TinyFPGA_B.v(345[10] 375[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1704.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1705 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2320 ), .I3(\data_out_frame[3] [1]), 
            .O(n52811));   // verilog/TinyFPGA_B.v(345[10] 375[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1705.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1706 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2320 ), .I3(\data_out_frame[3] [3]), 
            .O(n52810));   // verilog/TinyFPGA_B.v(345[10] 375[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1706.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1707 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2320 ), .I3(\data_out_frame[3] [4]), 
            .O(n52809));   // verilog/TinyFPGA_B.v(345[10] 375[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1707.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1708 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2320 ), .I3(\data_out_frame[3] [6]), 
            .O(n52808));   // verilog/TinyFPGA_B.v(345[10] 375[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1708.LUT_INIT = 16'h2300;
    SB_LUT4 n9409_bdd_4_lut_48777 (.I0(n9409), .I1(current[1]), .I2(duty[4]), 
            .I3(n9407), .O(n63521));
    defparam n9409_bdd_4_lut_48777.LUT_INIT = 16'he4aa;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1709 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2320 ), .I3(\data_out_frame[3] [7]), 
            .O(n52807));   // verilog/TinyFPGA_B.v(345[10] 375[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1709.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1710 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2320 ), .I3(\data_out_frame[10] [3]), 
            .O(n52713));   // verilog/TinyFPGA_B.v(345[10] 375[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1710.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1711 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2320 ), .I3(\data_out_frame[10] [4]), 
            .O(n52714));   // verilog/TinyFPGA_B.v(345[10] 375[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1711.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1712 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2320 ), .I3(\data_out_frame[10] [5]), 
            .O(n52715));   // verilog/TinyFPGA_B.v(345[10] 375[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1712.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1713 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2320 ), .I3(\data_out_frame[10] [6]), 
            .O(n52789));   // verilog/TinyFPGA_B.v(345[10] 375[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1713.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1714 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2320 ), .I3(\data_out_frame[10] [7]), 
            .O(n52716));   // verilog/TinyFPGA_B.v(345[10] 375[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1714.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1715 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2320 ), .I3(\data_out_frame[11] [0]), 
            .O(n52717));   // verilog/TinyFPGA_B.v(345[10] 375[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1715.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1716 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2320 ), .I3(\data_out_frame[11] [1]), 
            .O(n52718));   // verilog/TinyFPGA_B.v(345[10] 375[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1716.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1717 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2320 ), .I3(\data_out_frame[11] [2]), 
            .O(n52719));   // verilog/TinyFPGA_B.v(345[10] 375[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1717.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1718 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2320 ), .I3(\data_out_frame[11] [3]), 
            .O(n52720));   // verilog/TinyFPGA_B.v(345[10] 375[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1718.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1719 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2320 ), .I3(\data_out_frame[11] [4]), 
            .O(n52721));   // verilog/TinyFPGA_B.v(345[10] 375[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1719.LUT_INIT = 16'h2300;
    SB_LUT4 n63521_bdd_4_lut (.I0(n63521), .I1(duty[1]), .I2(n4550), .I3(n9407), 
            .O(pwm_setpoint_23__N_1[1]));
    defparam n63521_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1720 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2320 ), .I3(\data_out_frame[11] [5]), 
            .O(n52722));   // verilog/TinyFPGA_B.v(345[10] 375[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1720.LUT_INIT = 16'h2300;
    SB_LUT4 mux_1589_i5_3_lut (.I0(duty[7]), .I1(duty[4]), .I2(n259), 
            .I3(GND_net), .O(n9516));   // verilog/TinyFPGA_B.v(105[13] 116[7])
    defparam mux_1589_i5_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1721 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2320 ), .I3(\data_out_frame[11] [6]), 
            .O(n52723));   // verilog/TinyFPGA_B.v(345[10] 375[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1721.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1722 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2320 ), .I3(\data_out_frame[11] [7]), 
            .O(n52724));   // verilog/TinyFPGA_B.v(345[10] 375[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1722.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1723 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2320 ), .I3(\data_out_frame[4] [0]), 
            .O(n52806));   // verilog/TinyFPGA_B.v(345[10] 375[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1723.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1724 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2320 ), .I3(\data_out_frame[12] [0]), 
            .O(n52725));   // verilog/TinyFPGA_B.v(345[10] 375[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1724.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1725 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2320 ), .I3(\data_out_frame[12] [1]), 
            .O(n52726));   // verilog/TinyFPGA_B.v(345[10] 375[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1725.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1726 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2320 ), .I3(\data_out_frame[4] [1]), 
            .O(n52805));   // verilog/TinyFPGA_B.v(345[10] 375[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1726.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1727 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2320 ), .I3(\data_out_frame[4] [2]), 
            .O(n52796));   // verilog/TinyFPGA_B.v(345[10] 375[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1727.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1728 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2320 ), .I3(\data_out_frame[4] [3]), 
            .O(n52797));   // verilog/TinyFPGA_B.v(345[10] 375[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1728.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1729 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2320 ), .I3(\data_out_frame[4] [4]), 
            .O(n52798));   // verilog/TinyFPGA_B.v(345[10] 375[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1729.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1730 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2320 ), .I3(\data_out_frame[4] [5]), 
            .O(n52799));   // verilog/TinyFPGA_B.v(345[10] 375[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1730.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1731 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2320 ), .I3(\data_out_frame[4] [6]), 
            .O(n52800));   // verilog/TinyFPGA_B.v(345[10] 375[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1731.LUT_INIT = 16'h2300;
    SB_LUT4 mux_1589_i6_3_lut (.I0(duty[8]), .I1(duty[5]), .I2(n259), 
            .I3(GND_net), .O(n9514));   // verilog/TinyFPGA_B.v(105[13] 116[7])
    defparam mux_1589_i6_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1732 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2320 ), .I3(\data_out_frame[4] [7]), 
            .O(n52801));   // verilog/TinyFPGA_B.v(345[10] 375[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1732.LUT_INIT = 16'h2300;
    SB_LUT4 i12529_3_lut (.I0(\data_in_frame[11] [4]), .I1(rx_data[4]), 
            .I2(n25141), .I3(GND_net), .O(n26133));   // verilog/coms.v(128[12] 296[6])
    defparam i12529_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1733 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2320 ), .I3(\data_out_frame[5] [0]), 
            .O(n52802));   // verilog/TinyFPGA_B.v(345[10] 375[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1733.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1734 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2320 ), .I3(\data_out_frame[5] [1]), 
            .O(n52803));   // verilog/TinyFPGA_B.v(345[10] 375[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1734.LUT_INIT = 16'h2300;
    SB_LUT4 i39003_4_lut_4_lut_4_lut (.I0(hall1), .I1(commutation_state[2]), 
            .I2(hall2), .I3(hall3), .O(n53662));
    defparam i39003_4_lut_4_lut_4_lut.LUT_INIT = 16'hd504;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1735 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2320 ), .I3(\data_out_frame[5] [2]), 
            .O(n52804));   // verilog/TinyFPGA_B.v(345[10] 375[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1735.LUT_INIT = 16'h2300;
    SB_LUT4 mux_1589_i7_3_lut (.I0(duty[9]), .I1(duty[6]), .I2(n259), 
            .I3(GND_net), .O(n9512));   // verilog/TinyFPGA_B.v(105[13] 116[7])
    defparam mux_1589_i7_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1736 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2320 ), .I3(\data_out_frame[5] [3]), 
            .O(n52682));   // verilog/TinyFPGA_B.v(345[10] 375[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1736.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1737 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2320 ), .I3(\data_out_frame[5] [4]), 
            .O(n52681));   // verilog/TinyFPGA_B.v(345[10] 375[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1737.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1738 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2320 ), .I3(\data_out_frame[5] [5]), 
            .O(n52683));   // verilog/TinyFPGA_B.v(345[10] 375[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1738.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1739 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2320 ), .I3(\data_out_frame[5] [6]), 
            .O(n52684));   // verilog/TinyFPGA_B.v(345[10] 375[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1739.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1740 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2320 ), .I3(\data_out_frame[5] [7]), 
            .O(n52685));   // verilog/TinyFPGA_B.v(345[10] 375[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1740.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1741 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2320 ), .I3(\data_out_frame[6] [0]), 
            .O(n52686));   // verilog/TinyFPGA_B.v(345[10] 375[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1741.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1742 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2320 ), .I3(\data_out_frame[6] [1]), 
            .O(n52687));   // verilog/TinyFPGA_B.v(345[10] 375[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1742.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1743 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2320 ), .I3(\data_out_frame[12] [2]), 
            .O(n52727));   // verilog/TinyFPGA_B.v(345[10] 375[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1743.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1744 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2320 ), .I3(\data_out_frame[12] [3]), 
            .O(n52728));   // verilog/TinyFPGA_B.v(345[10] 375[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1744.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1745 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2320 ), .I3(\data_out_frame[6] [2]), 
            .O(n52688));   // verilog/TinyFPGA_B.v(345[10] 375[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1745.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1746 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2320 ), .I3(\data_out_frame[6] [3]), 
            .O(n52693));   // verilog/TinyFPGA_B.v(345[10] 375[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1746.LUT_INIT = 16'h2300;
    SB_LUT4 i12507_3_lut_4_lut (.I0(n1507), .I1(b_prev), .I2(a_new[1]), 
            .I3(position_31__N_3609), .O(n26111));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    defparam i12507_3_lut_4_lut.LUT_INIT = 16'h3caa;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1747 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2320 ), .I3(\data_out_frame[6] [4]), 
            .O(n52692));   // verilog/TinyFPGA_B.v(345[10] 375[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1747.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1748 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2320 ), .I3(\data_out_frame[6] [5]), 
            .O(n52691));   // verilog/TinyFPGA_B.v(345[10] 375[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1748.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1749 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2320 ), .I3(\data_out_frame[6] [6]), 
            .O(n52690));   // verilog/TinyFPGA_B.v(345[10] 375[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1749.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1750 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2320 ), .I3(\data_out_frame[6] [7]), 
            .O(n52689));   // verilog/TinyFPGA_B.v(345[10] 375[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1750.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1751 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2320 ), .I3(\data_out_frame[12] [4]), 
            .O(n52729));   // verilog/TinyFPGA_B.v(345[10] 375[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1751.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1752 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2320 ), .I3(\data_out_frame[12] [5]), 
            .O(n52730));   // verilog/TinyFPGA_B.v(345[10] 375[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1752.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1753 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2320 ), .I3(\data_out_frame[12] [6]), 
            .O(n52731));   // verilog/TinyFPGA_B.v(345[10] 375[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1753.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1754 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2320 ), .I3(\data_out_frame[12] [7]), 
            .O(n52732));   // verilog/TinyFPGA_B.v(345[10] 375[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1754.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1755 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2320 ), .I3(\data_out_frame[13] [0]), 
            .O(n52733));   // verilog/TinyFPGA_B.v(345[10] 375[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1755.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1756 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2320 ), .I3(\data_out_frame[13] [1]), 
            .O(n52680));   // verilog/TinyFPGA_B.v(345[10] 375[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1756.LUT_INIT = 16'h2300;
    SB_LUT4 i596_1_lut (.I0(reset), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n2568));   // verilog/TinyFPGA_B.v(345[10] 375[6])
    defparam i596_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1757 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2320 ), .I3(\data_out_frame[13] [2]), 
            .O(n52734));   // verilog/TinyFPGA_B.v(345[10] 375[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1757.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1758 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2320 ), .I3(\data_out_frame[13] [3]), 
            .O(n52735));   // verilog/TinyFPGA_B.v(345[10] 375[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1758.LUT_INIT = 16'h2300;
    SB_LUT4 i12927_3_lut (.I0(current[10]), .I1(data_adj_5634[10]), .I2(n24517), 
            .I3(GND_net), .O(n26531));   // verilog/tli4970.v(35[10] 68[6])
    defparam i12927_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_1759 (.I0(commutation_state[2]), .I1(commutation_state[1]), 
            .I2(commutation_state_prev[2]), .I3(commutation_state_prev[1]), 
            .O(n4_adj_5471));   // verilog/TinyFPGA_B.v(134[7:48])
    defparam i1_4_lut_adj_1759.LUT_INIT = 16'h7bde;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1760 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2320 ), .I3(\data_out_frame[13] [4]), 
            .O(n52736));   // verilog/TinyFPGA_B.v(345[10] 375[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1760.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1761 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2320 ), .I3(\data_out_frame[13] [5]), 
            .O(n52737));   // verilog/TinyFPGA_B.v(345[10] 375[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1761.LUT_INIT = 16'h2300;
    SB_LUT4 i4799_3_lut_4_lut (.I0(commutation_state[2]), .I1(commutation_state[1]), 
            .I2(commutation_state[0]), .I3(dir), .O(GLC_N_352));   // verilog/TinyFPGA_B.v(188[7] 207[14])
    defparam i4799_3_lut_4_lut.LUT_INIT = 16'hcc21;
    SB_LUT4 i2_2_lut_adj_1762 (.I0(dti_counter[1]), .I1(dti_counter[2]), 
            .I2(GND_net), .I3(GND_net), .O(n10_adj_5469));   // verilog/TinyFPGA_B.v(159[9:23])
    defparam i2_2_lut_adj_1762.LUT_INIT = 16'heeee;
    SB_LUT4 i4797_3_lut_4_lut (.I0(commutation_state[2]), .I1(commutation_state[1]), 
            .I2(commutation_state[0]), .I3(dir), .O(GHC_N_343));   // verilog/TinyFPGA_B.v(188[7] 207[14])
    defparam i4797_3_lut_4_lut.LUT_INIT = 16'h21cc;
    SB_LUT4 i6_4_lut_adj_1763 (.I0(dti_counter[7]), .I1(dti_counter[4]), 
            .I2(dti_counter[5]), .I3(dti_counter[6]), .O(n14_adj_5468));   // verilog/TinyFPGA_B.v(159[9:23])
    defparam i6_4_lut_adj_1763.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1764 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2320 ), .I3(\data_out_frame[13] [6]), 
            .O(n52738));   // verilog/TinyFPGA_B.v(345[10] 375[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1764.LUT_INIT = 16'h2300;
    SB_LUT4 i7_4_lut_adj_1765 (.I0(dti_counter[0]), .I1(n14_adj_5468), .I2(n10_adj_5469), 
            .I3(dti_counter[3]), .O(n19770));   // verilog/TinyFPGA_B.v(159[9:23])
    defparam i7_4_lut_adj_1765.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1766 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2320 ), .I3(\data_out_frame[13] [7]), 
            .O(n52739));   // verilog/TinyFPGA_B.v(345[10] 375[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1766.LUT_INIT = 16'h2300;
    SB_LUT4 i48443_2_lut (.I0(n19770), .I1(dti), .I2(GND_net), .I3(GND_net), 
            .O(dti_N_356));
    defparam i48443_2_lut.LUT_INIT = 16'hbbbb;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1767 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2320 ), .I3(\data_out_frame[14] [0]), 
            .O(n52740));   // verilog/TinyFPGA_B.v(345[10] 375[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1767.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1768 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2320 ), .I3(\data_out_frame[14] [1]), 
            .O(n52741));   // verilog/TinyFPGA_B.v(345[10] 375[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1768.LUT_INIT = 16'h2300;
    SB_LUT4 i12928_3_lut (.I0(current[9]), .I1(data_adj_5634[9]), .I2(n24517), 
            .I3(GND_net), .O(n26532));   // verilog/tli4970.v(35[10] 68[6])
    defparam i12928_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2_2_lut_3_lut (.I0(hall1), .I1(hall3), .I2(hall2), .I3(GND_net), 
            .O(commutation_state_7__N_168));   // verilog/TinyFPGA_B.v(154[7:32])
    defparam i2_2_lut_3_lut.LUT_INIT = 16'h0404;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1769 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2320 ), .I3(\data_out_frame[14] [2]), 
            .O(n25663));   // verilog/TinyFPGA_B.v(345[10] 375[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1769.LUT_INIT = 16'h2300;
    SB_LUT4 i12929_3_lut (.I0(current[8]), .I1(data_adj_5634[8]), .I2(n24517), 
            .I3(GND_net), .O(n26533));   // verilog/tli4970.v(35[10] 68[6])
    defparam i12929_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1770 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2320 ), .I3(\data_out_frame[14] [3]), 
            .O(n52742));   // verilog/TinyFPGA_B.v(345[10] 375[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1770.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1771 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2320 ), .I3(\data_out_frame[14] [4]), 
            .O(n52743));   // verilog/TinyFPGA_B.v(345[10] 375[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1771.LUT_INIT = 16'h2300;
    SB_LUT4 mux_1589_i8_3_lut (.I0(duty[10]), .I1(duty[7]), .I2(n259), 
            .I3(GND_net), .O(n9510));   // verilog/TinyFPGA_B.v(105[13] 116[7])
    defparam mux_1589_i8_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 i12526_3_lut (.I0(\data_in_frame[11] [3]), .I1(rx_data[3]), 
            .I2(n25141), .I3(GND_net), .O(n26130));   // verilog/coms.v(128[12] 296[6])
    defparam i12526_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1772 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2320 ), .I3(\data_out_frame[14] [5]), 
            .O(n52744));   // verilog/TinyFPGA_B.v(345[10] 375[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1772.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1773 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2320 ), .I3(\data_out_frame[14] [6]), 
            .O(n52745));   // verilog/TinyFPGA_B.v(345[10] 375[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1773.LUT_INIT = 16'h2300;
    SB_LUT4 i13106_3_lut (.I0(\data_in_frame[20] [7]), .I1(rx_data[7]), 
            .I2(n25123), .I3(GND_net), .O(n26710));   // verilog/coms.v(128[12] 296[6])
    defparam i13106_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i17855_3_lut (.I0(n25123), .I1(rx_data[6]), .I2(\data_in_frame[20] [6]), 
            .I3(GND_net), .O(n26709));   // verilog/coms.v(92[13:20])
    defparam i17855_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i12523_3_lut (.I0(\data_in_frame[11] [2]), .I1(rx_data[2]), 
            .I2(n25141), .I3(GND_net), .O(n26127));   // verilog/coms.v(128[12] 296[6])
    defparam i12523_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1774 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2320 ), .I3(\data_out_frame[14] [7]), 
            .O(n52746));   // verilog/TinyFPGA_B.v(345[10] 375[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1774.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1775 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2320 ), .I3(\data_out_frame[15] [0]), 
            .O(n52747));   // verilog/TinyFPGA_B.v(345[10] 375[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1775.LUT_INIT = 16'h2300;
    SB_LUT4 i13098_3_lut (.I0(\data_in_frame[20] [5]), .I1(rx_data[5]), 
            .I2(n25123), .I3(GND_net), .O(n26702));   // verilog/coms.v(128[12] 296[6])
    defparam i13098_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1776 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2320 ), .I3(\data_out_frame[15] [1]), 
            .O(n52748));   // verilog/TinyFPGA_B.v(345[10] 375[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1776.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1777 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2320 ), .I3(\data_out_frame[15] [2]), 
            .O(n52749));   // verilog/TinyFPGA_B.v(345[10] 375[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1777.LUT_INIT = 16'h2300;
    SB_LUT4 i17985_3_lut (.I0(n25141), .I1(rx_data[1]), .I2(\data_in_frame[11] [1]), 
            .I3(GND_net), .O(n26767));   // verilog/coms.v(92[13:20])
    defparam i17985_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i13095_3_lut (.I0(\data_in_frame[20] [4]), .I1(rx_data[4]), 
            .I2(n25123), .I3(GND_net), .O(n26699));   // verilog/coms.v(128[12] 296[6])
    defparam i13095_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13092_3_lut (.I0(\data_in_frame[20] [3]), .I1(rx_data[3]), 
            .I2(n25123), .I3(GND_net), .O(n26696));   // verilog/coms.v(128[12] 296[6])
    defparam i13092_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13089_3_lut (.I0(\data_in_frame[20] [2]), .I1(rx_data[2]), 
            .I2(n25123), .I3(GND_net), .O(n26693));   // verilog/coms.v(128[12] 296[6])
    defparam i13089_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_4_lut_adj_1778 (.I0(state_adj_5628[2]), .I1(n22361), 
            .I2(data_ready), .I3(n3), .O(n52313));   // verilog/eeprom.v(35[8] 81[4])
    defparam i1_4_lut_4_lut_adj_1778.LUT_INIT = 16'he2e0;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1779 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2320 ), .I3(\data_out_frame[15] [3]), 
            .O(n52750));   // verilog/TinyFPGA_B.v(345[10] 375[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1779.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1780 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2320 ), .I3(\data_out_frame[15] [4]), 
            .O(n52751));   // verilog/TinyFPGA_B.v(345[10] 375[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1780.LUT_INIT = 16'h2300;
    SB_LUT4 i3_4_lut (.I0(\ID_READOUT_FSM.state [1]), .I1(n62), .I2(delay_counter[31]), 
            .I3(\ID_READOUT_FSM.state [0]), .O(n55525));
    defparam i3_4_lut.LUT_INIT = 16'h0004;
    SB_LUT4 i12582_3_lut (.I0(a_prev_adj_5511), .I1(a_new_adj_5613[1]), 
            .I2(debounce_cnt_N_3606_adj_5513), .I3(GND_net), .O(n26186));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    defparam i12582_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1781 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2320 ), .I3(\data_out_frame[15] [5]), 
            .O(n52752));   // verilog/TinyFPGA_B.v(345[10] 375[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1781.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1782 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2320 ), .I3(\data_out_frame[15] [6]), 
            .O(n52753));   // verilog/TinyFPGA_B.v(345[10] 375[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1782.LUT_INIT = 16'h2300;
    SB_LUT4 i12607_3_lut (.I0(b_prev_adj_5512), .I1(b_new_adj_5614[1]), 
            .I2(debounce_cnt_N_3606_adj_5513), .I3(GND_net), .O(n26211));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    defparam i12607_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1783 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2320 ), .I3(\data_out_frame[15] [7]), 
            .O(n52754));   // verilog/TinyFPGA_B.v(345[10] 375[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1783.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1784 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2320 ), .I3(\data_out_frame[16] [0]), 
            .O(n52755));   // verilog/TinyFPGA_B.v(345[10] 375[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1784.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1785 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2320 ), .I3(\data_out_frame[16] [1]), 
            .O(n52756));   // verilog/TinyFPGA_B.v(345[10] 375[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1785.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1786 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2320 ), .I3(\data_out_frame[16] [2]), 
            .O(n52757));   // verilog/TinyFPGA_B.v(345[10] 375[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1786.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1787 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2320 ), .I3(\data_out_frame[16] [3]), 
            .O(n52758));   // verilog/TinyFPGA_B.v(345[10] 375[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1787.LUT_INIT = 16'h2300;
    \quadrature_decoder(0)_U0  quad_counter0 (.ENCODER0_B_N_keep(ENCODER0_B_N), 
            .n1543(clk16MHz), .ENCODER0_A_N_keep(ENCODER0_A_N), .encoder0_position({encoder0_position}), 
            .GND_net(GND_net), .VCC_net(VCC_net), .n26245(n26245), .a_prev(a_prev), 
            .n26244(n26244), .b_prev(b_prev), .position_31__N_3609(position_31__N_3609), 
            .\a_new[1] (a_new[1]), .\b_new[1] (b_new[1]), .n26111(n26111), 
            .n1507(n1507), .debounce_cnt_N_3606(debounce_cnt_N_3606)) /* synthesis lattice_noprune=1 */ ;   // verilog/TinyFPGA_B.v(291[27] 297[6])
    SB_LUT4 i12640_3_lut (.I0(b_prev), .I1(b_new[1]), .I2(debounce_cnt_N_3606), 
            .I3(GND_net), .O(n26244));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    defparam i12640_3_lut.LUT_INIT = 16'hacac;
    pll32MHz pll32MHz_inst (.GND_net(GND_net), .clk16MHz(clk16MHz), .VCC_net(VCC_net), 
            .clk32MHz(clk32MHz)) /* synthesis syn_module_defined=1 */ ;   // verilog/TinyFPGA_B.v(32[10] 36[2])
    SB_LUT4 i12641_3_lut (.I0(a_prev), .I1(a_new[1]), .I2(debounce_cnt_N_3606), 
            .I3(GND_net), .O(n26245));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    defparam i12641_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1788 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2320 ), .I3(\data_out_frame[16] [4]), 
            .O(n25620));   // verilog/TinyFPGA_B.v(345[10] 375[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1788.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1789 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2320 ), .I3(\data_out_frame[16] [5]), 
            .O(n52759));   // verilog/TinyFPGA_B.v(345[10] 375[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1789.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1790 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2320 ), .I3(\data_out_frame[16] [6]), 
            .O(n52760));   // verilog/TinyFPGA_B.v(345[10] 375[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1790.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1791 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2320 ), .I3(\data_out_frame[16] [7]), 
            .O(n52761));   // verilog/TinyFPGA_B.v(345[10] 375[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1791.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1792 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2320 ), .I3(\data_out_frame[17] [0]), 
            .O(n52762));   // verilog/TinyFPGA_B.v(345[10] 375[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1792.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1793 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2320 ), .I3(\data_out_frame[17] [1]), 
            .O(n52763));   // verilog/TinyFPGA_B.v(345[10] 375[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1793.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1794 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2320 ), .I3(\data_out_frame[17] [2]), 
            .O(n52764));   // verilog/TinyFPGA_B.v(345[10] 375[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1794.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1795 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2320 ), .I3(\data_out_frame[17] [3]), 
            .O(n52765));   // verilog/TinyFPGA_B.v(345[10] 375[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1795.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1796 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2320 ), .I3(\data_out_frame[17] [4]), 
            .O(n52766));   // verilog/TinyFPGA_B.v(345[10] 375[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1796.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1797 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2320 ), .I3(\data_out_frame[17] [5]), 
            .O(n52776));   // verilog/TinyFPGA_B.v(345[10] 375[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1797.LUT_INIT = 16'h2300;
    SB_LUT4 i1_4_lut_4_lut_adj_1798 (.I0(\ID_READOUT_FSM.state [0]), .I1(\ID_READOUT_FSM.state [1]), 
            .I2(reset), .I3(n35277), .O(n51303));   // verilog/TinyFPGA_B.v(345[10] 375[6])
    defparam i1_4_lut_4_lut_adj_1798.LUT_INIT = 16'hb1f1;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1799 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2320 ), .I3(\data_out_frame[17] [6]), 
            .O(n52767));   // verilog/TinyFPGA_B.v(345[10] 375[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1799.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1800 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2320 ), .I3(\data_out_frame[17] [7]), 
            .O(n52710));   // verilog/TinyFPGA_B.v(345[10] 375[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1800.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1801 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2320 ), .I3(\data_out_frame[21] [0]), 
            .O(n52769));   // verilog/TinyFPGA_B.v(345[10] 375[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1801.LUT_INIT = 16'h2300;
    SB_LUT4 mux_1589_i9_3_lut (.I0(duty[11]), .I1(duty[8]), .I2(n259), 
            .I3(GND_net), .O(n9508));   // verilog/TinyFPGA_B.v(105[13] 116[7])
    defparam mux_1589_i9_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1802 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2320 ), .I3(\data_out_frame[21] [1]), 
            .O(n52770));   // verilog/TinyFPGA_B.v(345[10] 375[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1802.LUT_INIT = 16'h2300;
    SB_LUT4 i11955_4_lut (.I0(n24501), .I1(n1159), .I2(n59865), .I3(n35374), 
            .O(n25559));   // verilog/TinyFPGA_B.v(345[10] 375[6])
    defparam i11955_4_lut.LUT_INIT = 16'ha088;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1803 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2320 ), .I3(\data_out_frame[21] [2]), 
            .O(n52771));   // verilog/TinyFPGA_B.v(345[10] 375[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1803.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1804 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2320 ), .I3(\data_out_frame[21] [3]), 
            .O(n52772));   // verilog/TinyFPGA_B.v(345[10] 375[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1804.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1805 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2320 ), .I3(\data_out_frame[21] [4]), 
            .O(n52773));   // verilog/TinyFPGA_B.v(345[10] 375[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1805.LUT_INIT = 16'h2300;
    SB_LUT4 i21748_2_lut (.I0(n19770), .I1(dti), .I2(GND_net), .I3(GND_net), 
            .O(n35258));
    defparam i21748_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1806 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2320 ), .I3(\data_out_frame[21] [5]), 
            .O(n52774));   // verilog/TinyFPGA_B.v(345[10] 375[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1806.LUT_INIT = 16'h2300;
    SB_LUT4 n9409_bdd_4_lut_48762 (.I0(n9409), .I1(current[0]), .I2(duty[3]), 
            .I3(n9407), .O(n63515));
    defparam n9409_bdd_4_lut_48762.LUT_INIT = 16'he4aa;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1807 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2320 ), .I3(\data_out_frame[21] [6]), 
            .O(n52777));   // verilog/TinyFPGA_B.v(345[10] 375[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1807.LUT_INIT = 16'h2300;
    SB_LUT4 n63515_bdd_4_lut (.I0(n63515), .I1(duty[0]), .I2(n4551), .I3(n9407), 
            .O(pwm_setpoint_23__N_1[0]));
    defparam n63515_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i2_3_lut_adj_1808 (.I0(n47777), .I1(n53474), .I2(\data_out_frame[22] [6]), 
            .I3(GND_net), .O(n53097));   // verilog/coms.v(98[12:26])
    defparam i2_3_lut_adj_1808.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1809 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2320 ), .I3(\data_out_frame[21] [7]), 
            .O(n52778));   // verilog/TinyFPGA_B.v(345[10] 375[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1809.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1810 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2320 ), .I3(\data_out_frame[22] [0]), 
            .O(n52779));   // verilog/TinyFPGA_B.v(345[10] 375[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1810.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1811 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2320 ), .I3(\data_out_frame[22] [1]), 
            .O(n52780));   // verilog/TinyFPGA_B.v(345[10] 375[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1811.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1812 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2320 ), .I3(\data_out_frame[22] [2]), 
            .O(n52781));   // verilog/TinyFPGA_B.v(345[10] 375[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1812.LUT_INIT = 16'h2300;
    SB_LUT4 mux_1589_i10_3_lut (.I0(duty[12]), .I1(duty[9]), .I2(n259), 
            .I3(GND_net), .O(n9506));   // verilog/TinyFPGA_B.v(105[13] 116[7])
    defparam mux_1589_i10_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1813 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2320 ), .I3(\data_out_frame[22] [3]), 
            .O(n52782));   // verilog/TinyFPGA_B.v(345[10] 375[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1813.LUT_INIT = 16'h2300;
    SB_LUT4 mux_1589_i11_3_lut (.I0(duty[13]), .I1(duty[10]), .I2(n259), 
            .I3(GND_net), .O(n9504));   // verilog/TinyFPGA_B.v(105[13] 116[7])
    defparam mux_1589_i11_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1814 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2320 ), .I3(\data_out_frame[22] [4]), 
            .O(n52783));   // verilog/TinyFPGA_B.v(345[10] 375[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1814.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1815 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2320 ), .I3(\data_out_frame[22] [5]), 
            .O(n52775));   // verilog/TinyFPGA_B.v(345[10] 375[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1815.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1816 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2320 ), .I3(\data_out_frame[22] [6]), 
            .O(n52795));   // verilog/TinyFPGA_B.v(345[10] 375[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1816.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1817 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2320 ), .I3(\data_out_frame[22] [7]), 
            .O(n52786));   // verilog/TinyFPGA_B.v(345[10] 375[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1817.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1818 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2320 ), .I3(\data_out_frame[7] [0]), 
            .O(n52700));   // verilog/TinyFPGA_B.v(345[10] 375[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1818.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1819 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2320 ), .I3(\data_out_frame[7] [1]), 
            .O(n52701));   // verilog/TinyFPGA_B.v(345[10] 375[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1819.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1820 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2320 ), .I3(\data_out_frame[7] [2]), 
            .O(n52793));   // verilog/TinyFPGA_B.v(345[10] 375[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1820.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1821 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2320 ), .I3(\data_out_frame[7] [3]), 
            .O(n52792));   // verilog/TinyFPGA_B.v(345[10] 375[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1821.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1822 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2320 ), .I3(\data_out_frame[7] [4]), 
            .O(n52784));   // verilog/TinyFPGA_B.v(345[10] 375[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1822.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1823 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2320 ), .I3(\data_out_frame[7] [5]), 
            .O(n52785));   // verilog/TinyFPGA_B.v(345[10] 375[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1823.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1824 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2320 ), .I3(\data_out_frame[7] [6]), 
            .O(n52787));   // verilog/TinyFPGA_B.v(345[10] 375[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1824.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1825 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2320 ), .I3(\data_out_frame[7] [7]), 
            .O(n52788));   // verilog/TinyFPGA_B.v(345[10] 375[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1825.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1826 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2320 ), .I3(\data_out_frame[8] [0]), 
            .O(n52790));   // verilog/TinyFPGA_B.v(345[10] 375[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1826.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1827 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2320 ), .I3(\data_out_frame[8] [1]), 
            .O(n52794));   // verilog/TinyFPGA_B.v(345[10] 375[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1827.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1828 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2320 ), .I3(\data_out_frame[8] [2]), 
            .O(n52791));   // verilog/TinyFPGA_B.v(345[10] 375[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1828.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1829 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2320 ), .I3(\data_out_frame[8] [3]), 
            .O(n52694));   // verilog/TinyFPGA_B.v(345[10] 375[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1829.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1830 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2320 ), .I3(\data_out_frame[8] [4]), 
            .O(n52695));   // verilog/TinyFPGA_B.v(345[10] 375[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1830.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1831 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2320 ), .I3(\data_out_frame[8] [5]), 
            .O(n52696));   // verilog/TinyFPGA_B.v(345[10] 375[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1831.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1832 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2320 ), .I3(\data_out_frame[8] [6]), 
            .O(n52697));   // verilog/TinyFPGA_B.v(345[10] 375[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1832.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1833 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2320 ), .I3(\data_out_frame[8] [7]), 
            .O(n52698));   // verilog/TinyFPGA_B.v(345[10] 375[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1833.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1834 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2320 ), .I3(\data_out_frame[9] [0]), 
            .O(n52699));   // verilog/TinyFPGA_B.v(345[10] 375[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1834.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1835 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2320 ), .I3(\data_out_frame[9] [1]), 
            .O(n52702));   // verilog/TinyFPGA_B.v(345[10] 375[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1835.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1836 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2320 ), .I3(\data_out_frame[9] [2]), 
            .O(n52703));   // verilog/TinyFPGA_B.v(345[10] 375[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1836.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1837 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2320 ), .I3(\data_out_frame[9] [3]), 
            .O(n52704));   // verilog/TinyFPGA_B.v(345[10] 375[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1837.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1838 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2320 ), .I3(\data_out_frame[9] [4]), 
            .O(n52705));   // verilog/TinyFPGA_B.v(345[10] 375[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1838.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1839 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2320 ), .I3(\data_out_frame[9] [5]), 
            .O(n52706));   // verilog/TinyFPGA_B.v(345[10] 375[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1839.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1840 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2320 ), .I3(\data_out_frame[9] [6]), 
            .O(n52707));   // verilog/TinyFPGA_B.v(345[10] 375[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1840.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1841 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2320 ), .I3(\data_out_frame[9] [7]), 
            .O(n52708));   // verilog/TinyFPGA_B.v(345[10] 375[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1841.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1842 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2320 ), .I3(\data_out_frame[10] [0]), 
            .O(n52709));   // verilog/TinyFPGA_B.v(345[10] 375[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1842.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1843 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2320 ), .I3(\data_out_frame[10] [1]), 
            .O(n52711));   // verilog/TinyFPGA_B.v(345[10] 375[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1843.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1844 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2320 ), .I3(\data_out_frame[10] [2]), 
            .O(n52712));   // verilog/TinyFPGA_B.v(345[10] 375[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1844.LUT_INIT = 16'h2300;
    SB_LUT4 i13086_3_lut (.I0(\data_in_frame[20] [1]), .I1(rx_data[1]), 
            .I2(n25123), .I3(GND_net), .O(n26690));   // verilog/coms.v(128[12] 296[6])
    defparam i13086_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13083_3_lut (.I0(\data_in_frame[20] [0]), .I1(rx_data[0]), 
            .I2(n25123), .I3(GND_net), .O(n26687));   // verilog/coms.v(128[12] 296[6])
    defparam i13083_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i42304_3_lut (.I0(n4531), .I1(duty[20]), .I2(n9409), .I3(GND_net), 
            .O(n57016));
    defparam i42304_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i42306_3_lut (.I0(n57016), .I1(n57014), .I2(n9407), .I3(GND_net), 
            .O(pwm_setpoint_23__N_1[20]));
    defparam i42306_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i42301_3_lut (.I0(n4530), .I1(duty[21]), .I2(n9409), .I3(GND_net), 
            .O(n57013));
    defparam i42301_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_1845 (.I0(o_Rx_DV_N_3261[12]), .I1(n4834), .I2(o_Rx_DV_N_3261[8]), 
            .I3(n55884), .O(n55890));
    defparam i1_4_lut_adj_1845.LUT_INIT = 16'hfffe;
    SB_LUT4 i42303_3_lut (.I0(n57013), .I1(n57014), .I2(n9407), .I3(GND_net), 
            .O(pwm_setpoint_23__N_1[21]));
    defparam i42303_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i42302_3_lut (.I0(current[15]), .I1(duty[23]), .I2(n9409), 
            .I3(GND_net), .O(n57014));
    defparam i42302_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_1091_i9_2_lut (.I0(r_Clock_Count[4]), .I1(o_Rx_DV_N_3261[4]), 
            .I2(GND_net), .I3(GND_net), .O(n9_adj_5546));   // verilog/uart_rx.v(119[17:57])
    defparam LessThan_1091_i9_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i42298_3_lut (.I0(n4529), .I1(duty[22]), .I2(n9409), .I3(GND_net), 
            .O(n57010));
    defparam i42298_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i42300_3_lut (.I0(n57010), .I1(n57014), .I2(n9407), .I3(GND_net), 
            .O(pwm_setpoint_23__N_1[22]));
    defparam i42300_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_1846 (.I0(o_Rx_DV_N_3261[24]), .I1(n29), .I2(n23_adj_5576), 
            .I3(n55890), .O(n55896));
    defparam i1_4_lut_adj_1846.LUT_INIT = 16'hfffe;
    SB_LUT4 i4925_3_lut (.I0(n4528), .I1(current[15]), .I2(n9407), .I3(GND_net), 
            .O(n18203));
    defparam i4925_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4926_3_lut (.I0(n18203), .I1(duty[23]), .I2(n9409), .I3(GND_net), 
            .O(pwm_setpoint_23__N_1[23]));
    defparam i4926_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_1589_i12_3_lut (.I0(duty[14]), .I1(duty[11]), .I2(n259), 
            .I3(GND_net), .O(n9502));   // verilog/TinyFPGA_B.v(105[13] 116[7])
    defparam mux_1589_i12_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 mux_1589_i13_3_lut (.I0(duty[15]), .I1(duty[12]), .I2(n259), 
            .I3(GND_net), .O(n9500));   // verilog/TinyFPGA_B.v(105[13] 116[7])
    defparam mux_1589_i13_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 i13176_3_lut (.I0(\PID_CONTROLLER.integral [23]), .I1(n336), 
            .I2(n24502), .I3(GND_net), .O(n26780));   // verilog/motorControl.v(42[14] 73[8])
    defparam i13176_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12912_4_lut (.I0(r_Rx_Data), .I1(rx_data[3]), .I2(n55896), 
            .I3(n27), .O(n26516));   // verilog/uart_rx.v(50[10] 145[8])
    defparam i12912_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 LessThan_1091_i4_4_lut (.I0(r_Clock_Count[0]), .I1(o_Rx_DV_N_3261[1]), 
            .I2(r_Clock_Count[1]), .I3(o_Rx_DV_N_3261[0]), .O(n4_adj_5543));   // verilog/uart_rx.v(119[17:57])
    defparam LessThan_1091_i4_4_lut.LUT_INIT = 16'h4d0c;
    SB_LUT4 mux_1589_i14_3_lut (.I0(duty[16]), .I1(duty[13]), .I2(n259), 
            .I3(GND_net), .O(n9498));   // verilog/TinyFPGA_B.v(105[13] 116[7])
    defparam mux_1589_i14_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 LessThan_1091_i8_3_lut (.I0(n6_adj_5544), .I1(o_Rx_DV_N_3261[4]), 
            .I2(n9_adj_5546), .I3(GND_net), .O(n8_adj_5545));   // verilog/uart_rx.v(119[17:57])
    defparam LessThan_1091_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i47874_4_lut (.I0(n8_adj_5545), .I1(n4_adj_5543), .I2(n9_adj_5546), 
            .I3(n60551), .O(n62587));   // verilog/uart_rx.v(119[17:57])
    defparam i47874_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 mux_1589_i15_3_lut (.I0(duty[17]), .I1(duty[14]), .I2(n259), 
            .I3(GND_net), .O(n9496));   // verilog/TinyFPGA_B.v(105[13] 116[7])
    defparam mux_1589_i15_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 i47875_3_lut (.I0(n62587), .I1(o_Rx_DV_N_3261[5]), .I2(r_Clock_Count[5]), 
            .I3(GND_net), .O(n62588));   // verilog/uart_rx.v(119[17:57])
    defparam i47875_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i47861_3_lut (.I0(n62588), .I1(o_Rx_DV_N_3261[6]), .I2(r_Clock_Count[6]), 
            .I3(GND_net), .O(n62574));   // verilog/uart_rx.v(119[17:57])
    defparam i47861_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 LessThan_1091_i6_3_lut_3_lut (.I0(r_Clock_Count[3]), .I1(o_Rx_DV_N_3261[3]), 
            .I2(o_Rx_DV_N_3261[2]), .I3(GND_net), .O(n6_adj_5544));   // verilog/uart_rx.v(119[17:57])
    defparam LessThan_1091_i6_3_lut_3_lut.LUT_INIT = 16'hd4d4;
    SB_LUT4 i45839_3_lut_4_lut (.I0(r_Clock_Count[3]), .I1(o_Rx_DV_N_3261[3]), 
            .I2(o_Rx_DV_N_3261[2]), .I3(r_Clock_Count[2]), .O(n60551));   // verilog/uart_rx.v(119[17:57])
    defparam i45839_3_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 i46504_3_lut (.I0(n62574), .I1(o_Rx_DV_N_3261[7]), .I2(r_Clock_Count[7]), 
            .I3(GND_net), .O(n4834));   // verilog/uart_rx.v(119[17:57])
    defparam i46504_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 mux_1589_i16_3_lut (.I0(duty[18]), .I1(duty[15]), .I2(n259), 
            .I3(GND_net), .O(n9494));   // verilog/TinyFPGA_B.v(105[13] 116[7])
    defparam mux_1589_i16_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 mux_1589_i17_3_lut (.I0(duty[19]), .I1(duty[16]), .I2(n259), 
            .I3(GND_net), .O(n9492));   // verilog/TinyFPGA_B.v(105[13] 116[7])
    defparam mux_1589_i17_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 mux_1589_i18_3_lut (.I0(duty[20]), .I1(duty[17]), .I2(n259), 
            .I3(GND_net), .O(n9490));   // verilog/TinyFPGA_B.v(105[13] 116[7])
    defparam mux_1589_i18_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 i45983_3_lut (.I0(state_7__N_3883[0]), .I1(n35402), .I2(enable_slow_N_3986), 
            .I3(GND_net), .O(n59914));   // verilog/i2c_controller.v(91[8] 173[6])
    defparam i45983_3_lut.LUT_INIT = 16'h4c4c;
    SB_LUT4 i16_4_lut (.I0(state_adj_5663[0]), .I1(n59914), .I2(n6319), 
            .I3(n6_adj_5560), .O(n8_adj_5572));   // verilog/i2c_controller.v(91[8] 173[6])
    defparam i16_4_lut.LUT_INIT = 16'h3afa;
    SB_LUT4 i21751_2_lut (.I0(pwm_out), .I1(GHC), .I2(GND_net), .I3(GND_net), 
            .O(INHC_c_0));   // verilog/TinyFPGA_B.v(80[16:31])
    defparam i21751_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i21750_2_lut (.I0(pwm_out), .I1(GHB), .I2(GND_net), .I3(GND_net), 
            .O(INHB_c_0));   // verilog/TinyFPGA_B.v(78[16:31])
    defparam i21750_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i21860_2_lut (.I0(pwm_out), .I1(GHA), .I2(GND_net), .I3(GND_net), 
            .O(INHA_c_0));   // verilog/TinyFPGA_B.v(76[16:31])
    defparam i21860_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_1589_i19_3_lut (.I0(duty[21]), .I1(duty[18]), .I2(n259), 
            .I3(GND_net), .O(n9488));   // verilog/TinyFPGA_B.v(105[13] 116[7])
    defparam mux_1589_i19_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 i13222_4_lut (.I0(state_7__N_3899[3]), .I1(data_adj_5627[0]), 
            .I2(n10_adj_5559), .I3(n22380), .O(n26826));   // verilog/i2c_controller.v(91[8] 173[6])
    defparam i13222_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i13225_3_lut (.I0(n47), .I1(r_Bit_Index_adj_5651[0]), .I2(n24612), 
            .I3(GND_net), .O(n26829));   // verilog/uart_tx.v(41[10] 144[8])
    defparam i13225_3_lut.LUT_INIT = 16'h1c1c;
    SB_LUT4 i13228_3_lut (.I0(n53789), .I1(r_Bit_Index[0]), .I2(n24621), 
            .I3(GND_net), .O(n26832));   // verilog/uart_rx.v(50[10] 145[8])
    defparam i13228_3_lut.LUT_INIT = 16'h1414;
    SB_LUT4 i1_4_lut_adj_1847 (.I0(o_Rx_DV_N_3261[12]), .I1(n4834), .I2(o_Rx_DV_N_3261[8]), 
            .I3(n55916), .O(n55922));
    defparam i1_4_lut_adj_1847.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1848 (.I0(o_Rx_DV_N_3261[24]), .I1(n29), .I2(n23_adj_5576), 
            .I3(n55922), .O(n55928));
    defparam i1_4_lut_adj_1848.LUT_INIT = 16'hfffe;
    SB_LUT4 i13232_4_lut (.I0(r_Rx_Data), .I1(rx_data[0]), .I2(n55928), 
            .I3(n27), .O(n26836));   // verilog/uart_rx.v(50[10] 145[8])
    defparam i13232_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i13233_4_lut (.I0(CS_MISO_c), .I1(data_adj_5634[0]), .I2(n11_adj_5516), 
            .I3(state_7__N_4092), .O(n26837));   // verilog/tli4970.v(35[10] 68[6])
    defparam i13233_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i13236_4_lut (.I0(n5_adj_5566), .I1(state_adj_5628[0]), .I2(n55082), 
            .I3(n4_adj_5474), .O(n26840));   // verilog/eeprom.v(35[8] 81[4])
    defparam i13236_4_lut.LUT_INIT = 16'h4144;
    SB_LUT4 i1_4_lut_adj_1849 (.I0(n23_adj_5576), .I1(o_Rx_DV_N_3261[12]), 
            .I2(n4834), .I3(o_Rx_DV_N_3261[8]), .O(n55718));
    defparam i1_4_lut_adj_1849.LUT_INIT = 16'hfffe;
    SB_LUT4 i45645_4_lut (.I0(data_ready), .I1(n6504), .I2(n24_adj_5562), 
            .I3(\ID_READOUT_FSM.state [0]), .O(n59888));   // verilog/TinyFPGA_B.v(345[10] 375[6])
    defparam i45645_4_lut.LUT_INIT = 16'hdccc;
    SB_LUT4 i46121_2_lut (.I0(n24_adj_5562), .I1(n6504), .I2(GND_net), 
            .I3(GND_net), .O(n59891));   // verilog/TinyFPGA_B.v(345[10] 375[6])
    defparam i46121_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i49_4_lut (.I0(n59891), .I1(n59888), .I2(\ID_READOUT_FSM.state [0]), 
            .I3(n6_adj_5561), .O(n51215));   // verilog/TinyFPGA_B.v(345[10] 375[6])
    defparam i49_4_lut.LUT_INIT = 16'hcac0;
    SB_LUT4 i6_4_lut_adj_1850 (.I0(ID[5]), .I1(ID[4]), .I2(ID[2]), .I3(ID[6]), 
            .O(n14_adj_5573));   // verilog/TinyFPGA_B.v(364[12:17])
    defparam i6_4_lut_adj_1850.LUT_INIT = 16'hfffe;
    SB_LUT4 i5_4_lut (.I0(ID[0]), .I1(ID[1]), .I2(ID[3]), .I3(ID[7]), 
            .O(n13_adj_5574));   // verilog/TinyFPGA_B.v(364[12:17])
    defparam i5_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i21767_4_lut (.I0(n13_adj_5574), .I1(n33), .I2(n14_adj_5573), 
            .I3(n34), .O(n35277));
    defparam i21767_4_lut.LUT_INIT = 16'hfac8;
    SB_LUT4 i1_2_lut_adj_1851 (.I0(delay_counter[12]), .I1(delay_counter[11]), 
            .I2(GND_net), .I3(GND_net), .O(n4_adj_5556));
    defparam i1_2_lut_adj_1851.LUT_INIT = 16'heeee;
    SB_LUT4 i2_4_lut (.I0(delay_counter[9]), .I1(n4_adj_5556), .I2(delay_counter[10]), 
            .I3(n22256), .O(n55221));
    defparam i2_4_lut.LUT_INIT = 16'hfcec;
    SB_LUT4 i2_4_lut_adj_1852 (.I0(n55221), .I1(n22269), .I2(delay_counter[13]), 
            .I3(delay_counter[14]), .O(n55183));
    defparam i2_4_lut_adj_1852.LUT_INIT = 16'hffec;
    SB_LUT4 i3_3_lut (.I0(delay_counter[20]), .I1(delay_counter[21]), .I2(delay_counter[23]), 
            .I3(GND_net), .O(n8_adj_5476));
    defparam i3_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 i1_4_lut_adj_1853 (.I0(o_Rx_DV_N_3261[24]), .I1(n27), .I2(n29), 
            .I3(n55718), .O(r_SM_Main_2__N_3219[1]));
    defparam i1_4_lut_adj_1853.LUT_INIT = 16'hfffe;
    SB_LUT4 i2_4_lut_adj_1854 (.I0(delay_counter[22]), .I1(n55183), .I2(delay_counter[19]), 
            .I3(delay_counter[18]), .O(n7_adj_5503));
    defparam i2_4_lut_adj_1854.LUT_INIT = 16'ha8a0;
    SB_LUT4 i21759_4_lut (.I0(n7_adj_5503), .I1(delay_counter[31]), .I2(n22253), 
            .I3(n8_adj_5476), .O(n1159));   // verilog/TinyFPGA_B.v(366[14:38])
    defparam i21759_4_lut.LUT_INIT = 16'h3230;
    SB_LUT4 i5_4_lut_adj_1855 (.I0(delay_counter[27]), .I1(delay_counter[29]), 
            .I2(delay_counter[24]), .I3(delay_counter[26]), .O(n12_adj_5542));
    defparam i5_4_lut_adj_1855.LUT_INIT = 16'hfffe;
    SB_LUT4 i6_4_lut_adj_1856 (.I0(delay_counter[28]), .I1(n12_adj_5542), 
            .I2(delay_counter[25]), .I3(delay_counter[30]), .O(n22253));
    defparam i6_4_lut_adj_1856.LUT_INIT = 16'hfffe;
    SB_LUT4 i2_3_lut_adj_1857 (.I0(delay_counter[17]), .I1(delay_counter[16]), 
            .I2(delay_counter[15]), .I3(GND_net), .O(n22269));
    defparam i2_3_lut_adj_1857.LUT_INIT = 16'hfefe;
    SB_LUT4 i5_3_lut (.I0(delay_counter[3]), .I1(delay_counter[5]), .I2(delay_counter[4]), 
            .I3(GND_net), .O(n14_adj_5473));
    defparam i5_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i6_4_lut_adj_1858 (.I0(delay_counter[8]), .I1(delay_counter[7]), 
            .I2(delay_counter[1]), .I3(delay_counter[0]), .O(n15_adj_5472));
    defparam i6_4_lut_adj_1858.LUT_INIT = 16'hfffe;
    SB_LUT4 i8_4_lut_adj_1859 (.I0(n15_adj_5472), .I1(delay_counter[2]), 
            .I2(n14_adj_5473), .I3(delay_counter[6]), .O(n22256));
    defparam i8_4_lut_adj_1859.LUT_INIT = 16'hfffe;
    SB_LUT4 i4086_4_lut (.I0(n22256), .I1(delay_counter[11]), .I2(delay_counter[10]), 
            .I3(delay_counter[9]), .O(n24_adj_5515));
    defparam i4086_4_lut.LUT_INIT = 16'hc8c0;
    SB_LUT4 i2_4_lut_adj_1860 (.I0(n24_adj_5515), .I1(delay_counter[14]), 
            .I2(delay_counter[12]), .I3(delay_counter[13]), .O(n55370));
    defparam i2_4_lut_adj_1860.LUT_INIT = 16'hc800;
    SB_LUT4 i1_2_lut_adj_1861 (.I0(delay_counter[22]), .I1(n22253), .I2(GND_net), 
            .I3(GND_net), .O(n6_adj_5540));
    defparam i1_2_lut_adj_1861.LUT_INIT = 16'heeee;
    SB_LUT4 i2_4_lut_adj_1862 (.I0(n55370), .I1(delay_counter[20]), .I2(n4_adj_5557), 
            .I3(delay_counter[19]), .O(n54628));
    defparam i2_4_lut_adj_1862.LUT_INIT = 16'hc800;
    SB_LUT4 i4_4_lut (.I0(delay_counter[23]), .I1(n54628), .I2(delay_counter[21]), 
            .I3(n6_adj_5540), .O(n62));
    defparam i4_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i21826_2_lut (.I0(n62), .I1(delay_counter[31]), .I2(GND_net), 
            .I3(GND_net), .O(read_N_361));   // verilog/TinyFPGA_B.v(352[12:35])
    defparam i21826_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i561_2_lut (.I0(n1159), .I1(n35277), .I2(GND_net), .I3(GND_net), 
            .O(n2533));   // verilog/TinyFPGA_B.v(370[18] 372[12])
    defparam i561_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i42023_2_lut (.I0(data_ready), .I1(\ID_READOUT_FSM.state [0]), 
            .I2(GND_net), .I3(GND_net), .O(n56726));
    defparam i42023_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i48514_4_lut (.I0(\ID_READOUT_FSM.state [1]), .I1(n6504), .I2(n56726), 
            .I3(n25_adj_5564), .O(n17_adj_5563));   // verilog/TinyFPGA_B.v(345[10] 375[6])
    defparam i48514_4_lut.LUT_INIT = 16'h88ba;
    SB_LUT4 i13245_3_lut (.I0(\PID_CONTROLLER.integral [22]), .I1(n337), 
            .I2(n24502), .I3(GND_net), .O(n26849));   // verilog/motorControl.v(42[14] 73[8])
    defparam i13245_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13246_3_lut (.I0(\PID_CONTROLLER.integral [21]), .I1(n338), 
            .I2(n24502), .I3(GND_net), .O(n26850));   // verilog/motorControl.v(42[14] 73[8])
    defparam i13246_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13247_3_lut (.I0(\PID_CONTROLLER.integral [20]), .I1(n339), 
            .I2(n24502), .I3(GND_net), .O(n26851));   // verilog/motorControl.v(42[14] 73[8])
    defparam i13247_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13248_3_lut (.I0(\PID_CONTROLLER.integral [19]), .I1(n340), 
            .I2(n24502), .I3(GND_net), .O(n26852));   // verilog/motorControl.v(42[14] 73[8])
    defparam i13248_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13249_3_lut (.I0(\PID_CONTROLLER.integral [18]), .I1(n341), 
            .I2(n24502), .I3(GND_net), .O(n26853));   // verilog/motorControl.v(42[14] 73[8])
    defparam i13249_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8_3_lut (.I0(\PID_CONTROLLER.integral [17]), .I1(n31535), .I2(n24502), 
            .I3(GND_net), .O(n26854));
    defparam i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13251_3_lut (.I0(\PID_CONTROLLER.integral [16]), .I1(n343), 
            .I2(n24502), .I3(GND_net), .O(n26855));   // verilog/motorControl.v(42[14] 73[8])
    defparam i13251_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13252_3_lut (.I0(\PID_CONTROLLER.integral [15]), .I1(n344), 
            .I2(n24502), .I3(GND_net), .O(n26856));   // verilog/motorControl.v(42[14] 73[8])
    defparam i13252_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13253_3_lut (.I0(\PID_CONTROLLER.integral [14]), .I1(n345), 
            .I2(n24502), .I3(GND_net), .O(n26857));   // verilog/motorControl.v(42[14] 73[8])
    defparam i13253_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13254_3_lut (.I0(\PID_CONTROLLER.integral [13]), .I1(n346), 
            .I2(n24502), .I3(GND_net), .O(n26858));   // verilog/motorControl.v(42[14] 73[8])
    defparam i13254_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13255_3_lut (.I0(\PID_CONTROLLER.integral [12]), .I1(n347), 
            .I2(n24502), .I3(GND_net), .O(n26859));   // verilog/motorControl.v(42[14] 73[8])
    defparam i13255_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13256_3_lut (.I0(\PID_CONTROLLER.integral [11]), .I1(n348), 
            .I2(n24502), .I3(GND_net), .O(n26860));   // verilog/motorControl.v(42[14] 73[8])
    defparam i13256_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13257_3_lut (.I0(\PID_CONTROLLER.integral [10]), .I1(n349), 
            .I2(n24502), .I3(GND_net), .O(n26861));   // verilog/motorControl.v(42[14] 73[8])
    defparam i13257_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13258_3_lut (.I0(\PID_CONTROLLER.integral [9]), .I1(n350), 
            .I2(n24502), .I3(GND_net), .O(n26862));   // verilog/motorControl.v(42[14] 73[8])
    defparam i13258_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13259_3_lut (.I0(\PID_CONTROLLER.integral [8]), .I1(n351), 
            .I2(n24502), .I3(GND_net), .O(n26863));   // verilog/motorControl.v(42[14] 73[8])
    defparam i13259_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13260_3_lut (.I0(\PID_CONTROLLER.integral [7]), .I1(n352), 
            .I2(n24502), .I3(GND_net), .O(n26864));   // verilog/motorControl.v(42[14] 73[8])
    defparam i13260_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13261_3_lut (.I0(\PID_CONTROLLER.integral [6]), .I1(n353), 
            .I2(n24502), .I3(GND_net), .O(n26865));   // verilog/motorControl.v(42[14] 73[8])
    defparam i13261_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13262_3_lut (.I0(\PID_CONTROLLER.integral [5]), .I1(n354), 
            .I2(n24502), .I3(GND_net), .O(n26866));   // verilog/motorControl.v(42[14] 73[8])
    defparam i13262_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13263_3_lut (.I0(\PID_CONTROLLER.integral [4]), .I1(n355), 
            .I2(n24502), .I3(GND_net), .O(n26867));   // verilog/motorControl.v(42[14] 73[8])
    defparam i13263_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13264_3_lut (.I0(\PID_CONTROLLER.integral [3]), .I1(n356), 
            .I2(n24502), .I3(GND_net), .O(n26868));   // verilog/motorControl.v(42[14] 73[8])
    defparam i13264_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13265_3_lut (.I0(\PID_CONTROLLER.integral [2]), .I1(n357), 
            .I2(n24502), .I3(GND_net), .O(n26869));   // verilog/motorControl.v(42[14] 73[8])
    defparam i13265_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_adj_1863 (.I0(control_mode[5]), .I1(control_mode[4]), 
            .I2(GND_net), .I3(GND_net), .O(n56512));   // verilog/TinyFPGA_B.v(272[5:22])
    defparam i1_2_lut_adj_1863.LUT_INIT = 16'heeee;
    SB_LUT4 i1_4_lut_adj_1864 (.I0(control_mode[7]), .I1(n1_adj_5541), .I2(n56512), 
            .I3(control_mode[6]), .O(n22431));   // verilog/TinyFPGA_B.v(272[5:22])
    defparam i1_4_lut_adj_1864.LUT_INIT = 16'hfffe;
    TLI4970 tli (.n26534(n26534), .\current[7] (current[7]), .n26533(n26533), 
            .\current[8] (current[8]), .n26532(n26532), .\current[9] (current[9]), 
            .n26531(n26531), .\current[10] (current[10]), .n26530(n26530), 
            .\current[11] (current[11]), .clk16MHz(clk16MHz), .n26439(n26439), 
            .\data[15] (data_adj_5634[15]), .n26437(n26437), .\data[12] (data_adj_5634[12]), 
            .n26435(n26435), .\data[11] (data_adj_5634[11]), .n26433(n26433), 
            .\data[10] (data_adj_5634[10]), .n26430(n26430), .\data[9] (data_adj_5634[9]), 
            .n26428(n26428), .\data[8] (data_adj_5634[8]), .n26427(n26427), 
            .\data[7] (data_adj_5634[7]), .n26424(n26424), .\data[6] (data_adj_5634[6]), 
            .n26422(n26422), .\data[5] (data_adj_5634[5]), .n26420(n26420), 
            .\data[4] (data_adj_5634[4]), .n26418(n26418), .\data[3] (data_adj_5634[3]), 
            .n26416(n26416), .\data[2] (data_adj_5634[2]), .GND_net(GND_net), 
            .VCC_net(VCC_net), .n26414(n26414), .\data[1] (data_adj_5634[1]), 
            .n6(n6_adj_5537), .n6_adj_14(n6_adj_5507), .n5(n5_adj_5508), 
            .n6_adj_15(n6_adj_5506), .n9(n9_adj_5517), .n35347(n35347), 
            .n35411(n35411), .n26837(n26837), .\data[0] (data_adj_5634[0]), 
            .n24517(n24517), .\current[15] (current[15]), .CS_c(CS_c), 
            .n26089(n26089), .\current[0] (current[0]), .n26540(n26540), 
            .\current[1] (current[1]), .n26539(n26539), .\current[2] (current[2]), 
            .n26538(n26538), .\current[3] (current[3]), .n26537(n26537), 
            .\current[4] (current[4]), .n26536(n26536), .\current[5] (current[5]), 
            .n26535(n26535), .\current[6] (current[6]), .n11(n11_adj_5516), 
            .state_7__N_4092(state_7__N_4092), .CS_CLK_c(CS_CLK_c), .n22373(n22373), 
            .n4(n4_adj_5470), .n22369(n22369), .n22357(n22357), .n22377(n22377), 
            .n4_adj_16(n4_adj_5565)) /* synthesis syn_noprune=1, syn_module_defined=1 */ ;   // verilog/TinyFPGA_B.v(391[11] 397[4])
    SB_LUT4 i13266_3_lut (.I0(\PID_CONTROLLER.integral [1]), .I1(n358), 
            .I2(n24502), .I3(GND_net), .O(n26870));   // verilog/motorControl.v(42[14] 73[8])
    defparam i13266_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_1094_i15_2_lut (.I0(r_Clock_Count_adj_5650[7]), .I1(o_Rx_DV_N_3261[7]), 
            .I2(GND_net), .I3(GND_net), .O(n15_adj_5553));   // verilog/uart_tx.v(117[17:57])
    defparam LessThan_1094_i15_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_1094_i13_2_lut (.I0(r_Clock_Count_adj_5650[6]), .I1(o_Rx_DV_N_3261[6]), 
            .I2(GND_net), .I3(GND_net), .O(n13_adj_5552));   // verilog/uart_tx.v(117[17:57])
    defparam LessThan_1094_i13_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_1094_i9_2_lut (.I0(r_Clock_Count_adj_5650[4]), .I1(o_Rx_DV_N_3261[4]), 
            .I2(GND_net), .I3(GND_net), .O(n9_adj_5550));   // verilog/uart_tx.v(117[17:57])
    defparam LessThan_1094_i9_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i13290_3_lut (.I0(current_limit[15]), .I1(\data_in_frame[20] [7]), 
            .I2(n19639), .I3(GND_net), .O(n26894));   // verilog/coms.v(128[12] 296[6])
    defparam i13290_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i17865_3_lut (.I0(current_limit[14]), .I1(\data_in_frame[20] [6]), 
            .I2(n19639), .I3(GND_net), .O(n26895));
    defparam i17865_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13292_3_lut (.I0(current_limit[13]), .I1(\data_in_frame[20] [5]), 
            .I2(n19639), .I3(GND_net), .O(n26896));   // verilog/coms.v(128[12] 296[6])
    defparam i13292_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13293_3_lut (.I0(current_limit[12]), .I1(\data_in_frame[20] [4]), 
            .I2(n19639), .I3(GND_net), .O(n26897));   // verilog/coms.v(128[12] 296[6])
    defparam i13293_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13294_3_lut (.I0(current_limit[11]), .I1(\data_in_frame[20] [3]), 
            .I2(n19639), .I3(GND_net), .O(n26898));   // verilog/coms.v(128[12] 296[6])
    defparam i13294_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13295_3_lut (.I0(current_limit[10]), .I1(\data_in_frame[20] [2]), 
            .I2(n19639), .I3(GND_net), .O(n26899));   // verilog/coms.v(128[12] 296[6])
    defparam i13295_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13296_3_lut (.I0(current_limit[9]), .I1(\data_in_frame[20] [1]), 
            .I2(n19639), .I3(GND_net), .O(n26900));   // verilog/coms.v(128[12] 296[6])
    defparam i13296_3_lut.LUT_INIT = 16'hcaca;
    coms setpoint_23__I_0 (.VCC_net(VCC_net), .clk16MHz(clk16MHz), .rx_data({rx_data}), 
         .\Kp[12] (Kp[12]), .IntegralLimit({IntegralLimit}), .\Kp[11] (Kp[11]), 
         .\Kp[10] (Kp[10]), .\Kp[9] (Kp[9]), .\Kp[5] (Kp[5]), .\Kp[4] (Kp[4]), 
         .\data_in_frame[3][3] (\data_in_frame[3] [3]), .\Kp[3] (Kp[3]), 
         .\data_in_frame[3][2] (\data_in_frame[3] [2]), .\Kp[2] (Kp[2]), 
         .\data_in_frame[3][1] (\data_in_frame[3] [1]), .\Kp[1] (Kp[1]), 
         .\data_in_frame[11] ({\data_in_frame[11] }), .rx_data_ready(rx_data_ready), 
         .\FRAME_MATCHER.rx_data_ready_prev (\FRAME_MATCHER.rx_data_ready_prev ), 
         .GND_net(GND_net), .deadband({deadband[23:3], Open_0, Open_1, 
         Open_2}), .\data_in_frame[3][6] (\data_in_frame[3] [6]), .\data_in_frame[3][7] (\data_in_frame[3] [7]), 
         .\data_in_frame[18] ({Open_3, Open_4, \data_in_frame[18] [5:0]}), 
         .n25157(n25157), .n2568(n2568), .\data_out_frame[0][2] (\data_out_frame[0] [2]), 
         .n52768(n52768), .\data_out_frame[0][3] (\data_out_frame[0] [3]), 
         .n52818(n52818), .\data_out_frame[0][4] (\data_out_frame[0] [4]), 
         .n52817(n52817), .\data_out_frame[1][0] (\data_out_frame[1] [0]), 
         .n52816(n52816), .\data_out_frame[1][1] (\data_out_frame[1] [1]), 
         .n52815(n52815), .\data_out_frame[1][3] (\data_out_frame[1] [3]), 
         .n52814(n52814), .\FRAME_MATCHER.state[3] (\FRAME_MATCHER.state [3]), 
         .\data_out_frame[1][5] (\data_out_frame[1] [5]), .n52819(n52819), 
         .\data_out_frame[1][6] (\data_out_frame[1] [6]), .n52813(n52813), 
         .\data_in_frame[18][7] (\data_in_frame[18] [7]), .\data_out_frame[1][7] (\data_out_frame[1] [7]), 
         .n52812(n52812), .\data_out_frame[6] ({\data_out_frame[6] }), .\FRAME_MATCHER.i_31__N_2320 (\FRAME_MATCHER.i_31__N_2320 ), 
         .encoder0_position({encoder0_position[23:0]}), .\data_out_frame[21] ({\data_out_frame[21] }), 
         .\data_out_frame[15] ({\data_out_frame[15] }), .reset(reset), .\data_out_frame[17] ({\data_out_frame[17] }), 
         .\data_in_frame[1][2] (\data_in_frame[1] [2]), .\data_out_frame[22] ({\data_out_frame[22] }), 
         .\data_in_frame[1][3] (\data_in_frame[1] [3]), .setpoint({setpoint}), 
         .\data_out_frame[13] ({\data_out_frame[13] }), .\data_in_frame[1][4] (\data_in_frame[1] [4]), 
         .\data_out_frame[11] ({\data_out_frame[11] }), .\data_out_frame[9] ({\data_out_frame[9] }), 
         .\data_out_frame[16] ({\data_out_frame[16] }), .byte_transmit_counter({Open_5, 
         Open_6, Open_7, Open_8, Open_9, Open_10, Open_11, byte_transmit_counter[0]}), 
         .\data_out_frame[14] ({\data_out_frame[14] }), .\data_out_frame[4] ({\data_out_frame[4] }), 
         .\data_out_frame[7] ({\data_out_frame[7] }), .\data_out_frame[8] ({\data_out_frame[8] }), 
         .\data_out_frame[12] ({\data_out_frame[12] }), .\data_in_frame[1][5] (\data_in_frame[1] [5]), 
         .\data_in_frame[1][6] (\data_in_frame[1] [6]), .\data_out_frame[3][1] (\data_out_frame[3] [1]), 
         .n52811(n52811), .n48858(n48858), .\data_out_frame[5] ({\data_out_frame[5] }), 
         .\data_out_frame[3][3] (\data_out_frame[3] [3]), .n52810(n52810), 
         .\data_out_frame[3][4] (\data_out_frame[3] [4]), .n52809(n52809), 
         .\data_out_frame[3][6] (\data_out_frame[3] [6]), .n52808(n52808), 
         .\data_out_frame[3][7] (\data_out_frame[3] [7]), .n52807(n52807), 
         .\data_out_frame[10] ({\data_out_frame[10] }), .n52713(n52713), 
         .n52714(n52714), .n52715(n52715), .n52789(n52789), .n52716(n52716), 
         .n52717(n52717), .n52718(n52718), .n52719(n52719), .n52720(n52720), 
         .n52721(n52721), .n52722(n52722), .n52723(n52723), .n52724(n52724), 
         .n52806(n52806), .n52725(n52725), .n52726(n52726), .n54590(n54590), 
         .n47777(n47777), .n52805(n52805), .n52796(n52796), .n26190(n26190), 
         .n26193(n26193), .n26196(n26196), .n52797(n52797), .n26199(n26199), 
         .n52798(n52798), .n26202(n26202), .n26205(n26205), .\data_in_frame[1][7] (\data_in_frame[1] [7]), 
         .n52799(n52799), .n52800(n52800), .n52801(n52801), .n52802(n52802), 
         .n52803(n52803), .n52804(n52804), .n52682(n52682), .control_mode({control_mode[7], 
         Open_12, Open_13, Open_14, Open_15, Open_16, Open_17, Open_18}), 
         .n26238(n26238), .n26250(n26250), .n26253(n26253), .n26262(n26262), 
         .n26265(n26265), .n26268(n26268), .\data_in_frame[4] ({Open_19, 
         Open_20, Open_21, Open_22, Open_23, \data_in_frame[4] [2:0]}), 
         .n26271(n26271), .n26274(n26274), .n26291(n26291), .\data_in_frame[4][6] (\data_in_frame[4] [6]), 
         .\control_mode[1] (control_mode[1]), .\control_mode[0] (control_mode[0]), 
         .n26294(n26294), .\data_in_frame[4][7] (\data_in_frame[4] [7]), 
         .n52681(n52681), .n52683(n52683), .n52684(n52684), .\byte_transmit_counter[2] (byte_transmit_counter[2]), 
         .n52685(n52685), .n52686(n52686), .\deadband[1] (deadband[1]), 
         .\Kp[8] (Kp[8]), .\Kp[7] (Kp[7]), .ID({ID}), .\Ki[15] (Ki[15]), 
         .\Ki[14] (Ki[14]), .\Ki[13] (Ki[13]), .n26634(n26634), .n27035(n27035), 
         .n26640(n26640), .n25161(n25161), .\control_mode[6] (control_mode[6]), 
         .\control_mode[5] (control_mode[5]), .n26643(n26643), .n26646(n26646), 
         .n26649(n26649), .n26655(n26655), .n26092(n26092), .\control_mode[4] (control_mode[4]), 
         .n26911(n26911), .n26910(n26910), .n26909(n26909), .n26908(n26908), 
         .current_limit({current_limit}), .n26907(n26907), .n26906(n26906), 
         .n26905(n26905), .n26904(n26904), .n26903(n26903), .n26902(n26902), 
         .n26901(n26901), .n26900(n26900), .n26899(n26899), .n26898(n26898), 
         .n26897(n26897), .n26896(n26896), .n26895(n26895), .n26894(n26894), 
         .PWMLimit({PWMLimit}), .\Ki[1] (Ki[1]), .\Ki[2] (Ki[2]), .\Ki[3] (Ki[3]), 
         .\Ki[4] (Ki[4]), .\Ki[5] (Ki[5]), .\Ki[6] (Ki[6]), .\Ki[7] (Ki[7]), 
         .\Ki[8] (Ki[8]), .\Ki[9] (Ki[9]), .\Ki[10] (Ki[10]), .\Ki[11] (Ki[11]), 
         .n52687(n52687), .n7(n7_adj_5575), .\Ki[12] (Ki[12]), .n26687(n26687), 
         .\data_in_frame[20] ({\data_in_frame[20] }), .n26690(n26690), .\data_out_frame[26][6] (\data_out_frame[26] [6]), 
         .\data_out_frame[27][6] (\data_out_frame[27] [6]), .encoder1_position({encoder1_position[23:0]}), 
         .n26243(n26243), .n52727(n52727), .n52728(n52728), .n26693(n26693), 
         .n26696(n26696), .n26699(n26699), .n26767(n26767), .n26702(n26702), 
         .n26127(n26127), .n26709(n26709), .n26710(n26710), .\Kp[13] (Kp[13]), 
         .n26130(n26130), .\data_in_frame[21] ({\data_in_frame[21] }), .n52688(n52688), 
         .n52693(n52693), .n52692(n52692), .\Kp[14] (Kp[14]), .n52691(n52691), 
         .n52690(n52690), .n52689(n52689), .n26133(n26133), .n52729(n52729), 
         .n52730(n52730), .n52731(n52731), .n52732(n52732), .n52733(n52733), 
         .n52680(n52680), .n52734(n52734), .n52735(n52735), .\Kp[15] (Kp[15]), 
         .n52736(n52736), .n52737(n52737), .n52738(n52738), .n52739(n52739), 
         .n52740(n52740), .n52741(n52741), .n25663(n25663), .n52742(n52742), 
         .n52743(n52743), .n52744(n52744), .n52745(n52745), .n52746(n52746), 
         .n52747(n52747), .n52748(n52748), .n52749(n52749), .n52750(n52750), 
         .n52751(n52751), .n52752(n52752), .n52753(n52753), .n52754(n52754), 
         .n52755(n52755), .n52756(n52756), .n52757(n52757), .n52758(n52758), 
         .n22431(n22431), .n15(n15_adj_5475), .control_update(control_update), 
         .n24502(n24502), .n25620(n25620), .n52759(n52759), .n52760(n52760), 
         .n52761(n52761), .n52762(n52762), .n26136(n26136), .n52763(n52763), 
         .n52764(n52764), .n52765(n52765), .n52766(n52766), .n52776(n52776), 
         .n52767(n52767), .n52710(n52710), .n52769(n52769), .n52770(n52770), 
         .n52771(n52771), .n52772(n52772), .n52773(n52773), .n52774(n52774), 
         .n52777(n52777), .n52778(n52778), .n52779(n52779), .n52780(n52780), 
         .n52781(n52781), .n52782(n52782), .n52783(n52783), .n52775(n52775), 
         .n52795(n52795), .n52786(n52786), .DE_c(DE_c), .n26139(n26139), 
         .n26142(n26142), .n52700(n52700), .n52701(n52701), .n52793(n52793), 
         .n52792(n52792), .n52784(n52784), .n52785(n52785), .n52787(n52787), 
         .n52788(n52788), .n52790(n52790), .n52794(n52794), .n52791(n52791), 
         .n52694(n52694), .n52695(n52695), .n52696(n52696), .n52697(n52697), 
         .n52698(n52698), .n52699(n52699), .n52702(n52702), .n52703(n52703), 
         .n52704(n52704), .n52705(n52705), .n52706(n52706), .n52707(n52707), 
         .n52708(n52708), .n52709(n52709), .n52711(n52711), .\Kp[6] (Kp[6]), 
         .n26083(n26083), .\Ki[0] (Ki[0]), .\Kp[0] (Kp[0]), .n52712(n52712), 
         .\deadband[0] (deadband[0]), .n25123(n25123), .n53097(n53097), 
         .n53474(n53474), .n59927(n59927), .n24840(n24840), .n15_adj_3(n15), 
         .n33792(n33792), .n1(n1_adj_5541), .n32007(n32007), .n19639(n19639), 
         .\current[7] (current[7]), .\current[6] (current[6]), .\current[5] (current[5]), 
         .\current[4] (current[4]), .n25127(n25127), .\current[3] (current[3]), 
         .\current[2] (current[2]), .\current[1] (current[1]), .\current[0] (current[0]), 
         .\current[15] (current[15]), .\current[11] (current[11]), .\current[10] (current[10]), 
         .\current[9] (current[9]), .\current[8] (current[8]), .pwm_setpoint({pwm_setpoint}), 
         .n52908(n52908), .n59928(n59928), .n25141(n25141), .r_Clock_Count({r_Clock_Count_adj_5650}), 
         .n24612(n24612), .n36763(n36763), .tx_o(tx_o), .n26829(n26829), 
         .\r_Bit_Index[0] (r_Bit_Index_adj_5651[0]), .\o_Rx_DV_N_3261[12] (o_Rx_DV_N_3261[12]), 
         .n4837(n4837), .\o_Rx_DV_N_3261[24] (o_Rx_DV_N_3261[24]), .n29(n29), 
         .n23(n23_adj_5576), .n27(n27), .n47(n47), .tx_enable(tx_enable), 
         .baudrate({baudrate}), .n24621(n24621), .n53789(n53789), .r_Clock_Count_adj_13({r_Clock_Count}), 
         .n26516(n26516), .\r_SM_Main[2] (r_SM_Main[2]), .r_Rx_Data(r_Rx_Data), 
         .RX_N_42(RX_N_42), .\r_Bit_Index[0]_adj_12 (r_Bit_Index[0]), .n55980(n55980), 
         .n55948(n55948), .n26445(n26445), .\o_Rx_DV_N_3261[8] (o_Rx_DV_N_3261[8]), 
         .n26443(n26443), .\o_Rx_DV_N_3261[7] (o_Rx_DV_N_3261[7]), .\o_Rx_DV_N_3261[6] (o_Rx_DV_N_3261[6]), 
         .\o_Rx_DV_N_3261[5] (o_Rx_DV_N_3261[5]), .n33(n33), .\o_Rx_DV_N_3261[4] (o_Rx_DV_N_3261[4]), 
         .\o_Rx_DV_N_3261[3] (o_Rx_DV_N_3261[3]), .\o_Rx_DV_N_3261[2] (o_Rx_DV_N_3261[2]), 
         .\o_Rx_DV_N_3261[1] (o_Rx_DV_N_3261[1]), .\o_Rx_DV_N_3261[0] (o_Rx_DV_N_3261[0]), 
         .n27051(n27051), .n26970(n26970), .n4834(n4834), .n52823(n52823), 
         .n26836(n26836), .n48959(n48959), .n26832(n26832), .n55964(n55964), 
         .n55996(n55996), .\r_SM_Main[1] (r_SM_Main[1]), .\r_SM_Main_2__N_3219[1] (r_SM_Main_2__N_3219[1]), 
         .n55461(n55461), .n26587(n26587), .n26062(n26062), .n55884(n55884), 
         .n55900(n55900), .n55916(n55916), .n55932(n55932), .n55814(n55814), 
         .n24535(n24535), .n34(n34)) /* synthesis syn_module_defined=1 */ ;   // verilog/TinyFPGA_B.v(243[22] 266[4])
    SB_LUT4 i13297_3_lut (.I0(current_limit[8]), .I1(\data_in_frame[20] [0]), 
            .I2(n19639), .I3(GND_net), .O(n26901));   // verilog/coms.v(128[12] 296[6])
    defparam i13297_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13298_3_lut (.I0(current_limit[7]), .I1(\data_in_frame[21] [7]), 
            .I2(n19639), .I3(GND_net), .O(n26902));   // verilog/coms.v(128[12] 296[6])
    defparam i13298_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13299_3_lut (.I0(current_limit[6]), .I1(\data_in_frame[21] [6]), 
            .I2(n19639), .I3(GND_net), .O(n26903));   // verilog/coms.v(128[12] 296[6])
    defparam i13299_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13300_3_lut (.I0(current_limit[5]), .I1(\data_in_frame[21] [5]), 
            .I2(n19639), .I3(GND_net), .O(n26904));   // verilog/coms.v(128[12] 296[6])
    defparam i13300_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13301_3_lut (.I0(current_limit[4]), .I1(\data_in_frame[21] [4]), 
            .I2(n19639), .I3(GND_net), .O(n26905));   // verilog/coms.v(128[12] 296[6])
    defparam i13301_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13302_3_lut (.I0(current_limit[3]), .I1(\data_in_frame[21] [3]), 
            .I2(n19639), .I3(GND_net), .O(n26906));   // verilog/coms.v(128[12] 296[6])
    defparam i13302_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12930_3_lut (.I0(current[7]), .I1(data_adj_5634[7]), .I2(n24517), 
            .I3(GND_net), .O(n26534));   // verilog/tli4970.v(35[10] 68[6])
    defparam i12930_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13303_3_lut (.I0(current_limit[2]), .I1(\data_in_frame[21] [2]), 
            .I2(n19639), .I3(GND_net), .O(n26907));   // verilog/coms.v(128[12] 296[6])
    defparam i13303_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13304_3_lut (.I0(current_limit[1]), .I1(\data_in_frame[21] [1]), 
            .I2(n19639), .I3(GND_net), .O(n26908));   // verilog/coms.v(128[12] 296[6])
    defparam i13304_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13305_3_lut (.I0(control_mode[7]), .I1(\data_in_frame[1] [7]), 
            .I2(n19639), .I3(GND_net), .O(n26909));   // verilog/coms.v(128[12] 296[6])
    defparam i13305_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13306_3_lut (.I0(control_mode[6]), .I1(\data_in_frame[1] [6]), 
            .I2(n19639), .I3(GND_net), .O(n26910));   // verilog/coms.v(128[12] 296[6])
    defparam i13306_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13307_3_lut (.I0(control_mode[5]), .I1(\data_in_frame[1] [5]), 
            .I2(n19639), .I3(GND_net), .O(n26911));   // verilog/coms.v(128[12] 296[6])
    defparam i13307_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_1094_i11_2_lut (.I0(r_Clock_Count_adj_5650[5]), .I1(o_Rx_DV_N_3261[5]), 
            .I2(GND_net), .I3(GND_net), .O(n11_adj_5551));   // verilog/uart_tx.v(117[17:57])
    defparam LessThan_1094_i11_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i12488_3_lut (.I0(\data_in_frame[11] [0]), .I1(rx_data[0]), 
            .I2(n25141), .I3(GND_net), .O(n26092));   // verilog/coms.v(128[12] 296[6])
    defparam i12488_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 LessThan_14_i6_3_lut_3_lut (.I0(current_limit[2]), .I1(current_limit[3]), 
            .I2(current[3]), .I3(GND_net), .O(n6_adj_5486));   // verilog/TinyFPGA_B.v(106[9:30])
    defparam LessThan_14_i6_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i45450_2_lut_4_lut (.I0(current[8]), .I1(current_limit[8]), 
            .I2(current[4]), .I3(current_limit[4]), .O(n60162));
    defparam i45450_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 LessThan_14_i8_3_lut_3_lut (.I0(current_limit[4]), .I1(current_limit[8]), 
            .I2(current[8]), .I3(GND_net), .O(n8_adj_5484));   // verilog/TinyFPGA_B.v(106[9:30])
    defparam LessThan_14_i8_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i13051_3_lut (.I0(\data_in_frame[18] [7]), .I1(rx_data[7]), 
            .I2(n25127), .I3(GND_net), .O(n26655));   // verilog/coms.v(128[12] 296[6])
    defparam i13051_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13045_3_lut (.I0(\data_in_frame[18] [5]), .I1(rx_data[5]), 
            .I2(n25127), .I3(GND_net), .O(n26649));   // verilog/coms.v(128[12] 296[6])
    defparam i13045_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13042_3_lut (.I0(\data_in_frame[18] [4]), .I1(rx_data[4]), 
            .I2(n25127), .I3(GND_net), .O(n26646));   // verilog/coms.v(128[12] 296[6])
    defparam i13042_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 unary_minus_15_inv_0_i24_1_lut (.I0(duty[23]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(pwm_setpoint_23__N_159));   // verilog/TinyFPGA_B.v(107[24:29])
    defparam unary_minus_15_inv_0_i24_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i13039_3_lut (.I0(\data_in_frame[18] [3]), .I1(rx_data[3]), 
            .I2(n25127), .I3(GND_net), .O(n26643));   // verilog/coms.v(128[12] 296[6])
    defparam i13039_3_lut.LUT_INIT = 16'hacac;
    \quadrature_decoder(0)  quad_counter1 (.ENCODER1_B_N_keep(ENCODER1_B_N), 
            .n1543(clk16MHz), .ENCODER1_A_N_keep(ENCODER1_A_N), .n26242(n26242), 
            .n1548(n1548), .n26211(n26211), .b_prev(b_prev_adj_5512), 
            .n26186(n26186), .a_prev(a_prev_adj_5511), .position_31__N_3609(position_31__N_3609_adj_5514), 
            .encoder1_position({encoder1_position}), .\a_new[1] (a_new_adj_5613[1]), 
            .\b_new[1] (b_new_adj_5614[1]), .GND_net(GND_net), .VCC_net(VCC_net), 
            .debounce_cnt_N_3606(debounce_cnt_N_3606_adj_5513)) /* synthesis lattice_noprune=1 */ ;   // verilog/TinyFPGA_B.v(299[27] 305[6])
    SB_LUT4 i1_2_lut_3_lut_adj_1865 (.I0(\data_out_frame[22] [4]), .I1(n48858), 
            .I2(n54590), .I3(GND_net), .O(n52908));   // verilog/coms.v(98[12:26])
    defparam i1_2_lut_3_lut_adj_1865.LUT_INIT = 16'h6969;
    SB_LUT4 LessThan_1094_i4_4_lut (.I0(r_Clock_Count_adj_5650[0]), .I1(o_Rx_DV_N_3261[1]), 
            .I2(r_Clock_Count_adj_5650[1]), .I3(o_Rx_DV_N_3261[0]), .O(n4_adj_5547));   // verilog/uart_tx.v(117[17:57])
    defparam LessThan_1094_i4_4_lut.LUT_INIT = 16'h4d0c;
    SB_LUT4 i1_4_lut_adj_1866 (.I0(o_Rx_DV_N_3261[12]), .I1(n4834), .I2(o_Rx_DV_N_3261[8]), 
            .I3(n55964), .O(n55970));
    defparam i1_4_lut_adj_1866.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1867 (.I0(o_Rx_DV_N_3261[24]), .I1(n29), .I2(n23_adj_5576), 
            .I3(n55970), .O(n55976));
    defparam i1_4_lut_adj_1867.LUT_INIT = 16'hfffe;
    SB_LUT4 i13366_4_lut (.I0(r_Rx_Data), .I1(rx_data[5]), .I2(n55976), 
            .I3(n27), .O(n26970));   // verilog/uart_rx.v(50[10] 145[8])
    defparam i13366_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 LessThan_11_i6_3_lut_3_lut (.I0(duty[2]), .I1(duty[3]), .I2(current[3]), 
            .I3(GND_net), .O(n6_adj_5501));   // verilog/TinyFPGA_B.v(98[10:22])
    defparam LessThan_11_i6_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 mux_1589_i20_3_lut (.I0(duty[22]), .I1(duty[19]), .I2(n259), 
            .I3(GND_net), .O(n9486));   // verilog/TinyFPGA_B.v(105[13] 116[7])
    defparam mux_1589_i20_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 LessThan_11_i10_3_lut_3_lut (.I0(duty[5]), .I1(duty[6]), .I2(current[6]), 
            .I3(GND_net), .O(n10_adj_5497));   // verilog/TinyFPGA_B.v(98[10:22])
    defparam LessThan_11_i10_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    pwm PWM (.n2568(n2568), .pwm_out(pwm_out), .clk32MHz(clk32MHz), .reset(reset), 
        .pwm_setpoint({pwm_setpoint}), .GND_net(GND_net), .VCC_net(VCC_net), 
        .\PWMLimit[7] (PWMLimit[7]), .\setpoint[7] (setpoint[7]), .n15(n15_adj_5538)) /* synthesis syn_module_defined=1 */ ;   // verilog/TinyFPGA_B.v(85[6] 90[3])
    SB_LUT4 LessThan_11_i8_3_lut_3_lut (.I0(duty[4]), .I1(duty[8]), .I2(current[8]), 
            .I3(GND_net), .O(n8_adj_5499));   // verilog/TinyFPGA_B.v(98[10:22])
    defparam LessThan_11_i8_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i45797_2_lut_4_lut (.I0(duty[6]), .I1(n303), .I2(duty[5]), 
            .I3(n304), .O(n60509));
    defparam i45797_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 i45787_2_lut_4_lut (.I0(duty[8]), .I1(n301), .I2(duty[4]), 
            .I3(n305), .O(n60499));
    defparam i45787_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    motorControl control (.GND_net(GND_net), .\Kp[12] (Kp[12]), .\Ki[3] (Ki[3]), 
            .n348(n348), .n32007(n32007), .\Kp[13] (Kp[13]), .VCC_net(VCC_net), 
            .\PID_CONTROLLER.integral ({\PID_CONTROLLER.integral }), .n292(n292), 
            .\Ki[4] (Ki[4]), .\Kp[6] (Kp[6]), .IntegralLimit({IntegralLimit}), 
            .\Ki[7] (Ki[7]), .n344(n344), .\Ki[0] (Ki[0]), .n341(n341), 
            .\Kp[1] (Kp[1]), .\Kp[0] (Kp[0]), .\Ki[5] (Ki[5]), .\Ki[6] (Ki[6]), 
            .\Kp[7] (Kp[7]), .\Ki[8] (Ki[8]), .\Kp[8] (Kp[8]), .\Ki[9] (Ki[9]), 
            .\Kp[9] (Kp[9]), .\Ki[10] (Ki[10]), .\Kp[10] (Kp[10]), .control_update(control_update), 
            .duty({duty}), .clk16MHz(clk16MHz), .reset(reset), .n240(n240), 
            .\Kp[2] (Kp[2]), .setpoint({setpoint}), .\Kp[3] (Kp[3]), .\Ki[11] (Ki[11]), 
            .\Ki[12] (Ki[12]), .n284(n284), .n258(n258), .\Kp[4] (Kp[4]), 
            .\Ki[1] (Ki[1]), .n349(n349), .n53(n53), .\Ki[2] (Ki[2]), 
            .\Kp[11] (Kp[11]), .\deadband[0] (deadband[0]), .n339(n339), 
            .n338(n338), .n336(n336), .n337(n337), .n340(n340), .\Kp[14] (Kp[14]), 
            .\Kp[5] (Kp[5]), .n490(n490), .n417(n417), .n344_adj_1(n344_adj_5558), 
            .n271(n271), .n198(n198), .n125(n125), .n35(n35), .n26870(n26870), 
            .n26869(n26869), .n26868(n26868), .n26867(n26867), .n26866(n26866), 
            .n26865(n26865), .n26864(n26864), .n26863(n26863), .n26862(n26862), 
            .n26861(n26861), .n26860(n26860), .n26859(n26859), .n26858(n26858), 
            .n26857(n26857), .n26856(n26856), .n26855(n26855), .n26854(n26854), 
            .n26853(n26853), .n26852(n26852), .n26851(n26851), .n26850(n26850), 
            .n26849(n26849), .n26780(n26780), .\Kp[15] (Kp[15]), .n343(n343), 
            .\deadband[1] (deadband[1]), .n26085(n26085), .\motor_state[23] (motor_state[23]), 
            .\motor_state[22] (motor_state[22]), .\motor_state[21] (motor_state[21]), 
            .\motor_state[20] (motor_state[20]), .\motor_state[19] (motor_state[19]), 
            .\motor_state[18] (motor_state[18]), .\motor_state[17] (motor_state[17]), 
            .\motor_state[16] (motor_state[16]), .\motor_state[15] (motor_state[15]), 
            .\motor_state[14] (motor_state[14]), .\motor_state[13] (motor_state[13]), 
            .\motor_state[12] (motor_state[12]), .n35211(n35211), .\motor_state[10] (motor_state[10]), 
            .\motor_state[9] (motor_state[9]), .\motor_state[8] (motor_state[8]), 
            .\motor_state[7] (motor_state[7]), .n33792(n33792), .\motor_state[5] (motor_state[5]), 
            .\motor_state[4] (motor_state[4]), .\motor_state[3] (motor_state[3]), 
            .\motor_state[2] (motor_state[2]), .n1(n1), .\motor_state[0] (motor_state[0]), 
            .n350(n350), .\Ki[13] (Ki[13]), .\Ki[14] (Ki[14]), .n351(n351), 
            .\deadband[5] (deadband[5]), .n345(n345), .\Ki[15] (Ki[15]), 
            .\deadband[6] (deadband[6]), .\deadband[7] (deadband[7]), .\deadband[8] (deadband[8]), 
            .\deadband[9] (deadband[9]), .\deadband[10] (deadband[10]), 
            .\deadband[11] (deadband[11]), .\deadband[12] (deadband[12]), 
            .\deadband[13] (deadband[13]), .\deadband[14] (deadband[14]), 
            .\deadband[15] (deadband[15]), .\deadband[16] (deadband[16]), 
            .n352(n352), .\deadband[17] (deadband[17]), .\deadband[18] (deadband[18]), 
            .PWMLimit({PWMLimit}), .\deadband[19] (deadband[19]), .\deadband[20] (deadband[20]), 
            .\deadband[21] (deadband[21]), .\deadband[22] (deadband[22]), 
            .\deadband[23] (deadband[23]), .n359(n359), .n353(n353), .n346(n346), 
            .n35713(n35713), .n354(n354), .\control_mode[0] (control_mode[0]), 
            .\control_mode[5] (control_mode[5]), .\control_mode[4] (control_mode[4]), 
            .n1_adj_2(n1_adj_5541), .n355(n355), .\control_mode[6] (control_mode[6]), 
            .\control_mode[7] (control_mode[7]), .\control_mode[1] (control_mode[1]), 
            .n19(n19_adj_5539), .n15(n15_adj_5538), .n356(n356), .\deadband[3] (deadband[3]), 
            .\deadband[4] (deadband[4]), .n357(n357), .n358(n358), .n347(n347)) /* synthesis syn_module_defined=1 */ ;   // verilog/TinyFPGA_B.v(276[16] 289[4])
    
endmodule
//
// Verilog Description of module EEPROM
//

module EEPROM (clk16MHz, enable_slow_N_3986, n5616, \state[2] , n52055, 
            n26840, VCC_net, \state[0] , \state[1] , GND_net, n3, 
            n55082, n26090, rw, n52313, data_ready, ID, baudrate, 
            n26567, n26566, n26565, n26564, n26563, n26562, n26561, 
            n26560, n35339, n55498, n4, \state[0]_adj_21 , n22361, 
            read, data, scl_enable, \state_7__N_3883[0] , n26826, 
            n8, n6319, sda_enable, n35402, n26091, \saved_addr[0] , 
            n26080, n26079, n26078, n26077, n26076, n26075, n26074, 
            n4_adj_22, n4_adj_23, n22404, n35435, n10, n52872, \state_7__N_3899[3] , 
            scl, sda_out, n6, n22380) /* synthesis syn_noprune=1, syn_module_defined=1 */ ;
    input clk16MHz;
    output enable_slow_N_3986;
    output [0:0]n5616;
    output \state[2] ;
    input n52055;
    input n26840;
    input VCC_net;
    output \state[0] ;
    output \state[1] ;
    input GND_net;
    output n3;
    output n55082;
    input n26090;
    output rw;
    input n52313;
    output data_ready;
    output [7:0]ID;
    output [31:0]baudrate;
    input n26567;
    input n26566;
    input n26565;
    input n26564;
    input n26563;
    input n26562;
    input n26561;
    input n26560;
    output n35339;
    output n55498;
    output n4;
    output \state[0]_adj_21 ;
    output n22361;
    input read;
    output [7:0]data;
    output scl_enable;
    output \state_7__N_3883[0] ;
    input n26826;
    input n8;
    output n6319;
    output sda_enable;
    output n35402;
    input n26091;
    output \saved_addr[0] ;
    input n26080;
    input n26079;
    input n26078;
    input n26077;
    input n26076;
    input n26075;
    input n26074;
    output n4_adj_22;
    output n4_adj_23;
    output n22404;
    output n35435;
    output n10;
    output n52872;
    input \state_7__N_3899[3] ;
    output scl;
    output sda_out;
    output n6;
    output n22380;
    
    wire clk16MHz /* synthesis SET_AS_NETWORK=clk16MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(31[6:14])
    
    wire n47941, n24676;
    wire [2:0]byte_counter;   // verilog/eeprom.v(30[11:23])
    
    wire n26045;
    wire [15:0]delay_counter_15__N_3729;
    
    wire n24562;
    wire [15:0]delay_counter;   // verilog/eeprom.v(28[12:25])
    
    wire n33079, n6527, n33075, n6529, n6530, n6531, n6532, n6533;
    wire [2:0]n17;
    
    wire ready_prev, enable;
    wire [7:0]state_7__N_3658;
    
    wire n55256, n33077, n47187, n52873;
    wire [15:0]n5010;
    
    wire n46276, n46275, n46274, n46273, n46272, n26087, n46271, 
        n26582, n26581, n26580, n26579, n26578, n26577, n26576, 
        n26575, n26574, n26573, n26572, n26571, n26570, n26569, 
        n26568, n26559, n26558, n26557, n26556, n26555, n26554, 
        n26553, n26552, n26551, n26550, n26549, n26548, n26547, 
        n46270, n26546, n26545, n26544, n46269, n46268, n46267, 
        n46266, n46265, n46264, n46263, n46262, n28, n26, n27, 
        n25, n22261, n52876;
    wire [7:0]state;   // verilog/i2c_controller.v(33[12:17])
    
    wire n7, n4_c, n56621, n4_adj_5460, n59921, n55087;
    
    SB_DFFESR byte_counter_1942__i0 (.Q(byte_counter[0]), .C(clk16MHz), 
            .E(n24676), .D(n47941), .R(n26045));   // verilog/eeprom.v(68[25:39])
    SB_DFFESR delay_counter_i0_i1 (.Q(delay_counter[1]), .C(clk16MHz), .E(n24562), 
            .D(delay_counter_15__N_3729[1]), .R(n33079));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFFESR delay_counter_i0_i2 (.Q(delay_counter[2]), .C(clk16MHz), .E(n24562), 
            .D(delay_counter_15__N_3729[2]), .R(n33079));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFFESR delay_counter_i0_i3 (.Q(delay_counter[3]), .C(clk16MHz), .E(n24562), 
            .D(delay_counter_15__N_3729[3]), .R(n33079));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFFESS delay_counter_i0_i4 (.Q(delay_counter[4]), .C(clk16MHz), .E(n24562), 
            .D(n6527), .S(n33075));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFFESR delay_counter_i0_i5 (.Q(delay_counter[5]), .C(clk16MHz), .E(n24562), 
            .D(delay_counter_15__N_3729[5]), .R(n33079));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFFESS delay_counter_i0_i6 (.Q(delay_counter[6]), .C(clk16MHz), .E(n24562), 
            .D(n6529), .S(n33075));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFFESS delay_counter_i0_i7 (.Q(delay_counter[7]), .C(clk16MHz), .E(n24562), 
            .D(n6530), .S(n33075));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFFESS delay_counter_i0_i8 (.Q(delay_counter[8]), .C(clk16MHz), .E(n24562), 
            .D(n6531), .S(n33075));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFFESS delay_counter_i0_i9 (.Q(delay_counter[9]), .C(clk16MHz), .E(n24562), 
            .D(n6532), .S(n33075));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFFESS delay_counter_i0_i10 (.Q(delay_counter[10]), .C(clk16MHz), 
            .E(n24562), .D(n6533), .S(n33075));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFFESR delay_counter_i0_i11 (.Q(delay_counter[11]), .C(clk16MHz), 
            .E(n24562), .D(delay_counter_15__N_3729[11]), .R(n33079));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFFESR delay_counter_i0_i12 (.Q(delay_counter[12]), .C(clk16MHz), 
            .E(n24562), .D(delay_counter_15__N_3729[12]), .R(n33079));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFFESR delay_counter_i0_i13 (.Q(delay_counter[13]), .C(clk16MHz), 
            .E(n24562), .D(delay_counter_15__N_3729[13]), .R(n33079));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFFESR delay_counter_i0_i14 (.Q(delay_counter[14]), .C(clk16MHz), 
            .E(n24562), .D(delay_counter_15__N_3729[14]), .R(n33079));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFFESR delay_counter_i0_i15 (.Q(delay_counter[15]), .C(clk16MHz), 
            .E(n24562), .D(delay_counter_15__N_3729[15]), .R(n33079));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFFESR byte_counter_1942__i2 (.Q(byte_counter[2]), .C(clk16MHz), 
            .E(n24676), .D(n17[2]), .R(n26045));   // verilog/eeprom.v(68[25:39])
    SB_DFFESR byte_counter_1942__i1 (.Q(byte_counter[1]), .C(clk16MHz), 
            .E(n24676), .D(n17[1]), .R(n26045));   // verilog/eeprom.v(68[25:39])
    SB_DFF ready_prev_59 (.Q(ready_prev), .C(clk16MHz), .D(enable_slow_N_3986));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFFSR enable_58 (.Q(enable), .C(clk16MHz), .D(n5616[0]), .R(\state[2] ));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF state_i2 (.Q(\state[2] ), .C(clk16MHz), .D(n52055));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFFE state_i0 (.Q(\state[0] ), .C(clk16MHz), .E(VCC_net), .D(n26840));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFFE state_i1 (.Q(\state[1] ), .C(clk16MHz), .E(n55256), .D(state_7__N_3658[1]));   // verilog/eeprom.v(35[8] 81[4])
    SB_LUT4 i1_2_lut_3_lut (.I0(\state[2] ), .I1(\state[0] ), .I2(n24562), 
            .I3(GND_net), .O(n33079));
    defparam i1_2_lut_3_lut.LUT_INIT = 16'he0e0;
    SB_LUT4 i9_1_lut_2_lut (.I0(\state[2] ), .I1(n3), .I2(GND_net), .I3(GND_net), 
            .O(n33077));
    defparam i9_1_lut_2_lut.LUT_INIT = 16'h7777;
    SB_LUT4 i2_2_lut_3_lut (.I0(byte_counter[0]), .I1(byte_counter[1]), 
            .I2(byte_counter[2]), .I3(GND_net), .O(n3));   // verilog/eeprom.v(68[25:39])
    defparam i2_2_lut_3_lut.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_2_lut_3_lut_adj_1664 (.I0(byte_counter[0]), .I1(byte_counter[1]), 
            .I2(n47187), .I3(GND_net), .O(n52873));   // verilog/eeprom.v(68[25:39])
    defparam i1_2_lut_3_lut_adj_1664.LUT_INIT = 16'hefef;
    SB_LUT4 add_1111_17_lut (.I0(GND_net), .I1(delay_counter[15]), .I2(n5010[13]), 
            .I3(n46276), .O(delay_counter_15__N_3729[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1111_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_1111_16_lut (.I0(GND_net), .I1(delay_counter[14]), .I2(n5010[13]), 
            .I3(n46275), .O(delay_counter_15__N_3729[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1111_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1111_16 (.CI(n46275), .I0(delay_counter[14]), .I1(n5010[13]), 
            .CO(n46276));
    SB_LUT4 add_1111_15_lut (.I0(GND_net), .I1(delay_counter[13]), .I2(n5010[13]), 
            .I3(n46274), .O(delay_counter_15__N_3729[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1111_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1111_15 (.CI(n46274), .I0(delay_counter[13]), .I1(n5010[13]), 
            .CO(n46275));
    SB_LUT4 i3_4_lut_4_lut_4_lut (.I0(\state[1] ), .I1(\state[0] ), .I2(enable_slow_N_3986), 
            .I3(ready_prev), .O(n55082));
    defparam i3_4_lut_4_lut_4_lut.LUT_INIT = 16'h8808;
    SB_LUT4 add_1111_14_lut (.I0(GND_net), .I1(delay_counter[12]), .I2(n5010[13]), 
            .I3(n46273), .O(delay_counter_15__N_3729[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1111_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1111_14 (.CI(n46273), .I0(delay_counter[12]), .I1(n5010[13]), 
            .CO(n46274));
    SB_DFFESR delay_counter_i0_i0 (.Q(delay_counter[0]), .C(clk16MHz), .E(n24562), 
            .D(delay_counter_15__N_3729[0]), .R(n33079));   // verilog/eeprom.v(35[8] 81[4])
    SB_LUT4 add_1111_13_lut (.I0(GND_net), .I1(delay_counter[11]), .I2(n5010[13]), 
            .I3(n46272), .O(delay_counter_15__N_3729[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1111_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1111_13 (.CI(n46272), .I0(delay_counter[11]), .I1(n5010[13]), 
            .CO(n46273));
    SB_DFF rw_64 (.Q(rw), .C(clk16MHz), .D(n26090));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF data_ready_61 (.Q(data_ready), .C(clk16MHz), .D(n52313));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i1 (.Q(ID[0]), .C(clk16MHz), .D(n26087));   // verilog/eeprom.v(35[8] 81[4])
    SB_LUT4 add_1111_12_lut (.I0(n33077), .I1(delay_counter[10]), .I2(n5010[13]), 
            .I3(n46271), .O(n6533)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1111_12_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_1111_12 (.CI(n46271), .I0(delay_counter[10]), .I1(n5010[13]), 
            .CO(n46272));
    SB_DFF bytes_0___i2 (.Q(ID[1]), .C(clk16MHz), .D(n26582));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i3 (.Q(ID[2]), .C(clk16MHz), .D(n26581));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i4 (.Q(ID[3]), .C(clk16MHz), .D(n26580));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i5 (.Q(ID[4]), .C(clk16MHz), .D(n26579));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i6 (.Q(ID[5]), .C(clk16MHz), .D(n26578));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i7 (.Q(ID[6]), .C(clk16MHz), .D(n26577));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i8 (.Q(ID[7]), .C(clk16MHz), .D(n26576));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i9 (.Q(baudrate[0]), .C(clk16MHz), .D(n26575));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i10 (.Q(baudrate[1]), .C(clk16MHz), .D(n26574));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i11 (.Q(baudrate[2]), .C(clk16MHz), .D(n26573));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i12 (.Q(baudrate[3]), .C(clk16MHz), .D(n26572));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i13 (.Q(baudrate[4]), .C(clk16MHz), .D(n26571));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i14 (.Q(baudrate[5]), .C(clk16MHz), .D(n26570));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i15 (.Q(baudrate[6]), .C(clk16MHz), .D(n26569));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i16 (.Q(baudrate[7]), .C(clk16MHz), .D(n26568));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i17 (.Q(baudrate[8]), .C(clk16MHz), .D(n26567));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i18 (.Q(baudrate[9]), .C(clk16MHz), .D(n26566));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i19 (.Q(baudrate[10]), .C(clk16MHz), .D(n26565));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i20 (.Q(baudrate[11]), .C(clk16MHz), .D(n26564));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i21 (.Q(baudrate[12]), .C(clk16MHz), .D(n26563));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i22 (.Q(baudrate[13]), .C(clk16MHz), .D(n26562));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i23 (.Q(baudrate[14]), .C(clk16MHz), .D(n26561));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i24 (.Q(baudrate[15]), .C(clk16MHz), .D(n26560));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i25 (.Q(baudrate[16]), .C(clk16MHz), .D(n26559));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i26 (.Q(baudrate[17]), .C(clk16MHz), .D(n26558));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i27 (.Q(baudrate[18]), .C(clk16MHz), .D(n26557));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i28 (.Q(baudrate[19]), .C(clk16MHz), .D(n26556));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i29 (.Q(baudrate[20]), .C(clk16MHz), .D(n26555));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i30 (.Q(baudrate[21]), .C(clk16MHz), .D(n26554));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i31 (.Q(baudrate[22]), .C(clk16MHz), .D(n26553));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i32 (.Q(baudrate[23]), .C(clk16MHz), .D(n26552));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i33 (.Q(baudrate[24]), .C(clk16MHz), .D(n26551));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i34 (.Q(baudrate[25]), .C(clk16MHz), .D(n26550));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i35 (.Q(baudrate[26]), .C(clk16MHz), .D(n26549));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i36 (.Q(baudrate[27]), .C(clk16MHz), .D(n26548));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i37 (.Q(baudrate[28]), .C(clk16MHz), .D(n26547));   // verilog/eeprom.v(35[8] 81[4])
    SB_LUT4 add_1111_11_lut (.I0(n33077), .I1(delay_counter[9]), .I2(n5010[13]), 
            .I3(n46270), .O(n6532)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1111_11_lut.LUT_INIT = 16'h8228;
    SB_DFF bytes_0___i38 (.Q(baudrate[29]), .C(clk16MHz), .D(n26546));   // verilog/eeprom.v(35[8] 81[4])
    SB_CARRY add_1111_11 (.CI(n46270), .I0(delay_counter[9]), .I1(n5010[13]), 
            .CO(n46271));
    SB_DFF bytes_0___i39 (.Q(baudrate[30]), .C(clk16MHz), .D(n26545));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i40 (.Q(baudrate[31]), .C(clk16MHz), .D(n26544));   // verilog/eeprom.v(35[8] 81[4])
    SB_LUT4 add_1111_10_lut (.I0(n33077), .I1(delay_counter[8]), .I2(n5010[13]), 
            .I3(n46269), .O(n6531)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1111_10_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_1111_10 (.CI(n46269), .I0(delay_counter[8]), .I1(n5010[13]), 
            .CO(n46270));
    SB_LUT4 add_1111_9_lut (.I0(n33077), .I1(delay_counter[7]), .I2(n5010[13]), 
            .I3(n46268), .O(n6530)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1111_9_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_1111_9 (.CI(n46268), .I0(delay_counter[7]), .I1(n5010[13]), 
            .CO(n46269));
    SB_LUT4 add_1111_8_lut (.I0(n33077), .I1(delay_counter[6]), .I2(n5010[13]), 
            .I3(n46267), .O(n6529)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1111_8_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_1111_8 (.CI(n46267), .I0(delay_counter[6]), .I1(n5010[13]), 
            .CO(n46268));
    SB_LUT4 add_1111_7_lut (.I0(GND_net), .I1(delay_counter[5]), .I2(n5010[13]), 
            .I3(n46266), .O(delay_counter_15__N_3729[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1111_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1111_7 (.CI(n46266), .I0(delay_counter[5]), .I1(n5010[13]), 
            .CO(n46267));
    SB_LUT4 add_1111_6_lut (.I0(n33077), .I1(delay_counter[4]), .I2(n5010[13]), 
            .I3(n46265), .O(n6527)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1111_6_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_1111_6 (.CI(n46265), .I0(delay_counter[4]), .I1(n5010[13]), 
            .CO(n46266));
    SB_LUT4 add_1111_5_lut (.I0(GND_net), .I1(delay_counter[3]), .I2(n5010[13]), 
            .I3(n46264), .O(delay_counter_15__N_3729[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1111_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1111_5 (.CI(n46264), .I0(delay_counter[3]), .I1(n5010[13]), 
            .CO(n46265));
    SB_LUT4 add_1111_4_lut (.I0(GND_net), .I1(delay_counter[2]), .I2(n5010[13]), 
            .I3(n46263), .O(delay_counter_15__N_3729[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1111_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1111_4 (.CI(n46263), .I0(delay_counter[2]), .I1(n5010[13]), 
            .CO(n46264));
    SB_LUT4 add_1111_3_lut (.I0(GND_net), .I1(delay_counter[1]), .I2(n5010[13]), 
            .I3(n46262), .O(delay_counter_15__N_3729[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1111_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1111_3 (.CI(n46262), .I0(delay_counter[1]), .I1(n5010[13]), 
            .CO(n46263));
    SB_LUT4 add_1111_2_lut (.I0(GND_net), .I1(delay_counter[0]), .I2(n5010[13]), 
            .I3(GND_net), .O(delay_counter_15__N_3729[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1111_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1111_2 (.CI(GND_net), .I0(delay_counter[0]), .I1(n5010[13]), 
            .CO(n46262));
    SB_LUT4 i32293_3_lut_4_lut (.I0(n35339), .I1(byte_counter[0]), .I2(byte_counter[1]), 
            .I3(byte_counter[2]), .O(n17[2]));   // verilog/eeprom.v(68[25:39])
    defparam i32293_3_lut_4_lut.LUT_INIT = 16'hbf40;
    SB_LUT4 i12_4_lut (.I0(delay_counter[6]), .I1(delay_counter[10]), .I2(delay_counter[12]), 
            .I3(delay_counter[8]), .O(n28));   // verilog/eeprom.v(55[12:28])
    defparam i12_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i10_4_lut (.I0(delay_counter[7]), .I1(delay_counter[14]), .I2(delay_counter[15]), 
            .I3(delay_counter[3]), .O(n26));   // verilog/eeprom.v(55[12:28])
    defparam i10_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i11_4_lut (.I0(delay_counter[1]), .I1(delay_counter[2]), .I2(delay_counter[0]), 
            .I3(delay_counter[5]), .O(n27));   // verilog/eeprom.v(55[12:28])
    defparam i11_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i9_4_lut (.I0(delay_counter[4]), .I1(delay_counter[9]), .I2(delay_counter[13]), 
            .I3(delay_counter[11]), .O(n25));   // verilog/eeprom.v(55[12:28])
    defparam i9_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i15_4_lut (.I0(n25), .I1(n27), .I2(n26), .I3(n28), .O(n22261));   // verilog/eeprom.v(55[12:28])
    defparam i15_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 mux_1437_Mux_0_i3_4_lut (.I0(\state[0] ), .I1(enable_slow_N_3986), 
            .I2(\state[1] ), .I3(n22261), .O(n5616[0]));   // verilog/eeprom.v(38[3] 80[10])
    defparam mux_1437_Mux_0_i3_4_lut.LUT_INIT = 16'h0a4a;
    SB_LUT4 i3_4_lut (.I0(byte_counter[1]), .I1(byte_counter[2]), .I2(byte_counter[0]), 
            .I3(n47187), .O(n55498));
    defparam i3_4_lut.LUT_INIT = 16'hfdff;
    SB_LUT4 i2_3_lut (.I0(byte_counter[2]), .I1(n47187), .I2(byte_counter[0]), 
            .I3(GND_net), .O(n52876));   // verilog/eeprom.v(68[25:39])
    defparam i2_3_lut.LUT_INIT = 16'hbfbf;
    SB_LUT4 i2_2_lut (.I0(state[1]), .I1(state[2]), .I2(GND_net), .I3(GND_net), 
            .O(n7));   // verilog/eeprom.v(55[12:28])
    defparam i2_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i1_2_lut_4_lut (.I0(\state[2] ), .I1(\state[0] ), .I2(\state[1] ), 
            .I3(n3), .O(n33075));
    defparam i1_2_lut_4_lut.LUT_INIT = 16'h0406;
    SB_LUT4 i1_4_lut_4_lut (.I0(\state[2] ), .I1(\state[0] ), .I2(\state[1] ), 
            .I3(n4_c), .O(n4));
    defparam i1_4_lut_4_lut.LUT_INIT = 16'h5702;
    SB_LUT4 i41920_2_lut_3_lut (.I0(\state[0]_adj_21 ), .I1(state[1]), .I2(state[2]), 
            .I3(GND_net), .O(n56621));
    defparam i41920_2_lut_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i48350_2_lut (.I0(n22261), .I1(enable_slow_N_3986), .I2(GND_net), 
            .I3(GND_net), .O(n5010[13]));   // verilog/eeprom.v(59[18] 61[12])
    defparam i48350_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i21829_2_lut (.I0(enable_slow_N_3986), .I1(ready_prev), .I2(GND_net), 
            .I3(GND_net), .O(n35339));
    defparam i21829_2_lut.LUT_INIT = 16'hdddd;
    SB_LUT4 i1_2_lut (.I0(\state[0] ), .I1(\state[1] ), .I2(GND_net), 
            .I3(GND_net), .O(n22361));   // verilog/eeprom.v(71[5:15])
    defparam i1_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i1_4_lut (.I0(\state[2] ), .I1(\state[0] ), .I2(\state[1] ), 
            .I3(read), .O(n24676));
    defparam i1_4_lut.LUT_INIT = 16'h4140;
    SB_LUT4 i1_2_lut_3_lut_adj_1665 (.I0(enable_slow_N_3986), .I1(ready_prev), 
            .I2(byte_counter[0]), .I3(GND_net), .O(n47941));
    defparam i1_2_lut_3_lut_adj_1665.LUT_INIT = 16'hd2d2;
    SB_LUT4 i1_4_lut_adj_1666 (.I0(\state[2] ), .I1(\state[1] ), .I2(read), 
            .I3(\state[0] ), .O(n4_adj_5460));
    defparam i1_4_lut_adj_1666.LUT_INIT = 16'hbbba;
    SB_LUT4 i45383_4_lut (.I0(n56621), .I1(n22261), .I2(\state[1] ), .I3(state[3]), 
            .O(n59921));
    defparam i45383_4_lut.LUT_INIT = 16'h0010;
    SB_LUT4 i2_4_lut (.I0(n59921), .I1(n4_adj_5460), .I2(n35339), .I3(\state[0] ), 
            .O(n55256));
    defparam i2_4_lut.LUT_INIT = 16'hcfee;
    SB_LUT4 i19542_4_lut (.I0(\state[1] ), .I1(n3), .I2(\state[2] ), .I3(\state[0] ), 
            .O(state_7__N_3658[1]));   // verilog/eeprom.v(27[11:16])
    defparam i19542_4_lut.LUT_INIT = 16'ha5ba;
    SB_LUT4 i2_2_lut_4_lut (.I0(read), .I1(\state[0] ), .I2(\state[1] ), 
            .I3(\state[2] ), .O(n26045));   // verilog/eeprom.v(68[25:39])
    defparam i2_2_lut_4_lut.LUT_INIT = 16'h0002;
    SB_LUT4 i12972_3_lut_4_lut (.I0(byte_counter[2]), .I1(n52873), .I2(data[7]), 
            .I3(ID[7]), .O(n26576));   // verilog/eeprom.v(35[8] 81[4])
    defparam i12972_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i12973_3_lut_4_lut (.I0(byte_counter[2]), .I1(n52873), .I2(data[6]), 
            .I3(ID[6]), .O(n26577));   // verilog/eeprom.v(35[8] 81[4])
    defparam i12973_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i12974_3_lut_4_lut (.I0(byte_counter[2]), .I1(n52873), .I2(data[5]), 
            .I3(ID[5]), .O(n26578));   // verilog/eeprom.v(35[8] 81[4])
    defparam i12974_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i12975_3_lut_4_lut (.I0(byte_counter[2]), .I1(n52873), .I2(data[4]), 
            .I3(ID[4]), .O(n26579));   // verilog/eeprom.v(35[8] 81[4])
    defparam i12975_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i12976_3_lut_4_lut (.I0(byte_counter[2]), .I1(n52873), .I2(data[3]), 
            .I3(ID[3]), .O(n26580));   // verilog/eeprom.v(35[8] 81[4])
    defparam i12976_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i12977_3_lut_4_lut (.I0(byte_counter[2]), .I1(n52873), .I2(data[2]), 
            .I3(ID[2]), .O(n26581));   // verilog/eeprom.v(35[8] 81[4])
    defparam i12977_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i12978_3_lut_4_lut (.I0(byte_counter[2]), .I1(n52873), .I2(data[1]), 
            .I3(ID[1]), .O(n26582));   // verilog/eeprom.v(35[8] 81[4])
    defparam i12978_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i12483_3_lut_4_lut (.I0(byte_counter[2]), .I1(n52873), .I2(data[0]), 
            .I3(ID[0]), .O(n26087));   // verilog/eeprom.v(35[8] 81[4])
    defparam i12483_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i12964_3_lut_4_lut (.I0(byte_counter[1]), .I1(n52876), .I2(data[7]), 
            .I3(baudrate[7]), .O(n26568));   // verilog/eeprom.v(35[8] 81[4])
    defparam i12964_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i12965_3_lut_4_lut (.I0(byte_counter[1]), .I1(n52876), .I2(data[6]), 
            .I3(baudrate[6]), .O(n26569));   // verilog/eeprom.v(35[8] 81[4])
    defparam i12965_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i12966_3_lut_4_lut (.I0(byte_counter[1]), .I1(n52876), .I2(data[5]), 
            .I3(baudrate[5]), .O(n26570));   // verilog/eeprom.v(35[8] 81[4])
    defparam i12966_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i12967_3_lut_4_lut (.I0(byte_counter[1]), .I1(n52876), .I2(data[4]), 
            .I3(baudrate[4]), .O(n26571));   // verilog/eeprom.v(35[8] 81[4])
    defparam i12967_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i12968_3_lut_4_lut (.I0(byte_counter[1]), .I1(n52876), .I2(data[3]), 
            .I3(baudrate[3]), .O(n26572));   // verilog/eeprom.v(35[8] 81[4])
    defparam i12968_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i12969_3_lut_4_lut (.I0(byte_counter[1]), .I1(n52876), .I2(data[2]), 
            .I3(baudrate[2]), .O(n26573));   // verilog/eeprom.v(35[8] 81[4])
    defparam i12969_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i12970_3_lut_4_lut (.I0(byte_counter[1]), .I1(n52876), .I2(data[1]), 
            .I3(baudrate[1]), .O(n26574));   // verilog/eeprom.v(35[8] 81[4])
    defparam i12970_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i12971_3_lut_4_lut (.I0(byte_counter[1]), .I1(n52876), .I2(data[0]), 
            .I3(baudrate[0]), .O(n26575));   // verilog/eeprom.v(35[8] 81[4])
    defparam i12971_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i12948_3_lut_4_lut (.I0(byte_counter[1]), .I1(n52876), .I2(data[7]), 
            .I3(baudrate[23]), .O(n26552));   // verilog/eeprom.v(35[8] 81[4])
    defparam i12948_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i12949_3_lut_4_lut (.I0(byte_counter[1]), .I1(n52876), .I2(data[6]), 
            .I3(baudrate[22]), .O(n26553));   // verilog/eeprom.v(35[8] 81[4])
    defparam i12949_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i12950_3_lut_4_lut (.I0(byte_counter[1]), .I1(n52876), .I2(data[5]), 
            .I3(baudrate[21]), .O(n26554));   // verilog/eeprom.v(35[8] 81[4])
    defparam i12950_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i12951_3_lut_4_lut (.I0(byte_counter[1]), .I1(n52876), .I2(data[4]), 
            .I3(baudrate[20]), .O(n26555));   // verilog/eeprom.v(35[8] 81[4])
    defparam i12951_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i12952_3_lut_4_lut (.I0(byte_counter[1]), .I1(n52876), .I2(data[3]), 
            .I3(baudrate[19]), .O(n26556));   // verilog/eeprom.v(35[8] 81[4])
    defparam i12952_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i12953_3_lut_4_lut (.I0(byte_counter[1]), .I1(n52876), .I2(data[2]), 
            .I3(baudrate[18]), .O(n26557));   // verilog/eeprom.v(35[8] 81[4])
    defparam i12953_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i12954_3_lut_4_lut (.I0(byte_counter[1]), .I1(n52876), .I2(data[1]), 
            .I3(baudrate[17]), .O(n26558));   // verilog/eeprom.v(35[8] 81[4])
    defparam i12954_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i12955_3_lut_4_lut (.I0(byte_counter[1]), .I1(n52876), .I2(data[0]), 
            .I3(baudrate[16]), .O(n26559));   // verilog/eeprom.v(35[8] 81[4])
    defparam i12955_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i12940_3_lut_4_lut (.I0(byte_counter[2]), .I1(n52873), .I2(data[7]), 
            .I3(baudrate[31]), .O(n26544));   // verilog/eeprom.v(35[8] 81[4])
    defparam i12940_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i12941_3_lut_4_lut (.I0(byte_counter[2]), .I1(n52873), .I2(data[6]), 
            .I3(baudrate[30]), .O(n26545));   // verilog/eeprom.v(35[8] 81[4])
    defparam i12941_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i12942_3_lut_4_lut (.I0(byte_counter[2]), .I1(n52873), .I2(data[5]), 
            .I3(baudrate[29]), .O(n26546));   // verilog/eeprom.v(35[8] 81[4])
    defparam i12942_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i12943_3_lut_4_lut (.I0(byte_counter[2]), .I1(n52873), .I2(data[4]), 
            .I3(baudrate[28]), .O(n26547));   // verilog/eeprom.v(35[8] 81[4])
    defparam i12943_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i12944_3_lut_4_lut (.I0(byte_counter[2]), .I1(n52873), .I2(data[3]), 
            .I3(baudrate[27]), .O(n26548));   // verilog/eeprom.v(35[8] 81[4])
    defparam i12944_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i12945_3_lut_4_lut (.I0(byte_counter[2]), .I1(n52873), .I2(data[2]), 
            .I3(baudrate[26]), .O(n26549));   // verilog/eeprom.v(35[8] 81[4])
    defparam i12945_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i12946_3_lut_4_lut (.I0(byte_counter[2]), .I1(n52873), .I2(data[1]), 
            .I3(baudrate[25]), .O(n26550));   // verilog/eeprom.v(35[8] 81[4])
    defparam i12946_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i12947_3_lut_4_lut (.I0(byte_counter[2]), .I1(n52873), .I2(data[0]), 
            .I3(baudrate[24]), .O(n26551));   // verilog/eeprom.v(35[8] 81[4])
    defparam i12947_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i32286_2_lut_3_lut_4_lut (.I0(enable_slow_N_3986), .I1(ready_prev), 
            .I2(byte_counter[0]), .I3(byte_counter[1]), .O(n17[1]));   // verilog/eeprom.v(68[25:39])
    defparam i32286_2_lut_3_lut_4_lut.LUT_INIT = 16'hdf20;
    SB_LUT4 i3_3_lut (.I0(n56621), .I1(state[3]), .I2(n22261), .I3(GND_net), 
            .O(n55087));
    defparam i3_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i1_4_lut_adj_1667 (.I0(\state[0] ), .I1(n55087), .I2(read), 
            .I3(\state[1] ), .O(n4_c));
    defparam i1_4_lut_adj_1667.LUT_INIT = 16'hbbfa;
    SB_LUT4 i48330_3_lut_4_lut_4_lut (.I0(\state[2] ), .I1(n3), .I2(\state[0] ), 
            .I3(\state[1] ), .O(n24562));
    defparam i48330_3_lut_4_lut_4_lut.LUT_INIT = 16'h0552;
    i2c_controller i2c (.clk16MHz(clk16MHz), .GND_net(GND_net), .VCC_net(VCC_net), 
            .scl_enable(scl_enable), .\state_7__N_3883[0] (\state_7__N_3883[0] ), 
            .n26826(n26826), .data({data}), .n8(n8), .\state[0] (\state[0]_adj_21 ), 
            .enable_slow_N_3986(enable_slow_N_3986), .n6319(n6319), .\state[1] (state[1]), 
            .\state[2] (state[2]), .\state[3] (state[3]), .sda_enable(sda_enable), 
            .n35402(n35402), .n26091(n26091), .\saved_addr[0] (\saved_addr[0] ), 
            .n26080(n26080), .n26079(n26079), .n26078(n26078), .n26077(n26077), 
            .n26076(n26076), .n26075(n26075), .n26074(n26074), .n4(n4_adj_22), 
            .n4_adj_17(n4_adj_23), .n22404(n22404), .n35435(n35435), .n10(n10), 
            .\state[0]_adj_18 (\state[0] ), .\state[1]_adj_19 (\state[1] ), 
            .ready_prev(ready_prev), .n52872(n52872), .\state[2]_adj_20 (\state[2] ), 
            .n47187(n47187), .n7(n7), .\state_7__N_3899[3] (\state_7__N_3899[3] ), 
            .scl(scl), .sda_out(sda_out), .enable(enable), .n6(n6), 
            .n22380(n22380)) /* synthesis syn_noprune=1, syn_module_defined=1 */ ;   // verilog/eeprom.v(83[16] 97[4])
    
endmodule
//
// Verilog Description of module i2c_controller
//

module i2c_controller (clk16MHz, GND_net, VCC_net, scl_enable, \state_7__N_3883[0] , 
            n26826, data, n8, \state[0] , enable_slow_N_3986, n6319, 
            \state[1] , \state[2] , \state[3] , sda_enable, n35402, 
            n26091, \saved_addr[0] , n26080, n26079, n26078, n26077, 
            n26076, n26075, n26074, n4, n4_adj_17, n22404, n35435, 
            n10, \state[0]_adj_18 , \state[1]_adj_19 , ready_prev, n52872, 
            \state[2]_adj_20 , n47187, n7, \state_7__N_3899[3] , scl, 
            sda_out, enable, n6, n22380) /* synthesis syn_noprune=1, syn_module_defined=1 */ ;
    input clk16MHz;
    input GND_net;
    input VCC_net;
    output scl_enable;
    output \state_7__N_3883[0] ;
    input n26826;
    output [7:0]data;
    input n8;
    output \state[0] ;
    output enable_slow_N_3986;
    output n6319;
    output \state[1] ;
    output \state[2] ;
    output \state[3] ;
    output sda_enable;
    output n35402;
    input n26091;
    output \saved_addr[0] ;
    input n26080;
    input n26079;
    input n26078;
    input n26077;
    input n26076;
    input n26075;
    input n26074;
    output n4;
    output n4_adj_17;
    output n22404;
    output n35435;
    output n10;
    input \state[0]_adj_18 ;
    input \state[1]_adj_19 ;
    input ready_prev;
    output n52872;
    input \state[2]_adj_20 ;
    output n47187;
    input n7;
    input \state_7__N_3899[3] ;
    output scl;
    output sda_out;
    input enable;
    output n6;
    output n22380;
    
    wire clk16MHz /* synthesis SET_AS_NETWORK=clk16MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(31[6:14])
    wire i2c_clk /* synthesis is_clock=1, SET_AS_NETWORK=\eeprom/i2c/i2c_clk */ ;   // verilog/i2c_controller.v(41[6:13])
    wire [5:0]n29;
    wire [7:0]counter2;   // verilog/i2c_controller.v(37[12:20])
    
    wire n25953;
    wire [7:0]n119;
    
    wire n24601;
    wire [7:0]counter;   // verilog/i2c_controller.v(36[12:19])
    
    wire n25932, n46689, n46688, n46687, n46686, n46685, n10_c, 
        i2c_clk_N_3972, scl_enable_N_3973, enable_slow_N_3985, n24565, 
        n5, n35464, n35559, n35719, n55496, n55420, n55253, n24561, 
        n52133, n55465, n24559, sda_out_adj_5442, n11, state_7__N_3882, 
        n11_adj_5443, n4_c, n9, n46261, n46260, n46259, n46258, 
        n46257, n46256, n46255, n15, n9_adj_5446, n12, n6_c, n6312, 
        n4_adj_5451, n59922, n6642, n28, n63023, n53714;
    wire [1:0]n6382;
    
    wire n11_adj_5452, n11_adj_5453, n11_adj_5454;
    
    SB_DFFSR counter2_1952_1953__i1 (.Q(counter2[0]), .C(clk16MHz), .D(n29[0]), 
            .R(n25953));   // verilog/i2c_controller.v(69[20:35])
    SB_DFFESS counter_i1 (.Q(counter[1]), .C(i2c_clk), .E(n24601), .D(n119[1]), 
            .S(n25932));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFFESS counter_i2 (.Q(counter[2]), .C(i2c_clk), .E(n24601), .D(n119[2]), 
            .S(n25932));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFFESR counter_i3 (.Q(counter[3]), .C(i2c_clk), .E(n24601), .D(n119[3]), 
            .R(n25932));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFFESR counter_i4 (.Q(counter[4]), .C(i2c_clk), .E(n24601), .D(n119[4]), 
            .R(n25932));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFFESR counter_i5 (.Q(counter[5]), .C(i2c_clk), .E(n24601), .D(n119[5]), 
            .R(n25932));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFFESR counter_i6 (.Q(counter[6]), .C(i2c_clk), .E(n24601), .D(n119[6]), 
            .R(n25932));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFFESR counter_i7 (.Q(counter[7]), .C(i2c_clk), .E(n24601), .D(n119[7]), 
            .R(n25932));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_LUT4 counter2_1952_1953_add_4_7_lut (.I0(GND_net), .I1(GND_net), 
            .I2(counter2[5]), .I3(n46689), .O(n29[5])) /* synthesis syn_instantiated=1 */ ;
    defparam counter2_1952_1953_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 counter2_1952_1953_add_4_6_lut (.I0(GND_net), .I1(GND_net), 
            .I2(counter2[4]), .I3(n46688), .O(n29[4])) /* synthesis syn_instantiated=1 */ ;
    defparam counter2_1952_1953_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter2_1952_1953_add_4_6 (.CI(n46688), .I0(GND_net), .I1(counter2[4]), 
            .CO(n46689));
    SB_LUT4 counter2_1952_1953_add_4_5_lut (.I0(GND_net), .I1(GND_net), 
            .I2(counter2[3]), .I3(n46687), .O(n29[3])) /* synthesis syn_instantiated=1 */ ;
    defparam counter2_1952_1953_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter2_1952_1953_add_4_5 (.CI(n46687), .I0(GND_net), .I1(counter2[3]), 
            .CO(n46688));
    SB_LUT4 counter2_1952_1953_add_4_4_lut (.I0(GND_net), .I1(GND_net), 
            .I2(counter2[2]), .I3(n46686), .O(n29[2])) /* synthesis syn_instantiated=1 */ ;
    defparam counter2_1952_1953_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter2_1952_1953_add_4_4 (.CI(n46686), .I0(GND_net), .I1(counter2[2]), 
            .CO(n46687));
    SB_LUT4 counter2_1952_1953_add_4_3_lut (.I0(GND_net), .I1(GND_net), 
            .I2(counter2[1]), .I3(n46685), .O(n29[1])) /* synthesis syn_instantiated=1 */ ;
    defparam counter2_1952_1953_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter2_1952_1953_add_4_3 (.CI(n46685), .I0(GND_net), .I1(counter2[1]), 
            .CO(n46686));
    SB_LUT4 counter2_1952_1953_add_4_2_lut (.I0(GND_net), .I1(GND_net), 
            .I2(counter2[0]), .I3(VCC_net), .O(n29[0])) /* synthesis syn_instantiated=1 */ ;
    defparam counter2_1952_1953_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter2_1952_1953_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(counter2[0]), 
            .CO(n46685));
    SB_LUT4 i4_4_lut (.I0(counter2[3]), .I1(counter2[5]), .I2(counter2[2]), 
            .I3(counter2[4]), .O(n10_c));
    defparam i4_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i5_3_lut (.I0(counter2[1]), .I1(n10_c), .I2(counter2[0]), 
            .I3(GND_net), .O(n25953));
    defparam i5_3_lut.LUT_INIT = 16'h8080;
    SB_DFF i2c_clk_122 (.Q(i2c_clk), .C(clk16MHz), .D(i2c_clk_N_3972));   // verilog/i2c_controller.v(58[9] 71[5])
    SB_DFFN i2c_scl_enable_124 (.Q(scl_enable), .C(i2c_clk), .D(scl_enable_N_3973));   // verilog/i2c_controller.v(76[12] 82[6])
    SB_DFFE enable_slow_121 (.Q(\state_7__N_3883[0] ), .C(clk16MHz), .E(n24565), 
            .D(enable_slow_N_3985));   // verilog/i2c_controller.v(58[9] 71[5])
    SB_DFF data_out_i0_i0 (.Q(data[0]), .C(i2c_clk), .D(n26826));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFFE state_i0_i0 (.Q(\state[0] ), .C(i2c_clk), .E(VCC_net), .D(n8));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_LUT4 i48341_2_lut (.I0(\state_7__N_3883[0] ), .I1(enable_slow_N_3986), 
            .I2(GND_net), .I3(GND_net), .O(enable_slow_N_3985));   // verilog/i2c_controller.v(62[6:32])
    defparam i48341_2_lut.LUT_INIT = 16'hdddd;
    SB_DFFESS state_i0_i1 (.Q(\state[1] ), .C(i2c_clk), .E(n6319), .D(n5), 
            .S(n35464));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFFESS state_i0_i2 (.Q(\state[2] ), .C(i2c_clk), .E(n6319), .D(n35559), 
            .S(n35719));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFFESS state_i0_i3 (.Q(\state[3] ), .C(i2c_clk), .E(n6319), .D(n55496), 
            .S(n55420));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFFNESS write_enable_132 (.Q(sda_enable), .C(i2c_clk), .E(n24561), 
            .D(n55253), .S(n52133));   // verilog/i2c_controller.v(180[12] 218[6])
    SB_DFFNESS sda_out_133 (.Q(sda_out_adj_5442), .C(i2c_clk), .E(n24559), 
            .D(n55465), .S(n52133));   // verilog/i2c_controller.v(180[12] 218[6])
    SB_DFFESS counter_i0 (.Q(counter[0]), .C(i2c_clk), .E(n24601), .D(n119[0]), 
            .S(n25932));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_LUT4 equal_1524_i11_2_lut_3_lut_4_lut (.I0(\state[2] ), .I1(\state[3] ), 
            .I2(\state[0] ), .I3(\state[1] ), .O(n11));   // verilog/i2c_controller.v(130[5:15])
    defparam equal_1524_i11_2_lut_3_lut_4_lut.LUT_INIT = 16'hdfff;
    SB_LUT4 i21890_2_lut_3_lut (.I0(\state[2] ), .I1(\state[3] ), .I2(\state[0] ), 
            .I3(GND_net), .O(n35402));   // verilog/i2c_controller.v(130[5:15])
    defparam i21890_2_lut_3_lut.LUT_INIT = 16'hfdfd;
    SB_LUT4 i48407_3_lut_4_lut (.I0(\state[2] ), .I1(\state[3] ), .I2(n6319), 
            .I3(\state[1] ), .O(n55420));   // verilog/i2c_controller.v(130[5:15])
    defparam i48407_3_lut_4_lut.LUT_INIT = 16'h0020;
    SB_LUT4 i22191_3_lut_4_lut (.I0(\state[1] ), .I1(\state[0] ), .I2(\state[2] ), 
            .I3(\state[3] ), .O(state_7__N_3882));
    defparam i22191_3_lut_4_lut.LUT_INIT = 16'hf800;
    SB_LUT4 state_7__I_0_140_i11_2_lut_3_lut_4_lut (.I0(\state[1] ), .I1(\state[0] ), 
            .I2(\state[3] ), .I3(\state[2] ), .O(n11_adj_5443));
    defparam state_7__I_0_140_i11_2_lut_3_lut_4_lut.LUT_INIT = 16'hfff7;
    SB_DFF saved_addr__i1 (.Q(\saved_addr[0] ), .C(i2c_clk), .D(n26091));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_LUT4 i2_3_lut_4_lut (.I0(\state[2] ), .I1(\state[3] ), .I2(n4_c), 
            .I3(n9), .O(n55496));   // verilog/i2c_controller.v(77[47:62])
    defparam i2_3_lut_4_lut.LUT_INIT = 16'hf0f4;
    SB_DFF data_out_i0_i7 (.Q(data[7]), .C(i2c_clk), .D(n26080));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFF data_out_i0_i6 (.Q(data[6]), .C(i2c_clk), .D(n26079));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFF data_out_i0_i5 (.Q(data[5]), .C(i2c_clk), .D(n26078));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFF data_out_i0_i4 (.Q(data[4]), .C(i2c_clk), .D(n26077));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFF data_out_i0_i3 (.Q(data[3]), .C(i2c_clk), .D(n26076));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFF data_out_i0_i2 (.Q(data[2]), .C(i2c_clk), .D(n26075));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFF data_out_i0_i1 (.Q(data[1]), .C(i2c_clk), .D(n26074));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFFSR counter2_1952_1953__i2 (.Q(counter2[1]), .C(clk16MHz), .D(n29[1]), 
            .R(n25953));   // verilog/i2c_controller.v(69[20:35])
    SB_DFFSR counter2_1952_1953__i3 (.Q(counter2[2]), .C(clk16MHz), .D(n29[2]), 
            .R(n25953));   // verilog/i2c_controller.v(69[20:35])
    SB_DFFSR counter2_1952_1953__i4 (.Q(counter2[3]), .C(clk16MHz), .D(n29[3]), 
            .R(n25953));   // verilog/i2c_controller.v(69[20:35])
    SB_DFFSR counter2_1952_1953__i5 (.Q(counter2[4]), .C(clk16MHz), .D(n29[4]), 
            .R(n25953));   // verilog/i2c_controller.v(69[20:35])
    SB_DFFSR counter2_1952_1953__i6 (.Q(counter2[5]), .C(clk16MHz), .D(n29[5]), 
            .R(n25953));   // verilog/i2c_controller.v(69[20:35])
    SB_LUT4 sub_39_add_2_9_lut (.I0(GND_net), .I1(counter[7]), .I2(VCC_net), 
            .I3(n46261), .O(n119[7])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_39_add_2_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_39_add_2_8_lut (.I0(GND_net), .I1(counter[6]), .I2(VCC_net), 
            .I3(n46260), .O(n119[6])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_39_add_2_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_39_add_2_8 (.CI(n46260), .I0(counter[6]), .I1(VCC_net), 
            .CO(n46261));
    SB_LUT4 sub_39_add_2_7_lut (.I0(GND_net), .I1(counter[5]), .I2(VCC_net), 
            .I3(n46259), .O(n119[5])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_39_add_2_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_39_add_2_7 (.CI(n46259), .I0(counter[5]), .I1(VCC_net), 
            .CO(n46260));
    SB_LUT4 sub_39_add_2_6_lut (.I0(GND_net), .I1(counter[4]), .I2(VCC_net), 
            .I3(n46258), .O(n119[4])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_39_add_2_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_39_add_2_6 (.CI(n46258), .I0(counter[4]), .I1(VCC_net), 
            .CO(n46259));
    SB_LUT4 sub_39_add_2_5_lut (.I0(GND_net), .I1(counter[3]), .I2(VCC_net), 
            .I3(n46257), .O(n119[3])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_39_add_2_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_39_add_2_5 (.CI(n46257), .I0(counter[3]), .I1(VCC_net), 
            .CO(n46258));
    SB_LUT4 sub_39_add_2_4_lut (.I0(GND_net), .I1(counter[2]), .I2(VCC_net), 
            .I3(n46256), .O(n119[2])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_39_add_2_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_39_add_2_4 (.CI(n46256), .I0(counter[2]), .I1(VCC_net), 
            .CO(n46257));
    SB_LUT4 sub_39_add_2_3_lut (.I0(GND_net), .I1(counter[1]), .I2(VCC_net), 
            .I3(n46255), .O(n119[1])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_39_add_2_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_39_add_2_3 (.CI(n46255), .I0(counter[1]), .I1(VCC_net), 
            .CO(n46256));
    SB_LUT4 sub_39_add_2_2_lut (.I0(GND_net), .I1(counter[0]), .I2(GND_net), 
            .I3(VCC_net), .O(n119[0])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_39_add_2_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_39_add_2_2 (.CI(VCC_net), .I0(counter[0]), .I1(GND_net), 
            .CO(n46255));
    SB_LUT4 i1_2_lut (.I0(i2c_clk), .I1(n25953), .I2(GND_net), .I3(GND_net), 
            .O(i2c_clk_N_3972));
    defparam i1_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 equal_339_i4_2_lut (.I0(counter[1]), .I1(counter[2]), .I2(GND_net), 
            .I3(GND_net), .O(n4));   // verilog/i2c_controller.v(153[6:23])
    defparam equal_339_i4_2_lut.LUT_INIT = 16'hdddd;
    SB_LUT4 equal_337_i4_2_lut (.I0(counter[1]), .I1(counter[2]), .I2(GND_net), 
            .I3(GND_net), .O(n4_adj_17));   // verilog/i2c_controller.v(153[6:23])
    defparam equal_337_i4_2_lut.LUT_INIT = 16'hbbbb;
    SB_LUT4 i1_2_lut_adj_1650 (.I0(n15), .I1(counter[0]), .I2(GND_net), 
            .I3(GND_net), .O(n22404));   // verilog/i2c_controller.v(91[8] 173[6])
    defparam i1_2_lut_adj_1650.LUT_INIT = 16'hbbbb;
    SB_LUT4 i21923_2_lut (.I0(counter[1]), .I1(counter[2]), .I2(GND_net), 
            .I3(GND_net), .O(n35435));
    defparam i21923_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 equal_262_i9_2_lut (.I0(\state[0] ), .I1(\state[1] ), .I2(GND_net), 
            .I3(GND_net), .O(n9_adj_5446));   // verilog/i2c_controller.v(77[27:43])
    defparam equal_262_i9_2_lut.LUT_INIT = 16'hdddd;
    SB_LUT4 i2_2_lut (.I0(counter[2]), .I1(counter[1]), .I2(GND_net), 
            .I3(GND_net), .O(n10));   // verilog/i2c_controller.v(110[10:22])
    defparam i2_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i5_4_lut (.I0(counter[3]), .I1(counter[5]), .I2(counter[0]), 
            .I3(counter[4]), .O(n12));   // verilog/i2c_controller.v(110[10:22])
    defparam i5_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_adj_1651 (.I0(\state[0]_adj_18 ), .I1(\state[1]_adj_19 ), 
            .I2(GND_net), .I3(GND_net), .O(n6_c));
    defparam i1_2_lut_adj_1651.LUT_INIT = 16'h8888;
    SB_LUT4 i4_4_lut_adj_1652 (.I0(ready_prev), .I1(n52872), .I2(\state[2]_adj_20 ), 
            .I3(n6_c), .O(n47187));
    defparam i4_4_lut_adj_1652.LUT_INIT = 16'h0100;
    SB_LUT4 i6_4_lut (.I0(counter[6]), .I1(n12), .I2(counter[7]), .I3(n10), 
            .O(n6312));   // verilog/i2c_controller.v(110[10:22])
    defparam i6_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_adj_1653 (.I0(\state[3] ), .I1(n6312), .I2(GND_net), 
            .I3(GND_net), .O(n4_adj_5451));
    defparam i1_2_lut_adj_1653.LUT_INIT = 16'hbbbb;
    SB_LUT4 i45782_4_lut (.I0(n7), .I1(n4_adj_5451), .I2(\state[2] ), 
            .I3(\state[0] ), .O(n59922));
    defparam i45782_4_lut.LUT_INIT = 16'hfcdd;
    SB_LUT4 i14_4_lut (.I0(n59922), .I1(n9_adj_5446), .I2(n6642), .I3(\state_7__N_3899[3] ), 
            .O(n24601));
    defparam i14_4_lut.LUT_INIT = 16'h35f5;
    SB_LUT4 i21846_2_lut (.I0(i2c_clk), .I1(scl_enable), .I2(GND_net), 
            .I3(GND_net), .O(scl));   // verilog/i2c_controller.v(45[19:61])
    defparam i21846_2_lut.LUT_INIT = 16'hbbbb;
    SB_LUT4 i1_4_lut (.I0(\state[3] ), .I1(\state[1] ), .I2(\state[0] ), 
            .I3(\state[2] ), .O(n28));
    defparam i1_4_lut.LUT_INIT = 16'h5110;
    SB_LUT4 i48310_2_lut (.I0(\state[3] ), .I1(\state[1] ), .I2(GND_net), 
            .I3(GND_net), .O(n63023));
    defparam i48310_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_4_lut_adj_1654 (.I0(n11), .I1(n63023), .I2(n28), .I3(n53714), 
            .O(n24559));
    defparam i1_4_lut_adj_1654.LUT_INIT = 16'ha0a8;
    SB_LUT4 mux_1734_Mux_1_i7_4_lut (.I0(counter[1]), .I1(counter[0]), .I2(counter[2]), 
            .I3(\saved_addr[0] ), .O(n6382[1]));   // verilog/i2c_controller.v(201[28:35])
    defparam mux_1734_Mux_1_i7_4_lut.LUT_INIT = 16'hc1c0;
    SB_LUT4 i2353_2_lut (.I0(sda_out_adj_5442), .I1(sda_enable), .I2(GND_net), 
            .I3(GND_net), .O(sda_out));   // verilog/i2c_controller.v(46[9:20])
    defparam i2353_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i39054_2_lut (.I0(\state[2] ), .I1(\state[0] ), .I2(GND_net), 
            .I3(GND_net), .O(n53714));
    defparam i39054_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i3_4_lut (.I0(\state[0] ), .I1(n7), .I2(\state[3] ), .I3(n11), 
            .O(n52133));
    defparam i3_4_lut.LUT_INIT = 16'h1000;
    SB_LUT4 i1_4_lut_adj_1655 (.I0(n11), .I1(\state[1] ), .I2(\state[3] ), 
            .I3(n53714), .O(n24561));
    defparam i1_4_lut_adj_1655.LUT_INIT = 16'h0a22;
    SB_LUT4 i1_4_lut_adj_1656 (.I0(\state_7__N_3899[3] ), .I1(n11_adj_5443), 
            .I2(n11), .I3(enable), .O(n4_c));
    defparam i1_4_lut_adj_1656.LUT_INIT = 16'h2a2f;
    SB_LUT4 i48409_3_lut (.I0(n6319), .I1(n15), .I2(n11_adj_5452), .I3(GND_net), 
            .O(n35719));
    defparam i48409_3_lut.LUT_INIT = 16'h2a2a;
    SB_LUT4 i48440_2_lut (.I0(\state_7__N_3899[3] ), .I1(n11_adj_5443), 
            .I2(GND_net), .I3(GND_net), .O(n35559));
    defparam i48440_2_lut.LUT_INIT = 16'h1111;
    SB_LUT4 i48410_4_lut (.I0(n6319), .I1(\state[0] ), .I2(n11_adj_5453), 
            .I3(n7), .O(n35464));
    defparam i48410_4_lut.LUT_INIT = 16'h0a8a;
    SB_LUT4 i1_4_lut_adj_1657 (.I0(n11_adj_5454), .I1(n11_adj_5443), .I2(\state_7__N_3899[3] ), 
            .I3(\saved_addr[0] ), .O(n5));   // verilog/i2c_controller.v(92[4] 172[11])
    defparam i1_4_lut_adj_1657.LUT_INIT = 16'h5755;
    SB_LUT4 state_7__I_0_139_i11_2_lut_3_lut_4_lut (.I0(\state[2] ), .I1(\state[3] ), 
            .I2(\state[0] ), .I3(\state[1] ), .O(n11_adj_5453));   // verilog/i2c_controller.v(44[32:47])
    defparam state_7__I_0_139_i11_2_lut_3_lut_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i48361_3_lut_4_lut (.I0(\state[2] ), .I1(\state[3] ), .I2(\state[0] ), 
            .I3(\state[1] ), .O(enable_slow_N_3986));   // verilog/i2c_controller.v(44[32:47])
    defparam i48361_3_lut_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 i2_3_lut_4_lut_adj_1658 (.I0(\state[3] ), .I1(\state[1] ), .I2(\state[2] ), 
            .I3(\state[0] ), .O(n55253));   // verilog/i2c_controller.v(181[4] 217[11])
    defparam i2_3_lut_4_lut_adj_1658.LUT_INIT = 16'h1110;
    SB_LUT4 i1_2_lut_3_lut (.I0(\state[2] ), .I1(\state[3] ), .I2(\state[0] ), 
            .I3(GND_net), .O(n6642));   // verilog/i2c_controller.v(44[32:47])
    defparam i1_2_lut_3_lut.LUT_INIT = 16'h1010;
    SB_LUT4 i2_3_lut_4_lut_adj_1659 (.I0(\state[2] ), .I1(\state[3] ), .I2(n6382[1]), 
            .I3(\state[1] ), .O(n55465));   // verilog/i2c_controller.v(44[32:47])
    defparam i2_3_lut_4_lut_adj_1659.LUT_INIT = 16'h1000;
    SB_LUT4 i2_3_lut_4_lut_adj_1660 (.I0(\state[1] ), .I1(\state[2] ), .I2(\state[0] ), 
            .I3(\state[3] ), .O(n52872));
    defparam i2_3_lut_4_lut_adj_1660.LUT_INIT = 16'hfffe;
    SB_LUT4 i12333_2_lut_4_lut (.I0(n24601), .I1(\state[2] ), .I2(\state[3] ), 
            .I3(\state[0] ), .O(n25932));   // verilog/i2c_controller.v(91[8] 173[6])
    defparam i12333_2_lut_4_lut.LUT_INIT = 16'h0200;
    SB_LUT4 i39145_3_lut_4_lut (.I0(\state[0] ), .I1(\state[1] ), .I2(\state[2] ), 
            .I3(\state[3] ), .O(scl_enable_N_3973));
    defparam i39145_3_lut_4_lut.LUT_INIT = 16'hfefc;
    SB_LUT4 state_7__I_0_142_i11_2_lut_3_lut_4_lut (.I0(\state[2] ), .I1(\state[3] ), 
            .I2(\state[0] ), .I3(\state[1] ), .O(n11_adj_5452));   // verilog/i2c_controller.v(77[47:62])
    defparam state_7__I_0_142_i11_2_lut_3_lut_4_lut.LUT_INIT = 16'hffbf;
    SB_LUT4 state_7__I_0_145_i11_2_lut_3_lut_4_lut (.I0(\state[2] ), .I1(\state[3] ), 
            .I2(\state[0] ), .I3(\state[1] ), .O(n11_adj_5454));   // verilog/i2c_controller.v(130[5:15])
    defparam state_7__I_0_145_i11_2_lut_3_lut_4_lut.LUT_INIT = 16'hffdf;
    SB_LUT4 state_7__I_0_144_i11_2_lut_3_lut_4_lut (.I0(\state[2] ), .I1(\state[3] ), 
            .I2(\state[0] ), .I3(\state[1] ), .O(n15));   // verilog/i2c_controller.v(130[5:15])
    defparam state_7__I_0_144_i11_2_lut_3_lut_4_lut.LUT_INIT = 16'hfdff;
    SB_LUT4 i48328_4_lut (.I0(state_7__N_3882), .I1(n6312), .I2(n11_adj_5453), 
            .I3(n35402), .O(n6319));
    defparam i48328_4_lut.LUT_INIT = 16'h5111;
    SB_LUT4 i2_2_lut_adj_1661 (.I0(n11_adj_5453), .I1(n11_adj_5452), .I2(GND_net), 
            .I3(GND_net), .O(n6));
    defparam i2_2_lut_adj_1661.LUT_INIT = 16'h8888;
    SB_LUT4 state_7__I_0_144_i9_2_lut (.I0(\state[0] ), .I1(\state[1] ), 
            .I2(GND_net), .I3(GND_net), .O(n9));   // verilog/i2c_controller.v(151[5:14])
    defparam state_7__I_0_144_i9_2_lut.LUT_INIT = 16'hbbbb;
    SB_LUT4 i1_2_lut_adj_1662 (.I0(counter[0]), .I1(n15), .I2(GND_net), 
            .I3(GND_net), .O(n22380));   // verilog/i2c_controller.v(91[8] 173[6])
    defparam i1_2_lut_adj_1662.LUT_INIT = 16'heeee;
    SB_LUT4 i1_2_lut_3_lut_adj_1663 (.I0(enable), .I1(\state_7__N_3883[0] ), 
            .I2(enable_slow_N_3986), .I3(GND_net), .O(n24565));
    defparam i1_2_lut_3_lut_adj_1663.LUT_INIT = 16'haeae;
    
endmodule
//
// Verilog Description of module \quadrature_decoder(0)_U0 
//

module \quadrature_decoder(0)_U0  (ENCODER0_B_N_keep, n1543, ENCODER0_A_N_keep, 
            encoder0_position, GND_net, VCC_net, n26245, a_prev, n26244, 
            b_prev, position_31__N_3609, \a_new[1] , \b_new[1] , n26111, 
            n1507, debounce_cnt_N_3606) /* synthesis lattice_noprune=1 */ ;
    input ENCODER0_B_N_keep;
    input n1543;
    input ENCODER0_A_N_keep;
    output [31:0]encoder0_position;
    input GND_net;
    input VCC_net;
    input n26245;
    output a_prev;
    input n26244;
    output b_prev;
    output position_31__N_3609;
    output \a_new[1] ;
    output \b_new[1] ;
    input n26111;
    output n1507;
    output debounce_cnt_N_3606;
    
    wire [1:0]b_new;   // vhdl/quadrature_decoder.vhd(40[9:14])
    wire [1:0]a_new;   // vhdl/quadrature_decoder.vhd(39[9:14])
    wire [31:0]n133;
    
    wire direction_N_3613, n46676, n46675, n46674, n46673, n46672, 
        n46671, n46670, n46669, n46668, n46667, n46666, n46665, 
        n46664, n46663, n46662, n46661, n46660, n46659, n46658, 
        n46657, n46656, n46655, n46654, n46653, n46652, n46651, 
        n46650, n46649, n46648, n46647, n46646;
    
    SB_DFF b_new_i0 (.Q(b_new[0]), .C(n1543), .D(ENCODER0_B_N_keep));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    SB_DFF a_new_i0 (.Q(a_new[0]), .C(n1543), .D(ENCODER0_A_N_keep));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    SB_LUT4 position_1949_add_4_33_lut (.I0(GND_net), .I1(direction_N_3613), 
            .I2(encoder0_position[31]), .I3(n46676), .O(n133[31])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1949_add_4_33_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 position_1949_add_4_32_lut (.I0(GND_net), .I1(direction_N_3613), 
            .I2(encoder0_position[30]), .I3(n46675), .O(n133[30])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1949_add_4_32_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1949_add_4_32 (.CI(n46675), .I0(direction_N_3613), 
            .I1(encoder0_position[30]), .CO(n46676));
    SB_LUT4 position_1949_add_4_31_lut (.I0(GND_net), .I1(direction_N_3613), 
            .I2(encoder0_position[29]), .I3(n46674), .O(n133[29])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1949_add_4_31_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1949_add_4_31 (.CI(n46674), .I0(direction_N_3613), 
            .I1(encoder0_position[29]), .CO(n46675));
    SB_LUT4 position_1949_add_4_30_lut (.I0(GND_net), .I1(direction_N_3613), 
            .I2(encoder0_position[28]), .I3(n46673), .O(n133[28])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1949_add_4_30_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1949_add_4_30 (.CI(n46673), .I0(direction_N_3613), 
            .I1(encoder0_position[28]), .CO(n46674));
    SB_LUT4 position_1949_add_4_29_lut (.I0(GND_net), .I1(direction_N_3613), 
            .I2(encoder0_position[27]), .I3(n46672), .O(n133[27])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1949_add_4_29_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1949_add_4_29 (.CI(n46672), .I0(direction_N_3613), 
            .I1(encoder0_position[27]), .CO(n46673));
    SB_LUT4 position_1949_add_4_28_lut (.I0(GND_net), .I1(direction_N_3613), 
            .I2(encoder0_position[26]), .I3(n46671), .O(n133[26])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1949_add_4_28_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1949_add_4_28 (.CI(n46671), .I0(direction_N_3613), 
            .I1(encoder0_position[26]), .CO(n46672));
    SB_LUT4 position_1949_add_4_27_lut (.I0(GND_net), .I1(direction_N_3613), 
            .I2(encoder0_position[25]), .I3(n46670), .O(n133[25])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1949_add_4_27_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1949_add_4_27 (.CI(n46670), .I0(direction_N_3613), 
            .I1(encoder0_position[25]), .CO(n46671));
    SB_LUT4 position_1949_add_4_26_lut (.I0(GND_net), .I1(direction_N_3613), 
            .I2(encoder0_position[24]), .I3(n46669), .O(n133[24])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1949_add_4_26_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1949_add_4_26 (.CI(n46669), .I0(direction_N_3613), 
            .I1(encoder0_position[24]), .CO(n46670));
    SB_LUT4 position_1949_add_4_25_lut (.I0(GND_net), .I1(direction_N_3613), 
            .I2(encoder0_position[23]), .I3(n46668), .O(n133[23])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1949_add_4_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1949_add_4_25 (.CI(n46668), .I0(direction_N_3613), 
            .I1(encoder0_position[23]), .CO(n46669));
    SB_LUT4 position_1949_add_4_24_lut (.I0(GND_net), .I1(direction_N_3613), 
            .I2(encoder0_position[22]), .I3(n46667), .O(n133[22])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1949_add_4_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1949_add_4_24 (.CI(n46667), .I0(direction_N_3613), 
            .I1(encoder0_position[22]), .CO(n46668));
    SB_LUT4 position_1949_add_4_23_lut (.I0(GND_net), .I1(direction_N_3613), 
            .I2(encoder0_position[21]), .I3(n46666), .O(n133[21])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1949_add_4_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1949_add_4_23 (.CI(n46666), .I0(direction_N_3613), 
            .I1(encoder0_position[21]), .CO(n46667));
    SB_LUT4 position_1949_add_4_22_lut (.I0(GND_net), .I1(direction_N_3613), 
            .I2(encoder0_position[20]), .I3(n46665), .O(n133[20])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1949_add_4_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1949_add_4_22 (.CI(n46665), .I0(direction_N_3613), 
            .I1(encoder0_position[20]), .CO(n46666));
    SB_LUT4 position_1949_add_4_21_lut (.I0(GND_net), .I1(direction_N_3613), 
            .I2(encoder0_position[19]), .I3(n46664), .O(n133[19])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1949_add_4_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1949_add_4_21 (.CI(n46664), .I0(direction_N_3613), 
            .I1(encoder0_position[19]), .CO(n46665));
    SB_LUT4 position_1949_add_4_20_lut (.I0(GND_net), .I1(direction_N_3613), 
            .I2(encoder0_position[18]), .I3(n46663), .O(n133[18])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1949_add_4_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1949_add_4_20 (.CI(n46663), .I0(direction_N_3613), 
            .I1(encoder0_position[18]), .CO(n46664));
    SB_LUT4 position_1949_add_4_19_lut (.I0(GND_net), .I1(direction_N_3613), 
            .I2(encoder0_position[17]), .I3(n46662), .O(n133[17])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1949_add_4_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1949_add_4_19 (.CI(n46662), .I0(direction_N_3613), 
            .I1(encoder0_position[17]), .CO(n46663));
    SB_LUT4 position_1949_add_4_18_lut (.I0(GND_net), .I1(direction_N_3613), 
            .I2(encoder0_position[16]), .I3(n46661), .O(n133[16])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1949_add_4_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1949_add_4_18 (.CI(n46661), .I0(direction_N_3613), 
            .I1(encoder0_position[16]), .CO(n46662));
    SB_LUT4 position_1949_add_4_17_lut (.I0(GND_net), .I1(direction_N_3613), 
            .I2(encoder0_position[15]), .I3(n46660), .O(n133[15])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1949_add_4_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1949_add_4_17 (.CI(n46660), .I0(direction_N_3613), 
            .I1(encoder0_position[15]), .CO(n46661));
    SB_LUT4 position_1949_add_4_16_lut (.I0(GND_net), .I1(direction_N_3613), 
            .I2(encoder0_position[14]), .I3(n46659), .O(n133[14])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1949_add_4_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1949_add_4_16 (.CI(n46659), .I0(direction_N_3613), 
            .I1(encoder0_position[14]), .CO(n46660));
    SB_LUT4 position_1949_add_4_15_lut (.I0(GND_net), .I1(direction_N_3613), 
            .I2(encoder0_position[13]), .I3(n46658), .O(n133[13])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1949_add_4_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1949_add_4_15 (.CI(n46658), .I0(direction_N_3613), 
            .I1(encoder0_position[13]), .CO(n46659));
    SB_LUT4 position_1949_add_4_14_lut (.I0(GND_net), .I1(direction_N_3613), 
            .I2(encoder0_position[12]), .I3(n46657), .O(n133[12])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1949_add_4_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1949_add_4_14 (.CI(n46657), .I0(direction_N_3613), 
            .I1(encoder0_position[12]), .CO(n46658));
    SB_LUT4 position_1949_add_4_13_lut (.I0(GND_net), .I1(direction_N_3613), 
            .I2(encoder0_position[11]), .I3(n46656), .O(n133[11])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1949_add_4_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1949_add_4_13 (.CI(n46656), .I0(direction_N_3613), 
            .I1(encoder0_position[11]), .CO(n46657));
    SB_LUT4 position_1949_add_4_12_lut (.I0(GND_net), .I1(direction_N_3613), 
            .I2(encoder0_position[10]), .I3(n46655), .O(n133[10])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1949_add_4_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1949_add_4_12 (.CI(n46655), .I0(direction_N_3613), 
            .I1(encoder0_position[10]), .CO(n46656));
    SB_LUT4 position_1949_add_4_11_lut (.I0(GND_net), .I1(direction_N_3613), 
            .I2(encoder0_position[9]), .I3(n46654), .O(n133[9])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1949_add_4_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1949_add_4_11 (.CI(n46654), .I0(direction_N_3613), 
            .I1(encoder0_position[9]), .CO(n46655));
    SB_LUT4 position_1949_add_4_10_lut (.I0(GND_net), .I1(direction_N_3613), 
            .I2(encoder0_position[8]), .I3(n46653), .O(n133[8])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1949_add_4_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1949_add_4_10 (.CI(n46653), .I0(direction_N_3613), 
            .I1(encoder0_position[8]), .CO(n46654));
    SB_LUT4 position_1949_add_4_9_lut (.I0(GND_net), .I1(direction_N_3613), 
            .I2(encoder0_position[7]), .I3(n46652), .O(n133[7])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1949_add_4_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1949_add_4_9 (.CI(n46652), .I0(direction_N_3613), 
            .I1(encoder0_position[7]), .CO(n46653));
    SB_LUT4 position_1949_add_4_8_lut (.I0(GND_net), .I1(direction_N_3613), 
            .I2(encoder0_position[6]), .I3(n46651), .O(n133[6])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1949_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1949_add_4_8 (.CI(n46651), .I0(direction_N_3613), 
            .I1(encoder0_position[6]), .CO(n46652));
    SB_LUT4 position_1949_add_4_7_lut (.I0(GND_net), .I1(direction_N_3613), 
            .I2(encoder0_position[5]), .I3(n46650), .O(n133[5])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1949_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1949_add_4_7 (.CI(n46650), .I0(direction_N_3613), 
            .I1(encoder0_position[5]), .CO(n46651));
    SB_LUT4 position_1949_add_4_6_lut (.I0(GND_net), .I1(direction_N_3613), 
            .I2(encoder0_position[4]), .I3(n46649), .O(n133[4])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1949_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1949_add_4_6 (.CI(n46649), .I0(direction_N_3613), 
            .I1(encoder0_position[4]), .CO(n46650));
    SB_LUT4 position_1949_add_4_5_lut (.I0(GND_net), .I1(direction_N_3613), 
            .I2(encoder0_position[3]), .I3(n46648), .O(n133[3])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1949_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1949_add_4_5 (.CI(n46648), .I0(direction_N_3613), 
            .I1(encoder0_position[3]), .CO(n46649));
    SB_LUT4 position_1949_add_4_4_lut (.I0(GND_net), .I1(direction_N_3613), 
            .I2(encoder0_position[2]), .I3(n46647), .O(n133[2])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1949_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1949_add_4_4 (.CI(n46647), .I0(direction_N_3613), 
            .I1(encoder0_position[2]), .CO(n46648));
    SB_LUT4 position_1949_add_4_3_lut (.I0(GND_net), .I1(direction_N_3613), 
            .I2(encoder0_position[1]), .I3(n46646), .O(n133[1])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1949_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1949_add_4_3 (.CI(n46646), .I0(direction_N_3613), 
            .I1(encoder0_position[1]), .CO(n46647));
    SB_LUT4 position_1949_add_4_2_lut (.I0(GND_net), .I1(GND_net), .I2(encoder0_position[0]), 
            .I3(VCC_net), .O(n133[0])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1949_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1949_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(encoder0_position[0]), 
            .CO(n46646));
    SB_DFF a_prev_40 (.Q(a_prev), .C(n1543), .D(n26245));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    SB_DFF b_prev_41 (.Q(b_prev), .C(n1543), .D(n26244));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    SB_DFFE position_1949__i0 (.Q(encoder0_position[0]), .C(n1543), .E(position_31__N_3609), 
            .D(n133[0]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFF a_new_i1 (.Q(\a_new[1] ), .C(n1543), .D(a_new[0]));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    SB_DFF b_new_i1 (.Q(\b_new[1] ), .C(n1543), .D(b_new[0]));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    SB_DFF direction_42 (.Q(n1507), .C(n1543), .D(n26111));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    SB_DFFE position_1949__i1 (.Q(encoder0_position[1]), .C(n1543), .E(position_31__N_3609), 
            .D(n133[1]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1949__i2 (.Q(encoder0_position[2]), .C(n1543), .E(position_31__N_3609), 
            .D(n133[2]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1949__i3 (.Q(encoder0_position[3]), .C(n1543), .E(position_31__N_3609), 
            .D(n133[3]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1949__i4 (.Q(encoder0_position[4]), .C(n1543), .E(position_31__N_3609), 
            .D(n133[4]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1949__i5 (.Q(encoder0_position[5]), .C(n1543), .E(position_31__N_3609), 
            .D(n133[5]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1949__i6 (.Q(encoder0_position[6]), .C(n1543), .E(position_31__N_3609), 
            .D(n133[6]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1949__i7 (.Q(encoder0_position[7]), .C(n1543), .E(position_31__N_3609), 
            .D(n133[7]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1949__i8 (.Q(encoder0_position[8]), .C(n1543), .E(position_31__N_3609), 
            .D(n133[8]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1949__i9 (.Q(encoder0_position[9]), .C(n1543), .E(position_31__N_3609), 
            .D(n133[9]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1949__i10 (.Q(encoder0_position[10]), .C(n1543), .E(position_31__N_3609), 
            .D(n133[10]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1949__i11 (.Q(encoder0_position[11]), .C(n1543), .E(position_31__N_3609), 
            .D(n133[11]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1949__i12 (.Q(encoder0_position[12]), .C(n1543), .E(position_31__N_3609), 
            .D(n133[12]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1949__i13 (.Q(encoder0_position[13]), .C(n1543), .E(position_31__N_3609), 
            .D(n133[13]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1949__i14 (.Q(encoder0_position[14]), .C(n1543), .E(position_31__N_3609), 
            .D(n133[14]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1949__i15 (.Q(encoder0_position[15]), .C(n1543), .E(position_31__N_3609), 
            .D(n133[15]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1949__i16 (.Q(encoder0_position[16]), .C(n1543), .E(position_31__N_3609), 
            .D(n133[16]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1949__i17 (.Q(encoder0_position[17]), .C(n1543), .E(position_31__N_3609), 
            .D(n133[17]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1949__i18 (.Q(encoder0_position[18]), .C(n1543), .E(position_31__N_3609), 
            .D(n133[18]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1949__i19 (.Q(encoder0_position[19]), .C(n1543), .E(position_31__N_3609), 
            .D(n133[19]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1949__i20 (.Q(encoder0_position[20]), .C(n1543), .E(position_31__N_3609), 
            .D(n133[20]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1949__i21 (.Q(encoder0_position[21]), .C(n1543), .E(position_31__N_3609), 
            .D(n133[21]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1949__i22 (.Q(encoder0_position[22]), .C(n1543), .E(position_31__N_3609), 
            .D(n133[22]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1949__i23 (.Q(encoder0_position[23]), .C(n1543), .E(position_31__N_3609), 
            .D(n133[23]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1949__i24 (.Q(encoder0_position[24]), .C(n1543), .E(position_31__N_3609), 
            .D(n133[24]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1949__i25 (.Q(encoder0_position[25]), .C(n1543), .E(position_31__N_3609), 
            .D(n133[25]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1949__i26 (.Q(encoder0_position[26]), .C(n1543), .E(position_31__N_3609), 
            .D(n133[26]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1949__i27 (.Q(encoder0_position[27]), .C(n1543), .E(position_31__N_3609), 
            .D(n133[27]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1949__i28 (.Q(encoder0_position[28]), .C(n1543), .E(position_31__N_3609), 
            .D(n133[28]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1949__i29 (.Q(encoder0_position[29]), .C(n1543), .E(position_31__N_3609), 
            .D(n133[29]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1949__i30 (.Q(encoder0_position[30]), .C(n1543), .E(position_31__N_3609), 
            .D(n133[30]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1949__i31 (.Q(encoder0_position[31]), .C(n1543), .E(position_31__N_3609), 
            .D(n133[31]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_LUT4 b_prev_I_0_48_2_lut (.I0(b_prev), .I1(\a_new[1] ), .I2(GND_net), 
            .I3(GND_net), .O(direction_N_3613));   // vhdl/quadrature_decoder.vhd(64[18:37])
    defparam b_prev_I_0_48_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 position_31__I_921_4_lut (.I0(a_prev), .I1(b_prev), .I2(\a_new[1] ), 
            .I3(\b_new[1] ), .O(position_31__N_3609));   // vhdl/quadrature_decoder.vhd(63[11:57])
    defparam position_31__I_921_4_lut.LUT_INIT = 16'h7bde;
    SB_LUT4 debounce_cnt_I_920_4_lut (.I0(a_new[0]), .I1(b_new[0]), .I2(\a_new[1] ), 
            .I3(\b_new[1] ), .O(debounce_cnt_N_3606));   // vhdl/quadrature_decoder.vhd(53[8:58])
    defparam debounce_cnt_I_920_4_lut.LUT_INIT = 16'h7bde;
    
endmodule
//
// Verilog Description of module pll32MHz
//

module pll32MHz (GND_net, clk16MHz, VCC_net, clk32MHz) /* synthesis syn_module_defined=1 */ ;
    input GND_net;
    input clk16MHz;
    input VCC_net;
    output clk32MHz;
    
    wire clk16MHz /* synthesis SET_AS_NETWORK=clk16MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(31[6:14])
    wire clk32MHz /* synthesis SET_AS_NETWORK=clk32MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(31[16:24])
    
    SB_PLL40_CORE pll32MHz_inst (.REFERENCECLK(clk16MHz), .PLLOUTCORE(clk32MHz), 
            .BYPASS(GND_net), .RESETB(VCC_net)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=51, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=32, LSE_RLINE=36 */ ;   // verilog/TinyFPGA_B.v(32[10] 36[2])
    defparam pll32MHz_inst.FEEDBACK_PATH = "PHASE_AND_DELAY";
    defparam pll32MHz_inst.DELAY_ADJUSTMENT_MODE_FEEDBACK = "FIXED";
    defparam pll32MHz_inst.DELAY_ADJUSTMENT_MODE_RELATIVE = "FIXED";
    defparam pll32MHz_inst.SHIFTREG_DIV_MODE = 2'b00;
    defparam pll32MHz_inst.FDA_FEEDBACK = 4'b0000;
    defparam pll32MHz_inst.FDA_RELATIVE = 4'b0000;
    defparam pll32MHz_inst.PLLOUT_SELECT = "SHIFTREG_0deg";
    defparam pll32MHz_inst.DIVR = 4'b0000;
    defparam pll32MHz_inst.DIVF = 7'b0000001;
    defparam pll32MHz_inst.DIVQ = 3'b011;
    defparam pll32MHz_inst.FILTER_RANGE = 3'b001;
    defparam pll32MHz_inst.ENABLE_ICEGATE = 1'b0;
    defparam pll32MHz_inst.TEST_MODE = 1'b0;
    defparam pll32MHz_inst.EXTERNAL_DIVIDE_FACTOR = 1;
    
endmodule
//
// Verilog Description of module TLI4970
//

module TLI4970 (n26534, \current[7] , n26533, \current[8] , n26532, 
            \current[9] , n26531, \current[10] , n26530, \current[11] , 
            clk16MHz, n26439, \data[15] , n26437, \data[12] , n26435, 
            \data[11] , n26433, \data[10] , n26430, \data[9] , n26428, 
            \data[8] , n26427, \data[7] , n26424, \data[6] , n26422, 
            \data[5] , n26420, \data[4] , n26418, \data[3] , n26416, 
            \data[2] , GND_net, VCC_net, n26414, \data[1] , n6, 
            n6_adj_14, n5, n6_adj_15, n9, n35347, n35411, n26837, 
            \data[0] , n24517, \current[15] , CS_c, n26089, \current[0] , 
            n26540, \current[1] , n26539, \current[2] , n26538, \current[3] , 
            n26537, \current[4] , n26536, \current[5] , n26535, \current[6] , 
            n11, state_7__N_4092, CS_CLK_c, n22373, n4, n22369, 
            n22357, n22377, n4_adj_16) /* synthesis syn_noprune=1, syn_module_defined=1 */ ;
    input n26534;
    output \current[7] ;
    input n26533;
    output \current[8] ;
    input n26532;
    output \current[9] ;
    input n26531;
    output \current[10] ;
    input n26530;
    output \current[11] ;
    input clk16MHz;
    input n26439;
    output \data[15] ;
    input n26437;
    output \data[12] ;
    input n26435;
    output \data[11] ;
    input n26433;
    output \data[10] ;
    input n26430;
    output \data[9] ;
    input n26428;
    output \data[8] ;
    input n26427;
    output \data[7] ;
    input n26424;
    output \data[6] ;
    input n26422;
    output \data[5] ;
    input n26420;
    output \data[4] ;
    input n26418;
    output \data[3] ;
    input n26416;
    output \data[2] ;
    input GND_net;
    input VCC_net;
    input n26414;
    output \data[1] ;
    output n6;
    output n6_adj_14;
    output n5;
    output n6_adj_15;
    output n9;
    output n35347;
    output n35411;
    input n26837;
    output \data[0] ;
    output n24517;
    output \current[15] ;
    output CS_c;
    input n26089;
    output \current[0] ;
    input n26540;
    output \current[1] ;
    input n26539;
    output \current[2] ;
    input n26538;
    output \current[3] ;
    input n26537;
    output \current[4] ;
    input n26536;
    output \current[5] ;
    input n26535;
    output \current[6] ;
    output n11;
    output state_7__N_4092;
    output CS_CLK_c;
    output n22373;
    output n4;
    output n22369;
    output n22357;
    output n22377;
    output n4_adj_16;
    
    wire clk_slow /* synthesis is_clock=1, SET_AS_NETWORK=\tli/clk_slow */ ;   // verilog/tli4970.v(11[7:15])
    wire clk16MHz /* synthesis SET_AS_NETWORK=clk16MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(31[6:14])
    wire [7:0]n37;
    
    wire n24610;
    wire [7:0]bit_counter;   // verilog/tli4970.v(26[13:24])
    
    wire n26041, clk_slow_N_4005;
    wire [2:0]n17;
    wire [7:0]counter;   // verilog/tli4970.v(12[13:20])
    
    wire n46638, n46637;
    wire [11:0]n1;
    wire [15:0]delay_counter;   // verilog/tli4970.v(28[14:27])
    
    wire n46636, n46635, n46634, n46633, n46632, n46631, n46630, 
        n46629, n46628, n46627, n46626, n9478, n24644;
    wire [7:0]state;   // verilog/tli4970.v(29[13:18])
    
    wire n25562, n19618, delay_counter_15__N_4087, clk_slow_N_4006;
    wire [13:0]n241;
    
    wire n46581, n46580, n46579, n46578, n46577, n46576, n46575, 
        n59852, n2, n35705, n9_adj_5438, clk_out, n26095;
    wire [7:0]n47;
    
    wire n15, n55407, n12, n10, n6_adj_5440;
    
    SB_DFFN current__i8 (.Q(\current[7] ), .C(clk_slow), .D(n26534));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN current__i9 (.Q(\current[8] ), .C(clk_slow), .D(n26533));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN current__i10 (.Q(\current[9] ), .C(clk_slow), .D(n26532));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN current__i11 (.Q(\current[10] ), .C(clk_slow), .D(n26531));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN current__i12 (.Q(\current[11] ), .C(clk_slow), .D(n26530));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFNESR bit_counter_1937__i7 (.Q(bit_counter[7]), .C(clk_slow), .E(n24610), 
            .D(n37[7]), .R(n26041));   // verilog/tli4970.v(55[24:39])
    SB_DFFNESR bit_counter_1937__i6 (.Q(bit_counter[6]), .C(clk_slow), .E(n24610), 
            .D(n37[6]), .R(n26041));   // verilog/tli4970.v(55[24:39])
    SB_DFF clk_slow_63 (.Q(clk_slow), .C(clk16MHz), .D(clk_slow_N_4005));   // verilog/tli4970.v(13[10] 19[6])
    SB_DFFNESR bit_counter_1937__i5 (.Q(bit_counter[5]), .C(clk_slow), .E(n24610), 
            .D(n37[5]), .R(n26041));   // verilog/tli4970.v(55[24:39])
    SB_DFFNESR bit_counter_1937__i4 (.Q(bit_counter[4]), .C(clk_slow), .E(n24610), 
            .D(n37[4]), .R(n26041));   // verilog/tli4970.v(55[24:39])
    SB_DFFN data_i15 (.Q(\data[15] ), .C(clk_slow), .D(n26439));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN data_i12 (.Q(\data[12] ), .C(clk_slow), .D(n26437));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN data_i11 (.Q(\data[11] ), .C(clk_slow), .D(n26435));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN data_i10 (.Q(\data[10] ), .C(clk_slow), .D(n26433));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN data_i9 (.Q(\data[9] ), .C(clk_slow), .D(n26430));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN data_i8 (.Q(\data[8] ), .C(clk_slow), .D(n26428));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN data_i7 (.Q(\data[7] ), .C(clk_slow), .D(n26427));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN data_i6 (.Q(\data[6] ), .C(clk_slow), .D(n26424));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN data_i5 (.Q(\data[5] ), .C(clk_slow), .D(n26422));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN data_i4 (.Q(\data[4] ), .C(clk_slow), .D(n26420));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN data_i3 (.Q(\data[3] ), .C(clk_slow), .D(n26418));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN data_i2 (.Q(\data[2] ), .C(clk_slow), .D(n26416));   // verilog/tli4970.v(35[10] 68[6])
    SB_LUT4 counter_1945_1946_add_4_4_lut (.I0(GND_net), .I1(GND_net), .I2(counter[2]), 
            .I3(n46638), .O(n17[2])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_1945_1946_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 counter_1945_1946_add_4_3_lut (.I0(GND_net), .I1(GND_net), .I2(counter[1]), 
            .I3(n46637), .O(n17[1])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_1945_1946_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_1945_1946_add_4_3 (.CI(n46637), .I0(GND_net), .I1(counter[1]), 
            .CO(n46638));
    SB_LUT4 counter_1945_1946_add_4_2_lut (.I0(GND_net), .I1(GND_net), .I2(counter[0]), 
            .I3(VCC_net), .O(n17[0])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_1945_1946_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_DFFN data_i1 (.Q(\data[1] ), .C(clk_slow), .D(n26414));   // verilog/tli4970.v(35[10] 68[6])
    SB_CARRY counter_1945_1946_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(counter[0]), 
            .CO(n46637));
    SB_LUT4 delay_counter_1943_1944_add_4_13_lut (.I0(GND_net), .I1(GND_net), 
            .I2(delay_counter[11]), .I3(n46636), .O(n1[11])) /* synthesis syn_instantiated=1 */ ;
    defparam delay_counter_1943_1944_add_4_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 delay_counter_1943_1944_add_4_12_lut (.I0(GND_net), .I1(GND_net), 
            .I2(delay_counter[10]), .I3(n46635), .O(n1[10])) /* synthesis syn_instantiated=1 */ ;
    defparam delay_counter_1943_1944_add_4_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY delay_counter_1943_1944_add_4_12 (.CI(n46635), .I0(GND_net), 
            .I1(delay_counter[10]), .CO(n46636));
    SB_LUT4 delay_counter_1943_1944_add_4_11_lut (.I0(GND_net), .I1(GND_net), 
            .I2(delay_counter[9]), .I3(n46634), .O(n1[9])) /* synthesis syn_instantiated=1 */ ;
    defparam delay_counter_1943_1944_add_4_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY delay_counter_1943_1944_add_4_11 (.CI(n46634), .I0(GND_net), 
            .I1(delay_counter[9]), .CO(n46635));
    SB_LUT4 delay_counter_1943_1944_add_4_10_lut (.I0(GND_net), .I1(GND_net), 
            .I2(delay_counter[8]), .I3(n46633), .O(n1[8])) /* synthesis syn_instantiated=1 */ ;
    defparam delay_counter_1943_1944_add_4_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY delay_counter_1943_1944_add_4_10 (.CI(n46633), .I0(GND_net), 
            .I1(delay_counter[8]), .CO(n46634));
    SB_LUT4 delay_counter_1943_1944_add_4_9_lut (.I0(GND_net), .I1(GND_net), 
            .I2(delay_counter[7]), .I3(n46632), .O(n1[7])) /* synthesis syn_instantiated=1 */ ;
    defparam delay_counter_1943_1944_add_4_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY delay_counter_1943_1944_add_4_9 (.CI(n46632), .I0(GND_net), 
            .I1(delay_counter[7]), .CO(n46633));
    SB_LUT4 delay_counter_1943_1944_add_4_8_lut (.I0(GND_net), .I1(GND_net), 
            .I2(delay_counter[6]), .I3(n46631), .O(n1[6])) /* synthesis syn_instantiated=1 */ ;
    defparam delay_counter_1943_1944_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY delay_counter_1943_1944_add_4_8 (.CI(n46631), .I0(GND_net), 
            .I1(delay_counter[6]), .CO(n46632));
    SB_LUT4 delay_counter_1943_1944_add_4_7_lut (.I0(GND_net), .I1(GND_net), 
            .I2(delay_counter[5]), .I3(n46630), .O(n1[5])) /* synthesis syn_instantiated=1 */ ;
    defparam delay_counter_1943_1944_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY delay_counter_1943_1944_add_4_7 (.CI(n46630), .I0(GND_net), 
            .I1(delay_counter[5]), .CO(n46631));
    SB_LUT4 delay_counter_1943_1944_add_4_6_lut (.I0(GND_net), .I1(GND_net), 
            .I2(delay_counter[4]), .I3(n46629), .O(n1[4])) /* synthesis syn_instantiated=1 */ ;
    defparam delay_counter_1943_1944_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY delay_counter_1943_1944_add_4_6 (.CI(n46629), .I0(GND_net), 
            .I1(delay_counter[4]), .CO(n46630));
    SB_LUT4 delay_counter_1943_1944_add_4_5_lut (.I0(GND_net), .I1(GND_net), 
            .I2(delay_counter[3]), .I3(n46628), .O(n1[3])) /* synthesis syn_instantiated=1 */ ;
    defparam delay_counter_1943_1944_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY delay_counter_1943_1944_add_4_5 (.CI(n46628), .I0(GND_net), 
            .I1(delay_counter[3]), .CO(n46629));
    SB_LUT4 delay_counter_1943_1944_add_4_4_lut (.I0(GND_net), .I1(GND_net), 
            .I2(delay_counter[2]), .I3(n46627), .O(n1[2])) /* synthesis syn_instantiated=1 */ ;
    defparam delay_counter_1943_1944_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY delay_counter_1943_1944_add_4_4 (.CI(n46627), .I0(GND_net), 
            .I1(delay_counter[2]), .CO(n46628));
    SB_LUT4 delay_counter_1943_1944_add_4_3_lut (.I0(GND_net), .I1(GND_net), 
            .I2(delay_counter[1]), .I3(n46626), .O(n1[1])) /* synthesis syn_instantiated=1 */ ;
    defparam delay_counter_1943_1944_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY delay_counter_1943_1944_add_4_3 (.CI(n46626), .I0(GND_net), 
            .I1(delay_counter[1]), .CO(n46627));
    SB_LUT4 delay_counter_1943_1944_add_4_2_lut (.I0(GND_net), .I1(GND_net), 
            .I2(delay_counter[0]), .I3(VCC_net), .O(n1[0])) /* synthesis syn_instantiated=1 */ ;
    defparam delay_counter_1943_1944_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY delay_counter_1943_1944_add_4_2 (.CI(VCC_net), .I0(GND_net), 
            .I1(delay_counter[0]), .CO(n46626));
    SB_LUT4 equal_323_i6_2_lut (.I0(bit_counter[2]), .I1(bit_counter[3]), 
            .I2(GND_net), .I3(GND_net), .O(n6));   // verilog/tli4970.v(54[9:26])
    defparam equal_323_i6_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 equal_321_i6_2_lut (.I0(bit_counter[2]), .I1(bit_counter[3]), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_14));   // verilog/tli4970.v(54[9:26])
    defparam equal_321_i6_2_lut.LUT_INIT = 16'hdddd;
    SB_LUT4 equal_313_i5_2_lut (.I0(bit_counter[0]), .I1(bit_counter[1]), 
            .I2(GND_net), .I3(GND_net), .O(n5));   // verilog/tli4970.v(54[9:26])
    defparam equal_313_i5_2_lut.LUT_INIT = 16'hdddd;
    SB_LUT4 equal_316_i6_2_lut (.I0(bit_counter[2]), .I1(bit_counter[3]), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_15));   // verilog/tli4970.v(54[9:26])
    defparam equal_316_i6_2_lut.LUT_INIT = 16'hbbbb;
    SB_LUT4 equal_254_i9_2_lut (.I0(bit_counter[0]), .I1(bit_counter[1]), 
            .I2(GND_net), .I3(GND_net), .O(n9));   // verilog/tli4970.v(56[12:26])
    defparam equal_254_i9_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i21837_2_lut (.I0(bit_counter[0]), .I1(bit_counter[1]), .I2(GND_net), 
            .I3(GND_net), .O(n35347));
    defparam i21837_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i21899_2_lut (.I0(bit_counter[2]), .I1(bit_counter[3]), .I2(GND_net), 
            .I3(GND_net), .O(n35411));
    defparam i21899_2_lut.LUT_INIT = 16'h8888;
    SB_DFFN data_i0 (.Q(\data[0] ), .C(clk_slow), .D(n26837));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFNESR state_i1 (.Q(state[1]), .C(clk_slow), .E(n24644), .D(n9478), 
            .R(n25562));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFNE bit_counter_1937__i0 (.Q(bit_counter[0]), .C(clk_slow), .E(n24610), 
            .D(n19618));   // verilog/tli4970.v(55[24:39])
    SB_DFFNSR delay_counter_1943_1944__i1 (.Q(delay_counter[0]), .C(clk_slow), 
            .D(n1[0]), .R(delay_counter_15__N_4087));   // verilog/tli4970.v(40[24:39])
    SB_DFFSR counter_1945_1946__i1 (.Q(counter[0]), .C(clk16MHz), .D(n17[0]), 
            .R(clk_slow_N_4006));   // verilog/tli4970.v(14[16:27])
    SB_DFFNE current__i13 (.Q(\current[15] ), .C(clk_slow), .E(n24517), 
            .D(n241[13]));   // verilog/tli4970.v(35[10] 68[6])
    SB_LUT4 bit_counter_1937_add_4_9_lut (.I0(GND_net), .I1(VCC_net), .I2(bit_counter[7]), 
            .I3(n46581), .O(n37[7])) /* synthesis syn_instantiated=1 */ ;
    defparam bit_counter_1937_add_4_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 bit_counter_1937_add_4_8_lut (.I0(GND_net), .I1(VCC_net), .I2(bit_counter[6]), 
            .I3(n46580), .O(n37[6])) /* synthesis syn_instantiated=1 */ ;
    defparam bit_counter_1937_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY bit_counter_1937_add_4_8 (.CI(n46580), .I0(VCC_net), .I1(bit_counter[6]), 
            .CO(n46581));
    SB_LUT4 bit_counter_1937_add_4_7_lut (.I0(GND_net), .I1(VCC_net), .I2(bit_counter[5]), 
            .I3(n46579), .O(n37[5])) /* synthesis syn_instantiated=1 */ ;
    defparam bit_counter_1937_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY bit_counter_1937_add_4_7 (.CI(n46579), .I0(VCC_net), .I1(bit_counter[5]), 
            .CO(n46580));
    SB_LUT4 bit_counter_1937_add_4_6_lut (.I0(GND_net), .I1(VCC_net), .I2(bit_counter[4]), 
            .I3(n46578), .O(n37[4])) /* synthesis syn_instantiated=1 */ ;
    defparam bit_counter_1937_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY bit_counter_1937_add_4_6 (.CI(n46578), .I0(VCC_net), .I1(bit_counter[4]), 
            .CO(n46579));
    SB_LUT4 bit_counter_1937_add_4_5_lut (.I0(GND_net), .I1(VCC_net), .I2(bit_counter[3]), 
            .I3(n46577), .O(n37[3])) /* synthesis syn_instantiated=1 */ ;
    defparam bit_counter_1937_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY bit_counter_1937_add_4_5 (.CI(n46577), .I0(VCC_net), .I1(bit_counter[3]), 
            .CO(n46578));
    SB_LUT4 bit_counter_1937_add_4_4_lut (.I0(GND_net), .I1(VCC_net), .I2(bit_counter[2]), 
            .I3(n46576), .O(n37[2])) /* synthesis syn_instantiated=1 */ ;
    defparam bit_counter_1937_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY bit_counter_1937_add_4_4 (.CI(n46576), .I0(VCC_net), .I1(bit_counter[2]), 
            .CO(n46577));
    SB_LUT4 bit_counter_1937_add_4_3_lut (.I0(GND_net), .I1(VCC_net), .I2(bit_counter[1]), 
            .I3(n46575), .O(n37[1])) /* synthesis syn_instantiated=1 */ ;
    defparam bit_counter_1937_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY bit_counter_1937_add_4_3 (.CI(n46575), .I0(VCC_net), .I1(bit_counter[1]), 
            .CO(n46576));
    SB_LUT4 bit_counter_1937_add_4_2_lut (.I0(n2), .I1(GND_net), .I2(bit_counter[0]), 
            .I3(VCC_net), .O(n59852)) /* synthesis syn_instantiated=1 */ ;
    defparam bit_counter_1937_add_4_2_lut.LUT_INIT = 16'h8228;
    SB_CARRY bit_counter_1937_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(bit_counter[0]), 
            .CO(n46575));
    SB_DFFNESS state_i0 (.Q(state[0]), .C(clk_slow), .E(n24644), .D(n35705), 
            .S(n25562));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN clk_out_67 (.Q(clk_out), .C(clk_slow), .D(n9_adj_5438));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN slave_select_66 (.Q(CS_c), .C(clk_slow), .D(n26095));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFNE bit_counter_1937__i1 (.Q(bit_counter[1]), .C(clk_slow), .E(n24610), 
            .D(n47[1]));   // verilog/tli4970.v(55[24:39])
    SB_DFFNE bit_counter_1937__i2 (.Q(bit_counter[2]), .C(clk_slow), .E(n24610), 
            .D(n47[2]));   // verilog/tli4970.v(55[24:39])
    SB_DFFNE bit_counter_1937__i3 (.Q(bit_counter[3]), .C(clk_slow), .E(n24610), 
            .D(n47[3]));   // verilog/tli4970.v(55[24:39])
    SB_DFFN current__i1 (.Q(\current[0] ), .C(clk_slow), .D(n26089));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFNSR delay_counter_1943_1944__i2 (.Q(delay_counter[1]), .C(clk_slow), 
            .D(n1[1]), .R(delay_counter_15__N_4087));   // verilog/tli4970.v(40[24:39])
    SB_DFFNSR delay_counter_1943_1944__i3 (.Q(delay_counter[2]), .C(clk_slow), 
            .D(n1[2]), .R(delay_counter_15__N_4087));   // verilog/tli4970.v(40[24:39])
    SB_DFFNSR delay_counter_1943_1944__i4 (.Q(delay_counter[3]), .C(clk_slow), 
            .D(n1[3]), .R(delay_counter_15__N_4087));   // verilog/tli4970.v(40[24:39])
    SB_DFFNSR delay_counter_1943_1944__i5 (.Q(delay_counter[4]), .C(clk_slow), 
            .D(n1[4]), .R(delay_counter_15__N_4087));   // verilog/tli4970.v(40[24:39])
    SB_DFFNSR delay_counter_1943_1944__i6 (.Q(delay_counter[5]), .C(clk_slow), 
            .D(n1[5]), .R(delay_counter_15__N_4087));   // verilog/tli4970.v(40[24:39])
    SB_DFFNSR delay_counter_1943_1944__i7 (.Q(delay_counter[6]), .C(clk_slow), 
            .D(n1[6]), .R(delay_counter_15__N_4087));   // verilog/tli4970.v(40[24:39])
    SB_DFFNSR delay_counter_1943_1944__i8 (.Q(delay_counter[7]), .C(clk_slow), 
            .D(n1[7]), .R(delay_counter_15__N_4087));   // verilog/tli4970.v(40[24:39])
    SB_DFFNSR delay_counter_1943_1944__i9 (.Q(delay_counter[8]), .C(clk_slow), 
            .D(n1[8]), .R(delay_counter_15__N_4087));   // verilog/tli4970.v(40[24:39])
    SB_DFFNSR delay_counter_1943_1944__i10 (.Q(delay_counter[9]), .C(clk_slow), 
            .D(n1[9]), .R(delay_counter_15__N_4087));   // verilog/tli4970.v(40[24:39])
    SB_DFFNSR delay_counter_1943_1944__i11 (.Q(delay_counter[10]), .C(clk_slow), 
            .D(n1[10]), .R(delay_counter_15__N_4087));   // verilog/tli4970.v(40[24:39])
    SB_DFFNSR delay_counter_1943_1944__i12 (.Q(delay_counter[11]), .C(clk_slow), 
            .D(n1[11]), .R(delay_counter_15__N_4087));   // verilog/tli4970.v(40[24:39])
    SB_DFFSR counter_1945_1946__i2 (.Q(counter[1]), .C(clk16MHz), .D(n17[1]), 
            .R(clk_slow_N_4006));   // verilog/tli4970.v(14[16:27])
    SB_DFFSR counter_1945_1946__i3 (.Q(counter[2]), .C(clk16MHz), .D(n17[2]), 
            .R(clk_slow_N_4006));   // verilog/tli4970.v(14[16:27])
    SB_DFFN current__i2 (.Q(\current[1] ), .C(clk_slow), .D(n26540));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN current__i3 (.Q(\current[2] ), .C(clk_slow), .D(n26539));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN current__i4 (.Q(\current[3] ), .C(clk_slow), .D(n26538));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN current__i5 (.Q(\current[4] ), .C(clk_slow), .D(n26537));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN current__i6 (.Q(\current[5] ), .C(clk_slow), .D(n26536));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN current__i7 (.Q(\current[6] ), .C(clk_slow), .D(n26535));   // verilog/tli4970.v(35[10] 68[6])
    SB_LUT4 i1_2_lut_4_lut (.I0(n15), .I1(state[0]), .I2(state[1]), .I3(delay_counter_15__N_4087), 
            .O(n24644));
    defparam i1_2_lut_4_lut.LUT_INIT = 16'hffdc;
    SB_LUT4 i11958_2_lut_4_lut (.I0(n15), .I1(state[0]), .I2(state[1]), 
            .I3(delay_counter_15__N_4087), .O(n25562));
    defparam i11958_2_lut_4_lut.LUT_INIT = 16'h2300;
    SB_LUT4 i2063_3_lut (.I0(counter[0]), .I1(counter[2]), .I2(counter[1]), 
            .I3(GND_net), .O(clk_slow_N_4006));
    defparam i2063_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 clk_slow_I_0_72_2_lut (.I0(clk_slow), .I1(clk_slow_N_4006), 
            .I2(GND_net), .I3(GND_net), .O(clk_slow_N_4005));   // verilog/tli4970.v(15[5] 18[8])
    defparam clk_slow_I_0_72_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i48353_2_lut (.I0(n15), .I1(state[0]), .I2(GND_net), .I3(GND_net), 
            .O(n35705));
    defparam i48353_2_lut.LUT_INIT = 16'h1111;
    SB_LUT4 equal_254_i11_2_lut_4_lut (.I0(bit_counter[0]), .I1(bit_counter[1]), 
            .I2(bit_counter[2]), .I3(bit_counter[3]), .O(n11));   // verilog/tli4970.v(56[12:26])
    defparam equal_254_i11_2_lut_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i2322_1_lut (.I0(state[0]), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n2));
    defparam i2322_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i12437_2_lut_2_lut (.I0(state[1]), .I1(state[0]), .I2(GND_net), 
            .I3(GND_net), .O(n26041));   // verilog/tli4970.v(55[24:39])
    defparam i12437_2_lut_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 state_7__I_0_77_i9_2_lut (.I0(state[0]), .I1(state[1]), .I2(GND_net), 
            .I3(GND_net), .O(state_7__N_4092));   // verilog/tli4970.v(53[7:17])
    defparam state_7__I_0_77_i9_2_lut.LUT_INIT = 16'hbbbb;
    SB_LUT4 i2151_1_lut (.I0(\data[12] ), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n241[13]));
    defparam i2151_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i11126_2_lut (.I0(state[1]), .I1(state[0]), .I2(GND_net), 
            .I3(GND_net), .O(n24610));
    defparam i11126_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i12491_3_lut_3_lut (.I0(state[0]), .I1(state[1]), .I2(CS_c), 
            .I3(GND_net), .O(n26095));
    defparam i12491_3_lut_3_lut.LUT_INIT = 16'hd1d1;
    SB_LUT4 i48546_4_lut_4_lut (.I0(state[0]), .I1(state[1]), .I2(clk_out), 
            .I3(n15), .O(n9_adj_5438));
    defparam i48546_4_lut_4_lut.LUT_INIT = 16'hf2b2;
    SB_LUT4 i6275_3_lut (.I0(state[0]), .I1(n59852), .I2(state[1]), .I3(GND_net), 
            .O(n19618));   // verilog/tli4970.v(55[24:39])
    defparam i6275_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 bit_counter_1937_mux_6_i4_3_lut_4_lut (.I0(state[1]), .I1(state[0]), 
            .I2(state_7__N_4092), .I3(n37[3]), .O(n47[3]));
    defparam bit_counter_1937_mux_6_i4_3_lut_4_lut.LUT_INIT = 16'h4f40;
    SB_LUT4 bit_counter_1937_mux_6_i3_3_lut_4_lut (.I0(state[1]), .I1(state[0]), 
            .I2(state_7__N_4092), .I3(n37[2]), .O(n47[2]));
    defparam bit_counter_1937_mux_6_i3_3_lut_4_lut.LUT_INIT = 16'h4f40;
    SB_LUT4 bit_counter_1937_mux_6_i2_3_lut_4_lut (.I0(state[1]), .I1(state[0]), 
            .I2(state_7__N_4092), .I3(n37[1]), .O(n47[1]));
    defparam bit_counter_1937_mux_6_i2_3_lut_4_lut.LUT_INIT = 16'h4f40;
    SB_LUT4 i2_3_lut (.I0(delay_counter[1]), .I1(delay_counter[4]), .I2(delay_counter[3]), 
            .I3(GND_net), .O(n55407));
    defparam i2_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i2064_4_lut (.I0(delay_counter[0]), .I1(delay_counter[5]), .I2(delay_counter[2]), 
            .I3(n55407), .O(n12));
    defparam i2064_4_lut.LUT_INIT = 16'hccc8;
    SB_LUT4 i4_4_lut (.I0(delay_counter[11]), .I1(delay_counter[7]), .I2(delay_counter[8]), 
            .I3(delay_counter[9]), .O(n10));
    defparam i4_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i5_4_lut (.I0(delay_counter[10]), .I1(n10), .I2(n12), .I3(delay_counter[6]), 
            .O(delay_counter_15__N_4087));
    defparam i5_4_lut.LUT_INIT = 16'h8880;
    SB_LUT4 i1_2_lut (.I0(bit_counter[5]), .I1(bit_counter[4]), .I2(GND_net), 
            .I3(GND_net), .O(n6_adj_5440));   // verilog/tli4970.v(56[12:26])
    defparam i1_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i4_4_lut_adj_1644 (.I0(bit_counter[6]), .I1(bit_counter[7]), 
            .I2(n11), .I3(n6_adj_5440), .O(n15));   // verilog/tli4970.v(56[12:26])
    defparam i4_4_lut_adj_1644.LUT_INIT = 16'hfffe;
    SB_LUT4 mux_2038_i2_3_lut (.I0(n15), .I1(state[1]), .I2(state[0]), 
            .I3(GND_net), .O(n9478));
    defparam mux_2038_i2_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 spi_clk_I_0_i1_3_lut (.I0(clk_slow), .I1(clk_out), .I2(CS_c), 
            .I3(GND_net), .O(CS_CLK_c));   // verilog/tli4970.v(23[20:53])
    defparam spi_clk_I_0_i1_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i1_2_lut_4_lut_adj_1645 (.I0(state[0]), .I1(state[1]), .I2(bit_counter[0]), 
            .I3(bit_counter[1]), .O(n22373));   // verilog/tli4970.v(43[5] 67[12])
    defparam i1_2_lut_4_lut_adj_1645.LUT_INIT = 16'hbfff;
    SB_LUT4 i1_2_lut_4_lut_adj_1646 (.I0(state[0]), .I1(state[1]), .I2(bit_counter[2]), 
            .I3(bit_counter[3]), .O(n4));   // verilog/tli4970.v(43[5] 67[12])
    defparam i1_2_lut_4_lut_adj_1646.LUT_INIT = 16'hbfff;
    SB_LUT4 i1_2_lut_4_lut_adj_1647 (.I0(state[0]), .I1(state[1]), .I2(bit_counter[2]), 
            .I3(bit_counter[3]), .O(n22369));   // verilog/tli4970.v(43[5] 67[12])
    defparam i1_2_lut_4_lut_adj_1647.LUT_INIT = 16'hfbff;
    SB_LUT4 i2_3_lut_4_lut (.I0(bit_counter[0]), .I1(bit_counter[1]), .I2(state[0]), 
            .I3(state[1]), .O(n22357));   // verilog/tli4970.v(43[5] 67[12])
    defparam i2_3_lut_4_lut.LUT_INIT = 16'hfbff;
    SB_LUT4 i1_2_lut_4_lut_adj_1648 (.I0(state[0]), .I1(state[1]), .I2(bit_counter[2]), 
            .I3(bit_counter[3]), .O(n22377));   // verilog/tli4970.v(43[5] 67[12])
    defparam i1_2_lut_4_lut_adj_1648.LUT_INIT = 16'hffbf;
    SB_LUT4 i1_2_lut_4_lut_adj_1649 (.I0(state[0]), .I1(state[1]), .I2(bit_counter[2]), 
            .I3(bit_counter[3]), .O(n4_adj_16));   // verilog/tli4970.v(43[5] 67[12])
    defparam i1_2_lut_4_lut_adj_1649.LUT_INIT = 16'hfffb;
    SB_LUT4 i48332_3_lut (.I0(\data[15] ), .I1(state[1]), .I2(state[0]), 
            .I3(GND_net), .O(n24517));
    defparam i48332_3_lut.LUT_INIT = 16'h4040;
    
endmodule
//
// Verilog Description of module coms
//

module coms (VCC_net, clk16MHz, rx_data, \Kp[12] , IntegralLimit, 
            \Kp[11] , \Kp[10] , \Kp[9] , \Kp[5] , \Kp[4] , \data_in_frame[3][3] , 
            \Kp[3] , \data_in_frame[3][2] , \Kp[2] , \data_in_frame[3][1] , 
            \Kp[1] , \data_in_frame[11] , rx_data_ready, \FRAME_MATCHER.rx_data_ready_prev , 
            GND_net, deadband, \data_in_frame[3][6] , \data_in_frame[3][7] , 
            \data_in_frame[18] , n25157, n2568, \data_out_frame[0][2] , 
            n52768, \data_out_frame[0][3] , n52818, \data_out_frame[0][4] , 
            n52817, \data_out_frame[1][0] , n52816, \data_out_frame[1][1] , 
            n52815, \data_out_frame[1][3] , n52814, \FRAME_MATCHER.state[3] , 
            \data_out_frame[1][5] , n52819, \data_out_frame[1][6] , n52813, 
            \data_in_frame[18][7] , \data_out_frame[1][7] , n52812, \data_out_frame[6] , 
            \FRAME_MATCHER.i_31__N_2320 , encoder0_position, \data_out_frame[21] , 
            \data_out_frame[15] , reset, \data_out_frame[17] , \data_in_frame[1][2] , 
            \data_out_frame[22] , \data_in_frame[1][3] , setpoint, \data_out_frame[13] , 
            \data_in_frame[1][4] , \data_out_frame[11] , \data_out_frame[9] , 
            \data_out_frame[16] , byte_transmit_counter, \data_out_frame[14] , 
            \data_out_frame[4] , \data_out_frame[7] , \data_out_frame[8] , 
            \data_out_frame[12] , \data_in_frame[1][5] , \data_in_frame[1][6] , 
            \data_out_frame[3][1] , n52811, n48858, \data_out_frame[5] , 
            \data_out_frame[3][3] , n52810, \data_out_frame[3][4] , n52809, 
            \data_out_frame[3][6] , n52808, \data_out_frame[3][7] , n52807, 
            \data_out_frame[10] , n52713, n52714, n52715, n52789, 
            n52716, n52717, n52718, n52719, n52720, n52721, n52722, 
            n52723, n52724, n52806, n52725, n52726, n54590, n47777, 
            n52805, n52796, n26190, n26193, n26196, n52797, n26199, 
            n52798, n26202, n26205, \data_in_frame[1][7] , n52799, 
            n52800, n52801, n52802, n52803, n52804, n52682, control_mode, 
            n26238, n26250, n26253, n26262, n26265, n26268, \data_in_frame[4] , 
            n26271, n26274, n26291, \data_in_frame[4][6] , \control_mode[1] , 
            \control_mode[0] , n26294, \data_in_frame[4][7] , n52681, 
            n52683, n52684, \byte_transmit_counter[2] , n52685, n52686, 
            \deadband[1] , \Kp[8] , \Kp[7] , ID, \Ki[15] , \Ki[14] , 
            \Ki[13] , n26634, n27035, n26640, n25161, \control_mode[6] , 
            \control_mode[5] , n26643, n26646, n26649, n26655, n26092, 
            \control_mode[4] , n26911, n26910, n26909, n26908, current_limit, 
            n26907, n26906, n26905, n26904, n26903, n26902, n26901, 
            n26900, n26899, n26898, n26897, n26896, n26895, n26894, 
            PWMLimit, \Ki[1] , \Ki[2] , \Ki[3] , \Ki[4] , \Ki[5] , 
            \Ki[6] , \Ki[7] , \Ki[8] , \Ki[9] , \Ki[10] , \Ki[11] , 
            n52687, n7, \Ki[12] , n26687, \data_in_frame[20] , n26690, 
            \data_out_frame[26][6] , \data_out_frame[27][6] , encoder1_position, 
            n26243, n52727, n52728, n26693, n26696, n26699, n26767, 
            n26702, n26127, n26709, n26710, \Kp[13] , n26130, \data_in_frame[21] , 
            n52688, n52693, n52692, \Kp[14] , n52691, n52690, n52689, 
            n26133, n52729, n52730, n52731, n52732, n52733, n52680, 
            n52734, n52735, \Kp[15] , n52736, n52737, n52738, n52739, 
            n52740, n52741, n25663, n52742, n52743, n52744, n52745, 
            n52746, n52747, n52748, n52749, n52750, n52751, n52752, 
            n52753, n52754, n52755, n52756, n52757, n52758, n22431, 
            n15, control_update, n24502, n25620, n52759, n52760, 
            n52761, n52762, n26136, n52763, n52764, n52765, n52766, 
            n52776, n52767, n52710, n52769, n52770, n52771, n52772, 
            n52773, n52774, n52777, n52778, n52779, n52780, n52781, 
            n52782, n52783, n52775, n52795, n52786, DE_c, n26139, 
            n26142, n52700, n52701, n52793, n52792, n52784, n52785, 
            n52787, n52788, n52790, n52794, n52791, n52694, n52695, 
            n52696, n52697, n52698, n52699, n52702, n52703, n52704, 
            n52705, n52706, n52707, n52708, n52709, n52711, \Kp[6] , 
            n26083, \Ki[0] , \Kp[0] , n52712, \deadband[0] , n25123, 
            n53097, n53474, n59927, n24840, n15_adj_3, n33792, n1, 
            n32007, n19639, \current[7] , \current[6] , \current[5] , 
            \current[4] , n25127, \current[3] , \current[2] , \current[1] , 
            \current[0] , \current[15] , \current[11] , \current[10] , 
            \current[9] , \current[8] , pwm_setpoint, n52908, n59928, 
            n25141, r_Clock_Count, n24612, n36763, tx_o, n26829, 
            \r_Bit_Index[0] , \o_Rx_DV_N_3261[12] , n4837, \o_Rx_DV_N_3261[24] , 
            n29, n23, n27, n47, tx_enable, baudrate, n24621, n53789, 
            r_Clock_Count_adj_13, n26516, \r_SM_Main[2] , r_Rx_Data, 
            RX_N_42, \r_Bit_Index[0]_adj_12 , n55980, n55948, n26445, 
            \o_Rx_DV_N_3261[8] , n26443, \o_Rx_DV_N_3261[7] , \o_Rx_DV_N_3261[6] , 
            \o_Rx_DV_N_3261[5] , n33, \o_Rx_DV_N_3261[4] , \o_Rx_DV_N_3261[3] , 
            \o_Rx_DV_N_3261[2] , \o_Rx_DV_N_3261[1] , \o_Rx_DV_N_3261[0] , 
            n27051, n26970, n4834, n52823, n26836, n48959, n26832, 
            n55964, n55996, \r_SM_Main[1] , \r_SM_Main_2__N_3219[1] , 
            n55461, n26587, n26062, n55884, n55900, n55916, n55932, 
            n55814, n24535, n34) /* synthesis syn_module_defined=1 */ ;
    input VCC_net;
    input clk16MHz;
    output [7:0]rx_data;
    output \Kp[12] ;
    output [23:0]IntegralLimit;
    output \Kp[11] ;
    output \Kp[10] ;
    output \Kp[9] ;
    output \Kp[5] ;
    output \Kp[4] ;
    output \data_in_frame[3][3] ;
    output \Kp[3] ;
    output \data_in_frame[3][2] ;
    output \Kp[2] ;
    output \data_in_frame[3][1] ;
    output \Kp[1] ;
    output [7:0]\data_in_frame[11] ;
    output rx_data_ready;
    output \FRAME_MATCHER.rx_data_ready_prev ;
    input GND_net;
    output [23:0]deadband;
    output \data_in_frame[3][6] ;
    output \data_in_frame[3][7] ;
    output [7:0]\data_in_frame[18] ;
    output n25157;
    input n2568;
    output \data_out_frame[0][2] ;
    input n52768;
    output \data_out_frame[0][3] ;
    input n52818;
    output \data_out_frame[0][4] ;
    input n52817;
    output \data_out_frame[1][0] ;
    input n52816;
    output \data_out_frame[1][1] ;
    input n52815;
    output \data_out_frame[1][3] ;
    input n52814;
    output \FRAME_MATCHER.state[3] ;
    output \data_out_frame[1][5] ;
    input n52819;
    output \data_out_frame[1][6] ;
    input n52813;
    output \data_in_frame[18][7] ;
    output \data_out_frame[1][7] ;
    input n52812;
    output [7:0]\data_out_frame[6] ;
    output \FRAME_MATCHER.i_31__N_2320 ;
    input [23:0]encoder0_position;
    output [7:0]\data_out_frame[21] ;
    output [7:0]\data_out_frame[15] ;
    input reset;
    output [7:0]\data_out_frame[17] ;
    output \data_in_frame[1][2] ;
    output [7:0]\data_out_frame[22] ;
    output \data_in_frame[1][3] ;
    output [23:0]setpoint;
    output [7:0]\data_out_frame[13] ;
    output \data_in_frame[1][4] ;
    output [7:0]\data_out_frame[11] ;
    output [7:0]\data_out_frame[9] ;
    output [7:0]\data_out_frame[16] ;
    output [7:0]byte_transmit_counter;
    output [7:0]\data_out_frame[14] ;
    output [7:0]\data_out_frame[4] ;
    output [7:0]\data_out_frame[7] ;
    output [7:0]\data_out_frame[8] ;
    output [7:0]\data_out_frame[12] ;
    output \data_in_frame[1][5] ;
    output \data_in_frame[1][6] ;
    output \data_out_frame[3][1] ;
    input n52811;
    output n48858;
    output [7:0]\data_out_frame[5] ;
    output \data_out_frame[3][3] ;
    input n52810;
    output \data_out_frame[3][4] ;
    input n52809;
    output \data_out_frame[3][6] ;
    input n52808;
    output \data_out_frame[3][7] ;
    input n52807;
    output [7:0]\data_out_frame[10] ;
    input n52713;
    input n52714;
    input n52715;
    input n52789;
    input n52716;
    input n52717;
    input n52718;
    input n52719;
    input n52720;
    input n52721;
    input n52722;
    input n52723;
    input n52724;
    input n52806;
    input n52725;
    input n52726;
    output n54590;
    output n47777;
    input n52805;
    input n52796;
    input n26190;
    input n26193;
    input n26196;
    input n52797;
    input n26199;
    input n52798;
    input n26202;
    input n26205;
    output \data_in_frame[1][7] ;
    input n52799;
    input n52800;
    input n52801;
    input n52802;
    input n52803;
    input n52804;
    input n52682;
    output [7:0]control_mode;
    input n26238;
    input n26250;
    input n26253;
    input n26262;
    input n26265;
    input n26268;
    output [7:0]\data_in_frame[4] ;
    input n26271;
    input n26274;
    input n26291;
    output \data_in_frame[4][6] ;
    output \control_mode[1] ;
    output \control_mode[0] ;
    input n26294;
    output \data_in_frame[4][7] ;
    input n52681;
    input n52683;
    input n52684;
    output \byte_transmit_counter[2] ;
    input n52685;
    input n52686;
    output \deadband[1] ;
    output \Kp[8] ;
    output \Kp[7] ;
    input [7:0]ID;
    output \Ki[15] ;
    output \Ki[14] ;
    output \Ki[13] ;
    input n26634;
    input n27035;
    input n26640;
    output n25161;
    output \control_mode[6] ;
    output \control_mode[5] ;
    input n26643;
    input n26646;
    input n26649;
    input n26655;
    input n26092;
    output \control_mode[4] ;
    input n26911;
    input n26910;
    input n26909;
    input n26908;
    output [15:0]current_limit;
    input n26907;
    input n26906;
    input n26905;
    input n26904;
    input n26903;
    input n26902;
    input n26901;
    input n26900;
    input n26899;
    input n26898;
    input n26897;
    input n26896;
    input n26895;
    input n26894;
    output [23:0]PWMLimit;
    output \Ki[1] ;
    output \Ki[2] ;
    output \Ki[3] ;
    output \Ki[4] ;
    output \Ki[5] ;
    output \Ki[6] ;
    output \Ki[7] ;
    output \Ki[8] ;
    output \Ki[9] ;
    output \Ki[10] ;
    output \Ki[11] ;
    input n52687;
    output n7;
    output \Ki[12] ;
    input n26687;
    output [7:0]\data_in_frame[20] ;
    input n26690;
    output \data_out_frame[26][6] ;
    output \data_out_frame[27][6] ;
    input [23:0]encoder1_position;
    input n26243;
    input n52727;
    input n52728;
    input n26693;
    input n26696;
    input n26699;
    input n26767;
    input n26702;
    input n26127;
    input n26709;
    input n26710;
    output \Kp[13] ;
    input n26130;
    output [7:0]\data_in_frame[21] ;
    input n52688;
    input n52693;
    input n52692;
    output \Kp[14] ;
    input n52691;
    input n52690;
    input n52689;
    input n26133;
    input n52729;
    input n52730;
    input n52731;
    input n52732;
    input n52733;
    input n52680;
    input n52734;
    input n52735;
    output \Kp[15] ;
    input n52736;
    input n52737;
    input n52738;
    input n52739;
    input n52740;
    input n52741;
    input n25663;
    input n52742;
    input n52743;
    input n52744;
    input n52745;
    input n52746;
    input n52747;
    input n52748;
    input n52749;
    input n52750;
    input n52751;
    input n52752;
    input n52753;
    input n52754;
    input n52755;
    input n52756;
    input n52757;
    input n52758;
    input n22431;
    output n15;
    input control_update;
    output n24502;
    input n25620;
    input n52759;
    input n52760;
    input n52761;
    input n52762;
    input n26136;
    input n52763;
    input n52764;
    input n52765;
    input n52766;
    input n52776;
    input n52767;
    input n52710;
    input n52769;
    input n52770;
    input n52771;
    input n52772;
    input n52773;
    input n52774;
    input n52777;
    input n52778;
    input n52779;
    input n52780;
    input n52781;
    input n52782;
    input n52783;
    input n52775;
    input n52795;
    input n52786;
    output DE_c;
    input n26139;
    input n26142;
    input n52700;
    input n52701;
    input n52793;
    input n52792;
    input n52784;
    input n52785;
    input n52787;
    input n52788;
    input n52790;
    input n52794;
    input n52791;
    input n52694;
    input n52695;
    input n52696;
    input n52697;
    input n52698;
    input n52699;
    input n52702;
    input n52703;
    input n52704;
    input n52705;
    input n52706;
    input n52707;
    input n52708;
    input n52709;
    input n52711;
    output \Kp[6] ;
    input n26083;
    output \Ki[0] ;
    output \Kp[0] ;
    input n52712;
    output \deadband[0] ;
    output n25123;
    input n53097;
    output n53474;
    input n59927;
    output n24840;
    output n15_adj_3;
    output n33792;
    output n1;
    output n32007;
    output n19639;
    input \current[7] ;
    input \current[6] ;
    input \current[5] ;
    input \current[4] ;
    output n25127;
    input \current[3] ;
    input \current[2] ;
    input \current[1] ;
    input \current[0] ;
    input \current[15] ;
    input \current[11] ;
    input \current[10] ;
    input \current[9] ;
    input \current[8] ;
    input [23:0]pwm_setpoint;
    input n52908;
    input n59928;
    output n25141;
    output [8:0]r_Clock_Count;
    output n24612;
    input n36763;
    output tx_o;
    input n26829;
    output \r_Bit_Index[0] ;
    output \o_Rx_DV_N_3261[12] ;
    input n4837;
    output \o_Rx_DV_N_3261[24] ;
    output n29;
    output n23;
    output n27;
    output n47;
    output tx_enable;
    input [31:0]baudrate;
    output n24621;
    output n53789;
    output [7:0]r_Clock_Count_adj_13;
    input n26516;
    output \r_SM_Main[2] ;
    output r_Rx_Data;
    input RX_N_42;
    output \r_Bit_Index[0]_adj_12 ;
    output n55980;
    output n55948;
    input n26445;
    output \o_Rx_DV_N_3261[8] ;
    input n26443;
    output \o_Rx_DV_N_3261[7] ;
    output \o_Rx_DV_N_3261[6] ;
    output \o_Rx_DV_N_3261[5] ;
    output n33;
    output \o_Rx_DV_N_3261[4] ;
    output \o_Rx_DV_N_3261[3] ;
    output \o_Rx_DV_N_3261[2] ;
    output \o_Rx_DV_N_3261[1] ;
    output \o_Rx_DV_N_3261[0] ;
    input n27051;
    input n26970;
    input n4834;
    input n52823;
    input n26836;
    input n48959;
    input n26832;
    output n55964;
    output n55996;
    output \r_SM_Main[1] ;
    input \r_SM_Main_2__N_3219[1] ;
    output n55461;
    input n26587;
    input n26062;
    output n55884;
    output n55900;
    output n55916;
    output n55932;
    input n55814;
    output n24535;
    output n34;
    
    wire clk16MHz /* synthesis SET_AS_NETWORK=clk16MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(31[6:14])
    
    wire n26527;
    wire [7:0]\data_in_frame[6] ;   // verilog/coms.v(97[12:25])
    
    wire n8, n52882;
    wire [7:0]\data_in_frame[10] ;   // verilog/coms.v(97[12:25])
    
    wire n26066, Kp_23__N_1583, n29100;
    wire [7:0]\data_in_frame[2] ;   // verilog/coms.v(97[12:25])
    
    wire n26762;
    wire [7:0]\data_in_frame[13] ;   // verilog/coms.v(97[12:25])
    
    wire n26763, n26765, n26766, n26771;
    wire [7:0]\data_in_frame[3] ;   // verilog/coms.v(97[12:25])
    
    wire n26230, n26237, n26241, n26246, n26247, n26524;
    wire [7:0]\data_in_frame[5] ;   // verilog/coms.v(97[12:25])
    
    wire n26521, n26248, n26518, n26166;
    wire [7:0]\data_in_frame[12] ;   // verilog/coms.v(97[12:25])
    
    wire n26249, n26169, n26172, n26175, n26510;
    wire [7:0]\data_in_frame[16] ;   // verilog/coms.v(97[12:25])
    
    wire n26280, n26281, n161, n26282, n26286;
    wire [7:0]\data_in_frame[14] ;   // verilog/coms.v(97[12:25])
    
    wire n26287, n26507, n26300, n26301, n26302, n26303;
    wire [7:0]\data_in_frame[19] ;   // verilog/coms.v(97[12:25])
    wire [23:0]n4553;
    
    wire n26504, n26501;
    wire [7:0]\data_in_frame[15] ;   // verilog/coms.v(97[12:25])
    
    wire n26498, n26495, n26492, n26489, n26486, n26483, n26480, 
        \FRAME_MATCHER.i_31__N_2325 , \FRAME_MATCHER.i_31__N_2323 , \FRAME_MATCHER.i_31__N_2319 , 
        n3133, n52227, n26477, n26256, n2, n2_adj_5052;
    wire [7:0]\data_in_frame[18]_c ;   // verilog/coms.v(97[12:25])
    
    wire n2_adj_5053, n2_adj_5054, n2_adj_5055, n26474, n2_adj_5056, 
        n5, n55477, n53279, n3, n2_adj_5057, n2_adj_5058;
    wire [7:0]\data_in_frame[1] ;   // verilog/coms.v(97[12:25])
    wire [7:0]\data_in_frame[17] ;   // verilog/coms.v(97[12:25])
    
    wire n2_adj_5059;
    wire [31:0]\FRAME_MATCHER.state_31__N_2423 ;
    
    wire n2_adj_5060, n53314, n53506, n23000, n48879, n23613, n2142, 
        n53339, n22958, n1816, n53305, n23361, n52927, n53082, 
        n52931, n24563, n53453, n52998, n53568, n10, n53131, n23110, 
        n22564, n47823, n53360, n53225, n23256, n53012, n26471, 
        n1129, n53153, n6, n23417, n47860, n48851, n23629, n53462, 
        n8_adj_5061, n53459, n53524, n33_c, n53357, n48777, n47766, 
        n47853;
    wire [7:0]byte_transmit_counter_c;   // verilog/coms.v(103[12:33])
    
    wire n63473, n53020, n10_adj_5062, n54765, n52912, n53160, n12, 
        n53544, n23635, n56886, n53189, n53237, n6_adj_5063, n48773, 
        n47956, n26468, n26304, n25077, n26631, n2_adj_5064, n26465, 
        n26462, n10_adj_5065, n14, n26305, n53324, n6_adj_5066, 
        n54577, n16, n2_adj_5067, n2_adj_5068, n53397, n15_c, n53204, 
        n53026, n24, n2_adj_5069, n2_adj_5070, n26459, n53100, n23083, 
        n53535, n23_c, n22526, n25, n52992, n13, n53037, n16_adj_5071, 
        n26306, n12_adj_5072, n55050, n26307, n53412, n24_adj_5073, 
        n1667, n53256, n22, n18, n26, n53103, n53273, n8_adj_5074;
    wire [7:0]\data_in_frame[9] ;   // verilog/coms.v(97[12:25])
    
    wire n27013, n27010, n53388, n53308, n2_adj_5075, n14_adj_5076, 
        n53518, n53332, n15_adj_5077, n22529, n6_adj_5078, n53150, 
        n6_adj_5079, n63021, n21977, n27007, n23720, n53216, n26308, 
        n26309, n26310, n26311, n2_adj_5080, n2_adj_5081, n2_adj_5082, 
        n2_adj_5083, n2_adj_5084, n2_adj_5085, n2_adj_5086, n2_adj_5087, 
        n2_adj_5088, n2_adj_5089, n2_adj_5090, n2_adj_5091, n2_adj_5092, 
        n22950, n22752, n6_adj_5093, n26628, n53226, n26312, n26313, 
        n2_adj_5094, n21993, n53068, n10_adj_5095, n26314, n14_adj_5096, 
        n53088, n48497, n48787, n26456, n2_adj_5097, n53219, n6_adj_5098, 
        n26315, n48885, n6_adj_5099, n55276, n47815, n2_adj_5100, 
        n26453, n54489, n2_adj_5101, n26450, n26447, n48809, n8_adj_5102, 
        n52932, n3_adj_5103, n26625, n26178, n26444, n52175, n26319, 
        n2_adj_5104, n2_adj_5105, n2_adj_5106, n2_adj_5107, n2_adj_5108, 
        n26208, n26212, n26215, n52143, n26221, n26224, n26227, 
        n2_adj_5109, n2_adj_5110, n2_adj_5111, n2_adj_5112, n26231, 
        n26413, n26320, n26321, n26322, n26323, n26324;
    wire [23:0]deadband_c;   // verilog/TinyFPGA_B.v(237[22:30])
    
    wire n26325, n26622, n2_adj_5113, n53023, n53415, n18_adj_5114;
    wire [7:0]control_mode_c;   // verilog/TinyFPGA_B.v(234[14:26])
    
    wire n52665, n46125, n52664, n16_adj_5115, n20, n52667, n46124, 
        n52668, n46123, n52223;
    wire [7:0]\data_in_frame[4]_c ;   // verilog/coms.v(97[12:25])
    
    wire n52221, n52215, n47750, n53436, n53094, n54719, n52669, 
        n46122, n52670, n46121, n26297, n2_adj_5116, n26392;
    wire [7:0]\data_in[0] ;   // verilog/coms.v(96[12:19])
    
    wire n2_adj_5117, n2_adj_5118, n52671, n46120, n3_adj_5119;
    wire [7:0]\data_out_frame[26] ;   // verilog/coms.v(98[12:26])
    
    wire n52841, n23134, n52672, n46119, n52666, tx_transmit_N_3189, 
        n26391, n52840, n26326, n26390, n52839, n26327, n52976, 
        n22519, n6_adj_5120, n26776, n23461, n22545, n26778, n23123, 
        n53342, n26340, n53439, n14_adj_5121, n10_adj_5122, n48764, 
        n26341, n53291, n4, n10_adj_5123, n53538, n4_adj_5124, n55268, 
        n53586, n12_adj_5125, n22533, n1521, n6_adj_5126, n53515, 
        n53043, n23077, n10_adj_5127, n14_adj_5128, n53559, n53109, 
        n53391, n26342, n23126, n26343, n10_adj_5129, n26389, n26344, 
        n53113, n7_c, n8_adj_5130, n53394, n52311, n22967, n26388, 
        n26387, n26584, n52961, n26593, n26596, n26599, n26602, 
        n26605, n52163, n52181, n26615, n26619, n27031, n10_adj_5131, 
        n26386, n26385;
    wire [7:0]\data_in[1] ;   // verilog/coms.v(96[12:19])
    
    wire n27028, n27025, n27022, n27019, n27016, n26384, n14_adj_5132, 
        n10_adj_5133, n53195, n26383, n26382, n26381, n26380, n26379, 
        n26378, n27004, n27001, n23375, n26998, n26995, n52968, 
        n26992, n53501, n26377;
    wire [7:0]\data_in[2] ;   // verilog/coms.v(96[12:19])
    
    wire n10_adj_5134, n26376, n26375, n53267, n26374, n26373, n26989;
    wire [7:0]\data_in_frame[8] ;   // verilog/coms.v(97[12:25])
    
    wire n26986, n26983, n26980, n10_adj_5135, n26977, n48833, n26372, 
        n26371, n53315, n26974, n26971, n26967, n26964;
    wire [7:0]\data_in_frame[7] ;   // verilog/coms.v(97[12:25])
    
    wire n26961, n26958, n26955, n26952, n26370, n26369;
    wire [7:0]\data_in[3] ;   // verilog/coms.v(96[12:19])
    
    wire n26368, n26367, n26366, n26949, n26946, n26943, n26940, 
        n26937, n26934, n26931, n26365, n26364, n26652, n52199, 
        n26662, n26665, n26671, n52233, n26677, n26917, n26915, 
        n26914, n26913, n26912, n24833, n63273;
    wire [31:0]\FRAME_MATCHER.i ;   // verilog/coms.v(116[11:12])
    
    wire n46612, n59781, n26893, n26892, n26891, n26363, n26362, 
        n26316, n26328, n26331, n26334, n26337, n26890, n26889, 
        n26888, n26887, n26886, n26885, n26884, n26883, n26882, 
        n26881, n26880, n26879, n26878, n26877, n26876, n26875, 
        n26874, n26356, n26355, n26354, n26353, n26352, n26351, 
        n26873, n26872, n26871, n26350, n26349, n26348, n26347, 
        n26346, n26842;
    wire [7:0]\data_in_frame[0] ;   // verilog/coms.v(97[12:25])
    
    wire n26102, n63653, n2_adj_5136, n26105, n26108, n26819;
    wire [7:0]\data_in_frame[23] ;   // verilog/coms.v(97[12:25])
    
    wire n26816, n26813, n26810, n26807, n26804, n24831, n46611, 
        n59793, n24829, n46610, n59807, n24827, n46609, n59808, 
        n26345, n26112, n26800, n26797, n26794;
    wire [7:0]\data_in_frame[22] ;   // verilog/coms.v(97[12:25])
    
    wire n26791, n24825, n46608, n59809, n26788, n26785, n26782, 
        n26115, n26118, n26681, n26684, n3_adj_5138, n52838, n56844, 
        n24823, n46607, n59810, n8_adj_5139, n24821, n46606, n59811, 
        n3_adj_5140, n52837, n3_adj_5141, n52836, n3_adj_5142, n52835, 
        n3_adj_5143, n52834, n3_adj_5144;
    wire [7:0]\data_out_frame[27] ;   // verilog/coms.v(98[12:26])
    
    wire n52833, n3_adj_5145, n52832, n3_adj_5146, n52831, n3_adj_5147, 
        n52830, n3_adj_5148, n52829, n3_adj_5149, n52828, n3_adj_5150, 
        n52827, n3_adj_5151, n52826, n1_c, n1_adj_5152, n1_adj_5153, 
        n1_adj_5154, n1_adj_5155, n1_adj_5156, n1_adj_5157, n24819, 
        n46605, n59812, n2_adj_5158, n2_adj_5159, n26121, n26756, 
        n26755, n26754, n26750, n63712, \FRAME_MATCHER.i_31__N_2318 , 
        n56605, n1796, n1797, n18192, \FRAME_MATCHER.i_31__N_2322 , 
        n51969, n26713, n1808, \FRAME_MATCHER.i_31__N_2324 , n2_adj_5160, 
        n23848, n24764, n2_adj_5161, n26746, n26743, n2_adj_5162, 
        n26740, n26739, n26738, n2_adj_5163, n2_adj_5164, n2_adj_5165, 
        n26737, n35372, n52895, n22_adj_5166, n59919, n63611, n14_adj_5167, 
        n7_adj_5168;
    wire [7:0]tx_data;   // verilog/coms.v(106[13:20])
    
    wire n63605, n56853, n26736, n25071, n24817, n46604, n59813, 
        n24815, n46603, n59814, n24813, n46602, n59815, n2_adj_5169, 
        n2_adj_5170, n2_adj_5171, n2_adj_5172, n2_adj_5173, n2_adj_5174, 
        n24811, n46601, n59816, n2_adj_5175, n2_adj_5176, n26732, 
        n24809, n46600, n59829, n26729, n24807, n46599, n59838, 
        n24805, n46598, n59840, n24803, n46597, n59841, n26728, 
        n24801, n46596, n59844, n24799, n46595, n59845, n24797, 
        n46594, n59846, n26725, n26722, n26719, n24795, n46593, 
        n59847, n24793, n46592, n59848, n2_adj_5177, n2_adj_5178, 
        n2_adj_5179, n2_adj_5180, n2_adj_5181, n2_adj_5182, n2_adj_5183, 
        n24791, n46591, n59849, n2_adj_5184, n2_adj_5185, n2_adj_5186, 
        n2_adj_5187, n2_adj_5188, n2_adj_5189, n2_adj_5190, n2_adj_5191, 
        n2_adj_5192, n2_adj_5193, n2_adj_5194, n2_adj_5195, n2_adj_5196, 
        n2_adj_5197, n2_adj_5198, n24789, n46590, n59850, n2_adj_5199, 
        n26716, n24787, n46589, n59853, n24785, n46588, n59855, 
        n2_adj_5200, n24783, n46587, n59856, n24781, n46586, n59857, 
        n24779, n46585, n59862, n24777, n46584, n59869, n24775, 
        n46583, n59870, n24773, n46582, n59871;
    wire [31:0]n133;
    
    wire n8_adj_5202, n53495, n53521, n7_adj_5203, n53492, n48923, 
        n53246, n54876, n55195, n52980, n2_adj_5204, n2_adj_5205, 
        n2_adj_5206, n22677, n2_adj_5207, n47932, n53163, n53321, 
        n52, n52921, n52995, n22631, n50, n22623, n53264, n48511, 
        n51, n49, n2_adj_5208, n26705, Kp_23__N_1224, n48800, n47783, 
        n56, n53298, n52940, n53249, Kp_23__N_902, n54, n2_adj_5209, 
        n48783, n55, n47756, n48785, n53512, n53, n62, n61, 
        n22_adj_5210, n53556, n28, n53409, n53222, n53234, n53079, 
        n36, n53583, n26_adj_5211, n34_c, n37, n53598, n39, n33_adj_5212, 
        n48295, n47898, n48794, n12_adj_5213, n22056, n53489, n53240, 
        n53228, n23039, n55031, n53370, n53366, n47764, n53091, 
        n47849, n53529, n23402, n23006, n48781, n53532, n18_adj_5214, 
        n48942, n52952, n24_adj_5215, n53375, n52937, n22_adj_5216, 
        n53468, n26_adj_5217, n22822, n23002, n53329, n48904, n52946, 
        n10_adj_5218, n54710, n22042, n53015, n47882, n10_adj_5219, 
        n48844, n53147, n48768, n8_adj_5220, n53363, n53085, n48813, 
        n22898, n23343, n53171, n48798, n48392, n53348, n53252, 
        n7_adj_5221, n54891, n53276, n63383, n23509, n53352, n2_adj_5222, 
        n2_adj_5223, n2_adj_5224, n2_adj_5225, n2_adj_5226, n2_adj_5227, 
        n2_adj_5228, n2_adj_5229, n2_adj_5230, n2_adj_5231, n2_adj_5232, 
        n2_adj_5233, n2_adj_5234, n2_adj_5235, n2_adj_5236, n2_adj_5237, 
        n2_adj_5238, n2_adj_5239, n2_adj_5240, n2_adj_5241, n2_adj_5242, 
        n2_adj_5243, n1_adj_5244;
    wire [2:0]r_SM_Main_2__N_3318;
    
    wire n25577, n23764, n25576, n53577, n1_adj_5245, n26101, n6_adj_5246, 
        n20730, n53509, n22837, n10_adj_5247, n26680, n26661, n2_adj_5248, 
        n2_adj_5249, n2_adj_5250, n2_adj_5251, n2_adj_5252, n2_adj_5253, 
        n2_adj_5254, n2_adj_5255, n2_adj_5256, n2_adj_5257, n2_adj_5258, 
        n2_adj_5259, n2_adj_5260, n2_adj_5261, n2_adj_5262, n2_adj_5263, 
        n2_adj_5264, n2_adj_5265, n2_adj_5266, n2_adj_5267, n2_adj_5268, 
        n2_adj_5269, n2_adj_5270, n2_adj_5271, n2_adj_5272, n2_adj_5273, 
        n26145, n26086, n26084, n26082, n26081, n3_adj_5274, n23288, 
        n52890, n48, n53607, n53592, n46, n26608, n26592, n53553, 
        n53125, n53288, n47_c, n53430, n53034, n45, n53285, n53595, 
        n44, n26148, n26151, n26589, n26154, n26583, n53571, n43, 
        n54_adj_5275, n48415, n49_adj_5276, n26157, n26072, n26160, 
        n26163, n7_adj_5277, n23201, n53004, n23152, n22610, n22828, 
        n23193, n23753, n22658, n22813, n23553, n53378, n26065, 
        n6_adj_5278, n53106, n53186, n23252, n53345, n52915, n22688, 
        n23479, n2_adj_5279, n26064, n10_adj_5280, n53712, n6_adj_5281, 
        n10_adj_5282, n23620, n48354, n53427, n53541, n6_adj_5283, 
        n6_adj_5284, Kp_23__N_1106, n53001, n23144, n22843, n6_adj_5285, 
        n20816, n52934, n47554, n47795, n8_adj_5286, n53168, n23221, 
        n53449, n10_adj_5287, n53565, n28_adj_5288, n32, n22594, 
        n53465, n30, n53403, n31, n23046, Kp_23__N_679, n29_c, 
        n6_adj_5289, n53550, n53424, n20672, n23506, n53471, n53135, 
        n23666, n53198, n22652, n6_adj_5290, Kp_23__N_550, n63386, 
        n53157, n23536, n52972, n53601, n6_adj_5291, n53243, n53073, 
        n33_adj_5292, n6_adj_5293, n53418, n53076, n53547, n53065, 
        Kp_23__N_704, Kp_23__N_710, n22713, n53007, n53116, n53192, 
        n6_adj_5294, n53406, n10_adj_5295, n52986, Kp_23__N_607, n53029, 
        n28_adj_5296, n26_adj_5297, n53318, n53058, n27_c, n53589, 
        n25_adj_5298, n53174, n20651, n53213, n16_adj_5299, n53141, 
        n53456, n17, n55110, n52989, n28_adj_5300, n53445, n26_adj_5301, 
        n27_adj_5302, n25_adj_5303, n47950, n16_adj_5304, n53183, 
        n22_adj_5305, n20_adj_5306, n24_adj_5307, Kp_23__N_915, n55472, 
        n16_adj_5308, n17_adj_5309, n22818, n6_adj_5310, Kp_23__N_602, 
        n53050, n21971, n47851, n53498, n48824, n6_adj_5311, n6_adj_5312, 
        n53458, Kp_23__N_920, n23741, n55482, n53207, n6_adj_5313, 
        n16_adj_5314, n17_adj_5315, n48239, n53253, n14_adj_5316, 
        n15_adj_5317, n10_adj_5318, n22021, n53311, n6_adj_5319, n47876, 
        n52924, n10_adj_5320, n8_adj_5321, n53400, n10_adj_5322, n12_adj_5323, 
        n54668, n54475, n6_adj_5324, n54715, n5_adj_5325, n10_adj_5326, 
        n55426, n18_adj_5327, n63878, n54852, n5_adj_5328, n6_adj_5329, 
        n54458, n54948, n54867, n54619, n12_adj_5330, n54950, n9, 
        n20_adj_5331, n54880, n28_adj_5332, n55002, n10_adj_5333, 
        n26_adj_5334, n56589, n8_adj_5335, n29_adj_5336, n31_adj_5337, 
        n25103, n56574, n10_adj_5338, n56576, n20820, n30_adj_5339, 
        n22_adj_5340, n56578, n32_adj_5341, n56724, n22333, n16_adj_5342, 
        n17_adj_5343, n55383, n55141, n55476, n29111, n4425, n1702, 
        n1705, n54660, n18_adj_5344, n16_adj_5345, n20_adj_5346, n4_adj_5347, 
        n54478, n22428, n56872, n21, n24742, n56927, n56928, n56926, 
        n63320, n14_adj_5348, n16_adj_5349, n61988, n61989, n56833, 
        n56834, n56945, n56944, n56941, n56942, n57008, n57007, 
        n56923, n56924, n59727, n59726, n24714, n56930, n56931, 
        n56929, n1_adj_5350, n56863, n59910, n21_adj_5351, n16_adj_5352, 
        n22_adj_5353, n56918, n24853, n56919, n56917, n59912, n21_adj_5354, 
        n16_adj_5355, n22_adj_5356, n63557, n63332, n7_adj_5358, n17_adj_5360, 
        n47634, n53144, n29098, n63302, n63371, n48790, n14_adj_5361, 
        n53574, n55349, n48259, n15_adj_5362, n63533, n56864, n63374, 
        n63326, n7_adj_5363, tx_active, n44_adj_5364, n22342, n5_adj_5365, 
        n52615, n3302, n771, n63527, n56597, Kp_23__N_583, n24_adj_5366, 
        n52983, n24745, n56933, n56934, n56932, n63338, n63284, 
        n53122, n21_adj_5367, n16_adj_5368, n53201, n33004, n16_adj_5369, 
        n61082, n56914, n12_adj_5370, n10_adj_5371, n56915, n56951, 
        n56916, n57324, n56952, n63296, n11, n21_adj_5372, n16_adj_5373, 
        n24_adj_5374, n22_adj_5375, n57080, n7_adj_5376, n21_adj_5377, 
        n9_adj_5378, n16_adj_5379, n24_adj_5380, n22_adj_5381, n56846, 
        n63290, n10_adj_5382, n52956, n33453, n56920, n56921, n56922, 
        n22_adj_5383, n27_adj_5384, n26_adj_5385, n29_adj_5386, n31_adj_5387, 
        n18187, n19648, n29112, n5_adj_5388, n1703, n22258, n30_adj_5389, 
        n52879, n54832, n10_adj_5390, n14_adj_5391, n22352, n20_adj_5392, 
        n22277, n19, n56728, n22425, n18_adj_5393, n22419, n20_adj_5394, 
        n15_adj_5395, n10_adj_5396, n56730, n15_adj_5397, n16_adj_5398, 
        n17_adj_5399, n16_adj_5400, n17_adj_5401, n4_adj_5402, n6_adj_5403, 
        n36757, n48758, n53335, n53477, n22_adj_5404, n24_adj_5405, 
        n20_adj_5406, n23272, n48935, n53282, n26_adj_5407, n53302, 
        n24_adj_5408, n25_adj_5409, n23712, n23_adj_5410, n18_adj_5411, 
        n19_adj_5412, n12_adj_5413, n23432, n13_adj_5414, n54606, 
        n12_adj_5415, n15_adj_5416, n8_adj_5417, n12_adj_5418, n63335, 
        n53580, n63497, n56873, n10_adj_5419, n63329, n63491, n63323, 
        n63317, n63311, n63305, n56961, n63299, n56877, n63293, 
        n63287, n63281;
    
    SB_DFFE data_in_frame_0___i49 (.Q(\data_in_frame[6] [0]), .C(clk16MHz), 
            .E(VCC_net), .D(n26527));   // verilog/coms.v(128[12] 296[6])
    SB_LUT4 i12462_3_lut_4_lut (.I0(n8), .I1(n52882), .I2(rx_data[6]), 
            .I3(\data_in_frame[10] [6]), .O(n26066));
    defparam i12462_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13158_3_lut_4_lut (.I0(Kp_23__N_1583), .I1(n29100), .I2(\data_in_frame[2] [4]), 
            .I3(\Kp[12] ), .O(n26762));
    defparam i13158_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i13159_3_lut_4_lut (.I0(Kp_23__N_1583), .I1(n29100), .I2(\data_in_frame[13] [1]), 
            .I3(IntegralLimit[1]), .O(n26763));
    defparam i13159_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i13161_3_lut_4_lut (.I0(Kp_23__N_1583), .I1(n29100), .I2(\data_in_frame[2] [3]), 
            .I3(\Kp[11] ), .O(n26765));
    defparam i13161_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i13162_3_lut_4_lut (.I0(Kp_23__N_1583), .I1(n29100), .I2(\data_in_frame[2] [2]), 
            .I3(\Kp[10] ), .O(n26766));
    defparam i13162_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i13167_3_lut_4_lut (.I0(Kp_23__N_1583), .I1(n29100), .I2(\data_in_frame[2] [1]), 
            .I3(\Kp[9] ), .O(n26771));
    defparam i13167_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i12626_3_lut_4_lut (.I0(Kp_23__N_1583), .I1(n29100), .I2(\data_in_frame[3] [5]), 
            .I3(\Kp[5] ), .O(n26230));
    defparam i12626_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i17222_3_lut_4_lut (.I0(Kp_23__N_1583), .I1(n29100), .I2(\data_in_frame[3] [4]), 
            .I3(\Kp[4] ), .O(n26237));
    defparam i17222_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i12637_3_lut_4_lut (.I0(Kp_23__N_1583), .I1(n29100), .I2(\data_in_frame[3][3] ), 
            .I3(\Kp[3] ), .O(n26241));
    defparam i12637_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i12642_3_lut_4_lut (.I0(Kp_23__N_1583), .I1(n29100), .I2(\data_in_frame[3][2] ), 
            .I3(\Kp[2] ), .O(n26246));
    defparam i12642_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i12643_3_lut_4_lut (.I0(Kp_23__N_1583), .I1(n29100), .I2(\data_in_frame[3][1] ), 
            .I3(\Kp[1] ), .O(n26247));
    defparam i12643_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFFE data_in_frame_0___i48 (.Q(\data_in_frame[5] [7]), .C(clk16MHz), 
            .E(VCC_net), .D(n26524));   // verilog/coms.v(128[12] 296[6])
    SB_DFFE data_in_frame_0___i47 (.Q(\data_in_frame[5] [6]), .C(clk16MHz), 
            .E(VCC_net), .D(n26521));   // verilog/coms.v(128[12] 296[6])
    SB_LUT4 i12644_3_lut_4_lut (.I0(Kp_23__N_1583), .I1(n29100), .I2(\data_in_frame[11] [7]), 
            .I3(IntegralLimit[23]), .O(n26248));
    defparam i12644_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFFE data_in_frame_0___i46 (.Q(\data_in_frame[5] [5]), .C(clk16MHz), 
            .E(VCC_net), .D(n26518));   // verilog/coms.v(128[12] 296[6])
    SB_DFF data_in_frame_0___i104 (.Q(\data_in_frame[12] [7]), .C(clk16MHz), 
           .D(n26166));   // verilog/coms.v(128[12] 296[6])
    SB_LUT4 i12645_3_lut_4_lut (.I0(Kp_23__N_1583), .I1(n29100), .I2(\data_in_frame[11] [6]), 
            .I3(IntegralLimit[22]), .O(n26249));
    defparam i12645_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFF data_in_frame_0___i105 (.Q(\data_in_frame[13] [0]), .C(clk16MHz), 
           .D(n26169));   // verilog/coms.v(128[12] 296[6])
    SB_DFF data_in_frame_0___i106 (.Q(\data_in_frame[13] [1]), .C(clk16MHz), 
           .D(n26172));   // verilog/coms.v(128[12] 296[6])
    SB_DFF data_in_frame_0___i107 (.Q(\data_in_frame[13] [2]), .C(clk16MHz), 
           .D(n26175));   // verilog/coms.v(128[12] 296[6])
    SB_DFFE data_in_frame_0___i131 (.Q(\data_in_frame[16] [2]), .C(clk16MHz), 
            .E(VCC_net), .D(n26510));   // verilog/coms.v(128[12] 296[6])
    SB_LUT4 i12676_3_lut_4_lut (.I0(Kp_23__N_1583), .I1(n29100), .I2(\data_in_frame[11] [5]), 
            .I3(IntegralLimit[21]), .O(n26280));
    defparam i12676_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i12677_3_lut_4_lut (.I0(Kp_23__N_1583), .I1(n29100), .I2(\data_in_frame[11] [4]), 
            .I3(IntegralLimit[20]), .O(n26281));
    defparam i12677_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i14_2_lut (.I0(rx_data_ready), .I1(\FRAME_MATCHER.rx_data_ready_prev ), 
            .I2(GND_net), .I3(GND_net), .O(n161));   // verilog/coms.v(153[9:50])
    defparam i14_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i12678_3_lut_4_lut (.I0(Kp_23__N_1583), .I1(n29100), .I2(\data_in_frame[11] [3]), 
            .I3(IntegralLimit[19]), .O(n26282));
    defparam i12678_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i12682_3_lut_4_lut (.I0(Kp_23__N_1583), .I1(n29100), .I2(\data_in_frame[11] [2]), 
            .I3(IntegralLimit[18]), .O(n26286));
    defparam i12682_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i12683_3_lut_4_lut (.I0(Kp_23__N_1583), .I1(n29100), .I2(\data_in_frame[14] [7]), 
            .I3(deadband[23]), .O(n26287));
    defparam i12683_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFFE data_in_frame_0___i130 (.Q(\data_in_frame[16] [1]), .C(clk16MHz), 
            .E(VCC_net), .D(n26507));   // verilog/coms.v(128[12] 296[6])
    SB_LUT4 i12696_3_lut_4_lut (.I0(Kp_23__N_1583), .I1(n29100), .I2(\data_in_frame[14] [6]), 
            .I3(deadband[22]), .O(n26300));
    defparam i12696_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i12697_3_lut_4_lut (.I0(Kp_23__N_1583), .I1(n29100), .I2(\data_in_frame[14] [5]), 
            .I3(deadband[21]), .O(n26301));
    defparam i12697_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i12698_3_lut_4_lut (.I0(Kp_23__N_1583), .I1(n29100), .I2(\data_in_frame[14] [4]), 
            .I3(deadband[20]), .O(n26302));
    defparam i12698_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i12699_3_lut_4_lut (.I0(Kp_23__N_1583), .I1(n29100), .I2(\data_in_frame[14] [3]), 
            .I3(deadband[19]), .O(n26303));
    defparam i12699_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 mux_1003_i2_3_lut_4_lut (.I0(Kp_23__N_1583), .I1(n29100), .I2(\data_in_frame[3][1] ), 
            .I3(\data_in_frame[19] [1]), .O(n4553[1]));
    defparam mux_1003_i2_3_lut_4_lut.LUT_INIT = 16'hf870;
    SB_DFFE data_in_frame_0___i129 (.Q(\data_in_frame[16] [0]), .C(clk16MHz), 
            .E(VCC_net), .D(n26504));   // verilog/coms.v(128[12] 296[6])
    SB_DFFE data_in_frame_0___i128 (.Q(\data_in_frame[15] [7]), .C(clk16MHz), 
            .E(VCC_net), .D(n26501));   // verilog/coms.v(128[12] 296[6])
    SB_DFFE data_in_frame_0___i127 (.Q(\data_in_frame[15] [6]), .C(clk16MHz), 
            .E(VCC_net), .D(n26498));   // verilog/coms.v(128[12] 296[6])
    SB_DFFE data_in_frame_0___i126 (.Q(\data_in_frame[15] [5]), .C(clk16MHz), 
            .E(VCC_net), .D(n26495));   // verilog/coms.v(128[12] 296[6])
    SB_DFFE data_in_frame_0___i125 (.Q(\data_in_frame[15] [4]), .C(clk16MHz), 
            .E(VCC_net), .D(n26492));   // verilog/coms.v(128[12] 296[6])
    SB_DFFE data_in_frame_0___i124 (.Q(\data_in_frame[15] [3]), .C(clk16MHz), 
            .E(VCC_net), .D(n26489));   // verilog/coms.v(128[12] 296[6])
    SB_DFFE data_in_frame_0___i123 (.Q(\data_in_frame[15] [2]), .C(clk16MHz), 
            .E(VCC_net), .D(n26486));   // verilog/coms.v(128[12] 296[6])
    SB_DFFE data_in_frame_0___i122 (.Q(\data_in_frame[15] [1]), .C(clk16MHz), 
            .E(VCC_net), .D(n26483));   // verilog/coms.v(128[12] 296[6])
    SB_LUT4 mux_1003_i3_3_lut_4_lut (.I0(Kp_23__N_1583), .I1(n29100), .I2(\data_in_frame[3][2] ), 
            .I3(\data_in_frame[19] [2]), .O(n4553[2]));
    defparam mux_1003_i3_3_lut_4_lut.LUT_INIT = 16'hf870;
    SB_LUT4 mux_1003_i4_3_lut_4_lut (.I0(Kp_23__N_1583), .I1(n29100), .I2(\data_in_frame[3][3] ), 
            .I3(\data_in_frame[19] [3]), .O(n4553[3]));
    defparam mux_1003_i4_3_lut_4_lut.LUT_INIT = 16'hf870;
    SB_LUT4 i17223_3_lut_4_lut (.I0(Kp_23__N_1583), .I1(n29100), .I2(\data_in_frame[3] [4]), 
            .I3(\data_in_frame[19] [4]), .O(n4553[4]));
    defparam i17223_3_lut_4_lut.LUT_INIT = 16'hf870;
    SB_DFFE data_in_frame_0___i121 (.Q(\data_in_frame[15] [0]), .C(clk16MHz), 
            .E(VCC_net), .D(n26480));   // verilog/coms.v(128[12] 296[6])
    SB_LUT4 mux_1003_i6_3_lut_4_lut (.I0(Kp_23__N_1583), .I1(n29100), .I2(\data_in_frame[3] [5]), 
            .I3(\data_in_frame[19] [5]), .O(n4553[5]));
    defparam mux_1003_i6_3_lut_4_lut.LUT_INIT = 16'hf870;
    SB_LUT4 mux_1003_i7_3_lut_4_lut (.I0(Kp_23__N_1583), .I1(n29100), .I2(\data_in_frame[3][6] ), 
            .I3(\data_in_frame[19] [6]), .O(n4553[6]));
    defparam mux_1003_i7_3_lut_4_lut.LUT_INIT = 16'hf870;
    SB_LUT4 mux_1003_i8_3_lut_4_lut (.I0(Kp_23__N_1583), .I1(n29100), .I2(\data_in_frame[3][7] ), 
            .I3(\data_in_frame[19] [7]), .O(n4553[7]));
    defparam mux_1003_i8_3_lut_4_lut.LUT_INIT = 16'hf870;
    SB_LUT4 mux_1003_i9_3_lut_4_lut (.I0(Kp_23__N_1583), .I1(n29100), .I2(\data_in_frame[2] [0]), 
            .I3(\data_in_frame[18] [0]), .O(n4553[8]));
    defparam mux_1003_i9_3_lut_4_lut.LUT_INIT = 16'hf870;
    SB_LUT4 i17864_3_lut_4_lut (.I0(Kp_23__N_1583), .I1(n29100), .I2(\data_in_frame[2] [1]), 
            .I3(\data_in_frame[18] [1]), .O(n4553[9]));
    defparam i17864_3_lut_4_lut.LUT_INIT = 16'hf870;
    SB_LUT4 mux_1003_i11_3_lut_4_lut (.I0(Kp_23__N_1583), .I1(n29100), .I2(\data_in_frame[2] [2]), 
            .I3(\data_in_frame[18] [2]), .O(n4553[10]));
    defparam mux_1003_i11_3_lut_4_lut.LUT_INIT = 16'hf870;
    SB_LUT4 i1_2_lut_3_lut (.I0(\FRAME_MATCHER.i_31__N_2325 ), .I1(\FRAME_MATCHER.i_31__N_2323 ), 
            .I2(\FRAME_MATCHER.i_31__N_2319 ), .I3(GND_net), .O(n3133));   // verilog/coms.v(146[4] 295[11])
    defparam i1_2_lut_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i17298_3_lut_4_lut (.I0(Kp_23__N_1583), .I1(n29100), .I2(\data_in_frame[2] [3]), 
            .I3(\data_in_frame[18] [3]), .O(n4553[11]));
    defparam i17298_3_lut_4_lut.LUT_INIT = 16'hf870;
    SB_LUT4 i11_3_lut (.I0(rx_data[5]), .I1(\data_in_frame[3] [5]), .I2(n25157), 
            .I3(GND_net), .O(n52227));   // verilog/coms.v(92[13:20])
    defparam i11_3_lut.LUT_INIT = 16'hcaca;
    SB_DFFE data_in_frame_0___i120 (.Q(\data_in_frame[14] [7]), .C(clk16MHz), 
            .E(VCC_net), .D(n26477));   // verilog/coms.v(128[12] 296[6])
    SB_LUT4 i12652_3_lut (.I0(\data_in_frame[3] [4]), .I1(rx_data[4]), .I2(n25157), 
            .I3(GND_net), .O(n26256));   // verilog/coms.v(128[12] 296[6])
    defparam i12652_3_lut.LUT_INIT = 16'hacac;
    SB_DFFESS data_out_frame_0___i3 (.Q(\data_out_frame[0][2] ), .C(clk16MHz), 
            .E(n2568), .D(n2), .S(n52768));   // verilog/coms.v(128[12] 296[6])
    SB_LUT4 mux_1003_i13_3_lut_4_lut (.I0(Kp_23__N_1583), .I1(n29100), .I2(\data_in_frame[2] [4]), 
            .I3(\data_in_frame[18] [4]), .O(n4553[12]));
    defparam mux_1003_i13_3_lut_4_lut.LUT_INIT = 16'hf870;
    SB_DFFESS data_out_frame_0___i4 (.Q(\data_out_frame[0][3] ), .C(clk16MHz), 
            .E(n2568), .D(n2_adj_5052), .S(n52818));   // verilog/coms.v(128[12] 296[6])
    SB_LUT4 mux_1003_i14_3_lut_4_lut (.I0(Kp_23__N_1583), .I1(n29100), .I2(\data_in_frame[2] [5]), 
            .I3(\data_in_frame[18] [5]), .O(n4553[13]));
    defparam mux_1003_i14_3_lut_4_lut.LUT_INIT = 16'hf870;
    SB_LUT4 i17260_3_lut_4_lut (.I0(Kp_23__N_1583), .I1(n29100), .I2(\data_in_frame[2] [6]), 
            .I3(\data_in_frame[18]_c [6]), .O(n4553[14]));
    defparam i17260_3_lut_4_lut.LUT_INIT = 16'hf870;
    SB_DFFESS data_out_frame_0___i5 (.Q(\data_out_frame[0][4] ), .C(clk16MHz), 
            .E(n2568), .D(n2_adj_5053), .S(n52817));   // verilog/coms.v(128[12] 296[6])
    SB_DFFESS data_out_frame_0___i9 (.Q(\data_out_frame[1][0] ), .C(clk16MHz), 
            .E(n2568), .D(n2_adj_5054), .S(n52816));   // verilog/coms.v(128[12] 296[6])
    SB_DFFESS data_out_frame_0___i10 (.Q(\data_out_frame[1][1] ), .C(clk16MHz), 
            .E(n2568), .D(n2_adj_5055), .S(n52815));   // verilog/coms.v(128[12] 296[6])
    SB_DFFE data_in_frame_0___i119 (.Q(\data_in_frame[14] [6]), .C(clk16MHz), 
            .E(VCC_net), .D(n26474));   // verilog/coms.v(128[12] 296[6])
    SB_DFFESS data_out_frame_0___i12 (.Q(\data_out_frame[1][3] ), .C(clk16MHz), 
            .E(n2568), .D(n2_adj_5056), .S(n52814));   // verilog/coms.v(128[12] 296[6])
    SB_LUT4 select_715_Select_210_i3_4_lut (.I0(n5), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(n55477), .I3(n53279), .O(n3));   // verilog/coms.v(146[4] 295[11])
    defparam select_715_Select_210_i3_4_lut.LUT_INIT = 16'h4884;
    SB_DFFESS data_out_frame_0___i14 (.Q(\data_out_frame[1][5] ), .C(clk16MHz), 
            .E(n2568), .D(n2_adj_5057), .S(n52819));   // verilog/coms.v(128[12] 296[6])
    SB_DFFESS data_out_frame_0___i15 (.Q(\data_out_frame[1][6] ), .C(clk16MHz), 
            .E(n2568), .D(n2_adj_5058), .S(n52813));   // verilog/coms.v(128[12] 296[6])
    SB_LUT4 mux_1003_i16_3_lut_4_lut (.I0(Kp_23__N_1583), .I1(n29100), .I2(\data_in_frame[2] [7]), 
            .I3(\data_in_frame[18][7] ), .O(n4553[15]));
    defparam mux_1003_i16_3_lut_4_lut.LUT_INIT = 16'hf870;
    SB_LUT4 i17424_3_lut_4_lut (.I0(Kp_23__N_1583), .I1(n29100), .I2(\data_in_frame[1] [0]), 
            .I3(\data_in_frame[17] [0]), .O(n4553[16]));
    defparam i17424_3_lut_4_lut.LUT_INIT = 16'hf870;
    SB_LUT4 i17378_3_lut_4_lut (.I0(Kp_23__N_1583), .I1(n29100), .I2(\data_in_frame[1] [1]), 
            .I3(\data_in_frame[17] [1]), .O(n4553[17]));
    defparam i17378_3_lut_4_lut.LUT_INIT = 16'hf870;
    SB_DFFESS data_out_frame_0___i16 (.Q(\data_out_frame[1][7] ), .C(clk16MHz), 
            .E(n2568), .D(n2_adj_5059), .S(n52812));   // verilog/coms.v(128[12] 296[6])
    SB_LUT4 select_715_Select_48_i2_4_lut (.I0(\data_out_frame[6] [0]), .I1(\FRAME_MATCHER.i_31__N_2320 ), 
            .I2(encoder0_position[16]), .I3(\FRAME_MATCHER.state_31__N_2423 [3]), 
            .O(n2_adj_5060));   // verilog/coms.v(146[4] 295[11])
    defparam select_715_Select_48_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut (.I0(\data_out_frame[21] [6]), .I1(n53314), .I2(GND_net), 
            .I3(GND_net), .O(n53506));
    defparam i1_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut (.I0(n23000), .I1(n48879), .I2(n23613), .I3(n2142), 
            .O(n53339));
    defparam i3_4_lut.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_adj_1044 (.I0(\data_out_frame[15] [4]), .I1(\data_out_frame[15] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n22958));
    defparam i1_2_lut_adj_1044.LUT_INIT = 16'h6666;
    SB_DFFR \FRAME_MATCHER.state_FSM_i1  (.Q(Kp_23__N_1583), .C(clk16MHz), 
            .D(n1816), .R(reset));   // verilog/coms.v(146[4] 295[11])
    SB_LUT4 i1_2_lut_adj_1045 (.I0(\data_out_frame[15] [5]), .I1(\data_out_frame[15] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n53305));
    defparam i1_2_lut_adj_1045.LUT_INIT = 16'h6666;
    SB_LUT4 i2_2_lut (.I0(\data_out_frame[17] [7]), .I1(n23361), .I2(GND_net), 
            .I3(GND_net), .O(n52927));
    defparam i2_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mux_1003_i19_3_lut_4_lut (.I0(Kp_23__N_1583), .I1(n29100), .I2(\data_in_frame[1][2] ), 
            .I3(\data_in_frame[17] [2]), .O(n4553[18]));
    defparam mux_1003_i19_3_lut_4_lut.LUT_INIT = 16'hf870;
    SB_LUT4 i3_4_lut_adj_1046 (.I0(\data_out_frame[17] [5]), .I1(n53305), 
            .I2(n53082), .I3(n52927), .O(n2142));
    defparam i3_4_lut_adj_1046.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut (.I0(n2142), .I1(\data_out_frame[22] [3]), .I2(\data_out_frame[22] [4]), 
            .I3(GND_net), .O(n52931));
    defparam i2_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 mux_1003_i20_3_lut_4_lut (.I0(Kp_23__N_1583), .I1(n29100), .I2(\data_in_frame[1][3] ), 
            .I3(\data_in_frame[17] [3]), .O(n4553[19]));
    defparam mux_1003_i20_3_lut_4_lut.LUT_INIT = 16'hf870;
    SB_DFFER setpoint_i0_i0 (.Q(setpoint[0]), .C(clk16MHz), .E(n24563), 
            .D(n4553[0]), .R(reset));   // verilog/coms.v(128[12] 296[6])
    SB_LUT4 i4_4_lut (.I0(n53453), .I1(n52998), .I2(\data_out_frame[13] [3]), 
            .I3(n53568), .O(n10));
    defparam i4_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 mux_1003_i21_3_lut_4_lut (.I0(Kp_23__N_1583), .I1(n29100), .I2(\data_in_frame[1][4] ), 
            .I3(\data_in_frame[17] [4]), .O(n4553[20]));
    defparam mux_1003_i21_3_lut_4_lut.LUT_INIT = 16'hf870;
    SB_LUT4 i5_3_lut (.I0(n53131), .I1(n10), .I2(\data_out_frame[11] [1]), 
            .I3(GND_net), .O(n23110));
    defparam i5_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_adj_1047 (.I0(n23110), .I1(n22564), .I2(n47823), 
            .I3(GND_net), .O(n53360));
    defparam i2_3_lut_adj_1047.LUT_INIT = 16'h9696;
    SB_LUT4 i3_4_lut_adj_1048 (.I0(n53225), .I1(n23256), .I2(\data_out_frame[13] [7]), 
            .I3(\data_out_frame[13] [6]), .O(n53012));   // verilog/coms.v(72[16:27])
    defparam i3_4_lut_adj_1048.LUT_INIT = 16'h6996;
    SB_DFFE data_in_frame_0___i118 (.Q(\data_in_frame[14] [5]), .C(clk16MHz), 
            .E(VCC_net), .D(n26471));   // verilog/coms.v(128[12] 296[6])
    SB_LUT4 i1_4_lut (.I0(n1129), .I1(\data_out_frame[6] [6]), .I2(n53153), 
            .I3(\data_out_frame[11] [4]), .O(n6));
    defparam i1_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_1049 (.I0(\data_out_frame[9] [2]), .I1(n53131), 
            .I2(n23417), .I3(n6), .O(n23256));
    defparam i4_4_lut_adj_1049.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1050 (.I0(n23256), .I1(n47860), .I2(\data_out_frame[13] [6]), 
            .I3(GND_net), .O(n48851));
    defparam i2_3_lut_adj_1050.LUT_INIT = 16'h9696;
    SB_LUT4 i3_3_lut (.I0(n23629), .I1(n52998), .I2(n53462), .I3(GND_net), 
            .O(n8_adj_5061));
    defparam i3_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 i1_4_lut_adj_1051 (.I0(\data_out_frame[13] [5]), .I1(\data_out_frame[11] [4]), 
            .I2(n8_adj_5061), .I3(n53459), .O(n23361));
    defparam i1_4_lut_adj_1051.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1052 (.I0(\data_out_frame[16] [1]), .I1(\data_out_frame[16] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n53524));
    defparam i1_2_lut_adj_1052.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_1053 (.I0(n33_c), .I1(n53524), .I2(n53357), .I3(n23361), 
            .O(n48777));
    defparam i3_4_lut_adj_1053.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1054 (.I0(\data_out_frame[16] [3]), .I1(n47766), 
            .I2(n53012), .I3(\data_out_frame[16] [2]), .O(n47853));
    defparam i3_4_lut_adj_1054.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1055 (.I0(n47853), .I1(n48777), .I2(GND_net), 
            .I3(GND_net), .O(n48879));
    defparam i1_2_lut_adj_1055.LUT_INIT = 16'h6666;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_48738 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[14] [2]), .I2(\data_out_frame[15] [2]), 
            .I3(byte_transmit_counter_c[1]), .O(n63473));
    defparam byte_transmit_counter_0__bdd_4_lut_48738.LUT_INIT = 16'he4aa;
    SB_LUT4 i4_4_lut_adj_1056 (.I0(n48777), .I1(n53020), .I2(n47823), 
            .I3(\data_out_frame[16] [0]), .O(n10_adj_5062));
    defparam i4_4_lut_adj_1056.LUT_INIT = 16'h9669;
    SB_LUT4 i5_3_lut_adj_1057 (.I0(n23361), .I1(n10_adj_5062), .I2(n48851), 
            .I3(GND_net), .O(n54765));
    defparam i5_3_lut_adj_1057.LUT_INIT = 16'h6969;
    SB_LUT4 i2_3_lut_adj_1058 (.I0(\data_out_frame[4] [6]), .I1(n52912), 
            .I2(\data_out_frame[7] [0]), .I3(GND_net), .O(n23417));   // verilog/coms.v(72[16:62])
    defparam i2_3_lut_adj_1058.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1059 (.I0(\data_out_frame[8] [7]), .I1(n23417), 
            .I2(GND_net), .I3(GND_net), .O(n53160));
    defparam i1_2_lut_adj_1059.LUT_INIT = 16'h6666;
    SB_LUT4 i5_4_lut (.I0(n53160), .I1(n53462), .I2(\data_out_frame[13] [4]), 
            .I3(\data_out_frame[11] [2]), .O(n12));
    defparam i5_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut (.I0(\data_out_frame[7] [1]), .I1(n12), .I2(n53544), 
            .I3(n23635), .O(n47823));
    defparam i6_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 n63473_bdd_4_lut (.I0(n63473), .I1(\data_out_frame[13] [2]), 
            .I2(\data_out_frame[12] [2]), .I3(byte_transmit_counter_c[1]), 
            .O(n56886));
    defparam n63473_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_2_lut_adj_1060 (.I0(\data_out_frame[15] [5]), .I1(n47823), 
            .I2(GND_net), .I3(GND_net), .O(n53189));
    defparam i1_2_lut_adj_1060.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1061 (.I0(\data_out_frame[17] [6]), .I1(\data_out_frame[17] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n53237));
    defparam i1_2_lut_adj_1061.LUT_INIT = 16'h6666;
    SB_LUT4 mux_1003_i22_3_lut_4_lut (.I0(Kp_23__N_1583), .I1(n29100), .I2(\data_in_frame[1][5] ), 
            .I3(\data_in_frame[17] [5]), .O(n4553[21]));
    defparam mux_1003_i22_3_lut_4_lut.LUT_INIT = 16'hf870;
    SB_LUT4 mux_1003_i23_3_lut_4_lut (.I0(Kp_23__N_1583), .I1(n29100), .I2(\data_in_frame[1][6] ), 
            .I3(\data_in_frame[17] [6]), .O(n4553[22]));
    defparam mux_1003_i23_3_lut_4_lut.LUT_INIT = 16'hf870;
    SB_LUT4 i4_4_lut_adj_1062 (.I0(\data_out_frame[22] [2]), .I1(\data_out_frame[15] [4]), 
            .I2(n53189), .I3(n6_adj_5063), .O(n48773));
    defparam i4_4_lut_adj_1062.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1063 (.I0(\data_out_frame[22] [1]), .I1(n47853), 
            .I2(n47956), .I3(GND_net), .O(n23613));
    defparam i2_3_lut_adj_1063.LUT_INIT = 16'h9696;
    SB_DFFE data_in_frame_0___i117 (.Q(\data_in_frame[14] [4]), .C(clk16MHz), 
            .E(VCC_net), .D(n26468));   // verilog/coms.v(128[12] 296[6])
    SB_LUT4 i12700_3_lut_4_lut (.I0(Kp_23__N_1583), .I1(n29100), .I2(\data_in_frame[14] [2]), 
            .I3(deadband[18]), .O(n26304));
    defparam i12700_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i13027_3_lut_4_lut (.I0(n25077), .I1(reset), .I2(rx_data[7]), 
            .I3(\data_in_frame[17] [7]), .O(n26631));
    defparam i13027_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFFESS data_out_frame_0___i26 (.Q(\data_out_frame[3][1] ), .C(clk16MHz), 
            .E(n2568), .D(n2_adj_5064), .S(n52811));   // verilog/coms.v(128[12] 296[6])
    SB_DFFE data_in_frame_0___i116 (.Q(\data_in_frame[14] [3]), .C(clk16MHz), 
            .E(VCC_net), .D(n26465));   // verilog/coms.v(128[12] 296[6])
    SB_DFFE data_in_frame_0___i115 (.Q(\data_in_frame[14] [2]), .C(clk16MHz), 
            .E(VCC_net), .D(n26462));   // verilog/coms.v(128[12] 296[6])
    SB_LUT4 i2_2_lut_adj_1064 (.I0(\data_out_frame[16] [0]), .I1(\data_out_frame[17] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n10_adj_5065));
    defparam i2_2_lut_adj_1064.LUT_INIT = 16'h6666;
    SB_LUT4 i6_4_lut_adj_1065 (.I0(n53360), .I1(\data_out_frame[15] [4]), 
            .I2(n53189), .I3(\data_out_frame[15] [6]), .O(n14));
    defparam i6_4_lut_adj_1065.LUT_INIT = 16'h6996;
    SB_LUT4 i12701_3_lut_4_lut (.I0(Kp_23__N_1583), .I1(n29100), .I2(\data_in_frame[14] [1]), 
            .I3(deadband[17]), .O(n26305));
    defparam i12701_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i7_4_lut (.I0(n23110), .I1(n14), .I2(n10_adj_5065), .I3(n53357), 
            .O(n48858));
    defparam i7_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1066 (.I0(\data_out_frame[9] [2]), .I1(\data_out_frame[9] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n53544));
    defparam i1_2_lut_adj_1066.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1067 (.I0(n23629), .I1(\data_out_frame[7] [5]), 
            .I2(n53324), .I3(n6_adj_5066), .O(n54577));
    defparam i4_4_lut_adj_1067.LUT_INIT = 16'h6996;
    SB_LUT4 i2_4_lut (.I0(\data_out_frame[7] [4]), .I1(\data_out_frame[7] [1]), 
            .I2(n54577), .I3(\data_out_frame[5] [3]), .O(n16));
    defparam i2_4_lut.LUT_INIT = 16'h9669;
    SB_DFFESS data_out_frame_0___i28 (.Q(\data_out_frame[3][3] ), .C(clk16MHz), 
            .E(n2568), .D(n2_adj_5067), .S(n52810));   // verilog/coms.v(128[12] 296[6])
    SB_DFFESS data_out_frame_0___i29 (.Q(\data_out_frame[3][4] ), .C(clk16MHz), 
            .E(n2568), .D(n2_adj_5068), .S(n52809));   // verilog/coms.v(128[12] 296[6])
    SB_LUT4 i1_2_lut_adj_1068 (.I0(n53397), .I1(\data_out_frame[4] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n15_c));
    defparam i1_2_lut_adj_1068.LUT_INIT = 16'h6666;
    SB_LUT4 i10_4_lut (.I0(n53204), .I1(\data_out_frame[6] [7]), .I2(n53026), 
            .I3(\data_out_frame[7] [0]), .O(n24));
    defparam i10_4_lut.LUT_INIT = 16'h6996;
    SB_DFFESS data_out_frame_0___i31 (.Q(\data_out_frame[3][6] ), .C(clk16MHz), 
            .E(n2568), .D(n2_adj_5069), .S(n52808));   // verilog/coms.v(128[12] 296[6])
    SB_DFFESS data_out_frame_0___i32 (.Q(\data_out_frame[3][7] ), .C(clk16MHz), 
            .E(n2568), .D(n2_adj_5070), .S(n52807));   // verilog/coms.v(128[12] 296[6])
    SB_DFFE data_in_frame_0___i114 (.Q(\data_in_frame[14] [1]), .C(clk16MHz), 
            .E(VCC_net), .D(n26459));   // verilog/coms.v(128[12] 296[6])
    SB_LUT4 i9_4_lut (.I0(n53100), .I1(n23083), .I2(\data_out_frame[6] [4]), 
            .I3(n53535), .O(n23_c));
    defparam i9_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i11_4_lut (.I0(n22526), .I1(n15_c), .I2(\data_out_frame[8] [0]), 
            .I3(n16), .O(n25));
    defparam i11_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_1069 (.I0(n52992), .I1(n25), .I2(n23_c), .I3(n24), 
            .O(n13));
    defparam i4_4_lut_adj_1069.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut_adj_1070 (.I0(n13), .I1(\data_out_frame[9] [1]), .I2(\data_out_frame[9] [3]), 
            .I3(n53037), .O(n16_adj_5071));
    defparam i7_4_lut_adj_1070.LUT_INIT = 16'h6996;
    SB_LUT4 i12702_3_lut_4_lut (.I0(Kp_23__N_1583), .I1(n29100), .I2(\data_in_frame[14] [0]), 
            .I3(deadband[16]), .O(n26306));
    defparam i12702_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i8_4_lut (.I0(n53544), .I1(n16_adj_5071), .I2(n12_adj_5072), 
            .I3(\data_out_frame[5] [4]), .O(n55050));
    defparam i8_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i12703_3_lut_4_lut (.I0(Kp_23__N_1583), .I1(n29100), .I2(\data_in_frame[15] [7]), 
            .I3(deadband[15]), .O(n26307));
    defparam i12703_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i10_4_lut_adj_1071 (.I0(n53412), .I1(\data_out_frame[10] [1]), 
            .I2(\data_out_frame[11] [3]), .I3(\data_out_frame[11] [6]), 
            .O(n24_adj_5073));   // verilog/coms.v(86[17:63])
    defparam i10_4_lut_adj_1071.LUT_INIT = 16'h6996;
    SB_LUT4 i8_4_lut_adj_1072 (.I0(n1667), .I1(n55050), .I2(n53256), .I3(\data_out_frame[11] [5]), 
            .O(n22));   // verilog/coms.v(86[17:63])
    defparam i8_4_lut_adj_1072.LUT_INIT = 16'h6996;
    SB_LUT4 i12_4_lut (.I0(n53453), .I1(n24_adj_5073), .I2(n18), .I3(\data_out_frame[10] [7]), 
            .O(n26));   // verilog/coms.v(86[17:63])
    defparam i12_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i13_4_lut (.I0(\data_out_frame[11] [4]), .I1(n26), .I2(n22), 
            .I3(n53103), .O(n53273));   // verilog/coms.v(86[17:63])
    defparam i13_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i13409_3_lut_4_lut (.I0(n8_adj_5074), .I1(n52882), .I2(rx_data[7]), 
            .I3(\data_in_frame[9] [7]), .O(n27013));
    defparam i13409_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13406_3_lut_4_lut (.I0(n8_adj_5074), .I1(n52882), .I2(rx_data[6]), 
            .I3(\data_in_frame[9] [6]), .O(n27010));
    defparam i13406_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i3_4_lut_adj_1073 (.I0(\data_out_frame[8] [2]), .I1(n53388), 
            .I2(\data_out_frame[7] [7]), .I3(\data_out_frame[10] [2]), .O(n53308));
    defparam i3_4_lut_adj_1073.LUT_INIT = 16'h6996;
    SB_DFFESS data_out_frame_0___i84 (.Q(\data_out_frame[10] [3]), .C(clk16MHz), 
            .E(n2568), .D(n2_adj_5075), .S(n52713));   // verilog/coms.v(128[12] 296[6])
    SB_LUT4 i5_3_lut_adj_1074 (.I0(\data_out_frame[12] [0]), .I1(n47860), 
            .I2(n53308), .I3(GND_net), .O(n14_adj_5076));
    defparam i5_3_lut_adj_1074.LUT_INIT = 16'h9696;
    SB_LUT4 i6_4_lut_adj_1075 (.I0(n53518), .I1(\data_out_frame[13] [7]), 
            .I2(n22526), .I3(n53332), .O(n15_adj_5077));
    defparam i6_4_lut_adj_1075.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1076 (.I0(\data_out_frame[14] [1]), .I1(n22529), 
            .I2(n6_adj_5078), .I3(n53150), .O(n6_adj_5079));   // verilog/coms.v(86[17:70])
    defparam i1_4_lut_adj_1076.LUT_INIT = 16'h6996;
    SB_LUT4 i48308_4_lut (.I0(n15_adj_5077), .I1(\data_out_frame[5] [3]), 
            .I2(n14_adj_5076), .I3(GND_net), .O(n63021));
    defparam i48308_4_lut.LUT_INIT = 16'h6969;
    SB_LUT4 i4_4_lut_adj_1077 (.I0(n21977), .I1(n63021), .I2(\data_out_frame[10] [4]), 
            .I3(n6_adj_5079), .O(n33_c));   // verilog/coms.v(86[17:70])
    defparam i4_4_lut_adj_1077.LUT_INIT = 16'h9669;
    SB_LUT4 i13403_3_lut_4_lut (.I0(n8_adj_5074), .I1(n52882), .I2(rx_data[5]), 
            .I3(\data_in_frame[9] [5]), .O(n27007));
    defparam i13403_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_1078 (.I0(\data_out_frame[9] [3]), .I1(n23720), 
            .I2(GND_net), .I3(GND_net), .O(n53153));
    defparam i1_2_lut_adj_1078.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_1079 (.I0(\data_out_frame[5] [4]), .I1(n53216), 
            .I2(\data_out_frame[5] [1]), .I3(\data_out_frame[5] [7]), .O(n23083));   // verilog/coms.v(74[16:34])
    defparam i3_4_lut_adj_1079.LUT_INIT = 16'h6996;
    SB_LUT4 i12704_3_lut_4_lut (.I0(Kp_23__N_1583), .I1(n29100), .I2(\data_in_frame[15] [6]), 
            .I3(deadband[14]), .O(n26308));
    defparam i12704_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i12705_3_lut_4_lut (.I0(Kp_23__N_1583), .I1(n29100), .I2(\data_in_frame[15] [5]), 
            .I3(deadband[13]), .O(n26309));
    defparam i12705_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i12706_3_lut_4_lut (.I0(Kp_23__N_1583), .I1(n29100), .I2(\data_in_frame[15] [4]), 
            .I3(deadband[12]), .O(n26310));
    defparam i12706_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i12707_3_lut_4_lut (.I0(Kp_23__N_1583), .I1(n29100), .I2(\data_in_frame[15] [3]), 
            .I3(deadband[11]), .O(n26311));
    defparam i12707_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2_3_lut_adj_1080 (.I0(n52912), .I1(\data_out_frame[6] [7]), 
            .I2(\data_out_frame[4] [5]), .I3(GND_net), .O(n53131));   // verilog/coms.v(72[16:62])
    defparam i2_3_lut_adj_1080.LUT_INIT = 16'h9696;
    SB_DFFESS data_out_frame_0___i85 (.Q(\data_out_frame[10] [4]), .C(clk16MHz), 
            .E(n2568), .D(n2_adj_5080), .S(n52714));   // verilog/coms.v(128[12] 296[6])
    SB_DFFESS data_out_frame_0___i86 (.Q(\data_out_frame[10] [5]), .C(clk16MHz), 
            .E(n2568), .D(n2_adj_5081), .S(n52715));   // verilog/coms.v(128[12] 296[6])
    SB_DFFESS data_out_frame_0___i87 (.Q(\data_out_frame[10] [6]), .C(clk16MHz), 
            .E(n2568), .D(n2_adj_5082), .S(n52789));   // verilog/coms.v(128[12] 296[6])
    SB_DFFESS data_out_frame_0___i88 (.Q(\data_out_frame[10] [7]), .C(clk16MHz), 
            .E(n2568), .D(n2_adj_5083), .S(n52716));   // verilog/coms.v(128[12] 296[6])
    SB_DFFESS data_out_frame_0___i89 (.Q(\data_out_frame[11] [0]), .C(clk16MHz), 
            .E(n2568), .D(n2_adj_5084), .S(n52717));   // verilog/coms.v(128[12] 296[6])
    SB_DFFESS data_out_frame_0___i90 (.Q(\data_out_frame[11] [1]), .C(clk16MHz), 
            .E(n2568), .D(n2_adj_5085), .S(n52718));   // verilog/coms.v(128[12] 296[6])
    SB_DFFESS data_out_frame_0___i91 (.Q(\data_out_frame[11] [2]), .C(clk16MHz), 
            .E(n2568), .D(n2_adj_5086), .S(n52719));   // verilog/coms.v(128[12] 296[6])
    SB_DFFESS data_out_frame_0___i92 (.Q(\data_out_frame[11] [3]), .C(clk16MHz), 
            .E(n2568), .D(n2_adj_5087), .S(n52720));   // verilog/coms.v(128[12] 296[6])
    SB_DFFESS data_out_frame_0___i93 (.Q(\data_out_frame[11] [4]), .C(clk16MHz), 
            .E(n2568), .D(n2_adj_5088), .S(n52721));   // verilog/coms.v(128[12] 296[6])
    SB_DFFESS data_out_frame_0___i94 (.Q(\data_out_frame[11] [5]), .C(clk16MHz), 
            .E(n2568), .D(n2_adj_5089), .S(n52722));   // verilog/coms.v(128[12] 296[6])
    SB_DFFESS data_out_frame_0___i95 (.Q(\data_out_frame[11] [6]), .C(clk16MHz), 
            .E(n2568), .D(n2_adj_5090), .S(n52723));   // verilog/coms.v(128[12] 296[6])
    SB_DFFESS data_out_frame_0___i96 (.Q(\data_out_frame[11] [7]), .C(clk16MHz), 
            .E(n2568), .D(n2_adj_5091), .S(n52724));   // verilog/coms.v(128[12] 296[6])
    SB_DFFESS data_out_frame_0___i33 (.Q(\data_out_frame[4] [0]), .C(clk16MHz), 
            .E(n2568), .D(n2_adj_5092), .S(n52806));   // verilog/coms.v(128[12] 296[6])
    SB_LUT4 i2_3_lut_adj_1081 (.I0(\data_out_frame[5] [2]), .I1(n53397), 
            .I2(\data_out_frame[9] [4]), .I3(GND_net), .O(n22950));   // verilog/coms.v(74[16:34])
    defparam i2_3_lut_adj_1081.LUT_INIT = 16'h9696;
    SB_LUT4 i3_4_lut_adj_1082 (.I0(\data_out_frame[11] [6]), .I1(n22950), 
            .I2(\data_out_frame[14] [0]), .I3(n22752), .O(n53225));
    defparam i3_4_lut_adj_1082.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1083 (.I0(\data_out_frame[11] [5]), .I1(n53459), 
            .I2(n6_adj_5093), .I3(n22950), .O(n47860));
    defparam i1_4_lut_adj_1083.LUT_INIT = 16'h6996;
    SB_LUT4 i13024_3_lut_4_lut (.I0(n25077), .I1(reset), .I2(rx_data[6]), 
            .I3(\data_in_frame[17] [6]), .O(n26628));
    defparam i13024_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_1084 (.I0(n47860), .I1(n53225), .I2(GND_net), 
            .I3(GND_net), .O(n53226));
    defparam i1_2_lut_adj_1084.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_1085 (.I0(\data_out_frame[15] [6]), .I1(n53226), 
            .I2(\data_out_frame[13] [7]), .I3(\data_out_frame[16] [1]), 
            .O(n53020));
    defparam i3_4_lut_adj_1085.LUT_INIT = 16'h9669;
    SB_LUT4 i12708_3_lut_4_lut (.I0(Kp_23__N_1583), .I1(n29100), .I2(\data_in_frame[15] [2]), 
            .I3(deadband[10]), .O(n26312));
    defparam i12708_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i341_2_lut (.I0(\data_out_frame[4] [5]), .I1(\data_out_frame[4] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n1129));   // verilog/coms.v(77[16:27])
    defparam i341_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1086 (.I0(\data_out_frame[11] [1]), .I1(\data_out_frame[11] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n53412));   // verilog/coms.v(75[16:43])
    defparam i1_2_lut_adj_1086.LUT_INIT = 16'h6666;
    SB_LUT4 i17986_3_lut_4_lut (.I0(Kp_23__N_1583), .I1(n29100), .I2(\data_in_frame[11] [1]), 
            .I3(IntegralLimit[17]), .O(n26313));
    defparam i17986_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i3_4_lut_adj_1087 (.I0(\data_out_frame[8] [7]), .I1(\data_out_frame[8] [6]), 
            .I2(\data_out_frame[6] [6]), .I3(\data_out_frame[8] [5]), .O(n53026));   // verilog/coms.v(75[16:43])
    defparam i3_4_lut_adj_1087.LUT_INIT = 16'h6996;
    SB_DFFESS data_out_frame_0___i97 (.Q(\data_out_frame[12] [0]), .C(clk16MHz), 
            .E(n2568), .D(n2_adj_5094), .S(n52725));   // verilog/coms.v(128[12] 296[6])
    SB_LUT4 i3_4_lut_adj_1088 (.I0(\data_out_frame[15] [2]), .I1(\data_out_frame[13] [0]), 
            .I2(\data_out_frame[15] [3]), .I3(n21993), .O(n53068));
    defparam i3_4_lut_adj_1088.LUT_INIT = 16'h6996;
    SB_LUT4 i2_2_lut_adj_1089 (.I0(n53026), .I1(\data_out_frame[10] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n10_adj_5095));   // verilog/coms.v(75[16:43])
    defparam i2_2_lut_adj_1089.LUT_INIT = 16'h6666;
    SB_LUT4 i12710_3_lut_4_lut (.I0(Kp_23__N_1583), .I1(n29100), .I2(\data_in_frame[11] [0]), 
            .I3(IntegralLimit[16]), .O(n26314));
    defparam i12710_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i6_4_lut_adj_1090 (.I0(n53412), .I1(\data_out_frame[13] [2]), 
            .I2(\data_out_frame[8] [4]), .I3(\data_out_frame[9] [0]), .O(n14_adj_5096));   // verilog/coms.v(75[16:43])
    defparam i6_4_lut_adj_1090.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut_adj_1091 (.I0(n22529), .I1(n14_adj_5096), .I2(n10_adj_5095), 
            .I3(n1129), .O(n22564));   // verilog/coms.v(75[16:43])
    defparam i7_4_lut_adj_1091.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1092 (.I0(\data_out_frame[17] [3]), .I1(n53088), 
            .I2(n48497), .I3(GND_net), .O(n48787));
    defparam i2_3_lut_adj_1092.LUT_INIT = 16'h9696;
    SB_DFFE data_in_frame_0___i113 (.Q(\data_in_frame[14] [0]), .C(clk16MHz), 
            .E(VCC_net), .D(n26456));   // verilog/coms.v(128[12] 296[6])
    SB_DFFESS data_out_frame_0___i98 (.Q(\data_out_frame[12] [1]), .C(clk16MHz), 
            .E(n2568), .D(n2_adj_5097), .S(n52726));   // verilog/coms.v(128[12] 296[6])
    SB_LUT4 i2_3_lut_adj_1093 (.I0(n47956), .I1(n48787), .I2(\data_out_frame[21] [7]), 
            .I3(GND_net), .O(n53219));
    defparam i2_3_lut_adj_1093.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1094 (.I0(\data_out_frame[15] [5]), .I1(n53020), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_5098));
    defparam i1_2_lut_adj_1094.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1095 (.I0(\data_out_frame[15] [7]), .I1(\data_out_frame[17] [7]), 
            .I2(n23110), .I3(n6_adj_5098), .O(n54590));
    defparam i4_4_lut_adj_1095.LUT_INIT = 16'h6996;
    SB_LUT4 i12711_3_lut_4_lut (.I0(Kp_23__N_1583), .I1(n29100), .I2(\data_in_frame[15] [1]), 
            .I3(deadband[9]), .O(n26315));
    defparam i12711_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4_4_lut_adj_1096 (.I0(n48858), .I1(n47777), .I2(n48885), 
            .I3(n6_adj_5099), .O(n55276));
    defparam i4_4_lut_adj_1096.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1097 (.I0(n48773), .I1(n48858), .I2(\data_out_frame[22] [3]), 
            .I3(GND_net), .O(n47815));
    defparam i2_3_lut_adj_1097.LUT_INIT = 16'h6969;
    SB_LUT4 i1_2_lut_adj_1098 (.I0(n48858), .I1(n54590), .I2(GND_net), 
            .I3(GND_net), .O(n23000));
    defparam i1_2_lut_adj_1098.LUT_INIT = 16'h9999;
    SB_DFFESS data_out_frame_0___i34 (.Q(\data_out_frame[4] [1]), .C(clk16MHz), 
            .E(n2568), .D(n2_adj_5100), .S(n52805));   // verilog/coms.v(128[12] 296[6])
    SB_DFFE data_in_frame_0___i112 (.Q(\data_in_frame[13] [7]), .C(clk16MHz), 
            .E(VCC_net), .D(n26453));   // verilog/coms.v(128[12] 296[6])
    SB_LUT4 i4_4_lut_adj_1099 (.I0(n54765), .I1(n47956), .I2(n53279), 
            .I3(n53339), .O(n54489));
    defparam i4_4_lut_adj_1099.LUT_INIT = 16'h9669;
    SB_DFFESS data_out_frame_0___i35 (.Q(\data_out_frame[4] [2]), .C(clk16MHz), 
            .E(n2568), .D(n2_adj_5101), .S(n52796));   // verilog/coms.v(128[12] 296[6])
    SB_DFFE data_in_frame_0___i111 (.Q(\data_in_frame[13] [6]), .C(clk16MHz), 
            .E(VCC_net), .D(n26450));   // verilog/coms.v(128[12] 296[6])
    SB_DFFE data_in_frame_0___i110 (.Q(\data_in_frame[13] [5]), .C(clk16MHz), 
            .E(VCC_net), .D(n26447));   // verilog/coms.v(128[12] 296[6])
    SB_LUT4 select_715_Select_209_i3_4_lut (.I0(n48809), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(n8_adj_5102), .I3(n52932), .O(n3_adj_5103));   // verilog/coms.v(146[4] 295[11])
    defparam select_715_Select_209_i3_4_lut.LUT_INIT = 16'h4884;
    SB_LUT4 i13021_3_lut_4_lut (.I0(n25077), .I1(reset), .I2(rx_data[5]), 
            .I3(\data_in_frame[17] [5]), .O(n26625));
    defparam i13021_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF data_in_frame_0___i108 (.Q(\data_in_frame[13] [3]), .C(clk16MHz), 
           .D(n26178));   // verilog/coms.v(128[12] 296[6])
    SB_DFF data_in_frame_0___i9 (.Q(\data_in_frame[1] [0]), .C(clk16MHz), 
           .D(n26444));   // verilog/coms.v(128[12] 296[6])
    SB_DFF data_in_frame_0___i10 (.Q(\data_in_frame[1] [1]), .C(clk16MHz), 
           .D(n52175));   // verilog/coms.v(128[12] 296[6])
    SB_DFF data_in_frame_0___i11 (.Q(\data_in_frame[1][2] ), .C(clk16MHz), 
           .D(n26190));   // verilog/coms.v(128[12] 296[6])
    SB_DFF data_in_frame_0___i12 (.Q(\data_in_frame[1][3] ), .C(clk16MHz), 
           .D(n26193));   // verilog/coms.v(128[12] 296[6])
    SB_DFF data_in_frame_0___i13 (.Q(\data_in_frame[1][4] ), .C(clk16MHz), 
           .D(n26196));   // verilog/coms.v(128[12] 296[6])
    SB_LUT4 i12715_3_lut_4_lut (.I0(Kp_23__N_1583), .I1(n29100), .I2(\data_in_frame[15] [0]), 
            .I3(deadband[8]), .O(n26319));
    defparam i12715_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFFESS data_out_frame_0___i36 (.Q(\data_out_frame[4] [3]), .C(clk16MHz), 
            .E(n2568), .D(n2_adj_5104), .S(n52797));   // verilog/coms.v(128[12] 296[6])
    SB_DFF data_in_frame_0___i14 (.Q(\data_in_frame[1][5] ), .C(clk16MHz), 
           .D(n26199));   // verilog/coms.v(128[12] 296[6])
    SB_DFFESS data_out_frame_0___i37 (.Q(\data_out_frame[4] [4]), .C(clk16MHz), 
            .E(n2568), .D(n2_adj_5105), .S(n52798));   // verilog/coms.v(128[12] 296[6])
    SB_DFF data_in_frame_0___i15 (.Q(\data_in_frame[1][6] ), .C(clk16MHz), 
           .D(n26202));   // verilog/coms.v(128[12] 296[6])
    SB_DFF data_in_frame_0___i16 (.Q(\data_in_frame[1][7] ), .C(clk16MHz), 
           .D(n26205));   // verilog/coms.v(128[12] 296[6])
    SB_DFFESS data_out_frame_0___i38 (.Q(\data_out_frame[4] [5]), .C(clk16MHz), 
            .E(n2568), .D(n2_adj_5106), .S(n52799));   // verilog/coms.v(128[12] 296[6])
    SB_DFFESS data_out_frame_0___i39 (.Q(\data_out_frame[4] [6]), .C(clk16MHz), 
            .E(n2568), .D(n2_adj_5107), .S(n52800));   // verilog/coms.v(128[12] 296[6])
    SB_DFFESS data_out_frame_0___i40 (.Q(\data_out_frame[4] [7]), .C(clk16MHz), 
            .E(n2568), .D(n2_adj_5108), .S(n52801));   // verilog/coms.v(128[12] 296[6])
    SB_DFF data_in_frame_0___i17 (.Q(\data_in_frame[2] [0]), .C(clk16MHz), 
           .D(n26208));   // verilog/coms.v(128[12] 296[6])
    SB_DFF data_in_frame_0___i18 (.Q(\data_in_frame[2] [1]), .C(clk16MHz), 
           .D(n26212));   // verilog/coms.v(128[12] 296[6])
    SB_DFF data_in_frame_0___i19 (.Q(\data_in_frame[2] [2]), .C(clk16MHz), 
           .D(n26215));   // verilog/coms.v(128[12] 296[6])
    SB_DFF data_in_frame_0___i20 (.Q(\data_in_frame[2] [3]), .C(clk16MHz), 
           .D(n52143));   // verilog/coms.v(128[12] 296[6])
    SB_DFF data_in_frame_0___i21 (.Q(\data_in_frame[2] [4]), .C(clk16MHz), 
           .D(n26221));   // verilog/coms.v(128[12] 296[6])
    SB_DFF data_in_frame_0___i22 (.Q(\data_in_frame[2] [5]), .C(clk16MHz), 
           .D(n26224));   // verilog/coms.v(128[12] 296[6])
    SB_DFF data_in_frame_0___i23 (.Q(\data_in_frame[2] [6]), .C(clk16MHz), 
           .D(n26227));   // verilog/coms.v(128[12] 296[6])
    SB_DFFESS data_out_frame_0___i41 (.Q(\data_out_frame[5] [0]), .C(clk16MHz), 
            .E(n2568), .D(n2_adj_5109), .S(n52802));   // verilog/coms.v(128[12] 296[6])
    SB_DFFESS data_out_frame_0___i42 (.Q(\data_out_frame[5] [1]), .C(clk16MHz), 
            .E(n2568), .D(n2_adj_5110), .S(n52803));   // verilog/coms.v(128[12] 296[6])
    SB_DFFESS data_out_frame_0___i43 (.Q(\data_out_frame[5] [2]), .C(clk16MHz), 
            .E(n2568), .D(n2_adj_5111), .S(n52804));   // verilog/coms.v(128[12] 296[6])
    SB_DFFESS data_out_frame_0___i44 (.Q(\data_out_frame[5] [3]), .C(clk16MHz), 
            .E(n2568), .D(n2_adj_5112), .S(n52682));   // verilog/coms.v(128[12] 296[6])
    SB_DFF data_in_frame_0___i24 (.Q(\data_in_frame[2] [7]), .C(clk16MHz), 
           .D(n26231));   // verilog/coms.v(128[12] 296[6])
    SB_DFF data_in_frame_0___i25 (.Q(\data_in_frame[3] [0]), .C(clk16MHz), 
           .D(n26413));   // verilog/coms.v(128[12] 296[6])
    SB_LUT4 i12716_3_lut_4_lut (.I0(Kp_23__N_1583), .I1(n29100), .I2(\data_in_frame[16] [7]), 
            .I3(deadband[7]), .O(n26320));
    defparam i12716_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i12717_3_lut_4_lut (.I0(Kp_23__N_1583), .I1(n29100), .I2(\data_in_frame[16] [6]), 
            .I3(deadband[6]), .O(n26321));
    defparam i12717_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i12718_3_lut_4_lut (.I0(Kp_23__N_1583), .I1(n29100), .I2(\data_in_frame[16] [5]), 
            .I3(deadband[5]), .O(n26322));
    defparam i12718_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i12719_3_lut_4_lut (.I0(Kp_23__N_1583), .I1(n29100), .I2(\data_in_frame[16] [4]), 
            .I3(deadband[4]), .O(n26323));
    defparam i12719_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i12720_3_lut_4_lut (.I0(Kp_23__N_1583), .I1(n29100), .I2(\data_in_frame[16] [3]), 
            .I3(deadband[3]), .O(n26324));
    defparam i12720_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i18451_3_lut_4_lut (.I0(Kp_23__N_1583), .I1(n29100), .I2(\data_in_frame[16] [2]), 
            .I3(deadband_c[2]), .O(n26325));
    defparam i18451_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i13018_3_lut_4_lut (.I0(n25077), .I1(reset), .I2(rx_data[4]), 
            .I3(\data_in_frame[17] [4]), .O(n26622));
    defparam i13018_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 select_715_Select_47_i2_4_lut (.I0(\data_out_frame[5] [7]), .I1(\FRAME_MATCHER.i_31__N_2320 ), 
            .I2(control_mode[7]), .I3(\FRAME_MATCHER.state_31__N_2423 [3]), 
            .O(n2_adj_5113));   // verilog/coms.v(146[4] 295[11])
    defparam select_715_Select_47_i2_4_lut.LUT_INIT = 16'hc088;
    SB_DFF data_in_frame_0___i26 (.Q(\data_in_frame[3][1] ), .C(clk16MHz), 
           .D(n26238));   // verilog/coms.v(128[12] 296[6])
    SB_LUT4 i17259_3_lut (.I0(n25157), .I1(rx_data[0]), .I2(\data_in_frame[3] [0]), 
            .I3(GND_net), .O(n26413));   // verilog/coms.v(92[13:20])
    defparam i17259_3_lut.LUT_INIT = 16'he4e4;
    SB_DFF data_in_frame_0___i27 (.Q(\data_in_frame[3][2] ), .C(clk16MHz), 
           .D(n26250));   // verilog/coms.v(128[12] 296[6])
    SB_DFF data_in_frame_0___i28 (.Q(\data_in_frame[3][3] ), .C(clk16MHz), 
           .D(n26253));   // verilog/coms.v(128[12] 296[6])
    SB_DFF data_in_frame_0___i29 (.Q(\data_in_frame[3] [4]), .C(clk16MHz), 
           .D(n26256));   // verilog/coms.v(128[12] 296[6])
    SB_DFF data_in_frame_0___i30 (.Q(\data_in_frame[3] [5]), .C(clk16MHz), 
           .D(n52227));   // verilog/coms.v(128[12] 296[6])
    SB_LUT4 i1_2_lut_adj_1100 (.I0(\data_out_frame[5] [5]), .I1(\data_out_frame[5] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n53023));   // verilog/coms.v(76[16:27])
    defparam i1_2_lut_adj_1100.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1101 (.I0(\data_out_frame[9] [4]), .I1(\data_out_frame[9] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n53415));   // verilog/coms.v(76[16:27])
    defparam i1_2_lut_adj_1101.LUT_INIT = 16'h6666;
    SB_DFF data_in_frame_0___i31 (.Q(\data_in_frame[3][6] ), .C(clk16MHz), 
           .D(n26262));   // verilog/coms.v(128[12] 296[6])
    SB_DFF data_in_frame_0___i32 (.Q(\data_in_frame[3][7] ), .C(clk16MHz), 
           .D(n26265));   // verilog/coms.v(128[12] 296[6])
    SB_DFF data_in_frame_0___i33 (.Q(\data_in_frame[4] [0]), .C(clk16MHz), 
           .D(n26268));   // verilog/coms.v(128[12] 296[6])
    SB_LUT4 i7_4_lut_adj_1102 (.I0(n23720), .I1(\data_out_frame[9] [6]), 
            .I2(\data_out_frame[7] [6]), .I3(\data_out_frame[12] [0]), .O(n18_adj_5114));   // verilog/coms.v(76[16:27])
    defparam i7_4_lut_adj_1102.LUT_INIT = 16'h6996;
    SB_LUT4 select_715_Select_43_i2_4_lut (.I0(\data_out_frame[5] [3]), .I1(\FRAME_MATCHER.i_31__N_2320 ), 
            .I2(control_mode_c[3]), .I3(\FRAME_MATCHER.state_31__N_2423 [3]), 
            .O(n2_adj_5112));   // verilog/coms.v(146[4] 295[11])
    defparam select_715_Select_43_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 add_1107_9_lut (.I0(n52664), .I1(byte_transmit_counter_c[7]), 
            .I2(GND_net), .I3(n46125), .O(n52665)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1107_9_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i5_2_lut (.I0(\data_out_frame[10] [0]), .I1(\data_out_frame[11] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n16_adj_5115));   // verilog/coms.v(76[16:27])
    defparam i5_2_lut.LUT_INIT = 16'h6666;
    SB_DFF data_in_frame_0___i34 (.Q(\data_in_frame[4] [1]), .C(clk16MHz), 
           .D(n26271));   // verilog/coms.v(128[12] 296[6])
    SB_DFF data_in_frame_0___i35 (.Q(\data_in_frame[4] [2]), .C(clk16MHz), 
           .D(n26274));   // verilog/coms.v(128[12] 296[6])
    SB_LUT4 i9_4_lut_adj_1103 (.I0(\data_out_frame[9] [5]), .I1(n18_adj_5114), 
            .I2(\data_out_frame[14] [2]), .I3(\data_out_frame[12] [1]), 
            .O(n20));   // verilog/coms.v(76[16:27])
    defparam i9_4_lut_adj_1103.LUT_INIT = 16'h6996;
    SB_LUT4 i10_4_lut_adj_1104 (.I0(n53415), .I1(n20), .I2(n16_adj_5115), 
            .I3(n53023), .O(n47766));   // verilog/coms.v(76[16:27])
    defparam i10_4_lut_adj_1104.LUT_INIT = 16'h6996;
    SB_LUT4 add_1107_8_lut (.I0(n52664), .I1(byte_transmit_counter_c[6]), 
            .I2(GND_net), .I3(n46124), .O(n52667)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1107_8_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_1107_8 (.CI(n46124), .I0(byte_transmit_counter_c[6]), .I1(GND_net), 
            .CO(n46125));
    SB_LUT4 add_1107_7_lut (.I0(n52664), .I1(byte_transmit_counter_c[5]), 
            .I2(GND_net), .I3(n46123), .O(n52668)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1107_7_lut.LUT_INIT = 16'h8228;
    SB_DFF data_in_frame_0___i36 (.Q(\data_in_frame[4]_c [3]), .C(clk16MHz), 
           .D(n52223));   // verilog/coms.v(128[12] 296[6])
    SB_LUT4 select_715_Select_42_i2_4_lut (.I0(\data_out_frame[5] [2]), .I1(\FRAME_MATCHER.i_31__N_2320 ), 
            .I2(control_mode_c[2]), .I3(\FRAME_MATCHER.state_31__N_2423 [3]), 
            .O(n2_adj_5111));   // verilog/coms.v(146[4] 295[11])
    defparam select_715_Select_42_i2_4_lut.LUT_INIT = 16'hc088;
    SB_DFF data_in_frame_0___i37 (.Q(\data_in_frame[4]_c [4]), .C(clk16MHz), 
           .D(n52221));   // verilog/coms.v(128[12] 296[6])
    SB_DFF data_in_frame_0___i38 (.Q(\data_in_frame[4]_c [5]), .C(clk16MHz), 
           .D(n52215));   // verilog/coms.v(128[12] 296[6])
    SB_DFF data_in_frame_0___i39 (.Q(\data_in_frame[4][6] ), .C(clk16MHz), 
           .D(n26291));   // verilog/coms.v(128[12] 296[6])
    SB_LUT4 i3_4_lut_adj_1105 (.I0(n47750), .I1(n53436), .I2(n53094), 
            .I3(\data_out_frame[16] [4]), .O(n54719));
    defparam i3_4_lut_adj_1105.LUT_INIT = 16'h6996;
    SB_CARRY add_1107_7 (.CI(n46123), .I0(byte_transmit_counter_c[5]), .I1(GND_net), 
            .CO(n46124));
    SB_LUT4 add_1107_6_lut (.I0(n52664), .I1(byte_transmit_counter_c[4]), 
            .I2(GND_net), .I3(n46122), .O(n52669)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1107_6_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_1107_6 (.CI(n46122), .I0(byte_transmit_counter_c[4]), .I1(GND_net), 
            .CO(n46123));
    SB_LUT4 i1_4_lut_adj_1106 (.I0(\FRAME_MATCHER.i_31__N_2320 ), .I1(\data_out_frame[5] [1]), 
            .I2(\control_mode[1] ), .I3(\FRAME_MATCHER.state_31__N_2423 [3]), 
            .O(n2_adj_5110));   // verilog/coms.v(146[4] 295[11])
    defparam i1_4_lut_adj_1106.LUT_INIT = 16'ha088;
    SB_LUT4 add_1107_5_lut (.I0(n52664), .I1(byte_transmit_counter_c[3]), 
            .I2(GND_net), .I3(n46121), .O(n52670)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1107_5_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i1_4_lut_adj_1107 (.I0(\FRAME_MATCHER.i_31__N_2320 ), .I1(\data_out_frame[5] [0]), 
            .I2(\control_mode[0] ), .I3(\FRAME_MATCHER.state_31__N_2423 [3]), 
            .O(n2_adj_5109));   // verilog/coms.v(146[4] 295[11])
    defparam i1_4_lut_adj_1107.LUT_INIT = 16'ha088;
    SB_DFF data_in_frame_0___i40 (.Q(\data_in_frame[4][7] ), .C(clk16MHz), 
           .D(n26294));   // verilog/coms.v(128[12] 296[6])
    SB_DFF data_in_frame_0___i41 (.Q(\data_in_frame[5] [0]), .C(clk16MHz), 
           .D(n26297));   // verilog/coms.v(128[12] 296[6])
    SB_DFFESS data_out_frame_0___i45 (.Q(\data_out_frame[5] [4]), .C(clk16MHz), 
            .E(n2568), .D(n2_adj_5116), .S(n52681));   // verilog/coms.v(128[12] 296[6])
    SB_DFF data_in_0___i2 (.Q(\data_in[0] [1]), .C(clk16MHz), .D(n26392));   // verilog/coms.v(128[12] 296[6])
    SB_DFFESS data_out_frame_0___i46 (.Q(\data_out_frame[5] [5]), .C(clk16MHz), 
            .E(n2568), .D(n2_adj_5117), .S(n52683));   // verilog/coms.v(128[12] 296[6])
    SB_DFFESS data_out_frame_0___i47 (.Q(\data_out_frame[5] [6]), .C(clk16MHz), 
            .E(n2568), .D(n2_adj_5118), .S(n52684));   // verilog/coms.v(128[12] 296[6])
    SB_CARRY add_1107_5 (.CI(n46121), .I0(byte_transmit_counter_c[3]), .I1(GND_net), 
            .CO(n46122));
    SB_LUT4 add_1107_4_lut (.I0(n52664), .I1(\byte_transmit_counter[2] ), 
            .I2(GND_net), .I3(n46120), .O(n52671)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1107_4_lut.LUT_INIT = 16'h8228;
    SB_DFFESS data_out_frame_0___i209 (.Q(\data_out_frame[26] [0]), .C(clk16MHz), 
            .E(n2568), .D(n3_adj_5119), .S(n52841));   // verilog/coms.v(128[12] 296[6])
    SB_CARRY add_1107_4 (.CI(n46120), .I0(\byte_transmit_counter[2] ), .I1(GND_net), 
            .CO(n46121));
    SB_LUT4 i1_2_lut_adj_1108 (.I0(\data_out_frame[17] [0]), .I1(n53094), 
            .I2(GND_net), .I3(GND_net), .O(n23134));
    defparam i1_2_lut_adj_1108.LUT_INIT = 16'h6666;
    SB_LUT4 add_1107_3_lut (.I0(n52664), .I1(byte_transmit_counter_c[1]), 
            .I2(GND_net), .I3(n46119), .O(n52672)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1107_3_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_1107_3 (.CI(n46119), .I0(byte_transmit_counter_c[1]), .I1(GND_net), 
            .CO(n46120));
    SB_LUT4 add_1107_2_lut (.I0(n52664), .I1(byte_transmit_counter[0]), 
            .I2(tx_transmit_N_3189), .I3(GND_net), .O(n52666)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1107_2_lut.LUT_INIT = 16'h8228;
    SB_DFFESS data_out_frame_0___i48 (.Q(\data_out_frame[5] [7]), .C(clk16MHz), 
            .E(n2568), .D(n2_adj_5113), .S(n52685));   // verilog/coms.v(128[12] 296[6])
    SB_CARRY add_1107_2 (.CI(GND_net), .I0(byte_transmit_counter[0]), .I1(tx_transmit_N_3189), 
            .CO(n46119));
    SB_DFF data_in_0___i3 (.Q(\data_in[0] [2]), .C(clk16MHz), .D(n26391));   // verilog/coms.v(128[12] 296[6])
    SB_DFFESS data_out_frame_0___i210 (.Q(\data_out_frame[26] [1]), .C(clk16MHz), 
            .E(n2568), .D(n3_adj_5103), .S(n52840));   // verilog/coms.v(128[12] 296[6])
    SB_DFFESS data_out_frame_0___i49 (.Q(\data_out_frame[6] [0]), .C(clk16MHz), 
            .E(n2568), .D(n2_adj_5060), .S(n52686));   // verilog/coms.v(128[12] 296[6])
    SB_LUT4 i12722_3_lut_4_lut (.I0(Kp_23__N_1583), .I1(n29100), .I2(\data_in_frame[16] [1]), 
            .I3(\deadband[1] ), .O(n26326));
    defparam i12722_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFF data_in_0___i4 (.Q(\data_in[0] [3]), .C(clk16MHz), .D(n26390));   // verilog/coms.v(128[12] 296[6])
    SB_DFFESS data_out_frame_0___i211 (.Q(\data_out_frame[26] [2]), .C(clk16MHz), 
            .E(n2568), .D(n3), .S(n52839));   // verilog/coms.v(128[12] 296[6])
    SB_LUT4 i12723_3_lut_4_lut (.I0(Kp_23__N_1583), .I1(n29100), .I2(\data_in_frame[12] [7]), 
            .I3(IntegralLimit[15]), .O(n26327));
    defparam i12723_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1_2_lut_adj_1109 (.I0(\data_out_frame[4] [7]), .I1(\data_out_frame[7] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n52976));   // verilog/coms.v(74[16:34])
    defparam i1_2_lut_adj_1109.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1110 (.I0(\data_out_frame[5] [3]), .I1(\data_out_frame[9] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n52992));
    defparam i1_2_lut_adj_1110.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_1111 (.I0(\data_out_frame[7] [4]), .I1(n52992), 
            .I2(n52976), .I3(\data_out_frame[5] [1]), .O(n22752));   // verilog/coms.v(74[16:34])
    defparam i3_4_lut_adj_1111.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1112 (.I0(\data_out_frame[5] [3]), .I1(\data_out_frame[5] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n22519));   // verilog/coms.v(72[16:62])
    defparam i1_2_lut_adj_1112.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1113 (.I0(\data_out_frame[10] [0]), .I1(\data_out_frame[11] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n53256));   // verilog/coms.v(77[16:43])
    defparam i1_2_lut_adj_1113.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1114 (.I0(\data_out_frame[7] [5]), .I1(\data_out_frame[9] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n53037));
    defparam i1_2_lut_adj_1114.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1115 (.I0(\data_out_frame[5] [6]), .I1(\data_out_frame[5] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n53216));   // verilog/coms.v(74[16:34])
    defparam i1_2_lut_adj_1115.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1116 (.I0(\data_out_frame[10] [0]), .I1(n53037), 
            .I2(\data_out_frame[10] [1]), .I3(n6_adj_5120), .O(n53150));
    defparam i4_4_lut_adj_1116.LUT_INIT = 16'h6996;
    SB_LUT4 mux_1003_i24_3_lut_4_lut (.I0(Kp_23__N_1583), .I1(n29100), .I2(\data_in_frame[1][7] ), 
            .I3(\data_in_frame[17] [7]), .O(n4553[23]));
    defparam mux_1003_i24_3_lut_4_lut.LUT_INIT = 16'hf870;
    SB_LUT4 i13172_3_lut_4_lut (.I0(Kp_23__N_1583), .I1(n29100), .I2(\data_in_frame[2] [0]), 
            .I3(\Kp[8] ), .O(n26776));
    defparam i13172_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2_3_lut_adj_1117 (.I0(n23461), .I1(n53150), .I2(\data_out_frame[12] [2]), 
            .I3(GND_net), .O(n22545));   // verilog/coms.v(75[16:27])
    defparam i2_3_lut_adj_1117.LUT_INIT = 16'h9696;
    SB_LUT4 i13174_3_lut_4_lut (.I0(Kp_23__N_1583), .I1(n29100), .I2(\data_in_frame[3][7] ), 
            .I3(\Kp[7] ), .O(n26778));
    defparam i13174_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i3_4_lut_adj_1118 (.I0(n23123), .I1(n53256), .I2(n22519), 
            .I3(n22752), .O(n21977));   // verilog/coms.v(77[16:43])
    defparam i3_4_lut_adj_1118.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1119 (.I0(\data_out_frame[14] [3]), .I1(n22545), 
            .I2(GND_net), .I3(GND_net), .O(n53342));
    defparam i1_2_lut_adj_1119.LUT_INIT = 16'h6666;
    SB_LUT4 i12736_3_lut_4_lut (.I0(Kp_23__N_1583), .I1(n29100), .I2(\data_in_frame[12] [6]), 
            .I3(IntegralLimit[14]), .O(n26340));
    defparam i12736_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i6_4_lut_adj_1120 (.I0(n53439), .I1(n47750), .I2(\data_out_frame[14] [7]), 
            .I3(\data_out_frame[17] [1]), .O(n14_adj_5121));
    defparam i6_4_lut_adj_1120.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut_adj_1121 (.I0(\data_out_frame[21] [3]), .I1(n14_adj_5121), 
            .I2(n10_adj_5122), .I3(n21993), .O(n48764));
    defparam i7_4_lut_adj_1121.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1122 (.I0(n55477), .I1(n48764), .I2(GND_net), 
            .I3(GND_net), .O(n48809));
    defparam i1_2_lut_adj_1122.LUT_INIT = 16'h6666;
    SB_LUT4 i12737_3_lut_4_lut (.I0(Kp_23__N_1583), .I1(n29100), .I2(\data_in_frame[12] [5]), 
            .I3(IntegralLimit[13]), .O(n26341));
    defparam i12737_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4_4_lut_adj_1123 (.I0(\data_out_frame[21] [2]), .I1(n53291), 
            .I2(n23134), .I3(n4), .O(n10_adj_5123));
    defparam i4_4_lut_adj_1123.LUT_INIT = 16'h6996;
    SB_LUT4 i5_4_lut_adj_1124 (.I0(\data_out_frame[16] [3]), .I1(n10_adj_5123), 
            .I2(n53538), .I3(n4_adj_5124), .O(n55268));
    defparam i5_4_lut_adj_1124.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1125 (.I0(\data_out_frame[10] [7]), .I1(n23635), 
            .I2(GND_net), .I3(GND_net), .O(n53568));
    defparam i1_2_lut_adj_1125.LUT_INIT = 16'h6666;
    SB_LUT4 i5_4_lut_adj_1126 (.I0(n53586), .I1(\data_out_frame[10] [5]), 
            .I2(\data_out_frame[6] [0]), .I3(\data_out_frame[8] [2]), .O(n12_adj_5125));   // verilog/coms.v(75[16:43])
    defparam i5_4_lut_adj_1126.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_1127 (.I0(n22533), .I1(n12_adj_5125), .I2(n53332), 
            .I3(\data_out_frame[8] [4]), .O(n1521));   // verilog/coms.v(75[16:43])
    defparam i6_4_lut_adj_1127.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1128 (.I0(\data_out_frame[4] [2]), .I1(\data_out_frame[6] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n53100));   // verilog/coms.v(76[16:43])
    defparam i1_2_lut_adj_1128.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_1129 (.I0(\data_out_frame[4] [4]), .I1(\data_out_frame[4] [3]), 
            .I2(\data_out_frame[6] [5]), .I3(GND_net), .O(n23629));
    defparam i2_3_lut_adj_1129.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1130 (.I0(\data_out_frame[6] [1]), .I1(\data_out_frame[5] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_5126));   // verilog/coms.v(75[16:27])
    defparam i1_2_lut_adj_1130.LUT_INIT = 16'h6666;
    SB_LUT4 select_715_Select_39_i2_4_lut (.I0(\data_out_frame[4] [7]), .I1(\FRAME_MATCHER.i_31__N_2320 ), 
            .I2(ID[7]), .I3(\FRAME_MATCHER.state_31__N_2423 [3]), .O(n2_adj_5108));   // verilog/coms.v(146[4] 295[11])
    defparam select_715_Select_39_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i4_4_lut_adj_1131 (.I0(n53324), .I1(n22533), .I2(\data_out_frame[4] [0]), 
            .I3(n6_adj_5126), .O(n53515));   // verilog/coms.v(75[16:27])
    defparam i4_4_lut_adj_1131.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1132 (.I0(n22533), .I1(n53043), .I2(GND_net), 
            .I3(GND_net), .O(n23077));   // verilog/coms.v(76[16:43])
    defparam i1_2_lut_adj_1132.LUT_INIT = 16'h6666;
    SB_LUT4 i2_2_lut_adj_1133 (.I0(\data_out_frame[11] [0]), .I1(\data_out_frame[10] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n10_adj_5127));   // verilog/coms.v(75[16:27])
    defparam i2_2_lut_adj_1133.LUT_INIT = 16'h6666;
    SB_LUT4 i6_4_lut_adj_1134 (.I0(\data_out_frame[12] [7]), .I1(n23077), 
            .I2(n53515), .I3(n23629), .O(n14_adj_5128));   // verilog/coms.v(75[16:27])
    defparam i6_4_lut_adj_1134.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut_adj_1135 (.I0(\data_out_frame[13] [1]), .I1(n14_adj_5128), 
            .I2(n10_adj_5127), .I3(n53568), .O(n53559));   // verilog/coms.v(75[16:27])
    defparam i7_4_lut_adj_1135.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1136 (.I0(\data_out_frame[12] [6]), .I1(n53109), 
            .I2(n1521), .I3(GND_net), .O(n53439));
    defparam i2_3_lut_adj_1136.LUT_INIT = 16'h9696;
    SB_LUT4 select_715_Select_38_i2_4_lut (.I0(\data_out_frame[4] [6]), .I1(\FRAME_MATCHER.i_31__N_2320 ), 
            .I2(ID[6]), .I3(\FRAME_MATCHER.state_31__N_2423 [3]), .O(n2_adj_5107));   // verilog/coms.v(146[4] 295[11])
    defparam select_715_Select_38_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_adj_1137 (.I0(\data_out_frame[15] [2]), .I1(\data_out_frame[15] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n53391));
    defparam i1_2_lut_adj_1137.LUT_INIT = 16'h6666;
    SB_LUT4 i12738_3_lut_4_lut (.I0(Kp_23__N_1583), .I1(n29100), .I2(\data_in_frame[4][7] ), 
            .I3(\Ki[15] ), .O(n26342));
    defparam i12738_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1_2_lut_adj_1138 (.I0(\data_out_frame[10] [4]), .I1(\data_out_frame[6] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n23126));   // verilog/coms.v(73[16:27])
    defparam i1_2_lut_adj_1138.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1139 (.I0(\data_out_frame[8] [3]), .I1(\data_out_frame[8] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n53388));   // verilog/coms.v(76[16:27])
    defparam i1_2_lut_adj_1139.LUT_INIT = 16'h6666;
    SB_LUT4 select_715_Select_37_i2_4_lut (.I0(\data_out_frame[4] [5]), .I1(\FRAME_MATCHER.i_31__N_2320 ), 
            .I2(ID[5]), .I3(\FRAME_MATCHER.state_31__N_2423 [3]), .O(n2_adj_5106));   // verilog/coms.v(146[4] 295[11])
    defparam select_715_Select_37_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_adj_1140 (.I0(\data_out_frame[4] [1]), .I1(\data_out_frame[6] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n53586));   // verilog/coms.v(76[16:27])
    defparam i1_2_lut_adj_1140.LUT_INIT = 16'h6666;
    SB_LUT4 i12739_3_lut_4_lut (.I0(Kp_23__N_1583), .I1(n29100), .I2(\data_in_frame[4][6] ), 
            .I3(\Ki[14] ), .O(n26343));
    defparam i12739_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4_4_lut_adj_1141 (.I0(\data_out_frame[12] [5]), .I1(n53586), 
            .I2(n53388), .I3(n23126), .O(n10_adj_5129));   // verilog/coms.v(76[16:27])
    defparam i4_4_lut_adj_1141.LUT_INIT = 16'h6996;
    SB_LUT4 select_715_Select_36_i2_4_lut (.I0(\data_out_frame[4] [4]), .I1(\FRAME_MATCHER.i_31__N_2320 ), 
            .I2(ID[4]), .I3(\FRAME_MATCHER.state_31__N_2423 [3]), .O(n2_adj_5105));   // verilog/coms.v(146[4] 295[11])
    defparam select_715_Select_36_i2_4_lut.LUT_INIT = 16'hc088;
    SB_DFF data_in_0___i5 (.Q(\data_in[0] [4]), .C(clk16MHz), .D(n26389));   // verilog/coms.v(128[12] 296[6])
    SB_LUT4 i5_3_lut_adj_1142 (.I0(n53535), .I1(n10_adj_5129), .I2(\data_out_frame[10] [3]), 
            .I3(GND_net), .O(n53109));   // verilog/coms.v(76[16:27])
    defparam i5_3_lut_adj_1142.LUT_INIT = 16'h9696;
    SB_LUT4 i12740_3_lut_4_lut (.I0(Kp_23__N_1583), .I1(n29100), .I2(\data_in_frame[4]_c [5]), 
            .I3(\Ki[13] ), .O(n26344));
    defparam i12740_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2_3_lut_adj_1143 (.I0(\data_out_frame[7] [6]), .I1(\data_out_frame[8] [0]), 
            .I2(\data_out_frame[7] [7]), .I3(GND_net), .O(n23461));   // verilog/coms.v(86[17:70])
    defparam i2_3_lut_adj_1143.LUT_INIT = 16'h9696;
    SB_DFF data_in_frame_0___i87 (.Q(\data_in_frame[10] [6]), .C(clk16MHz), 
           .D(n26066));   // verilog/coms.v(128[12] 296[6])
    SB_LUT4 i1_2_lut_adj_1144 (.I0(\data_out_frame[5] [4]), .I1(\data_out_frame[8] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n53113));   // verilog/coms.v(86[17:70])
    defparam i1_2_lut_adj_1144.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1145 (.I0(\data_out_frame[12] [4]), .I1(\data_out_frame[6] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n7_c));   // verilog/coms.v(86[17:70])
    defparam i1_2_lut_adj_1145.LUT_INIT = 16'h6666;
    SB_LUT4 i5_4_lut_adj_1146 (.I0(n53113), .I1(n7_c), .I2(n23461), .I3(n8_adj_5130), 
            .O(n53394));   // verilog/coms.v(86[17:70])
    defparam i5_4_lut_adj_1146.LUT_INIT = 16'h6996;
    SB_LUT4 select_715_Select_35_i2_4_lut (.I0(\data_out_frame[4] [3]), .I1(\FRAME_MATCHER.i_31__N_2320 ), 
            .I2(ID[3]), .I3(\FRAME_MATCHER.state_31__N_2423 [3]), .O(n2_adj_5104));   // verilog/coms.v(146[4] 295[11])
    defparam select_715_Select_35_i2_4_lut.LUT_INIT = 16'hc088;
    SB_DFF data_in_frame_0___i88 (.Q(\data_in_frame[10] [7]), .C(clk16MHz), 
           .D(n52311));   // verilog/coms.v(128[12] 296[6])
    SB_LUT4 i1_2_lut_adj_1147 (.I0(\data_out_frame[17] [2]), .I1(\data_out_frame[17] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n22967));
    defparam i1_2_lut_adj_1147.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1148 (.I0(\data_out_frame[7] [5]), .I1(\data_out_frame[7] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n53204));   // verilog/coms.v(76[16:27])
    defparam i1_2_lut_adj_1148.LUT_INIT = 16'h6666;
    SB_DFF data_in_0___i6 (.Q(\data_in[0] [5]), .C(clk16MHz), .D(n26388));   // verilog/coms.v(128[12] 296[6])
    SB_DFF data_in_0___i7 (.Q(\data_in[0] [6]), .C(clk16MHz), .D(n26387));   // verilog/coms.v(128[12] 296[6])
    SB_DFF data_in_frame_0___i50 (.Q(\data_in_frame[6] [1]), .C(clk16MHz), 
           .D(n26584));   // verilog/coms.v(128[12] 296[6])
    SB_LUT4 i1_2_lut_adj_1149 (.I0(\data_out_frame[7] [7]), .I1(\data_out_frame[6] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n52961));
    defparam i1_2_lut_adj_1149.LUT_INIT = 16'h6666;
    SB_DFF data_in_frame_0___i132 (.Q(\data_in_frame[16] [3]), .C(clk16MHz), 
           .D(n26593));   // verilog/coms.v(128[12] 296[6])
    SB_DFF data_in_frame_0___i133 (.Q(\data_in_frame[16] [4]), .C(clk16MHz), 
           .D(n26596));   // verilog/coms.v(128[12] 296[6])
    SB_DFF data_in_frame_0___i134 (.Q(\data_in_frame[16] [5]), .C(clk16MHz), 
           .D(n26599));   // verilog/coms.v(128[12] 296[6])
    SB_DFF data_in_frame_0___i135 (.Q(\data_in_frame[16] [6]), .C(clk16MHz), 
           .D(n26602));   // verilog/coms.v(128[12] 296[6])
    SB_DFF data_in_frame_0___i136 (.Q(\data_in_frame[16] [7]), .C(clk16MHz), 
           .D(n26605));   // verilog/coms.v(128[12] 296[6])
    SB_DFF data_in_frame_0___i137 (.Q(\data_in_frame[17] [0]), .C(clk16MHz), 
           .D(n52163));   // verilog/coms.v(128[12] 296[6])
    SB_DFF data_in_frame_0___i138 (.Q(\data_in_frame[17] [1]), .C(clk16MHz), 
           .D(n52181));   // verilog/coms.v(128[12] 296[6])
    SB_DFF data_in_frame_0___i139 (.Q(\data_in_frame[17] [2]), .C(clk16MHz), 
           .D(n26615));   // verilog/coms.v(128[12] 296[6])
    SB_DFF data_in_frame_0___i140 (.Q(\data_in_frame[17] [3]), .C(clk16MHz), 
           .D(n26619));   // verilog/coms.v(128[12] 296[6])
    SB_DFF data_in_frame_0___i141 (.Q(\data_in_frame[17] [4]), .C(clk16MHz), 
           .D(n26622));   // verilog/coms.v(128[12] 296[6])
    SB_DFF data_in_frame_0___i142 (.Q(\data_in_frame[17] [5]), .C(clk16MHz), 
           .D(n26625));   // verilog/coms.v(128[12] 296[6])
    SB_DFF data_in_frame_0___i143 (.Q(\data_in_frame[17] [6]), .C(clk16MHz), 
           .D(n26628));   // verilog/coms.v(128[12] 296[6])
    SB_DFF data_in_frame_0___i144 (.Q(\data_in_frame[17] [7]), .C(clk16MHz), 
           .D(n26631));   // verilog/coms.v(128[12] 296[6])
    SB_DFF data_in_frame_0___i145 (.Q(\data_in_frame[18] [0]), .C(clk16MHz), 
           .D(n26634));   // verilog/coms.v(128[12] 296[6])
    SB_DFF data_in_frame_0___i146 (.Q(\data_in_frame[18] [1]), .C(clk16MHz), 
           .D(n27035));   // verilog/coms.v(128[12] 296[6])
    SB_DFF data_in_frame_0___i147 (.Q(\data_in_frame[18] [2]), .C(clk16MHz), 
           .D(n26640));   // verilog/coms.v(128[12] 296[6])
    SB_DFFE data_in_frame_0___i86 (.Q(\data_in_frame[10] [5]), .C(clk16MHz), 
            .E(VCC_net), .D(n27031));   // verilog/coms.v(128[12] 296[6])
    SB_LUT4 i4_4_lut_adj_1150 (.I0(\data_out_frame[12] [3]), .I1(n53518), 
            .I2(n52961), .I3(\data_out_frame[10] [2]), .O(n10_adj_5131));   // verilog/coms.v(76[16:27])
    defparam i4_4_lut_adj_1150.LUT_INIT = 16'h6996;
    SB_LUT4 i879_2_lut (.I0(\data_out_frame[12] [7]), .I1(\data_out_frame[12] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n1667));   // verilog/coms.v(86[17:28])
    defparam i879_2_lut.LUT_INIT = 16'h6666;
    SB_DFF data_in_0___i8 (.Q(\data_in[0] [7]), .C(clk16MHz), .D(n26386));   // verilog/coms.v(128[12] 296[6])
    SB_DFF data_in_0___i9 (.Q(\data_in[1] [0]), .C(clk16MHz), .D(n26385));   // verilog/coms.v(128[12] 296[6])
    SB_DFFE data_in_frame_0___i85 (.Q(\data_in_frame[10] [4]), .C(clk16MHz), 
            .E(VCC_net), .D(n27028));   // verilog/coms.v(128[12] 296[6])
    SB_DFFE data_in_frame_0___i84 (.Q(\data_in_frame[10] [3]), .C(clk16MHz), 
            .E(VCC_net), .D(n27025));   // verilog/coms.v(128[12] 296[6])
    SB_DFFE data_in_frame_0___i83 (.Q(\data_in_frame[10] [2]), .C(clk16MHz), 
            .E(VCC_net), .D(n27022));   // verilog/coms.v(128[12] 296[6])
    SB_LUT4 i1_2_lut_adj_1151 (.I0(\data_out_frame[8] [3]), .I1(\data_out_frame[8] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n53324));   // verilog/coms.v(75[16:27])
    defparam i1_2_lut_adj_1151.LUT_INIT = 16'h6666;
    SB_DFFE data_in_frame_0___i82 (.Q(\data_in_frame[10] [1]), .C(clk16MHz), 
            .E(VCC_net), .D(n27019));   // verilog/coms.v(128[12] 296[6])
    SB_DFFE data_in_frame_0___i81 (.Q(\data_in_frame[10] [0]), .C(clk16MHz), 
            .E(VCC_net), .D(n27016));   // verilog/coms.v(128[12] 296[6])
    SB_DFFE data_in_frame_0___i80 (.Q(\data_in_frame[9] [7]), .C(clk16MHz), 
            .E(VCC_net), .D(n27013));   // verilog/coms.v(128[12] 296[6])
    SB_DFFE data_in_frame_0___i79 (.Q(\data_in_frame[9] [6]), .C(clk16MHz), 
            .E(VCC_net), .D(n27010));   // verilog/coms.v(128[12] 296[6])
    SB_DFF data_in_0___i10 (.Q(\data_in[1] [1]), .C(clk16MHz), .D(n26384));   // verilog/coms.v(128[12] 296[6])
    SB_LUT4 i1_2_lut_adj_1152 (.I0(\data_out_frame[10] [4]), .I1(\data_out_frame[10] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n53103));   // verilog/coms.v(86[17:63])
    defparam i1_2_lut_adj_1152.LUT_INIT = 16'h6666;
    SB_LUT4 i6_4_lut_adj_1153 (.I0(n53324), .I1(\data_out_frame[5] [6]), 
            .I2(n53043), .I3(\data_out_frame[5] [7]), .O(n14_adj_5132));   // verilog/coms.v(86[17:70])
    defparam i6_4_lut_adj_1153.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut_adj_1154 (.I0(n1667), .I1(n14_adj_5132), .I2(n10_adj_5133), 
            .I3(\data_out_frame[8] [2]), .O(n21993));   // verilog/coms.v(86[17:70])
    defparam i7_4_lut_adj_1154.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1155 (.I0(n21993), .I1(\data_out_frame[15] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n53195));
    defparam i1_2_lut_adj_1155.LUT_INIT = 16'h6666;
    SB_DFF data_in_0___i11 (.Q(\data_in[1] [2]), .C(clk16MHz), .D(n26383));   // verilog/coms.v(128[12] 296[6])
    SB_DFF data_in_0___i12 (.Q(\data_in[1] [3]), .C(clk16MHz), .D(n26382));   // verilog/coms.v(128[12] 296[6])
    SB_DFF data_in_0___i13 (.Q(\data_in[1] [4]), .C(clk16MHz), .D(n26381));   // verilog/coms.v(128[12] 296[6])
    SB_DFF data_in_0___i14 (.Q(\data_in[1] [5]), .C(clk16MHz), .D(n26380));   // verilog/coms.v(128[12] 296[6])
    SB_DFF data_in_0___i15 (.Q(\data_in[1] [6]), .C(clk16MHz), .D(n26379));   // verilog/coms.v(128[12] 296[6])
    SB_DFF data_in_0___i16 (.Q(\data_in[1] [7]), .C(clk16MHz), .D(n26378));   // verilog/coms.v(128[12] 296[6])
    SB_DFFE data_in_frame_0___i78 (.Q(\data_in_frame[9] [5]), .C(clk16MHz), 
            .E(VCC_net), .D(n27007));   // verilog/coms.v(128[12] 296[6])
    SB_DFFE data_in_frame_0___i77 (.Q(\data_in_frame[9] [4]), .C(clk16MHz), 
            .E(VCC_net), .D(n27004));   // verilog/coms.v(128[12] 296[6])
    SB_DFFE data_in_frame_0___i76 (.Q(\data_in_frame[9] [3]), .C(clk16MHz), 
            .E(VCC_net), .D(n27001));   // verilog/coms.v(128[12] 296[6])
    SB_LUT4 i1_2_lut_adj_1156 (.I0(\data_out_frame[13] [0]), .I1(\data_out_frame[15] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n23375));
    defparam i1_2_lut_adj_1156.LUT_INIT = 16'h6666;
    SB_DFFE data_in_frame_0___i75 (.Q(\data_in_frame[9] [2]), .C(clk16MHz), 
            .E(VCC_net), .D(n26998));   // verilog/coms.v(128[12] 296[6])
    SB_DFFE data_in_frame_0___i74 (.Q(\data_in_frame[9] [1]), .C(clk16MHz), 
            .E(VCC_net), .D(n26995));   // verilog/coms.v(128[12] 296[6])
    SB_LUT4 i1_2_lut_adj_1157 (.I0(\data_out_frame[14] [5]), .I1(n52968), 
            .I2(GND_net), .I3(GND_net), .O(n53538));   // verilog/coms.v(76[16:43])
    defparam i1_2_lut_adj_1157.LUT_INIT = 16'h6666;
    SB_DFFE data_in_frame_0___i73 (.Q(\data_in_frame[9] [0]), .C(clk16MHz), 
            .E(VCC_net), .D(n26992));   // verilog/coms.v(128[12] 296[6])
    SB_LUT4 i2_3_lut_adj_1158 (.I0(n1521), .I1(\data_out_frame[14] [6]), 
            .I2(\data_out_frame[14] [7]), .I3(GND_net), .O(n53501));
    defparam i2_3_lut_adj_1158.LUT_INIT = 16'h9696;
    SB_DFF data_in_0___i17 (.Q(\data_in[2] [0]), .C(clk16MHz), .D(n26377));   // verilog/coms.v(128[12] 296[6])
    SB_LUT4 i4_4_lut_adj_1159 (.I0(n53501), .I1(\data_out_frame[12] [6]), 
            .I2(\data_out_frame[15] [0]), .I3(n53538), .O(n10_adj_5134));
    defparam i4_4_lut_adj_1159.LUT_INIT = 16'h6996;
    SB_DFF data_in_0___i18 (.Q(\data_in[2] [1]), .C(clk16MHz), .D(n26376));   // verilog/coms.v(128[12] 296[6])
    SB_DFF data_in_0___i19 (.Q(\data_in[2] [2]), .C(clk16MHz), .D(n26375));   // verilog/coms.v(128[12] 296[6])
    SB_LUT4 i1_4_lut_adj_1160 (.I0(\data_out_frame[21] [5]), .I1(n53267), 
            .I2(n10_adj_5134), .I3(\data_out_frame[17] [1]), .O(n53314));
    defparam i1_4_lut_adj_1160.LUT_INIT = 16'h9669;
    SB_DFF data_in_0___i20 (.Q(\data_in[2] [3]), .C(clk16MHz), .D(n26374));   // verilog/coms.v(128[12] 296[6])
    SB_DFF data_in_0___i21 (.Q(\data_in[2] [4]), .C(clk16MHz), .D(n26373));   // verilog/coms.v(128[12] 296[6])
    SB_DFFE data_in_frame_0___i72 (.Q(\data_in_frame[8] [7]), .C(clk16MHz), 
            .E(VCC_net), .D(n26989));   // verilog/coms.v(128[12] 296[6])
    SB_DFFE data_in_frame_0___i71 (.Q(\data_in_frame[8] [6]), .C(clk16MHz), 
            .E(VCC_net), .D(n26986));   // verilog/coms.v(128[12] 296[6])
    SB_DFFE data_in_frame_0___i70 (.Q(\data_in_frame[8] [5]), .C(clk16MHz), 
            .E(VCC_net), .D(n26983));   // verilog/coms.v(128[12] 296[6])
    SB_DFFE data_in_frame_0___i69 (.Q(\data_in_frame[8] [4]), .C(clk16MHz), 
            .E(VCC_net), .D(n26980));   // verilog/coms.v(128[12] 296[6])
    SB_LUT4 i4_4_lut_adj_1161 (.I0(n23375), .I1(n22967), .I2(n53195), 
            .I3(n53394), .O(n10_adj_5135));   // verilog/coms.v(86[17:63])
    defparam i4_4_lut_adj_1161.LUT_INIT = 16'h6996;
    SB_DFFE data_in_frame_0___i68 (.Q(\data_in_frame[8] [3]), .C(clk16MHz), 
            .E(VCC_net), .D(n26977));   // verilog/coms.v(128[12] 296[6])
    SB_LUT4 i5_3_lut_adj_1162 (.I0(n48497), .I1(n10_adj_5135), .I2(n4), 
            .I3(GND_net), .O(n48833));   // verilog/coms.v(86[17:63])
    defparam i5_3_lut_adj_1162.LUT_INIT = 16'h9696;
    SB_DFF data_in_0___i22 (.Q(\data_in[2] [5]), .C(clk16MHz), .D(n26372));   // verilog/coms.v(128[12] 296[6])
    SB_LUT4 i11_3_lut_adj_1163 (.I0(rx_data[1]), .I1(\data_in_frame[1] [1]), 
            .I2(n25161), .I3(GND_net), .O(n52175));   // verilog/coms.v(92[13:20])
    defparam i11_3_lut_adj_1163.LUT_INIT = 16'hcaca;
    SB_DFF data_in_0___i23 (.Q(\data_in[2] [6]), .C(clk16MHz), .D(n26371));   // verilog/coms.v(128[12] 296[6])
    SB_LUT4 select_715_Select_208_i3_4_lut (.I0(n55268), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(n48809), .I3(n53315), .O(n3_adj_5119));   // verilog/coms.v(146[4] 295[11])
    defparam select_715_Select_208_i3_4_lut.LUT_INIT = 16'h8448;
    SB_DFFE data_in_frame_0___i67 (.Q(\data_in_frame[8] [2]), .C(clk16MHz), 
            .E(VCC_net), .D(n26974));   // verilog/coms.v(128[12] 296[6])
    SB_DFFE data_in_frame_0___i66 (.Q(\data_in_frame[8] [1]), .C(clk16MHz), 
            .E(VCC_net), .D(n26971));   // verilog/coms.v(128[12] 296[6])
    SB_DFFE data_in_frame_0___i65 (.Q(\data_in_frame[8] [0]), .C(clk16MHz), 
            .E(VCC_net), .D(n26967));   // verilog/coms.v(128[12] 296[6])
    SB_DFFE data_in_frame_0___i64 (.Q(\data_in_frame[7] [7]), .C(clk16MHz), 
            .E(VCC_net), .D(n26964));   // verilog/coms.v(128[12] 296[6])
    SB_DFFE data_in_frame_0___i63 (.Q(\data_in_frame[7] [6]), .C(clk16MHz), 
            .E(VCC_net), .D(n26961));   // verilog/coms.v(128[12] 296[6])
    SB_LUT4 select_715_Select_46_i2_4_lut (.I0(\data_out_frame[5] [6]), .I1(\FRAME_MATCHER.i_31__N_2320 ), 
            .I2(\control_mode[6] ), .I3(\FRAME_MATCHER.state_31__N_2423 [3]), 
            .O(n2_adj_5118));   // verilog/coms.v(146[4] 295[11])
    defparam select_715_Select_46_i2_4_lut.LUT_INIT = 16'hc088;
    SB_DFFE data_in_frame_0___i62 (.Q(\data_in_frame[7] [5]), .C(clk16MHz), 
            .E(VCC_net), .D(n26958));   // verilog/coms.v(128[12] 296[6])
    SB_DFFE data_in_frame_0___i61 (.Q(\data_in_frame[7] [4]), .C(clk16MHz), 
            .E(VCC_net), .D(n26955));   // verilog/coms.v(128[12] 296[6])
    SB_DFFE data_in_frame_0___i60 (.Q(\data_in_frame[7] [3]), .C(clk16MHz), 
            .E(VCC_net), .D(n26952));   // verilog/coms.v(128[12] 296[6])
    SB_DFF data_in_0___i24 (.Q(\data_in[2] [7]), .C(clk16MHz), .D(n26370));   // verilog/coms.v(128[12] 296[6])
    SB_LUT4 i17269_3_lut_4_lut (.I0(Kp_23__N_1583), .I1(n29100), .I2(\data_in_frame[3] [0]), 
            .I3(\data_in_frame[19] [0]), .O(n4553[0]));
    defparam i17269_3_lut_4_lut.LUT_INIT = 16'hf870;
    SB_DFF data_in_0___i25 (.Q(\data_in[3] [0]), .C(clk16MHz), .D(n26369));   // verilog/coms.v(128[12] 296[6])
    SB_DFF data_in_0___i26 (.Q(\data_in[3] [1]), .C(clk16MHz), .D(n26368));   // verilog/coms.v(128[12] 296[6])
    SB_DFF data_in_0___i27 (.Q(\data_in[3] [2]), .C(clk16MHz), .D(n26367));   // verilog/coms.v(128[12] 296[6])
    SB_DFF data_in_0___i28 (.Q(\data_in[3] [3]), .C(clk16MHz), .D(n26366));   // verilog/coms.v(128[12] 296[6])
    SB_DFFE data_in_frame_0___i59 (.Q(\data_in_frame[7] [2]), .C(clk16MHz), 
            .E(VCC_net), .D(n26949));   // verilog/coms.v(128[12] 296[6])
    SB_DFFE data_in_frame_0___i58 (.Q(\data_in_frame[7] [1]), .C(clk16MHz), 
            .E(VCC_net), .D(n26946));   // verilog/coms.v(128[12] 296[6])
    SB_DFFE data_in_frame_0___i57 (.Q(\data_in_frame[7] [0]), .C(clk16MHz), 
            .E(VCC_net), .D(n26943));   // verilog/coms.v(128[12] 296[6])
    SB_DFFE data_in_frame_0___i56 (.Q(\data_in_frame[6] [7]), .C(clk16MHz), 
            .E(VCC_net), .D(n26940));   // verilog/coms.v(128[12] 296[6])
    SB_DFFE data_in_frame_0___i55 (.Q(\data_in_frame[6] [6]), .C(clk16MHz), 
            .E(VCC_net), .D(n26937));   // verilog/coms.v(128[12] 296[6])
    SB_LUT4 select_715_Select_45_i2_4_lut (.I0(\data_out_frame[5] [5]), .I1(\FRAME_MATCHER.i_31__N_2320 ), 
            .I2(\control_mode[5] ), .I3(\FRAME_MATCHER.state_31__N_2423 [3]), 
            .O(n2_adj_5117));   // verilog/coms.v(146[4] 295[11])
    defparam select_715_Select_45_i2_4_lut.LUT_INIT = 16'hc088;
    SB_DFFE data_in_frame_0___i54 (.Q(\data_in_frame[6] [5]), .C(clk16MHz), 
            .E(VCC_net), .D(n26934));   // verilog/coms.v(128[12] 296[6])
    SB_DFFE data_in_frame_0___i53 (.Q(\data_in_frame[6] [4]), .C(clk16MHz), 
            .E(VCC_net), .D(n26931));   // verilog/coms.v(128[12] 296[6])
    SB_DFF data_in_0___i29 (.Q(\data_in[3] [4]), .C(clk16MHz), .D(n26365));   // verilog/coms.v(128[12] 296[6])
    SB_DFF data_in_0___i30 (.Q(\data_in[3] [5]), .C(clk16MHz), .D(n26364));   // verilog/coms.v(128[12] 296[6])
    SB_DFF data_in_frame_0___i148 (.Q(\data_in_frame[18] [3]), .C(clk16MHz), 
           .D(n26643));   // verilog/coms.v(128[12] 296[6])
    SB_DFF data_in_frame_0___i149 (.Q(\data_in_frame[18] [4]), .C(clk16MHz), 
           .D(n26646));   // verilog/coms.v(128[12] 296[6])
    SB_DFF data_in_frame_0___i150 (.Q(\data_in_frame[18] [5]), .C(clk16MHz), 
           .D(n26649));   // verilog/coms.v(128[12] 296[6])
    SB_DFF data_in_frame_0___i151 (.Q(\data_in_frame[18]_c [6]), .C(clk16MHz), 
           .D(n26652));   // verilog/coms.v(128[12] 296[6])
    SB_DFF data_in_frame_0___i152 (.Q(\data_in_frame[18][7] ), .C(clk16MHz), 
           .D(n26655));   // verilog/coms.v(128[12] 296[6])
    SB_DFF data_in_frame_0___i153 (.Q(\data_in_frame[19] [0]), .C(clk16MHz), 
           .D(n52199));   // verilog/coms.v(128[12] 296[6])
    SB_DFF data_in_frame_0___i154 (.Q(\data_in_frame[19] [1]), .C(clk16MHz), 
           .D(n26662));   // verilog/coms.v(128[12] 296[6])
    SB_DFF data_in_frame_0___i155 (.Q(\data_in_frame[19] [2]), .C(clk16MHz), 
           .D(n26665));   // verilog/coms.v(128[12] 296[6])
    SB_DFF data_in_frame_0___i156 (.Q(\data_in_frame[19] [3]), .C(clk16MHz), 
           .D(n26671));   // verilog/coms.v(128[12] 296[6])
    SB_DFF data_in_frame_0___i157 (.Q(\data_in_frame[19] [4]), .C(clk16MHz), 
           .D(n52233));   // verilog/coms.v(128[12] 296[6])
    SB_DFF data_in_frame_0___i158 (.Q(\data_in_frame[19] [5]), .C(clk16MHz), 
           .D(n26677));   // verilog/coms.v(128[12] 296[6])
    SB_DFFE data_in_frame_0___i52 (.Q(\data_in_frame[6] [3]), .C(clk16MHz), 
            .E(VCC_net), .D(n26917));   // verilog/coms.v(128[12] 296[6])
    SB_DFF data_in_frame_0___i89 (.Q(\data_in_frame[11] [0]), .C(clk16MHz), 
           .D(n26092));   // verilog/coms.v(128[12] 296[6])
    SB_DFF control_mode_i0_i1 (.Q(\control_mode[1] ), .C(clk16MHz), .D(n26915));   // verilog/coms.v(128[12] 296[6])
    SB_DFF control_mode_i0_i2 (.Q(control_mode_c[2]), .C(clk16MHz), .D(n26914));   // verilog/coms.v(128[12] 296[6])
    SB_DFF control_mode_i0_i3 (.Q(control_mode_c[3]), .C(clk16MHz), .D(n26913));   // verilog/coms.v(128[12] 296[6])
    SB_DFF control_mode_i0_i4 (.Q(\control_mode[4] ), .C(clk16MHz), .D(n26912));   // verilog/coms.v(128[12] 296[6])
    SB_DFF control_mode_i0_i5 (.Q(\control_mode[5] ), .C(clk16MHz), .D(n26911));   // verilog/coms.v(128[12] 296[6])
    SB_DFF control_mode_i0_i6 (.Q(\control_mode[6] ), .C(clk16MHz), .D(n26910));   // verilog/coms.v(128[12] 296[6])
    SB_DFF control_mode_i0_i7 (.Q(control_mode[7]), .C(clk16MHz), .D(n26909));   // verilog/coms.v(128[12] 296[6])
    SB_LUT4 select_715_Select_44_i2_4_lut (.I0(\data_out_frame[5] [4]), .I1(\FRAME_MATCHER.i_31__N_2320 ), 
            .I2(\control_mode[4] ), .I3(\FRAME_MATCHER.state_31__N_2423 [3]), 
            .O(n2_adj_5116));   // verilog/coms.v(146[4] 295[11])
    defparam select_715_Select_44_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 \FRAME_MATCHER.i_1939_add_4_33_lut  (.I0(n59781), .I1(n63273), 
            .I2(\FRAME_MATCHER.i [31]), .I3(n46612), .O(n24833)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_1939_add_4_33_lut .LUT_INIT = 16'h8BB8;
    SB_DFF current_limit_i0_i1 (.Q(current_limit[1]), .C(clk16MHz), .D(n26908));   // verilog/coms.v(128[12] 296[6])
    SB_DFF current_limit_i0_i2 (.Q(current_limit[2]), .C(clk16MHz), .D(n26907));   // verilog/coms.v(128[12] 296[6])
    SB_DFF current_limit_i0_i3 (.Q(current_limit[3]), .C(clk16MHz), .D(n26906));   // verilog/coms.v(128[12] 296[6])
    SB_DFF current_limit_i0_i4 (.Q(current_limit[4]), .C(clk16MHz), .D(n26905));   // verilog/coms.v(128[12] 296[6])
    SB_DFF current_limit_i0_i5 (.Q(current_limit[5]), .C(clk16MHz), .D(n26904));   // verilog/coms.v(128[12] 296[6])
    SB_DFF current_limit_i0_i6 (.Q(current_limit[6]), .C(clk16MHz), .D(n26903));   // verilog/coms.v(128[12] 296[6])
    SB_DFF current_limit_i0_i7 (.Q(current_limit[7]), .C(clk16MHz), .D(n26902));   // verilog/coms.v(128[12] 296[6])
    SB_DFF current_limit_i0_i8 (.Q(current_limit[8]), .C(clk16MHz), .D(n26901));   // verilog/coms.v(128[12] 296[6])
    SB_DFF current_limit_i0_i9 (.Q(current_limit[9]), .C(clk16MHz), .D(n26900));   // verilog/coms.v(128[12] 296[6])
    SB_DFF current_limit_i0_i10 (.Q(current_limit[10]), .C(clk16MHz), .D(n26899));   // verilog/coms.v(128[12] 296[6])
    SB_DFF current_limit_i0_i11 (.Q(current_limit[11]), .C(clk16MHz), .D(n26898));   // verilog/coms.v(128[12] 296[6])
    SB_DFF current_limit_i0_i12 (.Q(current_limit[12]), .C(clk16MHz), .D(n26897));   // verilog/coms.v(128[12] 296[6])
    SB_DFF current_limit_i0_i13 (.Q(current_limit[13]), .C(clk16MHz), .D(n26896));   // verilog/coms.v(128[12] 296[6])
    SB_DFF current_limit_i0_i14 (.Q(current_limit[14]), .C(clk16MHz), .D(n26895));   // verilog/coms.v(128[12] 296[6])
    SB_DFF current_limit_i0_i15 (.Q(current_limit[15]), .C(clk16MHz), .D(n26894));   // verilog/coms.v(128[12] 296[6])
    SB_DFFR PWMLimit_i0_i1 (.Q(PWMLimit[1]), .C(clk16MHz), .D(n26893), 
            .R(reset));   // verilog/coms.v(128[12] 296[6])
    SB_DFFS PWMLimit_i0_i2 (.Q(PWMLimit[2]), .C(clk16MHz), .D(n26892), 
            .S(reset));   // verilog/coms.v(128[12] 296[6])
    SB_DFFR PWMLimit_i0_i3 (.Q(PWMLimit[3]), .C(clk16MHz), .D(n26891), 
            .R(reset));   // verilog/coms.v(128[12] 296[6])
    SB_DFF data_in_0___i31 (.Q(\data_in[3] [6]), .C(clk16MHz), .D(n26363));   // verilog/coms.v(128[12] 296[6])
    SB_DFF data_in_0___i32 (.Q(\data_in[3] [7]), .C(clk16MHz), .D(n26362));   // verilog/coms.v(128[12] 296[6])
    SB_DFF data_in_frame_0___i42 (.Q(\data_in_frame[5] [1]), .C(clk16MHz), 
           .D(n26316));   // verilog/coms.v(128[12] 296[6])
    SB_DFF data_in_frame_0___i43 (.Q(\data_in_frame[5] [2]), .C(clk16MHz), 
           .D(n26328));   // verilog/coms.v(128[12] 296[6])
    SB_DFF data_in_frame_0___i44 (.Q(\data_in_frame[5] [3]), .C(clk16MHz), 
           .D(n26331));   // verilog/coms.v(128[12] 296[6])
    SB_DFF data_in_frame_0___i45 (.Q(\data_in_frame[5] [4]), .C(clk16MHz), 
           .D(n26334));   // verilog/coms.v(128[12] 296[6])
    SB_DFF data_in_frame_0___i109 (.Q(\data_in_frame[13] [4]), .C(clk16MHz), 
           .D(n26337));   // verilog/coms.v(128[12] 296[6])
    SB_DFFS PWMLimit_i0_i4 (.Q(PWMLimit[4]), .C(clk16MHz), .D(n26890), 
            .S(reset));   // verilog/coms.v(128[12] 296[6])
    SB_DFFS PWMLimit_i0_i5 (.Q(PWMLimit[5]), .C(clk16MHz), .D(n26889), 
            .S(reset));   // verilog/coms.v(128[12] 296[6])
    SB_DFFS PWMLimit_i0_i6 (.Q(PWMLimit[6]), .C(clk16MHz), .D(n26888), 
            .S(reset));   // verilog/coms.v(128[12] 296[6])
    SB_DFFS PWMLimit_i0_i7 (.Q(PWMLimit[7]), .C(clk16MHz), .D(n26887), 
            .S(reset));   // verilog/coms.v(128[12] 296[6])
    SB_DFFS PWMLimit_i0_i8 (.Q(PWMLimit[8]), .C(clk16MHz), .D(n26886), 
            .S(reset));   // verilog/coms.v(128[12] 296[6])
    SB_DFFR PWMLimit_i0_i9 (.Q(PWMLimit[9]), .C(clk16MHz), .D(n26885), 
            .R(reset));   // verilog/coms.v(128[12] 296[6])
    SB_DFFR PWMLimit_i0_i10 (.Q(PWMLimit[10]), .C(clk16MHz), .D(n26884), 
            .R(reset));   // verilog/coms.v(128[12] 296[6])
    SB_DFFR PWMLimit_i0_i11 (.Q(PWMLimit[11]), .C(clk16MHz), .D(n26883), 
            .R(reset));   // verilog/coms.v(128[12] 296[6])
    SB_DFFR PWMLimit_i0_i12 (.Q(PWMLimit[12]), .C(clk16MHz), .D(n26882), 
            .R(reset));   // verilog/coms.v(128[12] 296[6])
    SB_DFFR PWMLimit_i0_i13 (.Q(PWMLimit[13]), .C(clk16MHz), .D(n26881), 
            .R(reset));   // verilog/coms.v(128[12] 296[6])
    SB_DFFR PWMLimit_i0_i14 (.Q(PWMLimit[14]), .C(clk16MHz), .D(n26880), 
            .R(reset));   // verilog/coms.v(128[12] 296[6])
    SB_DFFR PWMLimit_i0_i15 (.Q(PWMLimit[15]), .C(clk16MHz), .D(n26879), 
            .R(reset));   // verilog/coms.v(128[12] 296[6])
    SB_DFFR PWMLimit_i0_i16 (.Q(PWMLimit[16]), .C(clk16MHz), .D(n26878), 
            .R(reset));   // verilog/coms.v(128[12] 296[6])
    SB_DFFR PWMLimit_i0_i17 (.Q(PWMLimit[17]), .C(clk16MHz), .D(n26877), 
            .R(reset));   // verilog/coms.v(128[12] 296[6])
    SB_DFFR PWMLimit_i0_i18 (.Q(PWMLimit[18]), .C(clk16MHz), .D(n26876), 
            .R(reset));   // verilog/coms.v(128[12] 296[6])
    SB_DFFR PWMLimit_i0_i19 (.Q(PWMLimit[19]), .C(clk16MHz), .D(n26875), 
            .R(reset));   // verilog/coms.v(128[12] 296[6])
    SB_DFFR PWMLimit_i0_i20 (.Q(PWMLimit[20]), .C(clk16MHz), .D(n26874), 
            .R(reset));   // verilog/coms.v(128[12] 296[6])
    SB_DFFR Ki_i1 (.Q(\Ki[1] ), .C(clk16MHz), .D(n26356), .R(reset));   // verilog/coms.v(128[12] 296[6])
    SB_DFFR Ki_i2 (.Q(\Ki[2] ), .C(clk16MHz), .D(n26355), .R(reset));   // verilog/coms.v(128[12] 296[6])
    SB_DFFR Ki_i3 (.Q(\Ki[3] ), .C(clk16MHz), .D(n26354), .R(reset));   // verilog/coms.v(128[12] 296[6])
    SB_DFFR Ki_i4 (.Q(\Ki[4] ), .C(clk16MHz), .D(n26353), .R(reset));   // verilog/coms.v(128[12] 296[6])
    SB_DFFR Ki_i5 (.Q(\Ki[5] ), .C(clk16MHz), .D(n26352), .R(reset));   // verilog/coms.v(128[12] 296[6])
    SB_DFFR Ki_i6 (.Q(\Ki[6] ), .C(clk16MHz), .D(n26351), .R(reset));   // verilog/coms.v(128[12] 296[6])
    SB_DFFR PWMLimit_i0_i21 (.Q(PWMLimit[21]), .C(clk16MHz), .D(n26873), 
            .R(reset));   // verilog/coms.v(128[12] 296[6])
    SB_DFFR PWMLimit_i0_i22 (.Q(PWMLimit[22]), .C(clk16MHz), .D(n26872), 
            .R(reset));   // verilog/coms.v(128[12] 296[6])
    SB_DFFR PWMLimit_i0_i23 (.Q(PWMLimit[23]), .C(clk16MHz), .D(n26871), 
            .R(reset));   // verilog/coms.v(128[12] 296[6])
    SB_DFFR Ki_i7 (.Q(\Ki[7] ), .C(clk16MHz), .D(n26350), .R(reset));   // verilog/coms.v(128[12] 296[6])
    SB_LUT4 i13289_3_lut_4_lut (.I0(Kp_23__N_1583), .I1(n29100), .I2(\data_in_frame[10] [1]), 
            .I3(PWMLimit[1]), .O(n26893));
    defparam i13289_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFFR Ki_i8 (.Q(\Ki[8] ), .C(clk16MHz), .D(n26349), .R(reset));   // verilog/coms.v(128[12] 296[6])
    SB_DFFR Ki_i9 (.Q(\Ki[9] ), .C(clk16MHz), .D(n26348), .R(reset));   // verilog/coms.v(128[12] 296[6])
    SB_DFFR Ki_i10 (.Q(\Ki[10] ), .C(clk16MHz), .D(n26347), .R(reset));   // verilog/coms.v(128[12] 296[6])
    SB_DFFR Ki_i11 (.Q(\Ki[11] ), .C(clk16MHz), .D(n26346), .R(reset));   // verilog/coms.v(128[12] 296[6])
    SB_DFFE data_in_frame_0___i1 (.Q(\data_in_frame[0] [0]), .C(clk16MHz), 
            .E(VCC_net), .D(n26842));   // verilog/coms.v(128[12] 296[6])
    SB_LUT4 i17413_3_lut (.I0(n25161), .I1(rx_data[0]), .I2(\data_in_frame[1] [0]), 
            .I3(GND_net), .O(n26444));   // verilog/coms.v(92[13:20])
    defparam i17413_3_lut.LUT_INIT = 16'he4e4;
    SB_DFF data_in_frame_0___i2 (.Q(\data_in_frame[0] [1]), .C(clk16MHz), 
           .D(n26102));   // verilog/coms.v(128[12] 296[6])
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[14] [3]), .I2(\data_out_frame[15] [3]), 
            .I3(byte_transmit_counter_c[1]), .O(n63653));
    defparam byte_transmit_counter_0__bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_DFFESS data_out_frame_0___i50 (.Q(\data_out_frame[6] [1]), .C(clk16MHz), 
            .E(n2568), .D(n2_adj_5136), .S(n52687));   // verilog/coms.v(128[12] 296[6])
    SB_DFF data_in_frame_0___i3 (.Q(\data_in_frame[0] [2]), .C(clk16MHz), 
           .D(n26105));   // verilog/coms.v(128[12] 296[6])
    SB_DFF data_in_frame_0___i4 (.Q(\data_in_frame[0] [3]), .C(clk16MHz), 
           .D(n26108));   // verilog/coms.v(128[12] 296[6])
    SB_DFFE data_in_frame_0___i192 (.Q(\data_in_frame[23] [7]), .C(clk16MHz), 
            .E(VCC_net), .D(n26819));   // verilog/coms.v(128[12] 296[6])
    SB_DFFE data_in_frame_0___i191 (.Q(\data_in_frame[23] [6]), .C(clk16MHz), 
            .E(VCC_net), .D(n26816));   // verilog/coms.v(128[12] 296[6])
    SB_DFFE data_in_frame_0___i190 (.Q(\data_in_frame[23] [5]), .C(clk16MHz), 
            .E(VCC_net), .D(n26813));   // verilog/coms.v(128[12] 296[6])
    SB_DFFE data_in_frame_0___i189 (.Q(\data_in_frame[23] [4]), .C(clk16MHz), 
            .E(VCC_net), .D(n26810));   // verilog/coms.v(128[12] 296[6])
    SB_DFFE data_in_frame_0___i188 (.Q(\data_in_frame[23] [3]), .C(clk16MHz), 
            .E(VCC_net), .D(n26807));   // verilog/coms.v(128[12] 296[6])
    SB_DFFE data_in_frame_0___i187 (.Q(\data_in_frame[23] [2]), .C(clk16MHz), 
            .E(VCC_net), .D(n26804));   // verilog/coms.v(128[12] 296[6])
    SB_LUT4 \FRAME_MATCHER.i_1939_add_4_32_lut  (.I0(n59793), .I1(n63273), 
            .I2(\FRAME_MATCHER.i [30]), .I3(n46611), .O(n24831)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_1939_add_4_32_lut .LUT_INIT = 16'h8BB8;
    SB_CARRY \FRAME_MATCHER.i_1939_add_4_32  (.CI(n46611), .I0(n63273), 
            .I1(\FRAME_MATCHER.i [30]), .CO(n46612));
    SB_LUT4 i13280_3_lut_4_lut (.I0(Kp_23__N_1583), .I1(n29100), .I2(\data_in_frame[9] [2]), 
            .I3(PWMLimit[10]), .O(n26884));
    defparam i13280_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i48301_3_lut (.I0(rx_data[5]), .I1(\data_in_frame[4]_c [5]), 
            .I2(n7), .I3(GND_net), .O(n52215));   // verilog/coms.v(92[13:20])
    defparam i48301_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 \FRAME_MATCHER.i_1939_add_4_31_lut  (.I0(n59807), .I1(n63273), 
            .I2(\FRAME_MATCHER.i [29]), .I3(n46610), .O(n24829)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_1939_add_4_31_lut .LUT_INIT = 16'h8BB8;
    SB_CARRY \FRAME_MATCHER.i_1939_add_4_31  (.CI(n46610), .I0(n63273), 
            .I1(\FRAME_MATCHER.i [29]), .CO(n46611));
    SB_LUT4 \FRAME_MATCHER.i_1939_add_4_30_lut  (.I0(n59808), .I1(n63273), 
            .I2(\FRAME_MATCHER.i [28]), .I3(n46609), .O(n24827)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_1939_add_4_30_lut .LUT_INIT = 16'h8BB8;
    SB_LUT4 i48302_3_lut (.I0(rx_data[4]), .I1(\data_in_frame[4]_c [4]), 
            .I2(n7), .I3(GND_net), .O(n52221));   // verilog/coms.v(92[13:20])
    defparam i48302_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i48303_3_lut (.I0(rx_data[3]), .I1(\data_in_frame[4]_c [3]), 
            .I2(n7), .I3(GND_net), .O(n52223));   // verilog/coms.v(92[13:20])
    defparam i48303_3_lut.LUT_INIT = 16'hcaca;
    SB_DFFR Ki_i12 (.Q(\Ki[12] ), .C(clk16MHz), .D(n26345), .R(reset));   // verilog/coms.v(128[12] 296[6])
    SB_DFFR Ki_i13 (.Q(\Ki[13] ), .C(clk16MHz), .D(n26344), .R(reset));   // verilog/coms.v(128[12] 296[6])
    SB_DFF data_in_frame_0___i5 (.Q(\data_in_frame[0] [4]), .C(clk16MHz), 
           .D(n26112));   // verilog/coms.v(128[12] 296[6])
    SB_DFFE data_in_frame_0___i186 (.Q(\data_in_frame[23] [1]), .C(clk16MHz), 
            .E(VCC_net), .D(n26800));   // verilog/coms.v(128[12] 296[6])
    SB_DFFR Ki_i14 (.Q(\Ki[14] ), .C(clk16MHz), .D(n26343), .R(reset));   // verilog/coms.v(128[12] 296[6])
    SB_DFFR Ki_i15 (.Q(\Ki[15] ), .C(clk16MHz), .D(n26342), .R(reset));   // verilog/coms.v(128[12] 296[6])
    SB_DFFE data_in_frame_0___i185 (.Q(\data_in_frame[23] [0]), .C(clk16MHz), 
            .E(VCC_net), .D(n26797));   // verilog/coms.v(128[12] 296[6])
    SB_DFFR IntegralLimit_i0_i13 (.Q(IntegralLimit[13]), .C(clk16MHz), .D(n26341), 
            .R(reset));   // verilog/coms.v(128[12] 296[6])
    SB_DFFE data_in_frame_0___i184 (.Q(\data_in_frame[22] [7]), .C(clk16MHz), 
            .E(VCC_net), .D(n26794));   // verilog/coms.v(128[12] 296[6])
    SB_DFFR IntegralLimit_i0_i14 (.Q(IntegralLimit[14]), .C(clk16MHz), .D(n26340), 
            .R(reset));   // verilog/coms.v(128[12] 296[6])
    SB_DFFE data_in_frame_0___i183 (.Q(\data_in_frame[22] [6]), .C(clk16MHz), 
            .E(VCC_net), .D(n26791));   // verilog/coms.v(128[12] 296[6])
    SB_CARRY \FRAME_MATCHER.i_1939_add_4_30  (.CI(n46609), .I0(n63273), 
            .I1(\FRAME_MATCHER.i [28]), .CO(n46610));
    SB_LUT4 select_715_Select_34_i2_4_lut (.I0(\data_out_frame[4] [2]), .I1(\FRAME_MATCHER.i_31__N_2320 ), 
            .I2(ID[2]), .I3(\FRAME_MATCHER.state_31__N_2423 [3]), .O(n2_adj_5101));   // verilog/coms.v(146[4] 295[11])
    defparam select_715_Select_34_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 \FRAME_MATCHER.i_1939_add_4_29_lut  (.I0(n59809), .I1(n63273), 
            .I2(\FRAME_MATCHER.i [27]), .I3(n46608), .O(n24825)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_1939_add_4_29_lut .LUT_INIT = 16'h8BB8;
    SB_DFFE data_in_frame_0___i182 (.Q(\data_in_frame[22] [5]), .C(clk16MHz), 
            .E(VCC_net), .D(n26788));   // verilog/coms.v(128[12] 296[6])
    SB_DFFE data_in_frame_0___i181 (.Q(\data_in_frame[22] [4]), .C(clk16MHz), 
            .E(VCC_net), .D(n26785));   // verilog/coms.v(128[12] 296[6])
    SB_DFFE data_in_frame_0___i51 (.Q(\data_in_frame[6] [2]), .C(clk16MHz), 
            .E(VCC_net), .D(n26782));   // verilog/coms.v(128[12] 296[6])
    SB_DFF data_in_frame_0___i6 (.Q(\data_in_frame[0] [5]), .C(clk16MHz), 
           .D(n26115));   // verilog/coms.v(128[12] 296[6])
    SB_DFF data_in_frame_0___i7 (.Q(\data_in_frame[0] [6]), .C(clk16MHz), 
           .D(n26118));   // verilog/coms.v(128[12] 296[6])
    SB_LUT4 select_715_Select_33_i2_4_lut (.I0(\data_out_frame[4] [1]), .I1(\FRAME_MATCHER.i_31__N_2320 ), 
            .I2(ID[1]), .I3(\FRAME_MATCHER.state_31__N_2423 [3]), .O(n2_adj_5100));   // verilog/coms.v(146[4] 295[11])
    defparam select_715_Select_33_i2_4_lut.LUT_INIT = 16'hc088;
    SB_CARRY \FRAME_MATCHER.i_1939_add_4_29  (.CI(n46608), .I0(n63273), 
            .I1(\FRAME_MATCHER.i [27]), .CO(n46609));
    SB_DFFR Kp_i7 (.Q(\Kp[7] ), .C(clk16MHz), .D(n26778), .R(reset));   // verilog/coms.v(128[12] 296[6])
    SB_DFF data_in_frame_0___i159 (.Q(\data_in_frame[19] [6]), .C(clk16MHz), 
           .D(n26681));   // verilog/coms.v(128[12] 296[6])
    SB_DFFR Kp_i8 (.Q(\Kp[8] ), .C(clk16MHz), .D(n26776), .R(reset));   // verilog/coms.v(128[12] 296[6])
    SB_DFF data_in_frame_0___i160 (.Q(\data_in_frame[19] [7]), .C(clk16MHz), 
           .D(n26684));   // verilog/coms.v(128[12] 296[6])
    SB_DFF data_in_frame_0___i161 (.Q(\data_in_frame[20] [0]), .C(clk16MHz), 
           .D(n26687));   // verilog/coms.v(128[12] 296[6])
    SB_DFF data_in_frame_0___i162 (.Q(\data_in_frame[20] [1]), .C(clk16MHz), 
           .D(n26690));   // verilog/coms.v(128[12] 296[6])
    SB_DFFESS data_out_frame_0___i212 (.Q(\data_out_frame[26] [3]), .C(clk16MHz), 
            .E(n2568), .D(n3_adj_5138), .S(n52838));   // verilog/coms.v(128[12] 296[6])
    SB_LUT4 n63653_bdd_4_lut (.I0(n63653), .I1(\data_out_frame[13] [3]), 
            .I2(\data_out_frame[12] [3]), .I3(byte_transmit_counter_c[1]), 
            .O(n56844));
    defparam n63653_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFFER setpoint_i0_i23 (.Q(setpoint[23]), .C(clk16MHz), .E(n24563), 
            .D(n4553[23]), .R(reset));   // verilog/coms.v(128[12] 296[6])
    SB_DFFR IntegralLimit_i0_i15 (.Q(IntegralLimit[15]), .C(clk16MHz), .D(n26327), 
            .R(reset));   // verilog/coms.v(128[12] 296[6])
    SB_DFFR deadband_i0_i1 (.Q(\deadband[1] ), .C(clk16MHz), .D(n26326), 
            .R(reset));   // verilog/coms.v(128[12] 296[6])
    SB_DFFR deadband_i0_i2 (.Q(deadband_c[2]), .C(clk16MHz), .D(n26325), 
            .R(reset));   // verilog/coms.v(128[12] 296[6])
    SB_DFFR deadband_i0_i3 (.Q(deadband[3]), .C(clk16MHz), .D(n26324), 
            .R(reset));   // verilog/coms.v(128[12] 296[6])
    SB_DFFR deadband_i0_i4 (.Q(deadband[4]), .C(clk16MHz), .D(n26323), 
            .R(reset));   // verilog/coms.v(128[12] 296[6])
    SB_DFFR deadband_i0_i5 (.Q(deadband[5]), .C(clk16MHz), .D(n26322), 
            .R(reset));   // verilog/coms.v(128[12] 296[6])
    SB_DFFR deadband_i0_i6 (.Q(deadband[6]), .C(clk16MHz), .D(n26321), 
            .R(reset));   // verilog/coms.v(128[12] 296[6])
    SB_DFFR deadband_i0_i7 (.Q(deadband[7]), .C(clk16MHz), .D(n26320), 
            .R(reset));   // verilog/coms.v(128[12] 296[6])
    SB_DFFR deadband_i0_i8 (.Q(deadband[8]), .C(clk16MHz), .D(n26319), 
            .R(reset));   // verilog/coms.v(128[12] 296[6])
    SB_DFFR deadband_i0_i9 (.Q(deadband[9]), .C(clk16MHz), .D(n26315), 
            .R(reset));   // verilog/coms.v(128[12] 296[6])
    SB_DFFR IntegralLimit_i0_i16 (.Q(IntegralLimit[16]), .C(clk16MHz), .D(n26314), 
            .R(reset));   // verilog/coms.v(128[12] 296[6])
    SB_DFFR IntegralLimit_i0_i17 (.Q(IntegralLimit[17]), .C(clk16MHz), .D(n26313), 
            .R(reset));   // verilog/coms.v(128[12] 296[6])
    SB_DFFR deadband_i0_i10 (.Q(deadband[10]), .C(clk16MHz), .D(n26312), 
            .R(reset));   // verilog/coms.v(128[12] 296[6])
    SB_DFFR deadband_i0_i11 (.Q(deadband[11]), .C(clk16MHz), .D(n26311), 
            .R(reset));   // verilog/coms.v(128[12] 296[6])
    SB_DFFR deadband_i0_i12 (.Q(deadband[12]), .C(clk16MHz), .D(n26310), 
            .R(reset));   // verilog/coms.v(128[12] 296[6])
    SB_DFFR deadband_i0_i13 (.Q(deadband[13]), .C(clk16MHz), .D(n26309), 
            .R(reset));   // verilog/coms.v(128[12] 296[6])
    SB_DFFR deadband_i0_i14 (.Q(deadband[14]), .C(clk16MHz), .D(n26308), 
            .R(reset));   // verilog/coms.v(128[12] 296[6])
    SB_DFFR deadband_i0_i15 (.Q(deadband[15]), .C(clk16MHz), .D(n26307), 
            .R(reset));   // verilog/coms.v(128[12] 296[6])
    SB_DFFR deadband_i0_i16 (.Q(deadband[16]), .C(clk16MHz), .D(n26306), 
            .R(reset));   // verilog/coms.v(128[12] 296[6])
    SB_DFFR deadband_i0_i17 (.Q(deadband[17]), .C(clk16MHz), .D(n26305), 
            .R(reset));   // verilog/coms.v(128[12] 296[6])
    SB_DFFR deadband_i0_i18 (.Q(deadband[18]), .C(clk16MHz), .D(n26304), 
            .R(reset));   // verilog/coms.v(128[12] 296[6])
    SB_LUT4 i13279_3_lut_4_lut (.I0(Kp_23__N_1583), .I1(n29100), .I2(\data_in_frame[9] [3]), 
            .I3(PWMLimit[11]), .O(n26883));
    defparam i13279_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFFER setpoint_i0_i22 (.Q(setpoint[22]), .C(clk16MHz), .E(n24563), 
            .D(n4553[22]), .R(reset));   // verilog/coms.v(128[12] 296[6])
    SB_DFFER setpoint_i0_i21 (.Q(setpoint[21]), .C(clk16MHz), .E(n24563), 
            .D(n4553[21]), .R(reset));   // verilog/coms.v(128[12] 296[6])
    SB_DFFER setpoint_i0_i20 (.Q(setpoint[20]), .C(clk16MHz), .E(n24563), 
            .D(n4553[20]), .R(reset));   // verilog/coms.v(128[12] 296[6])
    SB_DFFER setpoint_i0_i19 (.Q(setpoint[19]), .C(clk16MHz), .E(n24563), 
            .D(n4553[19]), .R(reset));   // verilog/coms.v(128[12] 296[6])
    SB_DFFER setpoint_i0_i18 (.Q(setpoint[18]), .C(clk16MHz), .E(n24563), 
            .D(n4553[18]), .R(reset));   // verilog/coms.v(128[12] 296[6])
    SB_DFFER setpoint_i0_i17 (.Q(setpoint[17]), .C(clk16MHz), .E(n24563), 
            .D(n4553[17]), .R(reset));   // verilog/coms.v(128[12] 296[6])
    SB_DFFER setpoint_i0_i16 (.Q(setpoint[16]), .C(clk16MHz), .E(n24563), 
            .D(n4553[16]), .R(reset));   // verilog/coms.v(128[12] 296[6])
    SB_DFFER setpoint_i0_i15 (.Q(setpoint[15]), .C(clk16MHz), .E(n24563), 
            .D(n4553[15]), .R(reset));   // verilog/coms.v(128[12] 296[6])
    SB_DFFER setpoint_i0_i14 (.Q(setpoint[14]), .C(clk16MHz), .E(n24563), 
            .D(n4553[14]), .R(reset));   // verilog/coms.v(128[12] 296[6])
    SB_DFFER setpoint_i0_i13 (.Q(setpoint[13]), .C(clk16MHz), .E(n24563), 
            .D(n4553[13]), .R(reset));   // verilog/coms.v(128[12] 296[6])
    SB_DFFER setpoint_i0_i12 (.Q(setpoint[12]), .C(clk16MHz), .E(n24563), 
            .D(n4553[12]), .R(reset));   // verilog/coms.v(128[12] 296[6])
    SB_DFFER setpoint_i0_i11 (.Q(setpoint[11]), .C(clk16MHz), .E(n24563), 
            .D(n4553[11]), .R(reset));   // verilog/coms.v(128[12] 296[6])
    SB_DFFER setpoint_i0_i10 (.Q(setpoint[10]), .C(clk16MHz), .E(n24563), 
            .D(n4553[10]), .R(reset));   // verilog/coms.v(128[12] 296[6])
    SB_DFFER setpoint_i0_i9 (.Q(setpoint[9]), .C(clk16MHz), .E(n24563), 
            .D(n4553[9]), .R(reset));   // verilog/coms.v(128[12] 296[6])
    SB_DFFER setpoint_i0_i8 (.Q(setpoint[8]), .C(clk16MHz), .E(n24563), 
            .D(n4553[8]), .R(reset));   // verilog/coms.v(128[12] 296[6])
    SB_DFFER setpoint_i0_i7 (.Q(setpoint[7]), .C(clk16MHz), .E(n24563), 
            .D(n4553[7]), .R(reset));   // verilog/coms.v(128[12] 296[6])
    SB_DFFER setpoint_i0_i6 (.Q(setpoint[6]), .C(clk16MHz), .E(n24563), 
            .D(n4553[6]), .R(reset));   // verilog/coms.v(128[12] 296[6])
    SB_DFFER setpoint_i0_i5 (.Q(setpoint[5]), .C(clk16MHz), .E(n24563), 
            .D(n4553[5]), .R(reset));   // verilog/coms.v(128[12] 296[6])
    SB_DFFER setpoint_i0_i4 (.Q(setpoint[4]), .C(clk16MHz), .E(n24563), 
            .D(n4553[4]), .R(reset));   // verilog/coms.v(128[12] 296[6])
    SB_DFFER setpoint_i0_i3 (.Q(setpoint[3]), .C(clk16MHz), .E(n24563), 
            .D(n4553[3]), .R(reset));   // verilog/coms.v(128[12] 296[6])
    SB_DFFER setpoint_i0_i2 (.Q(setpoint[2]), .C(clk16MHz), .E(n24563), 
            .D(n4553[2]), .R(reset));   // verilog/coms.v(128[12] 296[6])
    SB_DFFER setpoint_i0_i1 (.Q(setpoint[1]), .C(clk16MHz), .E(n24563), 
            .D(n4553[1]), .R(reset));   // verilog/coms.v(128[12] 296[6])
    SB_DFFR deadband_i0_i19 (.Q(deadband[19]), .C(clk16MHz), .D(n26303), 
            .R(reset));   // verilog/coms.v(128[12] 296[6])
    SB_LUT4 i13278_3_lut_4_lut (.I0(Kp_23__N_1583), .I1(n29100), .I2(\data_in_frame[9] [4]), 
            .I3(PWMLimit[12]), .O(n26882));
    defparam i13278_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 \FRAME_MATCHER.i_1939_add_4_28_lut  (.I0(n59810), .I1(n63273), 
            .I2(\FRAME_MATCHER.i [26]), .I3(n46607), .O(n24823)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_1939_add_4_28_lut .LUT_INIT = 16'h8BB8;
    SB_LUT4 i13363_3_lut_4_lut (.I0(n8_adj_5139), .I1(n52882), .I2(rx_data[0]), 
            .I3(\data_in_frame[8] [0]), .O(n26967));
    defparam i13363_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_CARRY \FRAME_MATCHER.i_1939_add_4_28  (.CI(n46607), .I0(n63273), 
            .I1(\FRAME_MATCHER.i [26]), .CO(n46608));
    SB_LUT4 \FRAME_MATCHER.i_1939_add_4_27_lut  (.I0(n59811), .I1(n63273), 
            .I2(\FRAME_MATCHER.i [25]), .I3(n46606), .O(n24821)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_1939_add_4_27_lut .LUT_INIT = 16'h8BB8;
    SB_CARRY \FRAME_MATCHER.i_1939_add_4_27  (.CI(n46606), .I0(n63273), 
            .I1(\FRAME_MATCHER.i [25]), .CO(n46607));
    SB_LUT4 select_715_Select_97_i2_4_lut (.I0(\data_out_frame[12] [1]), .I1(\FRAME_MATCHER.i_31__N_2320 ), 
            .I2(setpoint[17]), .I3(\FRAME_MATCHER.state_31__N_2423 [3]), 
            .O(n2_adj_5097));   // verilog/coms.v(146[4] 295[11])
    defparam select_715_Select_97_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_715_Select_96_i2_4_lut (.I0(\data_out_frame[12] [0]), .I1(\FRAME_MATCHER.i_31__N_2320 ), 
            .I2(setpoint[16]), .I3(\FRAME_MATCHER.state_31__N_2423 [3]), 
            .O(n2_adj_5094));   // verilog/coms.v(146[4] 295[11])
    defparam select_715_Select_96_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_715_Select_32_i2_4_lut (.I0(\data_out_frame[4] [0]), .I1(\FRAME_MATCHER.i_31__N_2320 ), 
            .I2(ID[0]), .I3(\FRAME_MATCHER.state_31__N_2423 [3]), .O(n2_adj_5092));   // verilog/coms.v(146[4] 295[11])
    defparam select_715_Select_32_i2_4_lut.LUT_INIT = 16'hc088;
    SB_DFFR deadband_i0_i20 (.Q(deadband[20]), .C(clk16MHz), .D(n26302), 
            .R(reset));   // verilog/coms.v(128[12] 296[6])
    SB_DFFESS data_out_frame_0___i213 (.Q(\data_out_frame[26] [4]), .C(clk16MHz), 
            .E(n2568), .D(n3_adj_5140), .S(n52837));   // verilog/coms.v(128[12] 296[6])
    SB_DFFR deadband_i0_i21 (.Q(deadband[21]), .C(clk16MHz), .D(n26301), 
            .R(reset));   // verilog/coms.v(128[12] 296[6])
    SB_DFFESS data_out_frame_0___i214 (.Q(\data_out_frame[26] [5]), .C(clk16MHz), 
            .E(n2568), .D(n3_adj_5141), .S(n52836));   // verilog/coms.v(128[12] 296[6])
    SB_DFFR deadband_i0_i22 (.Q(deadband[22]), .C(clk16MHz), .D(n26300), 
            .R(reset));   // verilog/coms.v(128[12] 296[6])
    SB_DFFESS data_out_frame_0___i215 (.Q(\data_out_frame[26][6] ), .C(clk16MHz), 
            .E(n2568), .D(n3_adj_5142), .S(n52835));   // verilog/coms.v(128[12] 296[6])
    SB_DFFESS data_out_frame_0___i216 (.Q(\data_out_frame[26] [7]), .C(clk16MHz), 
            .E(n2568), .D(n3_adj_5143), .S(n52834));   // verilog/coms.v(128[12] 296[6])
    SB_DFFESS data_out_frame_0___i217 (.Q(\data_out_frame[27] [0]), .C(clk16MHz), 
            .E(n2568), .D(n3_adj_5144), .S(n52833));   // verilog/coms.v(128[12] 296[6])
    SB_DFFESS data_out_frame_0___i218 (.Q(\data_out_frame[27] [1]), .C(clk16MHz), 
            .E(n2568), .D(n3_adj_5145), .S(n52832));   // verilog/coms.v(128[12] 296[6])
    SB_DFFESS data_out_frame_0___i219 (.Q(\data_out_frame[27] [2]), .C(clk16MHz), 
            .E(n2568), .D(n3_adj_5146), .S(n52831));   // verilog/coms.v(128[12] 296[6])
    SB_DFFESS data_out_frame_0___i220 (.Q(\data_out_frame[27] [3]), .C(clk16MHz), 
            .E(n2568), .D(n3_adj_5147), .S(n52830));   // verilog/coms.v(128[12] 296[6])
    SB_DFFESS data_out_frame_0___i221 (.Q(\data_out_frame[27] [4]), .C(clk16MHz), 
            .E(n2568), .D(n3_adj_5148), .S(n52829));   // verilog/coms.v(128[12] 296[6])
    SB_DFFESS data_out_frame_0___i222 (.Q(\data_out_frame[27] [5]), .C(clk16MHz), 
            .E(n2568), .D(n3_adj_5149), .S(n52828));   // verilog/coms.v(128[12] 296[6])
    SB_DFFESS data_out_frame_0___i223 (.Q(\data_out_frame[27][6] ), .C(clk16MHz), 
            .E(n2568), .D(n3_adj_5150), .S(n52827));   // verilog/coms.v(128[12] 296[6])
    SB_DFFESS data_out_frame_0___i224 (.Q(\data_out_frame[27] [7]), .C(clk16MHz), 
            .E(n2568), .D(n3_adj_5151), .S(n52826));   // verilog/coms.v(128[12] 296[6])
    SB_DFFR deadband_i0_i23 (.Q(deadband[23]), .C(clk16MHz), .D(n26287), 
            .R(reset));   // verilog/coms.v(128[12] 296[6])
    SB_DFFR IntegralLimit_i0_i18 (.Q(IntegralLimit[18]), .C(clk16MHz), .D(n26286), 
            .R(reset));   // verilog/coms.v(128[12] 296[6])
    SB_DFFR IntegralLimit_i0_i19 (.Q(IntegralLimit[19]), .C(clk16MHz), .D(n26282), 
            .R(reset));   // verilog/coms.v(128[12] 296[6])
    SB_DFFR IntegralLimit_i0_i20 (.Q(IntegralLimit[20]), .C(clk16MHz), .D(n26281), 
            .R(reset));   // verilog/coms.v(128[12] 296[6])
    SB_DFFR IntegralLimit_i0_i21 (.Q(IntegralLimit[21]), .C(clk16MHz), .D(n26280), 
            .R(reset));   // verilog/coms.v(128[12] 296[6])
    SB_LUT4 i13367_3_lut_4_lut (.I0(n8_adj_5139), .I1(n52882), .I2(rx_data[1]), 
            .I3(\data_in_frame[8] [1]), .O(n26971));
    defparam i13367_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 select_715_Select_95_i2_4_lut (.I0(\data_out_frame[11] [7]), .I1(\FRAME_MATCHER.i_31__N_2320 ), 
            .I2(encoder1_position[7]), .I3(\FRAME_MATCHER.state_31__N_2423 [3]), 
            .O(n2_adj_5091));   // verilog/coms.v(146[4] 295[11])
    defparam select_715_Select_95_i2_4_lut.LUT_INIT = 16'hc088;
    SB_DFFESS byte_transmit_counter_i0_i1 (.Q(byte_transmit_counter_c[1]), 
            .C(clk16MHz), .E(n2568), .D(n1_c), .S(n52672));   // verilog/coms.v(128[12] 296[6])
    SB_DFFESS byte_transmit_counter_i0_i2 (.Q(\byte_transmit_counter[2] ), 
            .C(clk16MHz), .E(n2568), .D(n1_adj_5152), .S(n52671));   // verilog/coms.v(128[12] 296[6])
    SB_DFFESS byte_transmit_counter_i0_i3 (.Q(byte_transmit_counter_c[3]), 
            .C(clk16MHz), .E(n2568), .D(n1_adj_5153), .S(n52670));   // verilog/coms.v(128[12] 296[6])
    SB_DFFESS byte_transmit_counter_i0_i4 (.Q(byte_transmit_counter_c[4]), 
            .C(clk16MHz), .E(n2568), .D(n1_adj_5154), .S(n52669));   // verilog/coms.v(128[12] 296[6])
    SB_DFFESS byte_transmit_counter_i0_i5 (.Q(byte_transmit_counter_c[5]), 
            .C(clk16MHz), .E(n2568), .D(n1_adj_5155), .S(n52668));   // verilog/coms.v(128[12] 296[6])
    SB_DFFESS byte_transmit_counter_i0_i6 (.Q(byte_transmit_counter_c[6]), 
            .C(clk16MHz), .E(n2568), .D(n1_adj_5156), .S(n52667));   // verilog/coms.v(128[12] 296[6])
    SB_DFFR IntegralLimit_i0_i22 (.Q(IntegralLimit[22]), .C(clk16MHz), .D(n26249), 
            .R(reset));   // verilog/coms.v(128[12] 296[6])
    SB_DFFR IntegralLimit_i0_i23 (.Q(IntegralLimit[23]), .C(clk16MHz), .D(n26248), 
            .R(reset));   // verilog/coms.v(128[12] 296[6])
    SB_DFFS Kp_i1 (.Q(\Kp[1] ), .C(clk16MHz), .D(n26247), .S(reset));   // verilog/coms.v(128[12] 296[6])
    SB_DFFR Kp_i2 (.Q(\Kp[2] ), .C(clk16MHz), .D(n26246), .R(reset));   // verilog/coms.v(128[12] 296[6])
    SB_DFFESS byte_transmit_counter_i0_i7 (.Q(byte_transmit_counter_c[7]), 
            .C(clk16MHz), .E(n2568), .D(n1_adj_5157), .S(n52665));   // verilog/coms.v(128[12] 296[6])
    SB_DFF \FRAME_MATCHER.rx_data_ready_prev_4001  (.Q(\FRAME_MATCHER.rx_data_ready_prev ), 
           .C(clk16MHz), .D(n26243));   // verilog/coms.v(128[12] 296[6])
    SB_DFFS Kp_i3 (.Q(\Kp[3] ), .C(clk16MHz), .D(n26241), .S(reset));   // verilog/coms.v(128[12] 296[6])
    SB_DFFR Kp_i4 (.Q(\Kp[4] ), .C(clk16MHz), .D(n26237), .R(reset));   // verilog/coms.v(128[12] 296[6])
    SB_DFFR Kp_i5 (.Q(\Kp[5] ), .C(clk16MHz), .D(n26230), .R(reset));   // verilog/coms.v(128[12] 296[6])
    SB_LUT4 i1_4_lut_adj_1164 (.I0(\FRAME_MATCHER.i_31__N_2320 ), .I1(\data_out_frame[11] [6]), 
            .I2(encoder1_position[6]), .I3(\FRAME_MATCHER.state_31__N_2423 [3]), 
            .O(n2_adj_5090));   // verilog/coms.v(146[4] 295[11])
    defparam i1_4_lut_adj_1164.LUT_INIT = 16'ha088;
    SB_LUT4 \FRAME_MATCHER.i_1939_add_4_26_lut  (.I0(n59812), .I1(n63273), 
            .I2(\FRAME_MATCHER.i [24]), .I3(n46605), .O(n24819)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_1939_add_4_26_lut .LUT_INIT = 16'h8BB8;
    SB_LUT4 select_715_Select_93_i2_4_lut (.I0(\data_out_frame[11] [5]), .I1(\FRAME_MATCHER.i_31__N_2320 ), 
            .I2(encoder1_position[5]), .I3(\FRAME_MATCHER.state_31__N_2423 [3]), 
            .O(n2_adj_5089));   // verilog/coms.v(146[4] 295[11])
    defparam select_715_Select_93_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i13370_3_lut_4_lut (.I0(n8_adj_5139), .I1(n52882), .I2(rx_data[2]), 
            .I3(\data_in_frame[8] [2]), .O(n26974));
    defparam i13370_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFFESS data_out_frame_0___i99 (.Q(\data_out_frame[12] [2]), .C(clk16MHz), 
            .E(n2568), .D(n2_adj_5158), .S(n52727));   // verilog/coms.v(128[12] 296[6])
    SB_LUT4 i13373_3_lut_4_lut (.I0(n8_adj_5139), .I1(n52882), .I2(rx_data[3]), 
            .I3(\data_in_frame[8] [3]), .O(n26977));
    defparam i13373_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13376_3_lut_4_lut (.I0(n8_adj_5139), .I1(n52882), .I2(rx_data[4]), 
            .I3(\data_in_frame[8] [4]), .O(n26980));
    defparam i13376_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13379_3_lut_4_lut (.I0(n8_adj_5139), .I1(n52882), .I2(rx_data[5]), 
            .I3(\data_in_frame[8] [5]), .O(n26983));
    defparam i13379_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 select_715_Select_92_i2_4_lut (.I0(\data_out_frame[11] [4]), .I1(\FRAME_MATCHER.i_31__N_2320 ), 
            .I2(encoder1_position[4]), .I3(\FRAME_MATCHER.state_31__N_2423 [3]), 
            .O(n2_adj_5088));   // verilog/coms.v(146[4] 295[11])
    defparam select_715_Select_92_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_715_Select_91_i2_4_lut (.I0(\data_out_frame[11] [3]), .I1(\FRAME_MATCHER.i_31__N_2320 ), 
            .I2(encoder1_position[3]), .I3(\FRAME_MATCHER.state_31__N_2423 [3]), 
            .O(n2_adj_5087));   // verilog/coms.v(146[4] 295[11])
    defparam select_715_Select_91_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i13382_3_lut_4_lut (.I0(n8_adj_5139), .I1(n52882), .I2(rx_data[6]), 
            .I3(\data_in_frame[8] [6]), .O(n26986));
    defparam i13382_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13385_3_lut_4_lut (.I0(n8_adj_5139), .I1(n52882), .I2(rx_data[7]), 
            .I3(\data_in_frame[8] [7]), .O(n26989));
    defparam i13385_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFFESS data_out_frame_0___i100 (.Q(\data_out_frame[12] [3]), .C(clk16MHz), 
            .E(n2568), .D(n2_adj_5159), .S(n52728));   // verilog/coms.v(128[12] 296[6])
    SB_DFF data_in_frame_0___i8 (.Q(\data_in_frame[0] [7]), .C(clk16MHz), 
           .D(n26121));   // verilog/coms.v(128[12] 296[6])
    SB_DFFR Kp_i9 (.Q(\Kp[9] ), .C(clk16MHz), .D(n26771), .R(reset));   // verilog/coms.v(128[12] 296[6])
    SB_DFF data_in_frame_0___i163 (.Q(\data_in_frame[20] [2]), .C(clk16MHz), 
           .D(n26693));   // verilog/coms.v(128[12] 296[6])
    SB_DFF data_in_frame_0___i164 (.Q(\data_in_frame[20] [3]), .C(clk16MHz), 
           .D(n26696));   // verilog/coms.v(128[12] 296[6])
    SB_DFF data_in_frame_0___i165 (.Q(\data_in_frame[20] [4]), .C(clk16MHz), 
           .D(n26699));   // verilog/coms.v(128[12] 296[6])
    SB_DFF data_in_frame_0___i90 (.Q(\data_in_frame[11] [1]), .C(clk16MHz), 
           .D(n26767));   // verilog/coms.v(128[12] 296[6])
    SB_DFFR Kp_i10 (.Q(\Kp[10] ), .C(clk16MHz), .D(n26766), .R(reset));   // verilog/coms.v(128[12] 296[6])
    SB_DFFR Kp_i11 (.Q(\Kp[11] ), .C(clk16MHz), .D(n26765), .R(reset));   // verilog/coms.v(128[12] 296[6])
    SB_DFF data_in_frame_0___i166 (.Q(\data_in_frame[20] [5]), .C(clk16MHz), 
           .D(n26702));   // verilog/coms.v(128[12] 296[6])
    SB_DFFS IntegralLimit_i0_i1 (.Q(IntegralLimit[1]), .C(clk16MHz), .D(n26763), 
            .S(reset));   // verilog/coms.v(128[12] 296[6])
    SB_DFFR Kp_i12 (.Q(\Kp[12] ), .C(clk16MHz), .D(n26762), .R(reset));   // verilog/coms.v(128[12] 296[6])
    SB_DFF data_in_frame_0___i91 (.Q(\data_in_frame[11] [2]), .C(clk16MHz), 
           .D(n26127));   // verilog/coms.v(128[12] 296[6])
    SB_DFF data_in_frame_0___i167 (.Q(\data_in_frame[20] [6]), .C(clk16MHz), 
           .D(n26709));   // verilog/coms.v(128[12] 296[6])
    SB_DFF data_in_frame_0___i168 (.Q(\data_in_frame[20] [7]), .C(clk16MHz), 
           .D(n26710));   // verilog/coms.v(128[12] 296[6])
    SB_DFFE data_in_frame_0___i180 (.Q(\data_in_frame[22] [3]), .C(clk16MHz), 
            .E(VCC_net), .D(n26756));   // verilog/coms.v(128[12] 296[6])
    SB_LUT4 select_715_Select_90_i2_4_lut (.I0(\data_out_frame[11] [2]), .I1(\FRAME_MATCHER.i_31__N_2320 ), 
            .I2(encoder1_position[2]), .I3(\FRAME_MATCHER.state_31__N_2423 [3]), 
            .O(n2_adj_5086));   // verilog/coms.v(146[4] 295[11])
    defparam select_715_Select_90_i2_4_lut.LUT_INIT = 16'hc088;
    SB_DFFR IntegralLimit_i0_i2 (.Q(IntegralLimit[2]), .C(clk16MHz), .D(n26755), 
            .R(reset));   // verilog/coms.v(128[12] 296[6])
    SB_DFFR Kp_i13 (.Q(\Kp[13] ), .C(clk16MHz), .D(n26754), .R(reset));   // verilog/coms.v(128[12] 296[6])
    SB_DFF data_in_frame_0___i92 (.Q(\data_in_frame[11] [3]), .C(clk16MHz), 
           .D(n26130));   // verilog/coms.v(128[12] 296[6])
    SB_DFFE data_in_frame_0___i179 (.Q(\data_in_frame[22] [2]), .C(clk16MHz), 
            .E(VCC_net), .D(n26750));   // verilog/coms.v(128[12] 296[6])
    SB_LUT4 select_715_Select_89_i2_4_lut (.I0(\data_out_frame[11] [1]), .I1(\FRAME_MATCHER.i_31__N_2320 ), 
            .I2(encoder1_position[1]), .I3(\FRAME_MATCHER.state_31__N_2423 [3]), 
            .O(n2_adj_5085));   // verilog/coms.v(146[4] 295[11])
    defparam select_715_Select_89_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i13277_3_lut_4_lut (.I0(Kp_23__N_1583), .I1(n29100), .I2(\data_in_frame[9] [5]), 
            .I3(PWMLimit[13]), .O(n26881));
    defparam i13277_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFFS \FRAME_MATCHER.state_FSM_i9  (.Q(\FRAME_MATCHER.i_31__N_2318 ), 
            .C(clk16MHz), .D(n63712), .S(reset));   // verilog/coms.v(146[4] 295[11])
    SB_DFFR \FRAME_MATCHER.state_FSM_i8  (.Q(\FRAME_MATCHER.i_31__N_2319 ), 
            .C(clk16MHz), .D(n56605), .R(reset));   // verilog/coms.v(146[4] 295[11])
    SB_DFFR \FRAME_MATCHER.state_FSM_i7  (.Q(\FRAME_MATCHER.i_31__N_2320 ), 
            .C(clk16MHz), .D(n1796), .R(reset));   // verilog/coms.v(146[4] 295[11])
    SB_DFFR \FRAME_MATCHER.state_FSM_i6  (.Q(\FRAME_MATCHER.state[3] ), .C(clk16MHz), 
            .D(n1797), .R(reset));   // verilog/coms.v(146[4] 295[11])
    SB_DFFR \FRAME_MATCHER.state_FSM_i5  (.Q(\FRAME_MATCHER.i_31__N_2322 ), 
            .C(clk16MHz), .D(n18192), .R(reset));   // verilog/coms.v(146[4] 295[11])
    SB_DFFR \FRAME_MATCHER.state_FSM_i4  (.Q(\FRAME_MATCHER.i_31__N_2323 ), 
            .C(clk16MHz), .D(n51969), .R(reset));   // verilog/coms.v(146[4] 295[11])
    SB_DFF data_in_frame_0___i169 (.Q(\data_in_frame[21] [0]), .C(clk16MHz), 
           .D(n26713));   // verilog/coms.v(128[12] 296[6])
    SB_DFFR \FRAME_MATCHER.state_FSM_i3  (.Q(\FRAME_MATCHER.i_31__N_2324 ), 
            .C(clk16MHz), .D(n1808), .R(reset));   // verilog/coms.v(146[4] 295[11])
    SB_DFFESS data_out_frame_0___i51 (.Q(\data_out_frame[6] [2]), .C(clk16MHz), 
            .E(n2568), .D(n2_adj_5160), .S(n52688));   // verilog/coms.v(128[12] 296[6])
    SB_DFFR \FRAME_MATCHER.state_FSM_i2  (.Q(\FRAME_MATCHER.i_31__N_2325 ), 
            .C(clk16MHz), .D(n23848), .R(reset));   // verilog/coms.v(146[4] 295[11])
    SB_DFFR \FRAME_MATCHER.i_1939__i0  (.Q(\FRAME_MATCHER.i [0]), .C(clk16MHz), 
            .D(n24764), .R(reset));   // verilog/coms.v(155[12:15])
    SB_DFFESS data_out_frame_0___i52 (.Q(\data_out_frame[6] [3]), .C(clk16MHz), 
            .E(n2568), .D(n2_adj_5161), .S(n52693));   // verilog/coms.v(128[12] 296[6])
    SB_DFFE data_in_frame_0___i178 (.Q(\data_in_frame[22] [1]), .C(clk16MHz), 
            .E(VCC_net), .D(n26746));   // verilog/coms.v(128[12] 296[6])
    SB_DFFE data_in_frame_0___i177 (.Q(\data_in_frame[22] [0]), .C(clk16MHz), 
            .E(VCC_net), .D(n26743));   // verilog/coms.v(128[12] 296[6])
    SB_DFFESS data_out_frame_0___i53 (.Q(\data_out_frame[6] [4]), .C(clk16MHz), 
            .E(n2568), .D(n2_adj_5162), .S(n52692));   // verilog/coms.v(128[12] 296[6])
    SB_DFFE data_in_frame_0___i176 (.Q(\data_in_frame[21] [7]), .C(clk16MHz), 
            .E(VCC_net), .D(n26740));   // verilog/coms.v(128[12] 296[6])
    SB_DFFR IntegralLimit_i0_i3 (.Q(IntegralLimit[3]), .C(clk16MHz), .D(n26739), 
            .R(reset));   // verilog/coms.v(128[12] 296[6])
    SB_DFFR Kp_i14 (.Q(\Kp[14] ), .C(clk16MHz), .D(n26738), .R(reset));   // verilog/coms.v(128[12] 296[6])
    SB_DFFESS data_out_frame_0___i54 (.Q(\data_out_frame[6] [5]), .C(clk16MHz), 
            .E(n2568), .D(n2_adj_5163), .S(n52691));   // verilog/coms.v(128[12] 296[6])
    SB_DFFESS data_out_frame_0___i55 (.Q(\data_out_frame[6] [6]), .C(clk16MHz), 
            .E(n2568), .D(n2_adj_5164), .S(n52690));   // verilog/coms.v(128[12] 296[6])
    SB_LUT4 select_715_Select_88_i2_4_lut (.I0(\data_out_frame[11] [0]), .I1(\FRAME_MATCHER.i_31__N_2320 ), 
            .I2(encoder1_position[0]), .I3(\FRAME_MATCHER.state_31__N_2423 [3]), 
            .O(n2_adj_5084));   // verilog/coms.v(146[4] 295[11])
    defparam select_715_Select_88_i2_4_lut.LUT_INIT = 16'hc088;
    SB_DFFESS data_out_frame_0___i56 (.Q(\data_out_frame[6] [7]), .C(clk16MHz), 
            .E(n2568), .D(n2_adj_5165), .S(n52689));   // verilog/coms.v(128[12] 296[6])
    SB_DFFS IntegralLimit_i0_i4 (.Q(IntegralLimit[4]), .C(clk16MHz), .D(n26737), 
            .S(reset));   // verilog/coms.v(128[12] 296[6])
    SB_LUT4 i13339_3_lut_4_lut (.I0(n35372), .I1(n52895), .I2(rx_data[0]), 
            .I3(\data_in_frame[7] [0]), .O(n26943));
    defparam i13339_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 select_715_Select_87_i2_4_lut (.I0(\data_out_frame[10] [7]), .I1(\FRAME_MATCHER.i_31__N_2320 ), 
            .I2(encoder1_position[15]), .I3(\FRAME_MATCHER.state_31__N_2423 [3]), 
            .O(n2_adj_5083));   // verilog/coms.v(146[4] 295[11])
    defparam select_715_Select_87_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i13342_3_lut_4_lut (.I0(n35372), .I1(n52895), .I2(rx_data[1]), 
            .I3(\data_in_frame[7] [1]), .O(n26946));
    defparam i13342_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 byte_transmit_counter_3__bdd_4_lut (.I0(byte_transmit_counter_c[3]), 
            .I1(n22_adj_5166), .I2(n59919), .I3(byte_transmit_counter_c[4]), 
            .O(n63611));
    defparam byte_transmit_counter_3__bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_LUT4 n63611_bdd_4_lut (.I0(n63611), .I1(n14_adj_5167), .I2(n7_adj_5168), 
            .I3(byte_transmit_counter_c[4]), .O(tx_data[7]));
    defparam n63611_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_48872 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[14] [4]), .I2(\data_out_frame[15] [4]), 
            .I3(byte_transmit_counter_c[1]), .O(n63605));
    defparam byte_transmit_counter_0__bdd_4_lut_48872.LUT_INIT = 16'he4aa;
    SB_LUT4 n63605_bdd_4_lut (.I0(n63605), .I1(\data_out_frame[13] [4]), 
            .I2(\data_out_frame[12] [4]), .I3(byte_transmit_counter_c[1]), 
            .O(n56853));
    defparam n63605_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_CARRY \FRAME_MATCHER.i_1939_add_4_26  (.CI(n46605), .I0(n63273), 
            .I1(\FRAME_MATCHER.i [24]), .CO(n46606));
    SB_LUT4 i13345_3_lut_4_lut (.I0(n35372), .I1(n52895), .I2(rx_data[2]), 
            .I3(\data_in_frame[7] [2]), .O(n26949));
    defparam i13345_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1_4_lut_adj_1165 (.I0(\FRAME_MATCHER.i_31__N_2320 ), .I1(\data_out_frame[10] [6]), 
            .I2(encoder1_position[14]), .I3(\FRAME_MATCHER.state_31__N_2423 [3]), 
            .O(n2_adj_5082));   // verilog/coms.v(146[4] 295[11])
    defparam i1_4_lut_adj_1165.LUT_INIT = 16'ha088;
    SB_LUT4 i13348_3_lut_4_lut (.I0(n35372), .I1(n52895), .I2(rx_data[3]), 
            .I3(\data_in_frame[7] [3]), .O(n26952));
    defparam i13348_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i13351_3_lut_4_lut (.I0(n35372), .I1(n52895), .I2(rx_data[4]), 
            .I3(\data_in_frame[7] [4]), .O(n26955));
    defparam i13351_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFFS IntegralLimit_i0_i5 (.Q(IntegralLimit[5]), .C(clk16MHz), .D(n26736), 
            .S(reset));   // verilog/coms.v(128[12] 296[6])
    SB_LUT4 select_715_Select_85_i2_4_lut (.I0(\data_out_frame[10] [5]), .I1(\FRAME_MATCHER.i_31__N_2320 ), 
            .I2(encoder1_position[13]), .I3(\FRAME_MATCHER.state_31__N_2423 [3]), 
            .O(n2_adj_5081));   // verilog/coms.v(146[4] 295[11])
    defparam select_715_Select_85_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i13354_3_lut_4_lut (.I0(n35372), .I1(n52895), .I2(rx_data[5]), 
            .I3(\data_in_frame[7] [5]), .O(n26958));
    defparam i13354_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i13357_3_lut_4_lut (.I0(n35372), .I1(n52895), .I2(rx_data[6]), 
            .I3(\data_in_frame[7] [6]), .O(n26961));
    defparam i13357_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 select_715_Select_84_i2_4_lut (.I0(\data_out_frame[10] [4]), .I1(\FRAME_MATCHER.i_31__N_2320 ), 
            .I2(encoder1_position[12]), .I3(\FRAME_MATCHER.state_31__N_2423 [3]), 
            .O(n2_adj_5080));   // verilog/coms.v(146[4] 295[11])
    defparam select_715_Select_84_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i13276_3_lut_4_lut (.I0(Kp_23__N_1583), .I1(n29100), .I2(\data_in_frame[9] [6]), 
            .I3(PWMLimit[14]), .O(n26880));
    defparam i13276_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i13275_3_lut_4_lut (.I0(Kp_23__N_1583), .I1(n29100), .I2(\data_in_frame[9] [7]), 
            .I3(PWMLimit[15]), .O(n26879));
    defparam i13275_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1_4_lut_adj_1166 (.I0(\FRAME_MATCHER.i_31__N_2320 ), .I1(\data_out_frame[10] [3]), 
            .I2(encoder1_position[11]), .I3(\FRAME_MATCHER.state_31__N_2423 [3]), 
            .O(n2_adj_5075));   // verilog/coms.v(146[4] 295[11])
    defparam i1_4_lut_adj_1166.LUT_INIT = 16'ha088;
    SB_LUT4 i13360_3_lut_4_lut (.I0(n35372), .I1(n52895), .I2(rx_data[7]), 
            .I3(\data_in_frame[7] [7]), .O(n26964));
    defparam i13360_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 select_715_Select_31_i2_3_lut (.I0(\data_out_frame[3][7] ), .I1(\FRAME_MATCHER.i_31__N_2320 ), 
            .I2(\FRAME_MATCHER.state_31__N_2423 [3]), .I3(GND_net), .O(n2_adj_5070));   // verilog/coms.v(146[4] 295[11])
    defparam select_715_Select_31_i2_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 select_715_Select_30_i2_3_lut (.I0(\data_out_frame[3][6] ), .I1(\FRAME_MATCHER.i_31__N_2320 ), 
            .I2(\FRAME_MATCHER.state_31__N_2423 [3]), .I3(GND_net), .O(n2_adj_5069));   // verilog/coms.v(146[4] 295[11])
    defparam select_715_Select_30_i2_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i13080_3_lut_4_lut (.I0(n25071), .I1(reset), .I2(rx_data[7]), 
            .I3(\data_in_frame[19] [7]), .O(n26684));
    defparam i13080_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13274_3_lut_4_lut (.I0(Kp_23__N_1583), .I1(n29100), .I2(\data_in_frame[8] [0]), 
            .I3(PWMLimit[16]), .O(n26878));
    defparam i13274_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 select_715_Select_28_i2_3_lut (.I0(\data_out_frame[3][4] ), .I1(\FRAME_MATCHER.i_31__N_2320 ), 
            .I2(\FRAME_MATCHER.state_31__N_2423 [3]), .I3(GND_net), .O(n2_adj_5068));   // verilog/coms.v(146[4] 295[11])
    defparam select_715_Select_28_i2_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 \FRAME_MATCHER.i_1939_add_4_25_lut  (.I0(n59813), .I1(n63273), 
            .I2(\FRAME_MATCHER.i [23]), .I3(n46604), .O(n24817)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_1939_add_4_25_lut .LUT_INIT = 16'h8BB8;
    SB_LUT4 select_715_Select_27_i2_3_lut (.I0(\data_out_frame[3][3] ), .I1(\FRAME_MATCHER.i_31__N_2320 ), 
            .I2(\FRAME_MATCHER.state_31__N_2423 [3]), .I3(GND_net), .O(n2_adj_5067));   // verilog/coms.v(146[4] 295[11])
    defparam select_715_Select_27_i2_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i13077_3_lut_4_lut (.I0(n25071), .I1(reset), .I2(rx_data[6]), 
            .I3(\data_in_frame[19] [6]), .O(n26681));
    defparam i13077_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF data_in_frame_0___i93 (.Q(\data_in_frame[11] [4]), .C(clk16MHz), 
           .D(n26133));   // verilog/coms.v(128[12] 296[6])
    SB_CARRY \FRAME_MATCHER.i_1939_add_4_25  (.CI(n46604), .I0(n63273), 
            .I1(\FRAME_MATCHER.i [23]), .CO(n46605));
    SB_LUT4 \FRAME_MATCHER.i_1939_add_4_24_lut  (.I0(n59814), .I1(n63273), 
            .I2(\FRAME_MATCHER.i [22]), .I3(n46603), .O(n24815)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_1939_add_4_24_lut .LUT_INIT = 16'h8BB8;
    SB_CARRY \FRAME_MATCHER.i_1939_add_4_24  (.CI(n46603), .I0(n63273), 
            .I1(\FRAME_MATCHER.i [22]), .CO(n46604));
    SB_LUT4 \FRAME_MATCHER.i_1939_add_4_23_lut  (.I0(n59815), .I1(n63273), 
            .I2(\FRAME_MATCHER.i [21]), .I3(n46602), .O(n24813)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_1939_add_4_23_lut .LUT_INIT = 16'h8BB8;
    SB_CARRY \FRAME_MATCHER.i_1939_add_4_23  (.CI(n46602), .I0(n63273), 
            .I1(\FRAME_MATCHER.i [21]), .CO(n46603));
    SB_LUT4 i13073_3_lut_4_lut (.I0(n25071), .I1(reset), .I2(rx_data[5]), 
            .I3(\data_in_frame[19] [5]), .O(n26677));
    defparam i13073_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFFESS data_out_frame_0___i101 (.Q(\data_out_frame[12] [4]), .C(clk16MHz), 
            .E(n2568), .D(n2_adj_5169), .S(n52729));   // verilog/coms.v(128[12] 296[6])
    SB_DFFESS data_out_frame_0___i102 (.Q(\data_out_frame[12] [5]), .C(clk16MHz), 
            .E(n2568), .D(n2_adj_5170), .S(n52730));   // verilog/coms.v(128[12] 296[6])
    SB_LUT4 i11_4_lut_4_lut (.I0(n25071), .I1(reset), .I2(rx_data[4]), 
            .I3(\data_in_frame[19] [4]), .O(n52233));
    defparam i11_4_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13273_3_lut_4_lut (.I0(Kp_23__N_1583), .I1(n29100), .I2(\data_in_frame[8] [1]), 
            .I3(PWMLimit[17]), .O(n26877));
    defparam i13273_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFFESS data_out_frame_0___i103 (.Q(\data_out_frame[12] [6]), .C(clk16MHz), 
            .E(n2568), .D(n2_adj_5171), .S(n52731));   // verilog/coms.v(128[12] 296[6])
    SB_LUT4 i13272_3_lut_4_lut (.I0(Kp_23__N_1583), .I1(n29100), .I2(\data_in_frame[8] [2]), 
            .I3(PWMLimit[18]), .O(n26876));
    defparam i13272_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i13288_3_lut_4_lut (.I0(Kp_23__N_1583), .I1(n29100), .I2(\data_in_frame[10] [2]), 
            .I3(PWMLimit[2]), .O(n26892));
    defparam i13288_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 select_715_Select_25_i2_3_lut (.I0(\data_out_frame[3][1] ), .I1(\FRAME_MATCHER.i_31__N_2320 ), 
            .I2(\FRAME_MATCHER.state_31__N_2423 [3]), .I3(GND_net), .O(n2_adj_5064));   // verilog/coms.v(146[4] 295[11])
    defparam select_715_Select_25_i2_3_lut.LUT_INIT = 16'hc8c8;
    SB_DFFESS data_out_frame_0___i104 (.Q(\data_out_frame[12] [7]), .C(clk16MHz), 
            .E(n2568), .D(n2_adj_5172), .S(n52732));   // verilog/coms.v(128[12] 296[6])
    SB_DFFESS data_out_frame_0___i105 (.Q(\data_out_frame[13] [0]), .C(clk16MHz), 
            .E(n2568), .D(n2_adj_5173), .S(n52733));   // verilog/coms.v(128[12] 296[6])
    SB_DFFESS data_out_frame_0___i106 (.Q(\data_out_frame[13] [1]), .C(clk16MHz), 
            .E(n2568), .D(n2_adj_5174), .S(n52680));   // verilog/coms.v(128[12] 296[6])
    SB_LUT4 \FRAME_MATCHER.i_1939_add_4_22_lut  (.I0(n59816), .I1(n63273), 
            .I2(\FRAME_MATCHER.i [20]), .I3(n46601), .O(n24811)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_1939_add_4_22_lut .LUT_INIT = 16'h8BB8;
    SB_DFFESS data_out_frame_0___i107 (.Q(\data_out_frame[13] [2]), .C(clk16MHz), 
            .E(n2568), .D(n2_adj_5175), .S(n52734));   // verilog/coms.v(128[12] 296[6])
    SB_DFFESS data_out_frame_0___i108 (.Q(\data_out_frame[13] [3]), .C(clk16MHz), 
            .E(n2568), .D(n2_adj_5176), .S(n52735));   // verilog/coms.v(128[12] 296[6])
    SB_DFFE data_in_frame_0___i175 (.Q(\data_in_frame[21] [6]), .C(clk16MHz), 
            .E(VCC_net), .D(n26732));   // verilog/coms.v(128[12] 296[6])
    SB_CARRY \FRAME_MATCHER.i_1939_add_4_22  (.CI(n46601), .I0(n63273), 
            .I1(\FRAME_MATCHER.i [20]), .CO(n46602));
    SB_LUT4 \FRAME_MATCHER.i_1939_add_4_21_lut  (.I0(n59829), .I1(n63273), 
            .I2(\FRAME_MATCHER.i [19]), .I3(n46600), .O(n24809)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_1939_add_4_21_lut .LUT_INIT = 16'h8BB8;
    SB_DFFE data_in_frame_0___i174 (.Q(\data_in_frame[21] [5]), .C(clk16MHz), 
            .E(VCC_net), .D(n26729));   // verilog/coms.v(128[12] 296[6])
    SB_LUT4 i13287_3_lut_4_lut (.I0(Kp_23__N_1583), .I1(n29100), .I2(\data_in_frame[10] [3]), 
            .I3(PWMLimit[3]), .O(n26891));
    defparam i13287_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i13271_3_lut_4_lut (.I0(Kp_23__N_1583), .I1(n29100), .I2(\data_in_frame[8] [3]), 
            .I3(PWMLimit[19]), .O(n26875));
    defparam i13271_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_CARRY \FRAME_MATCHER.i_1939_add_4_21  (.CI(n46600), .I0(n63273), 
            .I1(\FRAME_MATCHER.i [19]), .CO(n46601));
    SB_LUT4 \FRAME_MATCHER.i_1939_add_4_20_lut  (.I0(n59838), .I1(n63273), 
            .I2(\FRAME_MATCHER.i [18]), .I3(n46599), .O(n24807)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_1939_add_4_20_lut .LUT_INIT = 16'h8BB8;
    SB_LUT4 i13067_3_lut_4_lut (.I0(n25071), .I1(reset), .I2(rx_data[3]), 
            .I3(\data_in_frame[19] [3]), .O(n26671));
    defparam i13067_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13270_3_lut_4_lut (.I0(Kp_23__N_1583), .I1(n29100), .I2(\data_in_frame[8] [4]), 
            .I3(PWMLimit[20]), .O(n26874));
    defparam i13270_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i13015_3_lut_4_lut (.I0(n25077), .I1(reset), .I2(rx_data[3]), 
            .I3(\data_in_frame[17] [3]), .O(n26619));
    defparam i13015_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_CARRY \FRAME_MATCHER.i_1939_add_4_20  (.CI(n46599), .I0(n63273), 
            .I1(\FRAME_MATCHER.i [18]), .CO(n46600));
    SB_LUT4 \FRAME_MATCHER.i_1939_add_4_19_lut  (.I0(n59840), .I1(n63273), 
            .I2(\FRAME_MATCHER.i [17]), .I3(n46598), .O(n24805)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_1939_add_4_19_lut .LUT_INIT = 16'h8BB8;
    SB_CARRY \FRAME_MATCHER.i_1939_add_4_19  (.CI(n46598), .I0(n63273), 
            .I1(\FRAME_MATCHER.i [17]), .CO(n46599));
    SB_LUT4 \FRAME_MATCHER.i_1939_add_4_18_lut  (.I0(n59841), .I1(n63273), 
            .I2(\FRAME_MATCHER.i [16]), .I3(n46597), .O(n24803)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_1939_add_4_18_lut .LUT_INIT = 16'h8BB8;
    SB_DFFR Kp_i15 (.Q(\Kp[15] ), .C(clk16MHz), .D(n26728), .R(reset));   // verilog/coms.v(128[12] 296[6])
    SB_CARRY \FRAME_MATCHER.i_1939_add_4_18  (.CI(n46597), .I0(n63273), 
            .I1(\FRAME_MATCHER.i [16]), .CO(n46598));
    SB_LUT4 i13061_3_lut_4_lut (.I0(n25071), .I1(reset), .I2(rx_data[2]), 
            .I3(\data_in_frame[19] [2]), .O(n26665));
    defparam i13061_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 \FRAME_MATCHER.i_1939_add_4_17_lut  (.I0(n59844), .I1(n63273), 
            .I2(\FRAME_MATCHER.i [15]), .I3(n46596), .O(n24801)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_1939_add_4_17_lut .LUT_INIT = 16'h8BB8;
    SB_LUT4 i12752_3_lut_4_lut (.I0(Kp_23__N_1583), .I1(n29100), .I2(\data_in_frame[5] [1]), 
            .I3(\Ki[1] ), .O(n26356));
    defparam i12752_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_CARRY \FRAME_MATCHER.i_1939_add_4_17  (.CI(n46596), .I0(n63273), 
            .I1(\FRAME_MATCHER.i [15]), .CO(n46597));
    SB_LUT4 \FRAME_MATCHER.i_1939_add_4_16_lut  (.I0(n59845), .I1(n63273), 
            .I2(\FRAME_MATCHER.i [14]), .I3(n46595), .O(n24799)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_1939_add_4_16_lut .LUT_INIT = 16'h8BB8;
    SB_CARRY \FRAME_MATCHER.i_1939_add_4_16  (.CI(n46595), .I0(n63273), 
            .I1(\FRAME_MATCHER.i [14]), .CO(n46596));
    SB_LUT4 \FRAME_MATCHER.i_1939_add_4_15_lut  (.I0(n59846), .I1(n63273), 
            .I2(\FRAME_MATCHER.i [13]), .I3(n46594), .O(n24797)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_1939_add_4_15_lut .LUT_INIT = 16'h8BB8;
    SB_DFFE data_in_frame_0___i173 (.Q(\data_in_frame[21] [4]), .C(clk16MHz), 
            .E(VCC_net), .D(n26725));   // verilog/coms.v(128[12] 296[6])
    SB_DFFE data_in_frame_0___i172 (.Q(\data_in_frame[21] [3]), .C(clk16MHz), 
            .E(VCC_net), .D(n26722));   // verilog/coms.v(128[12] 296[6])
    SB_CARRY \FRAME_MATCHER.i_1939_add_4_15  (.CI(n46594), .I0(n63273), 
            .I1(\FRAME_MATCHER.i [13]), .CO(n46595));
    SB_DFFE data_in_frame_0___i171 (.Q(\data_in_frame[21] [2]), .C(clk16MHz), 
            .E(VCC_net), .D(n26719));   // verilog/coms.v(128[12] 296[6])
    SB_LUT4 \FRAME_MATCHER.i_1939_add_4_14_lut  (.I0(n59847), .I1(n63273), 
            .I2(\FRAME_MATCHER.i [12]), .I3(n46593), .O(n24795)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_1939_add_4_14_lut .LUT_INIT = 16'h8BB8;
    SB_CARRY \FRAME_MATCHER.i_1939_add_4_14  (.CI(n46593), .I0(n63273), 
            .I1(\FRAME_MATCHER.i [12]), .CO(n46594));
    SB_LUT4 \FRAME_MATCHER.i_1939_add_4_13_lut  (.I0(n59848), .I1(n63273), 
            .I2(\FRAME_MATCHER.i [11]), .I3(n46592), .O(n24793)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_1939_add_4_13_lut .LUT_INIT = 16'h8BB8;
    SB_LUT4 i13058_3_lut_4_lut (.I0(n25071), .I1(reset), .I2(rx_data[1]), 
            .I3(\data_in_frame[19] [1]), .O(n26662));
    defparam i13058_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFFESS data_out_frame_0___i109 (.Q(\data_out_frame[13] [4]), .C(clk16MHz), 
            .E(n2568), .D(n2_adj_5177), .S(n52736));   // verilog/coms.v(128[12] 296[6])
    SB_DFFESS data_out_frame_0___i110 (.Q(\data_out_frame[13] [5]), .C(clk16MHz), 
            .E(n2568), .D(n2_adj_5178), .S(n52737));   // verilog/coms.v(128[12] 296[6])
    SB_DFFESS data_out_frame_0___i111 (.Q(\data_out_frame[13] [6]), .C(clk16MHz), 
            .E(n2568), .D(n2_adj_5179), .S(n52738));   // verilog/coms.v(128[12] 296[6])
    SB_DFFESS data_out_frame_0___i112 (.Q(\data_out_frame[13] [7]), .C(clk16MHz), 
            .E(n2568), .D(n2_adj_5180), .S(n52739));   // verilog/coms.v(128[12] 296[6])
    SB_DFFESS data_out_frame_0___i113 (.Q(\data_out_frame[14] [0]), .C(clk16MHz), 
            .E(n2568), .D(n2_adj_5181), .S(n52740));   // verilog/coms.v(128[12] 296[6])
    SB_DFFESS data_out_frame_0___i114 (.Q(\data_out_frame[14] [1]), .C(clk16MHz), 
            .E(n2568), .D(n2_adj_5182), .S(n52741));   // verilog/coms.v(128[12] 296[6])
    SB_DFFESS data_out_frame_0___i115 (.Q(\data_out_frame[14] [2]), .C(clk16MHz), 
            .E(n2568), .D(n2_adj_5183), .S(n25663));   // verilog/coms.v(128[12] 296[6])
    SB_CARRY \FRAME_MATCHER.i_1939_add_4_13  (.CI(n46592), .I0(n63273), 
            .I1(\FRAME_MATCHER.i [11]), .CO(n46593));
    SB_LUT4 i11_3_lut_4_lut (.I0(n25071), .I1(reset), .I2(\data_in_frame[19] [0]), 
            .I3(rx_data[0]), .O(n52199));
    defparam i11_3_lut_4_lut.LUT_INIT = 16'hf1e0;
    SB_LUT4 \FRAME_MATCHER.i_1939_add_4_12_lut  (.I0(n59849), .I1(n63273), 
            .I2(\FRAME_MATCHER.i [10]), .I3(n46591), .O(n24791)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_1939_add_4_12_lut .LUT_INIT = 16'h8BB8;
    SB_DFFESS data_out_frame_0___i116 (.Q(\data_out_frame[14] [3]), .C(clk16MHz), 
            .E(n2568), .D(n2_adj_5184), .S(n52742));   // verilog/coms.v(128[12] 296[6])
    SB_DFFESS data_out_frame_0___i117 (.Q(\data_out_frame[14] [4]), .C(clk16MHz), 
            .E(n2568), .D(n2_adj_5185), .S(n52743));   // verilog/coms.v(128[12] 296[6])
    SB_DFFESS data_out_frame_0___i118 (.Q(\data_out_frame[14] [5]), .C(clk16MHz), 
            .E(n2568), .D(n2_adj_5186), .S(n52744));   // verilog/coms.v(128[12] 296[6])
    SB_DFFESS data_out_frame_0___i119 (.Q(\data_out_frame[14] [6]), .C(clk16MHz), 
            .E(n2568), .D(n2_adj_5187), .S(n52745));   // verilog/coms.v(128[12] 296[6])
    SB_DFFESS data_out_frame_0___i120 (.Q(\data_out_frame[14] [7]), .C(clk16MHz), 
            .E(n2568), .D(n2_adj_5188), .S(n52746));   // verilog/coms.v(128[12] 296[6])
    SB_DFFESS data_out_frame_0___i121 (.Q(\data_out_frame[15] [0]), .C(clk16MHz), 
            .E(n2568), .D(n2_adj_5189), .S(n52747));   // verilog/coms.v(128[12] 296[6])
    SB_DFFESS data_out_frame_0___i122 (.Q(\data_out_frame[15] [1]), .C(clk16MHz), 
            .E(n2568), .D(n2_adj_5190), .S(n52748));   // verilog/coms.v(128[12] 296[6])
    SB_DFFESS data_out_frame_0___i123 (.Q(\data_out_frame[15] [2]), .C(clk16MHz), 
            .E(n2568), .D(n2_adj_5191), .S(n52749));   // verilog/coms.v(128[12] 296[6])
    SB_DFFESS data_out_frame_0___i124 (.Q(\data_out_frame[15] [3]), .C(clk16MHz), 
            .E(n2568), .D(n2_adj_5192), .S(n52750));   // verilog/coms.v(128[12] 296[6])
    SB_DFFESS data_out_frame_0___i125 (.Q(\data_out_frame[15] [4]), .C(clk16MHz), 
            .E(n2568), .D(n2_adj_5193), .S(n52751));   // verilog/coms.v(128[12] 296[6])
    SB_DFFESS data_out_frame_0___i126 (.Q(\data_out_frame[15] [5]), .C(clk16MHz), 
            .E(n2568), .D(n2_adj_5194), .S(n52752));   // verilog/coms.v(128[12] 296[6])
    SB_CARRY \FRAME_MATCHER.i_1939_add_4_12  (.CI(n46591), .I0(n63273), 
            .I1(\FRAME_MATCHER.i [10]), .CO(n46592));
    SB_DFFESS data_out_frame_0___i127 (.Q(\data_out_frame[15] [6]), .C(clk16MHz), 
            .E(n2568), .D(n2_adj_5195), .S(n52753));   // verilog/coms.v(128[12] 296[6])
    SB_DFFESS data_out_frame_0___i128 (.Q(\data_out_frame[15] [7]), .C(clk16MHz), 
            .E(n2568), .D(n2_adj_5196), .S(n52754));   // verilog/coms.v(128[12] 296[6])
    SB_DFFESS data_out_frame_0___i129 (.Q(\data_out_frame[16] [0]), .C(clk16MHz), 
            .E(n2568), .D(n2_adj_5197), .S(n52755));   // verilog/coms.v(128[12] 296[6])
    SB_DFFESS data_out_frame_0___i130 (.Q(\data_out_frame[16] [1]), .C(clk16MHz), 
            .E(n2568), .D(n2_adj_5198), .S(n52756));   // verilog/coms.v(128[12] 296[6])
    SB_LUT4 \FRAME_MATCHER.i_1939_add_4_11_lut  (.I0(n59850), .I1(n63273), 
            .I2(\FRAME_MATCHER.i [9]), .I3(n46590), .O(n24789)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_1939_add_4_11_lut .LUT_INIT = 16'h8BB8;
    SB_DFFESS data_out_frame_0___i131 (.Q(\data_out_frame[16] [2]), .C(clk16MHz), 
            .E(n2568), .D(n2_adj_5199), .S(n52757));   // verilog/coms.v(128[12] 296[6])
    SB_DFFE data_in_frame_0___i170 (.Q(\data_in_frame[21] [1]), .C(clk16MHz), 
            .E(VCC_net), .D(n26716));   // verilog/coms.v(128[12] 296[6])
    SB_LUT4 i12751_3_lut_4_lut (.I0(Kp_23__N_1583), .I1(n29100), .I2(\data_in_frame[5] [2]), 
            .I3(\Ki[2] ), .O(n26355));
    defparam i12751_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_CARRY \FRAME_MATCHER.i_1939_add_4_11  (.CI(n46590), .I0(n63273), 
            .I1(\FRAME_MATCHER.i [9]), .CO(n46591));
    SB_LUT4 \FRAME_MATCHER.i_1939_add_4_10_lut  (.I0(n59853), .I1(n63273), 
            .I2(\FRAME_MATCHER.i [8]), .I3(n46589), .O(n24787)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_1939_add_4_10_lut .LUT_INIT = 16'h8BB8;
    SB_CARRY \FRAME_MATCHER.i_1939_add_4_10  (.CI(n46589), .I0(n63273), 
            .I1(\FRAME_MATCHER.i [8]), .CO(n46590));
    SB_LUT4 \FRAME_MATCHER.i_1939_add_4_9_lut  (.I0(n59855), .I1(n63273), 
            .I2(\FRAME_MATCHER.i [7]), .I3(n46588), .O(n24785)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_1939_add_4_9_lut .LUT_INIT = 16'h8BB8;
    SB_CARRY \FRAME_MATCHER.i_1939_add_4_9  (.CI(n46588), .I0(n63273), .I1(\FRAME_MATCHER.i [7]), 
            .CO(n46589));
    SB_DFFESS data_out_frame_0___i132 (.Q(\data_out_frame[16] [3]), .C(clk16MHz), 
            .E(n2568), .D(n2_adj_5200), .S(n52758));   // verilog/coms.v(128[12] 296[6])
    SB_LUT4 \FRAME_MATCHER.i_1939_add_4_8_lut  (.I0(n59856), .I1(n63273), 
            .I2(\FRAME_MATCHER.i [6]), .I3(n46587), .O(n24783)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_1939_add_4_8_lut .LUT_INIT = 16'h8BB8;
    SB_CARRY \FRAME_MATCHER.i_1939_add_4_8  (.CI(n46587), .I0(n63273), .I1(\FRAME_MATCHER.i [6]), 
            .CO(n46588));
    SB_LUT4 \FRAME_MATCHER.i_1939_add_4_7_lut  (.I0(n59857), .I1(n63273), 
            .I2(\FRAME_MATCHER.i [5]), .I3(n46586), .O(n24781)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_1939_add_4_7_lut .LUT_INIT = 16'h8BB8;
    SB_CARRY \FRAME_MATCHER.i_1939_add_4_7  (.CI(n46586), .I0(n63273), .I1(\FRAME_MATCHER.i [5]), 
            .CO(n46587));
    SB_LUT4 \FRAME_MATCHER.i_1939_add_4_6_lut  (.I0(n59862), .I1(n63273), 
            .I2(\FRAME_MATCHER.i [4]), .I3(n46585), .O(n24779)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_1939_add_4_6_lut .LUT_INIT = 16'h8BB8;
    SB_CARRY \FRAME_MATCHER.i_1939_add_4_6  (.CI(n46585), .I0(n63273), .I1(\FRAME_MATCHER.i [4]), 
            .CO(n46586));
    SB_LUT4 \FRAME_MATCHER.i_1939_add_4_5_lut  (.I0(n59869), .I1(n63273), 
            .I2(\FRAME_MATCHER.i [3]), .I3(n46584), .O(n24777)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_1939_add_4_5_lut .LUT_INIT = 16'h8BB8;
    SB_CARRY \FRAME_MATCHER.i_1939_add_4_5  (.CI(n46584), .I0(n63273), .I1(\FRAME_MATCHER.i [3]), 
            .CO(n46585));
    SB_LUT4 \FRAME_MATCHER.i_1939_add_4_4_lut  (.I0(n59870), .I1(n63273), 
            .I2(\FRAME_MATCHER.i [2]), .I3(n46583), .O(n24775)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_1939_add_4_4_lut .LUT_INIT = 16'h8BB8;
    SB_CARRY \FRAME_MATCHER.i_1939_add_4_4  (.CI(n46583), .I0(n63273), .I1(\FRAME_MATCHER.i [2]), 
            .CO(n46584));
    SB_LUT4 \FRAME_MATCHER.i_1939_add_4_3_lut  (.I0(n59871), .I1(n63273), 
            .I2(\FRAME_MATCHER.i [1]), .I3(n46582), .O(n24773)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_1939_add_4_3_lut .LUT_INIT = 16'h8BB8;
    SB_CARRY \FRAME_MATCHER.i_1939_add_4_3  (.CI(n46582), .I0(n63273), .I1(\FRAME_MATCHER.i [1]), 
            .CO(n46583));
    SB_LUT4 \FRAME_MATCHER.i_1939_add_4_2_lut  (.I0(GND_net), .I1(n161), 
            .I2(\FRAME_MATCHER.i [0]), .I3(GND_net), .O(n133[0])) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_1939_add_4_2_lut .LUT_INIT = 16'hC33C;
    SB_LUT4 i1_2_lut_3_lut_adj_1167 (.I0(\control_mode[0] ), .I1(n22431), 
            .I2(\control_mode[1] ), .I3(GND_net), .O(n15));   // verilog/coms.v(128[12] 296[6])
    defparam i1_2_lut_3_lut_adj_1167.LUT_INIT = 16'hfdfd;
    SB_CARRY \FRAME_MATCHER.i_1939_add_4_2  (.CI(GND_net), .I0(n161), .I1(\FRAME_MATCHER.i [0]), 
            .CO(n46582));
    SB_LUT4 i21853_3_lut_4_lut (.I0(\control_mode[0] ), .I1(n22431), .I2(control_update), 
            .I3(\control_mode[1] ), .O(n24502));   // verilog/coms.v(128[12] 296[6])
    defparam i21853_3_lut_4_lut.LUT_INIT = 16'hd0f0;
    SB_LUT4 i12730_3_lut_4_lut (.I0(n8_adj_5202), .I1(n52895), .I2(rx_data[4]), 
            .I3(\data_in_frame[5] [4]), .O(n26334));
    defparam i12730_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_2_lut_adj_1168 (.I0(n53495), .I1(n53521), .I2(GND_net), 
            .I3(GND_net), .O(n7_adj_5203));
    defparam i2_2_lut_adj_1168.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1169 (.I0(n7_adj_5203), .I1(n53492), .I2(n48923), 
            .I3(n53246), .O(n54876));
    defparam i4_4_lut_adj_1169.LUT_INIT = 16'h9669;
    SB_LUT4 i2_3_lut_adj_1170 (.I0(\data_in_frame[20] [4]), .I1(\data_in_frame[20] [3]), 
            .I2(n55195), .I3(GND_net), .O(n52980));
    defparam i2_3_lut_adj_1170.LUT_INIT = 16'h6969;
    SB_LUT4 i12750_3_lut_4_lut (.I0(Kp_23__N_1583), .I1(n29100), .I2(\data_in_frame[5] [3]), 
            .I3(\Ki[3] ), .O(n26354));
    defparam i12750_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFFESS data_out_frame_0___i133 (.Q(\data_out_frame[16] [4]), .C(clk16MHz), 
            .E(n2568), .D(n2_adj_5204), .S(n25620));   // verilog/coms.v(128[12] 296[6])
    SB_DFFESS data_out_frame_0___i134 (.Q(\data_out_frame[16] [5]), .C(clk16MHz), 
            .E(n2568), .D(n2_adj_5205), .S(n52759));   // verilog/coms.v(128[12] 296[6])
    SB_DFFESS data_out_frame_0___i135 (.Q(\data_out_frame[16] [6]), .C(clk16MHz), 
            .E(n2568), .D(n2_adj_5206), .S(n52760));   // verilog/coms.v(128[12] 296[6])
    SB_LUT4 i1_2_lut_adj_1171 (.I0(\data_in_frame[18] [3]), .I1(\data_in_frame[18] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n22677));
    defparam i1_2_lut_adj_1171.LUT_INIT = 16'h6666;
    SB_DFFESS data_out_frame_0___i136 (.Q(\data_out_frame[16] [7]), .C(clk16MHz), 
            .E(n2568), .D(n2_adj_5207), .S(n52761));   // verilog/coms.v(128[12] 296[6])
    SB_LUT4 i20_4_lut (.I0(n47932), .I1(n53163), .I2(n53321), .I3(\data_in_frame[16] [7]), 
            .O(n52));
    defparam i20_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i18_4_lut (.I0(n52921), .I1(\data_in_frame[18][7] ), .I2(n52995), 
            .I3(n22631), .O(n50));
    defparam i18_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i19_4_lut (.I0(n22623), .I1(n53264), .I2(\data_in_frame[15] [4]), 
            .I3(n48511), .O(n51));
    defparam i19_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i17_4_lut (.I0(\data_in_frame[18] [1]), .I1(\data_in_frame[20] [7]), 
            .I2(\data_in_frame[16] [3]), .I3(n22677), .O(n49));
    defparam i17_4_lut.LUT_INIT = 16'h6996;
    SB_DFFESS data_out_frame_0___i137 (.Q(\data_out_frame[17] [0]), .C(clk16MHz), 
            .E(n2568), .D(n2_adj_5208), .S(n52762));   // verilog/coms.v(128[12] 296[6])
    SB_DFF data_in_frame_0___i94 (.Q(\data_in_frame[11] [5]), .C(clk16MHz), 
           .D(n26136));   // verilog/coms.v(128[12] 296[6])
    SB_DFFR IntegralLimit_i0_i6 (.Q(IntegralLimit[6]), .C(clk16MHz), .D(n26705), 
            .R(reset));   // verilog/coms.v(128[12] 296[6])
    SB_LUT4 i24_4_lut (.I0(Kp_23__N_1224), .I1(n48800), .I2(n47783), .I3(\data_in_frame[21] [7]), 
            .O(n56));
    defparam i24_4_lut.LUT_INIT = 16'h9669;
    SB_LUT4 i22_4_lut (.I0(n53298), .I1(n52940), .I2(n53249), .I3(Kp_23__N_902), 
            .O(n54));
    defparam i22_4_lut.LUT_INIT = 16'h6996;
    SB_DFFESS data_out_frame_0___i138 (.Q(\data_out_frame[17] [1]), .C(clk16MHz), 
            .E(n2568), .D(n2_adj_5209), .S(n52763));   // verilog/coms.v(128[12] 296[6])
    SB_LUT4 i12749_3_lut_4_lut (.I0(Kp_23__N_1583), .I1(n29100), .I2(\data_in_frame[5] [4]), 
            .I3(\Ki[4] ), .O(n26353));
    defparam i12749_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i23_4_lut (.I0(n48783), .I1(\data_in_frame[15] [1]), .I2(\data_in_frame[15] [6]), 
            .I3(\data_in_frame[10] [6]), .O(n55));
    defparam i23_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i21_4_lut (.I0(n47756), .I1(n48785), .I2(\data_in_frame[16] [5]), 
            .I3(n53512), .O(n53));
    defparam i21_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i30_4_lut (.I0(n53), .I1(n55), .I2(n54), .I3(n56), .O(n62));
    defparam i30_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i29_4_lut (.I0(n49), .I1(n51), .I2(n50), .I3(n52), .O(n61));
    defparam i29_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1172 (.I0(\data_in_frame[20] [1]), .I1(n61), .I2(\data_in_frame[20] [2]), 
            .I3(n62), .O(n22_adj_5210));
    defparam i1_4_lut_adj_1172.LUT_INIT = 16'h6996;
    SB_LUT4 i7_3_lut (.I0(n53556), .I1(\data_in_frame[19] [7]), .I2(\data_in_frame[19] [5]), 
            .I3(GND_net), .O(n28));
    defparam i7_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 i15_4_lut (.I0(n53409), .I1(n53222), .I2(n53234), .I3(n53079), 
            .O(n36));
    defparam i15_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i13_4_lut_adj_1173 (.I0(n53583), .I1(n26_adj_5211), .I2(\data_in_frame[19] [6]), 
            .I3(\data_in_frame[21] [6]), .O(n34_c));
    defparam i13_4_lut_adj_1173.LUT_INIT = 16'h6996;
    SB_LUT4 i16_4_lut (.I0(n52980), .I1(\data_in_frame[21] [2]), .I2(\data_in_frame[15] [7]), 
            .I3(n22_adj_5210), .O(n37));
    defparam i16_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i12727_3_lut_4_lut (.I0(n8_adj_5202), .I1(n52895), .I2(rx_data[3]), 
            .I3(\data_in_frame[5] [3]), .O(n26331));
    defparam i12727_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i18_4_lut_adj_1174 (.I0(\data_in_frame[20] [0]), .I1(n36), .I2(n28), 
            .I3(n53598), .O(n39));
    defparam i18_4_lut_adj_1174.LUT_INIT = 16'h6996;
    SB_LUT4 i12724_3_lut_4_lut (.I0(n8_adj_5202), .I1(n52895), .I2(rx_data[2]), 
            .I3(\data_in_frame[5] [2]), .O(n26328));
    defparam i12724_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i20_4_lut_adj_1175 (.I0(n39), .I1(n37), .I2(n33_adj_5212), 
            .I3(n34_c), .O(n48923));
    defparam i20_4_lut_adj_1175.LUT_INIT = 16'h6996;
    SB_LUT4 i5_4_lut_adj_1176 (.I0(n48295), .I1(n47898), .I2(n48794), 
            .I3(\data_in_frame[20] [7]), .O(n12_adj_5213));
    defparam i5_4_lut_adj_1176.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_1177 (.I0(n22056), .I1(n12_adj_5213), .I2(n53489), 
            .I3(\data_in_frame[18] [5]), .O(n53240));
    defparam i6_4_lut_adj_1177.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1178 (.I0(\data_in_frame[21] [7]), .I1(n48785), 
            .I2(GND_net), .I3(GND_net), .O(n53228));
    defparam i1_2_lut_adj_1178.LUT_INIT = 16'h6666;
    SB_LUT4 i3_3_lut_adj_1179 (.I0(\data_in_frame[16] [5]), .I1(n23039), 
            .I2(\data_in_frame[16] [6]), .I3(GND_net), .O(n47932));
    defparam i3_3_lut_adj_1179.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_adj_1180 (.I0(\data_in_frame[19] [1]), .I1(n55031), 
            .I2(n47932), .I3(GND_net), .O(n53492));
    defparam i2_3_lut_adj_1180.LUT_INIT = 16'h6969;
    SB_LUT4 i12712_3_lut_4_lut (.I0(n8_adj_5202), .I1(n52895), .I2(rx_data[1]), 
            .I3(\data_in_frame[5] [1]), .O(n26316));
    defparam i12712_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i12693_3_lut_4_lut (.I0(n8_adj_5202), .I1(n52895), .I2(rx_data[0]), 
            .I3(\data_in_frame[5] [0]), .O(n26297));
    defparam i12693_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i3_4_lut_adj_1181 (.I0(\data_in_frame[17] [3]), .I1(n53370), 
            .I2(n53366), .I3(n47764), .O(n53583));
    defparam i3_4_lut_adj_1181.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1182 (.I0(\data_in_frame[13] [4]), .I1(n53091), 
            .I2(GND_net), .I3(GND_net), .O(n47849));   // verilog/coms.v(86[17:63])
    defparam i1_2_lut_adj_1182.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_1183 (.I0(n47849), .I1(n53583), .I2(n53529), 
            .I3(n23402), .O(n23006));
    defparam i3_4_lut_adj_1183.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1184 (.I0(n23006), .I1(n48781), .I2(GND_net), 
            .I3(GND_net), .O(n48800));
    defparam i1_2_lut_adj_1184.LUT_INIT = 16'h9999;
    SB_LUT4 i1_2_lut_adj_1185 (.I0(\data_in_frame[17] [0]), .I1(\data_in_frame[17] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n53264));
    defparam i1_2_lut_adj_1185.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1186 (.I0(\data_in_frame[15] [1]), .I1(\data_in_frame[14] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n53366));
    defparam i1_2_lut_adj_1186.LUT_INIT = 16'h6666;
    SB_LUT4 i12748_3_lut_4_lut (.I0(Kp_23__N_1583), .I1(n29100), .I2(\data_in_frame[5] [5]), 
            .I3(\Ki[5] ), .O(n26352));
    defparam i12748_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i12914_3_lut_4_lut (.I0(n8_adj_5202), .I1(n52895), .I2(rx_data[5]), 
            .I3(\data_in_frame[5] [5]), .O(n26518));
    defparam i12914_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i4_2_lut (.I0(\data_in_frame[14] [6]), .I1(n53532), .I2(GND_net), 
            .I3(GND_net), .O(n18_adj_5214));
    defparam i4_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i10_4_lut_adj_1187 (.I0(\data_in_frame[14] [7]), .I1(n48942), 
            .I2(n48511), .I3(n52952), .O(n24_adj_5215));
    defparam i10_4_lut_adj_1187.LUT_INIT = 16'h6996;
    SB_LUT4 i8_4_lut_adj_1188 (.I0(\data_in_frame[17] [2]), .I1(n53375), 
            .I2(n52937), .I3(\data_in_frame[12] [6]), .O(n22_adj_5216));
    defparam i8_4_lut_adj_1188.LUT_INIT = 16'h6996;
    SB_LUT4 i12_4_lut_adj_1189 (.I0(n53468), .I1(n24_adj_5215), .I2(n18_adj_5214), 
            .I3(n53366), .O(n26_adj_5217));
    defparam i12_4_lut_adj_1189.LUT_INIT = 16'h6996;
    SB_LUT4 i13_4_lut_adj_1190 (.I0(n22822), .I1(n26_adj_5217), .I2(n22_adj_5216), 
            .I3(n23002), .O(n48781));
    defparam i13_4_lut_adj_1190.LUT_INIT = 16'h6996;
    SB_LUT4 i1_3_lut (.I0(\data_in_frame[19] [3]), .I1(n48781), .I2(n53329), 
            .I3(GND_net), .O(n48904));
    defparam i1_3_lut.LUT_INIT = 16'h6969;
    SB_LUT4 i4_4_lut_adj_1191 (.I0(n52946), .I1(\data_in_frame[14] [7]), 
            .I2(\data_in_frame[16] [7]), .I3(n53375), .O(n10_adj_5218));   // verilog/coms.v(72[16:27])
    defparam i4_4_lut_adj_1191.LUT_INIT = 16'h6996;
    SB_LUT4 i5_3_lut_adj_1192 (.I0(n54710), .I1(n10_adj_5218), .I2(\data_in_frame[14] [5]), 
            .I3(GND_net), .O(n22042));   // verilog/coms.v(72[16:27])
    defparam i5_3_lut_adj_1192.LUT_INIT = 16'h6969;
    SB_LUT4 i1_2_lut_adj_1193 (.I0(\data_in_frame[21] [5]), .I1(n48904), 
            .I2(GND_net), .I3(GND_net), .O(n53015));
    defparam i1_2_lut_adj_1193.LUT_INIT = 16'h9999;
    SB_LUT4 i4_4_lut_adj_1194 (.I0(n47882), .I1(n48904), .I2(n53264), 
            .I3(\data_in_frame[19] [2]), .O(n10_adj_5219));
    defparam i4_4_lut_adj_1194.LUT_INIT = 16'h9669;
    SB_LUT4 i12917_3_lut_4_lut (.I0(n8_adj_5202), .I1(n52895), .I2(rx_data[6]), 
            .I3(\data_in_frame[5] [6]), .O(n26521));
    defparam i12917_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i5_3_lut_adj_1195 (.I0(n22042), .I1(n10_adj_5219), .I2(n48844), 
            .I3(GND_net), .O(n53409));
    defparam i5_3_lut_adj_1195.LUT_INIT = 16'h9696;
    SB_LUT4 i12920_3_lut_4_lut (.I0(n8_adj_5202), .I1(n52895), .I2(rx_data[7]), 
            .I3(\data_in_frame[5] [7]), .O(n26524));
    defparam i12920_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_1196 (.I0(\data_in_frame[18] [2]), .I1(\data_in_frame[18] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n22631));
    defparam i1_2_lut_adj_1196.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_1197 (.I0(n22056), .I1(\data_in_frame[17] [0]), 
            .I2(\data_in_frame[19] [0]), .I3(GND_net), .O(n53246));
    defparam i2_3_lut_adj_1197.LUT_INIT = 16'h9696;
    SB_LUT4 equal_292_i8_2_lut_3_lut (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(\FRAME_MATCHER.i [0]), .I3(GND_net), .O(n8_adj_5202));   // verilog/coms.v(154[7:23])
    defparam equal_292_i8_2_lut_3_lut.LUT_INIT = 16'hbfbf;
    SB_LUT4 i2_3_lut_adj_1198 (.I0(\data_in_frame[9] [7]), .I1(n53147), 
            .I2(n48768), .I3(GND_net), .O(n54710));
    defparam i2_3_lut_adj_1198.LUT_INIT = 16'h9696;
    SB_LUT4 equal_293_i8_2_lut_3_lut (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(\FRAME_MATCHER.i [0]), .I3(GND_net), .O(n8_adj_5220));   // verilog/coms.v(154[7:23])
    defparam equal_293_i8_2_lut_3_lut.LUT_INIT = 16'hfbfb;
    SB_LUT4 i3_4_lut_adj_1199 (.I0(\data_in_frame[14] [5]), .I1(n54710), 
            .I2(n53363), .I3(n52937), .O(n47783));
    defparam i3_4_lut_adj_1199.LUT_INIT = 16'h9669;
    SB_LUT4 i2_3_lut_adj_1200 (.I0(\data_in_frame[16] [6]), .I1(n53085), 
            .I2(n48813), .I3(GND_net), .O(n48844));
    defparam i2_3_lut_adj_1200.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1201 (.I0(n22898), .I1(n23343), .I2(GND_net), 
            .I3(GND_net), .O(n53468));
    defparam i1_2_lut_adj_1201.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_1202 (.I0(n53171), .I1(\data_in_frame[14] [6]), 
            .I2(\data_in_frame[16] [7]), .I3(n53468), .O(n53085));
    defparam i3_4_lut_adj_1202.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1203 (.I0(\data_in_frame[18][7] ), .I1(n48844), 
            .I2(n47783), .I3(GND_net), .O(n55031));
    defparam i2_3_lut_adj_1203.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1204 (.I0(n55031), .I1(n53085), .I2(GND_net), 
            .I3(GND_net), .O(n48295));   // verilog/coms.v(71[16:69])
    defparam i1_2_lut_adj_1204.LUT_INIT = 16'h9999;
    SB_LUT4 i1_2_lut_adj_1205 (.I0(n48798), .I1(n48392), .I2(GND_net), 
            .I3(GND_net), .O(n48783));
    defparam i1_2_lut_adj_1205.LUT_INIT = 16'h9999;
    SB_LUT4 i12747_3_lut_4_lut (.I0(Kp_23__N_1583), .I1(n29100), .I2(\data_in_frame[5] [6]), 
            .I3(\Ki[6] ), .O(n26351));
    defparam i12747_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i3_4_lut_adj_1206 (.I0(n48783), .I1(n53348), .I2(\data_in_frame[20] [6]), 
            .I3(\data_in_frame[19] [0]), .O(n53521));
    defparam i3_4_lut_adj_1206.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1207 (.I0(\data_in_frame[18] [5]), .I1(n53252), 
            .I2(\data_in_frame[21] [0]), .I3(\data_in_frame[18] [4]), .O(n53495));
    defparam i3_4_lut_adj_1207.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1208 (.I0(\data_in_frame[21] [1]), .I1(n53521), 
            .I2(GND_net), .I3(GND_net), .O(n53222));
    defparam i1_2_lut_adj_1208.LUT_INIT = 16'h6666;
    SB_LUT4 data_in_frame_17__7__I_0_4027_2_lut (.I0(\data_in_frame[17] [7]), 
            .I1(\data_in_frame[17] [6]), .I2(GND_net), .I3(GND_net), .O(Kp_23__N_1224));   // verilog/coms.v(71[16:27])
    defparam data_in_frame_17__7__I_0_4027_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i13269_3_lut_4_lut (.I0(Kp_23__N_1583), .I1(n29100), .I2(\data_in_frame[8] [5]), 
            .I3(PWMLimit[21]), .O(n26873));
    defparam i13269_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4_4_lut_adj_1209 (.I0(n7_adj_5221), .I1(n53079), .I2(n54891), 
            .I3(Kp_23__N_1224), .O(n53276));   // verilog/coms.v(77[16:43])
    defparam i4_4_lut_adj_1209.LUT_INIT = 16'h9669;
    SB_LUT4 i13268_3_lut_4_lut (.I0(Kp_23__N_1583), .I1(n29100), .I2(\data_in_frame[8] [6]), 
            .I3(PWMLimit[22]), .O(n26872));
    defparam i13268_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_48673 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[14] [6]), .I2(\data_out_frame[15] [6]), 
            .I3(byte_transmit_counter_c[1]), .O(n63383));
    defparam byte_transmit_counter_0__bdd_4_lut_48673.LUT_INIT = 16'he4aa;
    SB_LUT4 i3_4_lut_adj_1210 (.I0(\data_in_frame[13] [2]), .I1(\data_in_frame[15] [2]), 
            .I2(\data_in_frame[12] [7]), .I3(\data_in_frame[12] [6]), .O(n52921));   // verilog/coms.v(77[16:43])
    defparam i3_4_lut_adj_1210.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1211 (.I0(n23509), .I1(n53352), .I2(n52921), 
            .I3(\data_in_frame[13] [0]), .O(n47764));   // verilog/coms.v(77[16:43])
    defparam i3_4_lut_adj_1211.LUT_INIT = 16'h6996;
    SB_DFFESS data_out_frame_0___i139 (.Q(\data_out_frame[17] [2]), .C(clk16MHz), 
            .E(n2568), .D(n2_adj_5222), .S(n52764));   // verilog/coms.v(128[12] 296[6])
    SB_DFFESS data_out_frame_0___i140 (.Q(\data_out_frame[17] [3]), .C(clk16MHz), 
            .E(n2568), .D(n2_adj_5223), .S(n52765));   // verilog/coms.v(128[12] 296[6])
    SB_DFFESS data_out_frame_0___i141 (.Q(\data_out_frame[17] [4]), .C(clk16MHz), 
            .E(n2568), .D(n2_adj_5224), .S(n52766));   // verilog/coms.v(128[12] 296[6])
    SB_DFFESS data_out_frame_0___i142 (.Q(\data_out_frame[17] [5]), .C(clk16MHz), 
            .E(n2568), .D(n2_adj_5225), .S(n52776));   // verilog/coms.v(128[12] 296[6])
    SB_DFFESS data_out_frame_0___i143 (.Q(\data_out_frame[17] [6]), .C(clk16MHz), 
            .E(n2568), .D(n2_adj_5226), .S(n52767));   // verilog/coms.v(128[12] 296[6])
    SB_DFFESS data_out_frame_0___i144 (.Q(\data_out_frame[17] [7]), .C(clk16MHz), 
            .E(n2568), .D(n2_adj_5227), .S(n52710));   // verilog/coms.v(128[12] 296[6])
    SB_LUT4 i1_2_lut_adj_1212 (.I0(\data_in_frame[15] [7]), .I1(\data_in_frame[16] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n53321));   // verilog/coms.v(86[17:28])
    defparam i1_2_lut_adj_1212.LUT_INIT = 16'h6666;
    SB_DFFESS data_out_frame_0___i169 (.Q(\data_out_frame[21] [0]), .C(clk16MHz), 
            .E(n2568), .D(n2_adj_5228), .S(n52769));   // verilog/coms.v(128[12] 296[6])
    SB_DFFESS data_out_frame_0___i170 (.Q(\data_out_frame[21] [1]), .C(clk16MHz), 
            .E(n2568), .D(n2_adj_5229), .S(n52770));   // verilog/coms.v(128[12] 296[6])
    SB_DFFESS data_out_frame_0___i171 (.Q(\data_out_frame[21] [2]), .C(clk16MHz), 
            .E(n2568), .D(n2_adj_5230), .S(n52771));   // verilog/coms.v(128[12] 296[6])
    SB_DFFESS data_out_frame_0___i172 (.Q(\data_out_frame[21] [3]), .C(clk16MHz), 
            .E(n2568), .D(n2_adj_5231), .S(n52772));   // verilog/coms.v(128[12] 296[6])
    SB_DFFESS data_out_frame_0___i173 (.Q(\data_out_frame[21] [4]), .C(clk16MHz), 
            .E(n2568), .D(n2_adj_5232), .S(n52773));   // verilog/coms.v(128[12] 296[6])
    SB_DFFESS data_out_frame_0___i174 (.Q(\data_out_frame[21] [5]), .C(clk16MHz), 
            .E(n2568), .D(n2_adj_5233), .S(n52774));   // verilog/coms.v(128[12] 296[6])
    SB_DFFESS data_out_frame_0___i175 (.Q(\data_out_frame[21] [6]), .C(clk16MHz), 
            .E(n2568), .D(n2_adj_5234), .S(n52777));   // verilog/coms.v(128[12] 296[6])
    SB_DFFESS data_out_frame_0___i176 (.Q(\data_out_frame[21] [7]), .C(clk16MHz), 
            .E(n2568), .D(n2_adj_5235), .S(n52778));   // verilog/coms.v(128[12] 296[6])
    SB_DFFESS data_out_frame_0___i177 (.Q(\data_out_frame[22] [0]), .C(clk16MHz), 
            .E(n2568), .D(n2_adj_5236), .S(n52779));   // verilog/coms.v(128[12] 296[6])
    SB_DFFESS data_out_frame_0___i178 (.Q(\data_out_frame[22] [1]), .C(clk16MHz), 
            .E(n2568), .D(n2_adj_5237), .S(n52780));   // verilog/coms.v(128[12] 296[6])
    SB_DFFESS data_out_frame_0___i179 (.Q(\data_out_frame[22] [2]), .C(clk16MHz), 
            .E(n2568), .D(n2_adj_5238), .S(n52781));   // verilog/coms.v(128[12] 296[6])
    SB_DFFESS data_out_frame_0___i180 (.Q(\data_out_frame[22] [3]), .C(clk16MHz), 
            .E(n2568), .D(n2_adj_5239), .S(n52782));   // verilog/coms.v(128[12] 296[6])
    SB_DFFESS data_out_frame_0___i181 (.Q(\data_out_frame[22] [4]), .C(clk16MHz), 
            .E(n2568), .D(n2_adj_5240), .S(n52783));   // verilog/coms.v(128[12] 296[6])
    SB_DFFESS data_out_frame_0___i182 (.Q(\data_out_frame[22] [5]), .C(clk16MHz), 
            .E(n2568), .D(n2_adj_5241), .S(n52775));   // verilog/coms.v(128[12] 296[6])
    SB_DFFESS data_out_frame_0___i183 (.Q(\data_out_frame[22] [6]), .C(clk16MHz), 
            .E(n2568), .D(n2_adj_5242), .S(n52795));   // verilog/coms.v(128[12] 296[6])
    SB_DFFESS data_out_frame_0___i184 (.Q(\data_out_frame[22] [7]), .C(clk16MHz), 
            .E(n2568), .D(n2_adj_5243), .S(n52786));   // verilog/coms.v(128[12] 296[6])
    SB_DFFESS tx_transmit_4000 (.Q(r_SM_Main_2__N_3318[0]), .C(clk16MHz), 
            .E(n2568), .D(n1_adj_5244), .S(n25577));   // verilog/coms.v(128[12] 296[6])
    SB_LUT4 i2_3_lut_adj_1213 (.I0(\data_in_frame[16] [1]), .I1(n53163), 
            .I2(\data_in_frame[13] [7]), .I3(GND_net), .O(n53556));
    defparam i2_3_lut_adj_1213.LUT_INIT = 16'h9696;
    SB_DFFESS driver_enable_4003 (.Q(DE_c), .C(clk16MHz), .E(n2568), .D(n23764), 
            .S(n25576));   // verilog/coms.v(128[12] 296[6])
    SB_LUT4 i1_2_lut_adj_1214 (.I0(\data_in_frame[13] [5]), .I1(\data_in_frame[13] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n53577));   // verilog/coms.v(86[17:28])
    defparam i1_2_lut_adj_1214.LUT_INIT = 16'h6666;
    SB_LUT4 i12517_3_lut_4_lut (.I0(n8_adj_5139), .I1(n52895), .I2(rx_data[7]), 
            .I3(\data_in_frame[0] [7]), .O(n26121));
    defparam i12517_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFFESS byte_transmit_counter_i0_i0 (.Q(byte_transmit_counter[0]), .C(clk16MHz), 
            .E(n2568), .D(n1_adj_5245), .S(n52666));   // verilog/coms.v(128[12] 296[6])
    SB_LUT4 i12514_3_lut_4_lut (.I0(n8_adj_5139), .I1(n52895), .I2(rx_data[6]), 
            .I3(\data_in_frame[0] [6]), .O(n26118));
    defparam i12514_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i12511_3_lut_4_lut (.I0(n8_adj_5139), .I1(n52895), .I2(rx_data[5]), 
            .I3(\data_in_frame[0] [5]), .O(n26115));
    defparam i12511_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF data_in_0___i1 (.Q(\data_in[0] [0]), .C(clk16MHz), .D(n26101));   // verilog/coms.v(128[12] 296[6])
    SB_LUT4 i12508_3_lut_4_lut (.I0(n8_adj_5139), .I1(n52895), .I2(rx_data[4]), 
            .I3(\data_in_frame[0] [4]), .O(n26112));
    defparam i12508_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i12504_3_lut_4_lut (.I0(n8_adj_5139), .I1(n52895), .I2(rx_data[3]), 
            .I3(\data_in_frame[0] [3]), .O(n26108));
    defparam i12504_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i12501_3_lut_4_lut (.I0(n8_adj_5139), .I1(n52895), .I2(rx_data[2]), 
            .I3(\data_in_frame[0] [2]), .O(n26105));
    defparam i12501_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i12498_3_lut_4_lut (.I0(n8_adj_5139), .I1(n52895), .I2(rx_data[1]), 
            .I3(\data_in_frame[0] [1]), .O(n26102));
    defparam i12498_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13238_3_lut_4_lut (.I0(n8_adj_5139), .I1(n52895), .I2(rx_data[0]), 
            .I3(\data_in_frame[0] [0]), .O(n26842));
    defparam i13238_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13011_3_lut_4_lut (.I0(n25077), .I1(reset), .I2(rx_data[2]), 
            .I3(\data_in_frame[17] [2]), .O(n26615));
    defparam i13011_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13267_3_lut_4_lut (.I0(Kp_23__N_1583), .I1(n29100), .I2(\data_in_frame[8] [7]), 
            .I3(PWMLimit[23]), .O(n26871));
    defparam i13267_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i11_4_lut_4_lut_adj_1215 (.I0(n25077), .I1(reset), .I2(rx_data[1]), 
            .I3(\data_in_frame[17] [1]), .O(n52181));
    defparam i11_4_lut_4_lut_adj_1215.LUT_INIT = 16'hfe10;
    SB_LUT4 i12746_3_lut_4_lut (.I0(Kp_23__N_1583), .I1(n29100), .I2(\data_in_frame[5] [7]), 
            .I3(\Ki[7] ), .O(n26350));
    defparam i12746_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4_4_lut_adj_1216 (.I0(n23402), .I1(\data_in_frame[16] [0]), 
            .I2(n53556), .I3(n6_adj_5246), .O(n20730));
    defparam i4_4_lut_adj_1216.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_1217 (.I0(n53509), .I1(n22837), .I2(\data_in_frame[15] [5]), 
            .I3(n53577), .O(n10_adj_5247));   // verilog/coms.v(86[17:28])
    defparam i4_4_lut_adj_1217.LUT_INIT = 16'h6996;
    SB_DFFR IntegralLimit_i0_i7 (.Q(IntegralLimit[7]), .C(clk16MHz), .D(n26680), 
            .R(reset));   // verilog/coms.v(128[12] 296[6])
    SB_DFF data_in_frame_0___i95 (.Q(\data_in_frame[11] [6]), .C(clk16MHz), 
           .D(n26139));   // verilog/coms.v(128[12] 296[6])
    SB_DFF data_in_frame_0___i96 (.Q(\data_in_frame[11] [7]), .C(clk16MHz), 
           .D(n26142));   // verilog/coms.v(128[12] 296[6])
    SB_DFFR IntegralLimit_i0_i8 (.Q(IntegralLimit[8]), .C(clk16MHz), .D(n26661), 
            .R(reset));   // verilog/coms.v(128[12] 296[6])
    SB_LUT4 i1_2_lut_adj_1218 (.I0(\data_in_frame[13] [3]), .I1(\data_in_frame[13] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n22837));   // verilog/coms.v(86[17:63])
    defparam i1_2_lut_adj_1218.LUT_INIT = 16'h6666;
    SB_LUT4 i12745_3_lut_4_lut (.I0(Kp_23__N_1583), .I1(n29100), .I2(\data_in_frame[4] [0]), 
            .I3(\Ki[8] ), .O(n26349));
    defparam i12745_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFFR \FRAME_MATCHER.i_1939__i1  (.Q(\FRAME_MATCHER.i [1]), .C(clk16MHz), 
            .D(n24773), .R(reset));   // verilog/coms.v(155[12:15])
    SB_DFFESS data_out_frame_0___i57 (.Q(\data_out_frame[7] [0]), .C(clk16MHz), 
            .E(n2568), .D(n2_adj_5248), .S(n52700));   // verilog/coms.v(128[12] 296[6])
    SB_DFFESS data_out_frame_0___i58 (.Q(\data_out_frame[7] [1]), .C(clk16MHz), 
            .E(n2568), .D(n2_adj_5249), .S(n52701));   // verilog/coms.v(128[12] 296[6])
    SB_DFFESS data_out_frame_0___i59 (.Q(\data_out_frame[7] [2]), .C(clk16MHz), 
            .E(n2568), .D(n2_adj_5250), .S(n52793));   // verilog/coms.v(128[12] 296[6])
    SB_DFFESS data_out_frame_0___i60 (.Q(\data_out_frame[7] [3]), .C(clk16MHz), 
            .E(n2568), .D(n2_adj_5251), .S(n52792));   // verilog/coms.v(128[12] 296[6])
    SB_DFFESS data_out_frame_0___i61 (.Q(\data_out_frame[7] [4]), .C(clk16MHz), 
            .E(n2568), .D(n2_adj_5252), .S(n52784));   // verilog/coms.v(128[12] 296[6])
    SB_DFFESS data_out_frame_0___i62 (.Q(\data_out_frame[7] [5]), .C(clk16MHz), 
            .E(n2568), .D(n2_adj_5253), .S(n52785));   // verilog/coms.v(128[12] 296[6])
    SB_DFFESS data_out_frame_0___i63 (.Q(\data_out_frame[7] [6]), .C(clk16MHz), 
            .E(n2568), .D(n2_adj_5254), .S(n52787));   // verilog/coms.v(128[12] 296[6])
    SB_DFFESS data_out_frame_0___i64 (.Q(\data_out_frame[7] [7]), .C(clk16MHz), 
            .E(n2568), .D(n2_adj_5255), .S(n52788));   // verilog/coms.v(128[12] 296[6])
    SB_DFFESS data_out_frame_0___i65 (.Q(\data_out_frame[8] [0]), .C(clk16MHz), 
            .E(n2568), .D(n2_adj_5256), .S(n52790));   // verilog/coms.v(128[12] 296[6])
    SB_DFFESS data_out_frame_0___i66 (.Q(\data_out_frame[8] [1]), .C(clk16MHz), 
            .E(n2568), .D(n2_adj_5257), .S(n52794));   // verilog/coms.v(128[12] 296[6])
    SB_DFFESS data_out_frame_0___i67 (.Q(\data_out_frame[8] [2]), .C(clk16MHz), 
            .E(n2568), .D(n2_adj_5258), .S(n52791));   // verilog/coms.v(128[12] 296[6])
    SB_DFFESS data_out_frame_0___i68 (.Q(\data_out_frame[8] [3]), .C(clk16MHz), 
            .E(n2568), .D(n2_adj_5259), .S(n52694));   // verilog/coms.v(128[12] 296[6])
    SB_DFFESS data_out_frame_0___i69 (.Q(\data_out_frame[8] [4]), .C(clk16MHz), 
            .E(n2568), .D(n2_adj_5260), .S(n52695));   // verilog/coms.v(128[12] 296[6])
    SB_DFFESS data_out_frame_0___i70 (.Q(\data_out_frame[8] [5]), .C(clk16MHz), 
            .E(n2568), .D(n2_adj_5261), .S(n52696));   // verilog/coms.v(128[12] 296[6])
    SB_DFFESS data_out_frame_0___i71 (.Q(\data_out_frame[8] [6]), .C(clk16MHz), 
            .E(n2568), .D(n2_adj_5262), .S(n52697));   // verilog/coms.v(128[12] 296[6])
    SB_DFFESS data_out_frame_0___i72 (.Q(\data_out_frame[8] [7]), .C(clk16MHz), 
            .E(n2568), .D(n2_adj_5263), .S(n52698));   // verilog/coms.v(128[12] 296[6])
    SB_DFFESS data_out_frame_0___i73 (.Q(\data_out_frame[9] [0]), .C(clk16MHz), 
            .E(n2568), .D(n2_adj_5264), .S(n52699));   // verilog/coms.v(128[12] 296[6])
    SB_DFFESS data_out_frame_0___i74 (.Q(\data_out_frame[9] [1]), .C(clk16MHz), 
            .E(n2568), .D(n2_adj_5265), .S(n52702));   // verilog/coms.v(128[12] 296[6])
    SB_DFFESS data_out_frame_0___i75 (.Q(\data_out_frame[9] [2]), .C(clk16MHz), 
            .E(n2568), .D(n2_adj_5266), .S(n52703));   // verilog/coms.v(128[12] 296[6])
    SB_DFFESS data_out_frame_0___i76 (.Q(\data_out_frame[9] [3]), .C(clk16MHz), 
            .E(n2568), .D(n2_adj_5267), .S(n52704));   // verilog/coms.v(128[12] 296[6])
    SB_DFFESS data_out_frame_0___i77 (.Q(\data_out_frame[9] [4]), .C(clk16MHz), 
            .E(n2568), .D(n2_adj_5268), .S(n52705));   // verilog/coms.v(128[12] 296[6])
    SB_DFFESS data_out_frame_0___i78 (.Q(\data_out_frame[9] [5]), .C(clk16MHz), 
            .E(n2568), .D(n2_adj_5269), .S(n52706));   // verilog/coms.v(128[12] 296[6])
    SB_DFFESS data_out_frame_0___i79 (.Q(\data_out_frame[9] [6]), .C(clk16MHz), 
            .E(n2568), .D(n2_adj_5270), .S(n52707));   // verilog/coms.v(128[12] 296[6])
    SB_DFFESS data_out_frame_0___i80 (.Q(\data_out_frame[9] [7]), .C(clk16MHz), 
            .E(n2568), .D(n2_adj_5271), .S(n52708));   // verilog/coms.v(128[12] 296[6])
    SB_DFFESS data_out_frame_0___i81 (.Q(\data_out_frame[10] [0]), .C(clk16MHz), 
            .E(n2568), .D(n2_adj_5272), .S(n52709));   // verilog/coms.v(128[12] 296[6])
    SB_DFFESS data_out_frame_0___i82 (.Q(\data_out_frame[10] [1]), .C(clk16MHz), 
            .E(n2568), .D(n2_adj_5273), .S(n52711));   // verilog/coms.v(128[12] 296[6])
    SB_DFFR \FRAME_MATCHER.i_1939__i2  (.Q(\FRAME_MATCHER.i [2]), .C(clk16MHz), 
            .D(n24775), .R(reset));   // verilog/coms.v(155[12:15])
    SB_DFFR \FRAME_MATCHER.i_1939__i3  (.Q(\FRAME_MATCHER.i [3]), .C(clk16MHz), 
            .D(n24777), .R(reset));   // verilog/coms.v(155[12:15])
    SB_DFFR \FRAME_MATCHER.i_1939__i4  (.Q(\FRAME_MATCHER.i [4]), .C(clk16MHz), 
            .D(n24779), .R(reset));   // verilog/coms.v(155[12:15])
    SB_DFFR \FRAME_MATCHER.i_1939__i5  (.Q(\FRAME_MATCHER.i [5]), .C(clk16MHz), 
            .D(n24781), .R(reset));   // verilog/coms.v(155[12:15])
    SB_DFFR \FRAME_MATCHER.i_1939__i6  (.Q(\FRAME_MATCHER.i [6]), .C(clk16MHz), 
            .D(n24783), .R(reset));   // verilog/coms.v(155[12:15])
    SB_DFFR \FRAME_MATCHER.i_1939__i7  (.Q(\FRAME_MATCHER.i [7]), .C(clk16MHz), 
            .D(n24785), .R(reset));   // verilog/coms.v(155[12:15])
    SB_DFFR \FRAME_MATCHER.i_1939__i8  (.Q(\FRAME_MATCHER.i [8]), .C(clk16MHz), 
            .D(n24787), .R(reset));   // verilog/coms.v(155[12:15])
    SB_DFFR \FRAME_MATCHER.i_1939__i9  (.Q(\FRAME_MATCHER.i [9]), .C(clk16MHz), 
            .D(n24789), .R(reset));   // verilog/coms.v(155[12:15])
    SB_DFFR \FRAME_MATCHER.i_1939__i10  (.Q(\FRAME_MATCHER.i [10]), .C(clk16MHz), 
            .D(n24791), .R(reset));   // verilog/coms.v(155[12:15])
    SB_DFFR \FRAME_MATCHER.i_1939__i11  (.Q(\FRAME_MATCHER.i [11]), .C(clk16MHz), 
            .D(n24793), .R(reset));   // verilog/coms.v(155[12:15])
    SB_DFFR \FRAME_MATCHER.i_1939__i12  (.Q(\FRAME_MATCHER.i [12]), .C(clk16MHz), 
            .D(n24795), .R(reset));   // verilog/coms.v(155[12:15])
    SB_DFFR \FRAME_MATCHER.i_1939__i13  (.Q(\FRAME_MATCHER.i [13]), .C(clk16MHz), 
            .D(n24797), .R(reset));   // verilog/coms.v(155[12:15])
    SB_DFFR \FRAME_MATCHER.i_1939__i14  (.Q(\FRAME_MATCHER.i [14]), .C(clk16MHz), 
            .D(n24799), .R(reset));   // verilog/coms.v(155[12:15])
    SB_DFFR \FRAME_MATCHER.i_1939__i15  (.Q(\FRAME_MATCHER.i [15]), .C(clk16MHz), 
            .D(n24801), .R(reset));   // verilog/coms.v(155[12:15])
    SB_DFFR \FRAME_MATCHER.i_1939__i16  (.Q(\FRAME_MATCHER.i [16]), .C(clk16MHz), 
            .D(n24803), .R(reset));   // verilog/coms.v(155[12:15])
    SB_DFFR \FRAME_MATCHER.i_1939__i17  (.Q(\FRAME_MATCHER.i [17]), .C(clk16MHz), 
            .D(n24805), .R(reset));   // verilog/coms.v(155[12:15])
    SB_DFFR \FRAME_MATCHER.i_1939__i18  (.Q(\FRAME_MATCHER.i [18]), .C(clk16MHz), 
            .D(n24807), .R(reset));   // verilog/coms.v(155[12:15])
    SB_DFFR \FRAME_MATCHER.i_1939__i19  (.Q(\FRAME_MATCHER.i [19]), .C(clk16MHz), 
            .D(n24809), .R(reset));   // verilog/coms.v(155[12:15])
    SB_DFFR \FRAME_MATCHER.i_1939__i20  (.Q(\FRAME_MATCHER.i [20]), .C(clk16MHz), 
            .D(n24811), .R(reset));   // verilog/coms.v(155[12:15])
    SB_DFFR \FRAME_MATCHER.i_1939__i21  (.Q(\FRAME_MATCHER.i [21]), .C(clk16MHz), 
            .D(n24813), .R(reset));   // verilog/coms.v(155[12:15])
    SB_DFFR \FRAME_MATCHER.i_1939__i22  (.Q(\FRAME_MATCHER.i [22]), .C(clk16MHz), 
            .D(n24815), .R(reset));   // verilog/coms.v(155[12:15])
    SB_DFFR \FRAME_MATCHER.i_1939__i23  (.Q(\FRAME_MATCHER.i [23]), .C(clk16MHz), 
            .D(n24817), .R(reset));   // verilog/coms.v(155[12:15])
    SB_DFFR \FRAME_MATCHER.i_1939__i24  (.Q(\FRAME_MATCHER.i [24]), .C(clk16MHz), 
            .D(n24819), .R(reset));   // verilog/coms.v(155[12:15])
    SB_DFFR \FRAME_MATCHER.i_1939__i25  (.Q(\FRAME_MATCHER.i [25]), .C(clk16MHz), 
            .D(n24821), .R(reset));   // verilog/coms.v(155[12:15])
    SB_DFFR \FRAME_MATCHER.i_1939__i26  (.Q(\FRAME_MATCHER.i [26]), .C(clk16MHz), 
            .D(n24823), .R(reset));   // verilog/coms.v(155[12:15])
    SB_DFFR \FRAME_MATCHER.i_1939__i27  (.Q(\FRAME_MATCHER.i [27]), .C(clk16MHz), 
            .D(n24825), .R(reset));   // verilog/coms.v(155[12:15])
    SB_DFFR \FRAME_MATCHER.i_1939__i28  (.Q(\FRAME_MATCHER.i [28]), .C(clk16MHz), 
            .D(n24827), .R(reset));   // verilog/coms.v(155[12:15])
    SB_DFFR \FRAME_MATCHER.i_1939__i29  (.Q(\FRAME_MATCHER.i [29]), .C(clk16MHz), 
            .D(n24829), .R(reset));   // verilog/coms.v(155[12:15])
    SB_DFFR \FRAME_MATCHER.i_1939__i30  (.Q(\FRAME_MATCHER.i [30]), .C(clk16MHz), 
            .D(n24831), .R(reset));   // verilog/coms.v(155[12:15])
    SB_DFFR \FRAME_MATCHER.i_1939__i31  (.Q(\FRAME_MATCHER.i [31]), .C(clk16MHz), 
            .D(n24833), .R(reset));   // verilog/coms.v(155[12:15])
    SB_LUT4 i1_2_lut_adj_1219 (.I0(\data_in_frame[10] [1]), .I1(\data_in_frame[12] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n53363));
    defparam i1_2_lut_adj_1219.LUT_INIT = 16'h6666;
    SB_DFF data_in_frame_0___i97 (.Q(\data_in_frame[12] [0]), .C(clk16MHz), 
           .D(n26145));   // verilog/coms.v(128[12] 296[6])
    SB_LUT4 i12744_3_lut_4_lut (.I0(Kp_23__N_1583), .I1(n29100), .I2(\data_in_frame[4] [1]), 
            .I3(\Ki[9] ), .O(n26348));
    defparam i12744_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1_2_lut_adj_1220 (.I0(\data_in_frame[12] [5]), .I1(\data_in_frame[12] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n53171));
    defparam i1_2_lut_adj_1220.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_1221 (.I0(n53171), .I1(n53363), .I2(\data_in_frame[12] [6]), 
            .I3(GND_net), .O(n52946));   // verilog/coms.v(72[16:27])
    defparam i2_3_lut_adj_1221.LUT_INIT = 16'h9696;
    SB_DFFR Kp_i6 (.Q(\Kp[6] ), .C(clk16MHz), .D(n26086), .R(reset));   // verilog/coms.v(128[12] 296[6])
    SB_DFFR PWMLimit_i0_i0 (.Q(PWMLimit[0]), .C(clk16MHz), .D(n26084), 
            .R(reset));   // verilog/coms.v(128[12] 296[6])
    SB_DFF current_limit_i0_i0 (.Q(current_limit[0]), .C(clk16MHz), .D(n26083));   // verilog/coms.v(128[12] 296[6])
    SB_DFF control_mode_i0_i0 (.Q(\control_mode[0] ), .C(clk16MHz), .D(n26082));   // verilog/coms.v(128[12] 296[6])
    SB_DFFR Ki_i0 (.Q(\Ki[0] ), .C(clk16MHz), .D(n26081), .R(reset));   // verilog/coms.v(128[12] 296[6])
    SB_LUT4 i2_3_lut_adj_1222 (.I0(n3_adj_5274), .I1(n23288), .I2(\data_in_frame[10] [4]), 
            .I3(GND_net), .O(n22898));   // verilog/coms.v(75[16:43])
    defparam i2_3_lut_adj_1222.LUT_INIT = 16'h9696;
    SB_LUT4 i13193_3_lut_4_lut (.I0(n35372), .I1(n52890), .I2(rx_data[0]), 
            .I3(\data_in_frame[23] [0]), .O(n26797));
    defparam i13193_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i13196_3_lut_4_lut (.I0(n35372), .I1(n52890), .I2(rx_data[1]), 
            .I3(\data_in_frame[23] [1]), .O(n26800));
    defparam i13196_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i20_4_lut_adj_1223 (.I0(\data_in_frame[3] [4]), .I1(\data_in_frame[10] [3]), 
            .I2(\data_in_frame[10] [6]), .I3(\data_in_frame[9] [5]), .O(n48));
    defparam i20_4_lut_adj_1223.LUT_INIT = 16'h6996;
    SB_LUT4 i18_4_lut_adj_1224 (.I0(\data_in_frame[7] [6]), .I1(n53607), 
            .I2(\data_in_frame[11] [2]), .I3(n53592), .O(n46));
    defparam i18_4_lut_adj_1224.LUT_INIT = 16'h6996;
    SB_DFFR IntegralLimit_i0_i9 (.Q(IntegralLimit[9]), .C(clk16MHz), .D(n26608), 
            .R(reset));   // verilog/coms.v(128[12] 296[6])
    SB_DFFR IntegralLimit_i0_i10 (.Q(IntegralLimit[10]), .C(clk16MHz), .D(n26592), 
            .R(reset));   // verilog/coms.v(128[12] 296[6])
    SB_LUT4 i19_4_lut_adj_1225 (.I0(n53553), .I1(n53125), .I2(n53288), 
            .I3(n52946), .O(n47_c));
    defparam i19_4_lut_adj_1225.LUT_INIT = 16'h6996;
    SB_LUT4 i13200_3_lut_4_lut (.I0(n35372), .I1(n52890), .I2(rx_data[2]), 
            .I3(\data_in_frame[23] [2]), .O(n26804));
    defparam i13200_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i17_4_lut_adj_1226 (.I0(n53430), .I1(\data_in_frame[10] [5]), 
            .I2(n53034), .I3(\data_in_frame[10] [7]), .O(n45));
    defparam i17_4_lut_adj_1226.LUT_INIT = 16'h6996;
    SB_LUT4 i16_4_lut_adj_1227 (.I0(n53285), .I1(\data_in_frame[11] [4]), 
            .I2(\data_in_frame[10] [4]), .I3(n53595), .O(n44));
    defparam i16_4_lut_adj_1227.LUT_INIT = 16'h6996;
    SB_LUT4 i11_3_lut_4_lut_adj_1228 (.I0(n25077), .I1(reset), .I2(\data_in_frame[17] [0]), 
            .I3(rx_data[0]), .O(n52163));
    defparam i11_3_lut_4_lut_adj_1228.LUT_INIT = 16'hf1e0;
    SB_DFF data_in_frame_0___i98 (.Q(\data_in_frame[12] [1]), .C(clk16MHz), 
           .D(n26148));   // verilog/coms.v(128[12] 296[6])
    SB_DFF data_in_frame_0___i99 (.Q(\data_in_frame[12] [2]), .C(clk16MHz), 
           .D(n26151));   // verilog/coms.v(128[12] 296[6])
    SB_DFFR IntegralLimit_i0_i11 (.Q(IntegralLimit[11]), .C(clk16MHz), .D(n26589), 
            .R(reset));   // verilog/coms.v(128[12] 296[6])
    SB_DFF data_in_frame_0___i100 (.Q(\data_in_frame[12] [3]), .C(clk16MHz), 
           .D(n26154));   // verilog/coms.v(128[12] 296[6])
    SB_DFFR IntegralLimit_i0_i12 (.Q(IntegralLimit[12]), .C(clk16MHz), .D(n26583), 
            .R(reset));   // verilog/coms.v(128[12] 296[6])
    SB_LUT4 i15_4_lut_adj_1229 (.I0(n53571), .I1(\data_in_frame[1][4] ), 
            .I2(\data_in_frame[11] [1]), .I3(\data_in_frame[12] [0]), .O(n43));
    defparam i15_4_lut_adj_1229.LUT_INIT = 16'h6996;
    SB_LUT4 i26_4_lut (.I0(n45), .I1(n47_c), .I2(n46), .I3(n48), .O(n54_adj_5275));
    defparam i26_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i21_4_lut_adj_1230 (.I0(n48415), .I1(\data_in_frame[11] [7]), 
            .I2(\data_in_frame[11] [0]), .I3(\data_in_frame[12] [7]), .O(n49_adj_5276));
    defparam i21_4_lut_adj_1230.LUT_INIT = 16'h6996;
    SB_LUT4 i27_4_lut (.I0(n49_adj_5276), .I1(n54_adj_5275), .I2(n43), 
            .I3(n44), .O(n48942));
    defparam i27_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1231 (.I0(\data_in_frame[13] [0]), .I1(n52940), 
            .I2(GND_net), .I3(GND_net), .O(n53370));
    defparam i1_2_lut_adj_1231.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1232 (.I0(\data_in_frame[16] [1]), .I1(\data_in_frame[16] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n53249));
    defparam i1_2_lut_adj_1232.LUT_INIT = 16'h6666;
    SB_LUT4 i13286_3_lut_4_lut (.I0(Kp_23__N_1583), .I1(n29100), .I2(\data_in_frame[10] [4]), 
            .I3(PWMLimit[4]), .O(n26890));
    defparam i13286_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i13203_3_lut_4_lut (.I0(n35372), .I1(n52890), .I2(rx_data[3]), 
            .I3(\data_in_frame[23] [3]), .O(n26807));
    defparam i13203_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF data_in_frame_0___i101 (.Q(\data_in_frame[12] [4]), .C(clk16MHz), 
           .D(n26157));   // verilog/coms.v(128[12] 296[6])
    SB_DFFR Kp_i0 (.Q(\Kp[0] ), .C(clk16MHz), .D(n26072), .R(reset));   // verilog/coms.v(128[12] 296[6])
    SB_DFF data_in_frame_0___i102 (.Q(\data_in_frame[12] [5]), .C(clk16MHz), 
           .D(n26160));   // verilog/coms.v(128[12] 296[6])
    SB_DFF data_in_frame_0___i103 (.Q(\data_in_frame[12] [6]), .C(clk16MHz), 
           .D(n26163));   // verilog/coms.v(128[12] 296[6])
    SB_LUT4 i3_4_lut_adj_1233 (.I0(n53607), .I1(n7_adj_5277), .I2(n23201), 
            .I3(n53004), .O(n23152));   // verilog/coms.v(71[16:27])
    defparam i3_4_lut_adj_1233.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1234 (.I0(n22610), .I1(n23152), .I2(\data_in_frame[11] [5]), 
            .I3(GND_net), .O(n22828));   // verilog/coms.v(77[16:43])
    defparam i2_3_lut_adj_1234.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1235 (.I0(\data_in_frame[11] [0]), .I1(n23193), 
            .I2(GND_net), .I3(GND_net), .O(n23509));
    defparam i1_2_lut_adj_1235.LUT_INIT = 16'h6666;
    SB_LUT4 i13206_3_lut_4_lut (.I0(n35372), .I1(n52890), .I2(rx_data[4]), 
            .I3(\data_in_frame[23] [4]), .O(n26810));
    defparam i13206_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1_2_lut_adj_1236 (.I0(\data_in_frame[9] [0]), .I1(n23753), 
            .I2(GND_net), .I3(GND_net), .O(n22658));   // verilog/coms.v(72[16:27])
    defparam i1_2_lut_adj_1236.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_1237 (.I0(\data_in_frame[11] [2]), .I1(n22658), 
            .I2(\data_in_frame[9] [1]), .I3(n23193), .O(n23402));
    defparam i3_4_lut_adj_1237.LUT_INIT = 16'h6996;
    SB_LUT4 i1_3_lut_adj_1238 (.I0(\data_in_frame[13] [3]), .I1(n23002), 
            .I2(n23402), .I3(GND_net), .O(n53091));
    defparam i1_3_lut_adj_1238.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_adj_1239 (.I0(n22813), .I1(n23288), .I2(\data_in_frame[10] [5]), 
            .I3(GND_net), .O(n23553));
    defparam i2_3_lut_adj_1239.LUT_INIT = 16'h9696;
    SB_LUT4 i13209_3_lut_4_lut (.I0(n35372), .I1(n52890), .I2(rx_data[5]), 
            .I3(\data_in_frame[23] [5]), .O(n26813));
    defparam i13209_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1_2_lut_adj_1240 (.I0(\data_in_frame[10] [6]), .I1(n22813), 
            .I2(GND_net), .I3(GND_net), .O(n53378));
    defparam i1_2_lut_adj_1240.LUT_INIT = 16'h6666;
    SB_DFFR IntegralLimit_i0_i0 (.Q(IntegralLimit[0]), .C(clk16MHz), .D(n26065), 
            .R(reset));   // verilog/coms.v(128[12] 296[6])
    SB_LUT4 i1_2_lut_adj_1241 (.I0(\data_in_frame[6] [5]), .I1(\data_in_frame[2] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_5278));   // verilog/coms.v(97[12:25])
    defparam i1_2_lut_adj_1241.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1242 (.I0(n53106), .I1(n53186), .I2(n23252), 
            .I3(n6_adj_5278), .O(n53345));   // verilog/coms.v(97[12:25])
    defparam i4_4_lut_adj_1242.LUT_INIT = 16'h6996;
    SB_LUT4 i13285_3_lut_4_lut (.I0(Kp_23__N_1583), .I1(n29100), .I2(\data_in_frame[10] [5]), 
            .I3(PWMLimit[5]), .O(n26889));
    defparam i13285_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i3_4_lut_adj_1243 (.I0(\data_in_frame[6] [6]), .I1(n53345), 
            .I2(n52915), .I3(n22688), .O(n23479));   // verilog/coms.v(77[16:43])
    defparam i3_4_lut_adj_1243.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1244 (.I0(n23479), .I1(\data_in_frame[11] [1]), 
            .I2(\data_in_frame[9] [0]), .I3(GND_net), .O(n53352));   // verilog/coms.v(77[16:43])
    defparam i2_3_lut_adj_1244.LUT_INIT = 16'h9696;
    SB_DFFESS data_out_frame_0___i83 (.Q(\data_out_frame[10] [2]), .C(clk16MHz), 
            .E(n2568), .D(n2_adj_5279), .S(n52712));   // verilog/coms.v(128[12] 296[6])
    SB_DFFR deadband_i0_i0 (.Q(\deadband[0] ), .C(clk16MHz), .D(n26064), 
            .R(reset));   // verilog/coms.v(128[12] 296[6])
    SB_LUT4 i13212_3_lut_4_lut (.I0(n35372), .I1(n52890), .I2(rx_data[6]), 
            .I3(\data_in_frame[23] [6]), .O(n26816));
    defparam i13212_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i11520_3_lut_4_lut (.I0(n10_adj_5280), .I1(n53712), .I2(reset), 
            .I3(n8_adj_5220), .O(n25123));
    defparam i11520_3_lut_4_lut.LUT_INIT = 16'hfffb;
    SB_LUT4 i1_2_lut_adj_1245 (.I0(\data_in_frame[10] [7]), .I1(n53352), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_5281));
    defparam i1_2_lut_adj_1245.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1246 (.I0(\data_in_frame[12] [7]), .I1(n53378), 
            .I2(n23553), .I3(n6_adj_5281), .O(n53532));
    defparam i4_4_lut_adj_1246.LUT_INIT = 16'h6996;
    SB_LUT4 i13215_3_lut_4_lut (.I0(n35372), .I1(n52890), .I2(rx_data[7]), 
            .I3(\data_in_frame[23] [7]), .O(n26819));
    defparam i13215_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4_4_lut_adj_1247 (.I0(\data_in_frame[15] [4]), .I1(\data_in_frame[13] [2]), 
            .I2(n53091), .I3(n53378), .O(n10_adj_5282));
    defparam i4_4_lut_adj_1247.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1248 (.I0(n54891), .I1(n47756), .I2(\data_in_frame[17] [5]), 
            .I3(GND_net), .O(n23620));
    defparam i2_3_lut_adj_1248.LUT_INIT = 16'h6969;
    SB_LUT4 i1_2_lut_adj_1249 (.I0(\data_in_frame[10] [2]), .I1(n48354), 
            .I2(GND_net), .I3(GND_net), .O(n53592));
    defparam i1_2_lut_adj_1249.LUT_INIT = 16'h6666;
    SB_LUT4 i12559_3_lut_4_lut (.I0(n8_adj_5220), .I1(n52882), .I2(rx_data[6]), 
            .I3(\data_in_frame[12] [6]), .O(n26163));
    defparam i12559_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13284_3_lut_4_lut (.I0(Kp_23__N_1583), .I1(n29100), .I2(\data_in_frame[10] [6]), 
            .I3(PWMLimit[6]), .O(n26888));
    defparam i13284_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4_4_lut_adj_1250 (.I0(\data_in_frame[8] [1]), .I1(n53427), 
            .I2(n53541), .I3(n6_adj_5283), .O(n23343));
    defparam i4_4_lut_adj_1250.LUT_INIT = 16'h6996;
    SB_LUT4 i12556_3_lut_4_lut (.I0(n8_adj_5220), .I1(n52882), .I2(rx_data[5]), 
            .I3(\data_in_frame[12] [5]), .O(n26160));
    defparam i12556_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i3_4_lut_adj_1251 (.I0(\data_in_frame[14] [4]), .I1(n53288), 
            .I2(\data_in_frame[12] [3]), .I3(n23343), .O(n48813));
    defparam i3_4_lut_adj_1251.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1252 (.I0(n48813), .I1(\data_in_frame[16] [5]), 
            .I2(n23039), .I3(GND_net), .O(n47898));
    defparam i2_3_lut_adj_1252.LUT_INIT = 16'h6969;
    SB_LUT4 i12553_3_lut_4_lut (.I0(n8_adj_5220), .I1(n52882), .I2(rx_data[4]), 
            .I3(\data_in_frame[12] [4]), .O(n26157));
    defparam i12553_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i4_4_lut_adj_1253 (.I0(\data_in_frame[16] [5]), .I1(n23620), 
            .I2(n48813), .I3(n6_adj_5284), .O(n53598));
    defparam i4_4_lut_adj_1253.LUT_INIT = 16'h6996;
    SB_LUT4 data_in_frame_13__7__I_0_2_lut (.I0(\data_in_frame[13] [7]), .I1(\data_in_frame[13] [6]), 
            .I2(GND_net), .I3(GND_net), .O(Kp_23__N_1106));   // verilog/coms.v(86[17:28])
    defparam data_in_frame_13__7__I_0_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_1254 (.I0(\data_in_frame[11] [4]), .I1(n53001), 
            .I2(\data_in_frame[9] [2]), .I3(n23144), .O(n22843));   // verilog/coms.v(74[16:42])
    defparam i3_4_lut_adj_1254.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1255 (.I0(\data_in_frame[14] [0]), .I1(\data_in_frame[11] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_5285));
    defparam i1_2_lut_adj_1255.LUT_INIT = 16'h6666;
    SB_LUT4 i12550_3_lut_4_lut (.I0(n8_adj_5220), .I1(n52882), .I2(rx_data[3]), 
            .I3(\data_in_frame[12] [3]), .O(n26154));
    defparam i12550_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i4_4_lut_adj_1256 (.I0(n23144), .I1(n20816), .I2(n52934), 
            .I3(n6_adj_5285), .O(n53163));
    defparam i4_4_lut_adj_1256.LUT_INIT = 16'h6996;
    SB_LUT4 i12547_3_lut_4_lut (.I0(n8_adj_5220), .I1(n52882), .I2(rx_data[2]), 
            .I3(\data_in_frame[12] [2]), .O(n26151));
    defparam i12547_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_1257 (.I0(n47554), .I1(\data_in_frame[10] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n47795));
    defparam i1_2_lut_adj_1257.LUT_INIT = 16'h6666;
    SB_LUT4 i18499_3_lut_4_lut (.I0(Kp_23__N_1583), .I1(n29100), .I2(\data_in_frame[10] [7]), 
            .I3(PWMLimit[7]), .O(n26887));
    defparam i18499_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i12544_3_lut_4_lut (.I0(n8_adj_5220), .I1(n52882), .I2(rx_data[1]), 
            .I3(\data_in_frame[12] [1]), .O(n26148));
    defparam i12544_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_3_lut_adj_1258 (.I0(\data_in_frame[12] [1]), .I1(\data_in_frame[11] [6]), 
            .I2(\data_in_frame[7] [3]), .I3(GND_net), .O(n53595));   // verilog/coms.v(166[9:87])
    defparam i2_3_lut_adj_1258.LUT_INIT = 16'h9696;
    SB_LUT4 i12541_3_lut_4_lut (.I0(n8_adj_5220), .I1(n52882), .I2(rx_data[0]), 
            .I3(\data_in_frame[12] [0]), .O(n26145));
    defparam i12541_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i12562_3_lut_4_lut (.I0(n8_adj_5220), .I1(n52882), .I2(rx_data[7]), 
            .I3(\data_in_frame[12] [7]), .O(n26166));
    defparam i12562_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13139_3_lut_4_lut (.I0(n8_adj_5286), .I1(n52890), .I2(rx_data[0]), 
            .I3(\data_in_frame[22] [0]), .O(n26743));
    defparam i13139_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13142_3_lut_4_lut (.I0(n8_adj_5286), .I1(n52890), .I2(rx_data[1]), 
            .I3(\data_in_frame[22] [1]), .O(n26746));
    defparam i13142_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i4_4_lut_adj_1259 (.I0(n53168), .I1(n23221), .I2(\data_in_frame[7] [0]), 
            .I3(n53449), .O(n10_adj_5287));   // verilog/coms.v(75[16:43])
    defparam i4_4_lut_adj_1259.LUT_INIT = 16'h6996;
    SB_LUT4 i13146_3_lut_4_lut (.I0(n8_adj_5286), .I1(n52890), .I2(rx_data[2]), 
            .I3(\data_in_frame[22] [2]), .O(n26750));
    defparam i13146_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_1260 (.I0(\data_in_frame[9] [3]), .I1(n23753), 
            .I2(GND_net), .I3(GND_net), .O(n53001));   // verilog/coms.v(74[16:42])
    defparam i1_2_lut_adj_1260.LUT_INIT = 16'h6666;
    SB_LUT4 i10_4_lut_adj_1261 (.I0(\data_in_frame[14] [2]), .I1(n53001), 
            .I2(\data_in_frame[5] [0]), .I3(n53565), .O(n28_adj_5288));   // verilog/coms.v(166[9:87])
    defparam i10_4_lut_adj_1261.LUT_INIT = 16'h6996;
    SB_LUT4 i14_3_lut (.I0(n22688), .I1(n28_adj_5288), .I2(\data_in_frame[3][2] ), 
            .I3(GND_net), .O(n32));   // verilog/coms.v(166[9:87])
    defparam i14_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 i13282_3_lut_4_lut (.I0(Kp_23__N_1583), .I1(n29100), .I2(\data_in_frame[9] [0]), 
            .I3(PWMLimit[8]), .O(n26886));
    defparam i13282_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i12_4_lut_adj_1262 (.I0(n22594), .I1(n53595), .I2(n47795), 
            .I3(n53465), .O(n30));   // verilog/coms.v(166[9:87])
    defparam i12_4_lut_adj_1262.LUT_INIT = 16'h6996;
    SB_LUT4 i13_4_lut_adj_1263 (.I0(n53403), .I1(\data_in_frame[7] [5]), 
            .I2(\data_in_frame[1][3] ), .I3(\data_in_frame[9] [0]), .O(n31));   // verilog/coms.v(166[9:87])
    defparam i13_4_lut_adj_1263.LUT_INIT = 16'h6996;
    SB_LUT4 i11_4_lut_adj_1264 (.I0(n23046), .I1(Kp_23__N_679), .I2(n7_adj_5277), 
            .I3(\data_in_frame[9] [6]), .O(n29_c));   // verilog/coms.v(166[9:87])
    defparam i11_4_lut_adj_1264.LUT_INIT = 16'h6996;
    SB_LUT4 i17_4_lut_adj_1265 (.I0(n29_c), .I1(n31), .I2(n30), .I3(n32), 
            .O(n48798));   // verilog/coms.v(166[9:87])
    defparam i17_4_lut_adj_1265.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1266 (.I0(n48798), .I1(\data_in_frame[16] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_5289));   // verilog/coms.v(77[16:43])
    defparam i1_2_lut_adj_1266.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1267 (.I0(n53163), .I1(n22843), .I2(Kp_23__N_1106), 
            .I3(n6_adj_5289), .O(n53252));   // verilog/coms.v(77[16:43])
    defparam i4_4_lut_adj_1267.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1268 (.I0(\data_in_frame[5] [5]), .I1(n53550), 
            .I2(n53424), .I3(\data_in_frame[7] [7]), .O(n20672));
    defparam i3_4_lut_adj_1268.LUT_INIT = 16'h6996;
    SB_LUT4 i13152_3_lut_4_lut (.I0(n8_adj_5286), .I1(n52890), .I2(rx_data[3]), 
            .I3(\data_in_frame[22] [3]), .O(n26756));
    defparam i13152_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_3_lut_adj_1269 (.I0(n20672), .I1(n23506), .I2(\data_in_frame[8] [0]), 
            .I3(GND_net), .O(n53147));
    defparam i2_3_lut_adj_1269.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1270 (.I0(\data_in_frame[1][2] ), .I1(\data_in_frame[7] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n53553));
    defparam i1_2_lut_adj_1270.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_1271 (.I0(\data_in_frame[5] [0]), .I1(n53471), 
            .I2(\data_in_frame[5] [1]), .I3(GND_net), .O(n53125));
    defparam i2_3_lut_adj_1271.LUT_INIT = 16'h9696;
    SB_LUT4 i3_4_lut_adj_1272 (.I0(\data_in_frame[2] [6]), .I1(\data_in_frame[3] [0]), 
            .I2(n53135), .I3(\data_in_frame[0] [6]), .O(n53471));   // verilog/coms.v(78[16:27])
    defparam i3_4_lut_adj_1272.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1273 (.I0(n23666), .I1(n53571), .I2(n53471), 
            .I3(n53198), .O(n20816));   // verilog/coms.v(86[17:70])
    defparam i3_4_lut_adj_1273.LUT_INIT = 16'h6996;
    SB_LUT4 i13181_3_lut_4_lut (.I0(n8_adj_5286), .I1(n52890), .I2(rx_data[4]), 
            .I3(\data_in_frame[22] [4]), .O(n26785));
    defparam i13181_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13281_3_lut_4_lut (.I0(Kp_23__N_1583), .I1(n29100), .I2(\data_in_frame[9] [1]), 
            .I3(PWMLimit[9]), .O(n26885));
    defparam i13281_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4_4_lut_adj_1274 (.I0(\data_in_frame[3][6] ), .I1(\data_in_frame[5] [7]), 
            .I2(n22652), .I3(n6_adj_5290), .O(n23506));   // verilog/coms.v(77[16:43])
    defparam i4_4_lut_adj_1274.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1275 (.I0(n23506), .I1(Kp_23__N_550), .I2(\data_in_frame[6] [1]), 
            .I3(\data_in_frame[8] [2]), .O(n3_adj_5274));   // verilog/coms.v(235[9:81])
    defparam i3_4_lut_adj_1275.LUT_INIT = 16'h6996;
    SB_LUT4 n63383_bdd_4_lut (.I0(n63383), .I1(\data_out_frame[13] [6]), 
            .I2(\data_out_frame[12] [6]), .I3(byte_transmit_counter_c[1]), 
            .O(n63386));
    defparam n63383_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_2_lut_adj_1276 (.I0(\data_in_frame[8] [1]), .I1(n3_adj_5274), 
            .I2(GND_net), .I3(GND_net), .O(n53157));
    defparam i1_2_lut_adj_1276.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1277 (.I0(n23536), .I1(\data_in_frame[4]_c [5]), 
            .I2(GND_net), .I3(GND_net), .O(n52972));   // verilog/coms.v(97[12:25])
    defparam i1_2_lut_adj_1277.LUT_INIT = 16'h6666;
    SB_LUT4 i13184_3_lut_4_lut (.I0(n8_adj_5286), .I1(n52890), .I2(rx_data[5]), 
            .I3(\data_in_frame[22] [5]), .O(n26788));
    defparam i13184_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i12741_3_lut_4_lut (.I0(Kp_23__N_1583), .I1(n29100), .I2(\data_in_frame[4]_c [4]), 
            .I3(\Ki[12] ), .O(n26345));
    defparam i12741_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1_2_lut_adj_1278 (.I0(\data_in_frame[6] [6]), .I1(n53601), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_5291));
    defparam i1_2_lut_adj_1278.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1279 (.I0(\data_in_frame[6] [7]), .I1(\data_in_frame[6] [4]), 
            .I2(\data_in_frame[6] [3]), .I3(n6_adj_5291), .O(n53243));
    defparam i4_4_lut_adj_1279.LUT_INIT = 16'h6996;
    SB_LUT4 i13187_3_lut_4_lut (.I0(n8_adj_5286), .I1(n52890), .I2(rx_data[6]), 
            .I3(\data_in_frame[22] [6]), .O(n26791));
    defparam i13187_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_1280 (.I0(\data_in_frame[3] [5]), .I1(\data_in_frame[5] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n53034));   // verilog/coms.v(97[12:25])
    defparam i1_2_lut_adj_1280.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_1281 (.I0(n22652), .I1(n53073), .I2(n53034), 
            .I3(n33_adj_5292), .O(n48415));   // verilog/coms.v(97[12:25])
    defparam i3_4_lut_adj_1281.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1282 (.I0(\data_in_frame[6] [3]), .I1(\data_in_frame[3][7] ), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_5293));   // verilog/coms.v(71[16:69])
    defparam i1_2_lut_adj_1282.LUT_INIT = 16'h6666;
    SB_LUT4 i13190_3_lut_4_lut (.I0(n8_adj_5286), .I1(n52890), .I2(rx_data[7]), 
            .I3(\data_in_frame[22] [7]), .O(n26794));
    defparam i13190_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i4_4_lut_adj_1283 (.I0(n53418), .I1(n53076), .I2(n53547), 
            .I3(n6_adj_5293), .O(n53065));   // verilog/coms.v(71[16:69])
    defparam i4_4_lut_adj_1283.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1284 (.I0(\data_in_frame[8] [4]), .I1(n53065), 
            .I2(\data_in_frame[6] [2]), .I3(Kp_23__N_704), .O(n22813));   // verilog/coms.v(75[16:43])
    defparam i3_4_lut_adj_1284.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1285 (.I0(\data_in_frame[8] [5]), .I1(n53065), 
            .I2(Kp_23__N_710), .I3(\data_in_frame[6] [4]), .O(n22713));   // verilog/coms.v(76[16:43])
    defparam i3_4_lut_adj_1285.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1286 (.I0(n53007), .I1(n53116), .I2(\data_in_frame[6] [0]), 
            .I3(GND_net), .O(n53550));
    defparam i2_3_lut_adj_1286.LUT_INIT = 16'h9696;
    SB_LUT4 i12743_3_lut_4_lut (.I0(Kp_23__N_1583), .I1(n29100), .I2(\data_in_frame[4] [2]), 
            .I3(\Ki[10] ), .O(n26347));
    defparam i12743_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1_2_lut_adj_1287 (.I0(\data_in_frame[8] [0]), .I1(n48415), 
            .I2(GND_net), .I3(GND_net), .O(n53192));
    defparam i1_2_lut_adj_1287.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1288 (.I0(n22713), .I1(n22813), .I2(GND_net), 
            .I3(GND_net), .O(Kp_23__N_902));   // verilog/coms.v(77[16:43])
    defparam i1_2_lut_adj_1288.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1289 (.I0(\data_in_frame[1][5] ), .I1(\data_in_frame[3][6] ), 
            .I2(GND_net), .I3(GND_net), .O(n53007));   // verilog/coms.v(79[16:27])
    defparam i1_2_lut_adj_1289.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1290 (.I0(\data_in_frame[4] [0]), .I1(\data_in_frame[1][5] ), 
            .I2(n53116), .I3(n6_adj_5294), .O(Kp_23__N_550));   // verilog/coms.v(76[16:27])
    defparam i4_4_lut_adj_1290.LUT_INIT = 16'h6996;
    SB_LUT4 i12733_3_lut_4_lut (.I0(n8_adj_5202), .I1(n52882), .I2(rx_data[4]), 
            .I3(\data_in_frame[13] [4]), .O(n26337));
    defparam i12733_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i12574_3_lut_4_lut (.I0(n8_adj_5202), .I1(n52882), .I2(rx_data[3]), 
            .I3(\data_in_frame[13] [3]), .O(n26178));
    defparam i12574_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i4_4_lut_adj_1291 (.I0(n53007), .I1(\data_in_frame[1][7] ), 
            .I2(\data_in_frame[2] [0]), .I3(n53406), .O(n10_adj_5295));   // verilog/coms.v(79[16:27])
    defparam i4_4_lut_adj_1291.LUT_INIT = 16'h6996;
    SB_LUT4 i5_3_lut_adj_1292 (.I0(\data_in_frame[1][6] ), .I1(n10_adj_5295), 
            .I2(\data_in_frame[1][4] ), .I3(GND_net), .O(Kp_23__N_704));   // verilog/coms.v(79[16:27])
    defparam i5_3_lut_adj_1292.LUT_INIT = 16'h9696;
    SB_LUT4 i3_4_lut_adj_1293 (.I0(\data_in_frame[8] [3]), .I1(n52986), 
            .I2(Kp_23__N_704), .I3(Kp_23__N_550), .O(n23288));
    defparam i3_4_lut_adj_1293.LUT_INIT = 16'h6996;
    SB_LUT4 i12843_3_lut_4_lut (.I0(n8_adj_5202), .I1(n52882), .I2(rx_data[5]), 
            .I3(\data_in_frame[13] [5]), .O(n26447));
    defparam i12843_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i3_4_lut_adj_1294 (.I0(\data_in_frame[5] [4]), .I1(Kp_23__N_607), 
            .I2(\data_in_frame[7] [1]), .I3(\data_in_frame[7] [4]), .O(n53403));   // verilog/coms.v(166[9:87])
    defparam i3_4_lut_adj_1294.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1295 (.I0(\data_in_frame[6] [4]), .I1(\data_in_frame[8] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n53029));   // verilog/coms.v(77[16:43])
    defparam i1_2_lut_adj_1295.LUT_INIT = 16'h6666;
    SB_LUT4 i12846_3_lut_4_lut (.I0(n8_adj_5202), .I1(n52882), .I2(rx_data[6]), 
            .I3(\data_in_frame[13] [6]), .O(n26450));
    defparam i12846_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i12849_3_lut_4_lut (.I0(n8_adj_5202), .I1(n52882), .I2(rx_data[7]), 
            .I3(\data_in_frame[13] [7]), .O(n26453));
    defparam i12849_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i12571_3_lut_4_lut (.I0(n8_adj_5202), .I1(n52882), .I2(rx_data[2]), 
            .I3(\data_in_frame[13] [2]), .O(n26175));
    defparam i12571_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_1296 (.I0(n23221), .I1(\data_in_frame[8] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n52915));   // verilog/coms.v(77[16:43])
    defparam i1_2_lut_adj_1296.LUT_INIT = 16'h6666;
    SB_LUT4 i12_4_lut_adj_1297 (.I0(n52915), .I1(\data_in_frame[4] [2]), 
            .I2(\data_in_frame[5] [3]), .I3(\data_in_frame[7] [6]), .O(n28_adj_5296));
    defparam i12_4_lut_adj_1297.LUT_INIT = 16'h6996;
    SB_LUT4 i10_4_lut_adj_1298 (.I0(\data_in_frame[7] [0]), .I1(n53029), 
            .I2(n53403), .I3(n23288), .O(n26_adj_5297));
    defparam i10_4_lut_adj_1298.LUT_INIT = 16'h6996;
    SB_LUT4 i11_4_lut_adj_1299 (.I0(Kp_23__N_902), .I1(n53318), .I2(n53541), 
            .I3(n53058), .O(n27_c));
    defparam i11_4_lut_adj_1299.LUT_INIT = 16'h6996;
    SB_LUT4 i9_4_lut_adj_1300 (.I0(\data_in_frame[9] [0]), .I1(\data_in_frame[7] [2]), 
            .I2(n53589), .I3(n53157), .O(n25_adj_5298));
    defparam i9_4_lut_adj_1300.LUT_INIT = 16'h6996;
    SB_LUT4 i15_4_lut_adj_1301 (.I0(n25_adj_5298), .I1(n27_c), .I2(n26_adj_5297), 
            .I3(n28_adj_5296), .O(n53285));
    defparam i15_4_lut_adj_1301.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1302 (.I0(\data_in_frame[1] [1]), .I1(\data_in_frame[3][2] ), 
            .I2(GND_net), .I3(GND_net), .O(n53174));   // verilog/coms.v(71[16:27])
    defparam i1_2_lut_adj_1302.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1303 (.I0(\data_in_frame[6] [1]), .I1(\data_in_frame[6] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n52986));   // verilog/coms.v(86[17:28])
    defparam i1_2_lut_adj_1303.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1304 (.I0(\data_in_frame[4] [1]), .I1(\data_in_frame[4] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n53406));   // verilog/coms.v(79[16:27])
    defparam i1_2_lut_adj_1304.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1305 (.I0(\data_in_frame[1][3] ), .I1(n53424), 
            .I2(GND_net), .I3(GND_net), .O(n20651));
    defparam i1_2_lut_adj_1305.LUT_INIT = 16'h6666;
    SB_LUT4 i12568_3_lut_4_lut (.I0(n8_adj_5202), .I1(n52882), .I2(rx_data[1]), 
            .I3(\data_in_frame[13] [1]), .O(n26172));
    defparam i12568_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_1306 (.I0(n23536), .I1(\data_in_frame[4][6] ), 
            .I2(GND_net), .I3(GND_net), .O(n53449));
    defparam i1_2_lut_adj_1306.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1307 (.I0(\data_in_frame[5] [0]), .I1(\data_in_frame[4][7] ), 
            .I2(GND_net), .I3(GND_net), .O(n53004));   // verilog/coms.v(71[16:27])
    defparam i1_2_lut_adj_1307.LUT_INIT = 16'h6666;
    SB_LUT4 i12565_3_lut_4_lut (.I0(n8_adj_5202), .I1(n52882), .I2(rx_data[0]), 
            .I3(\data_in_frame[13] [0]), .O(n26169));
    defparam i12565_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_1308 (.I0(\data_in_frame[3] [5]), .I1(\data_in_frame[5] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n53116));   // verilog/coms.v(76[16:27])
    defparam i1_2_lut_adj_1308.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1309 (.I0(\data_in_frame[4]_c [3]), .I1(\data_in_frame[4]_c [4]), 
            .I2(GND_net), .I3(GND_net), .O(n53106));   // verilog/coms.v(97[12:25])
    defparam i1_2_lut_adj_1309.LUT_INIT = 16'h6666;
    SB_LUT4 i13001_3_lut_4_lut (.I0(n8_adj_5139), .I1(n52890), .I2(rx_data[7]), 
            .I3(\data_in_frame[16] [7]), .O(n26605));
    defparam i13001_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_1310 (.I0(\data_in_frame[5] [3]), .I1(\data_in_frame[5] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n53198));   // verilog/coms.v(86[17:70])
    defparam i1_2_lut_adj_1310.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1311 (.I0(\data_in_frame[1][5] ), .I1(\data_in_frame[2] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n53076));
    defparam i1_2_lut_adj_1311.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1312 (.I0(\data_in_frame[5] [4]), .I1(\data_in_frame[5] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n53213));
    defparam i1_2_lut_adj_1312.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1313 (.I0(\data_in_frame[5] [1]), .I1(\data_in_frame[3] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n53565));   // verilog/coms.v(79[16:27])
    defparam i1_2_lut_adj_1313.LUT_INIT = 16'h6666;
    SB_LUT4 i12742_3_lut_4_lut (.I0(Kp_23__N_1583), .I1(n29100), .I2(\data_in_frame[4]_c [3]), 
            .I3(\Ki[11] ), .O(n26346));
    defparam i12742_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i6_4_lut_adj_1314 (.I0(n23046), .I1(\data_in_frame[3][1] ), 
            .I2(Kp_23__N_679), .I3(n23536), .O(n16_adj_5299));   // verilog/coms.v(79[16:27])
    defparam i6_4_lut_adj_1314.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut_adj_1315 (.I0(n53141), .I1(n53456), .I2(n23221), 
            .I3(n53076), .O(n17));   // verilog/coms.v(79[16:27])
    defparam i7_4_lut_adj_1315.LUT_INIT = 16'h6996;
    SB_LUT4 i9_4_lut_adj_1316 (.I0(n17), .I1(n23252), .I2(n16_adj_5299), 
            .I3(\data_in_frame[0] [7]), .O(n55110));   // verilog/coms.v(79[16:27])
    defparam i9_4_lut_adj_1316.LUT_INIT = 16'h6996;
    SB_LUT4 i12998_3_lut_4_lut (.I0(n8_adj_5139), .I1(n52890), .I2(rx_data[6]), 
            .I3(\data_in_frame[16] [6]), .O(n26602));
    defparam i12998_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i12_4_lut_adj_1317 (.I0(n53198), .I1(n52989), .I2(n53106), 
            .I3(\data_in_frame[4] [2]), .O(n28_adj_5300));   // verilog/coms.v(79[16:27])
    defparam i12_4_lut_adj_1317.LUT_INIT = 16'h6996;
    SB_LUT4 i10_4_lut_adj_1318 (.I0(n53445), .I1(n53565), .I2(\data_in_frame[5] [6]), 
            .I3(n53213), .O(n26_adj_5301));   // verilog/coms.v(79[16:27])
    defparam i10_4_lut_adj_1318.LUT_INIT = 16'h6996;
    SB_LUT4 i11_4_lut_adj_1319 (.I0(n53004), .I1(n53449), .I2(n20651), 
            .I3(n53406), .O(n27_adj_5302));   // verilog/coms.v(79[16:27])
    defparam i11_4_lut_adj_1319.LUT_INIT = 16'h6996;
    SB_LUT4 i12995_3_lut_4_lut (.I0(n8_adj_5139), .I1(n52890), .I2(rx_data[5]), 
            .I3(\data_in_frame[16] [5]), .O(n26599));
    defparam i12995_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i9_4_lut_adj_1320 (.I0(\data_in_frame[6] [5]), .I1(n52986), 
            .I2(n55110), .I3(n53174), .O(n25_adj_5303));   // verilog/coms.v(79[16:27])
    defparam i9_4_lut_adj_1320.LUT_INIT = 16'h6996;
    SB_LUT4 i15_4_lut_adj_1321 (.I0(n25_adj_5303), .I1(n27_adj_5302), .I2(n26_adj_5301), 
            .I3(n28_adj_5300), .O(n53601));   // verilog/coms.v(79[16:27])
    defparam i15_4_lut_adj_1321.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1322 (.I0(\data_in_frame[1][4] ), .I1(\data_in_frame[1][3] ), 
            .I2(GND_net), .I3(GND_net), .O(n33_adj_5292));   // verilog/coms.v(97[12:25])
    defparam i1_2_lut_adj_1322.LUT_INIT = 16'h6666;
    SB_LUT4 data_in_frame_1__5__I_0_2_lut (.I0(\data_in_frame[1][5] ), .I1(\data_in_frame[1][4] ), 
            .I2(GND_net), .I3(GND_net), .O(Kp_23__N_679));   // verilog/coms.v(77[16:27])
    defparam data_in_frame_1__5__I_0_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1323 (.I0(\data_in_frame[4] [1]), .I1(\data_in_frame[0] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n53547));   // verilog/coms.v(71[16:69])
    defparam i1_2_lut_adj_1323.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_1324 (.I0(n47950), .I1(n53553), .I2(n53427), 
            .I3(\data_in_frame[5] [3]), .O(n48768));
    defparam i3_4_lut_adj_1324.LUT_INIT = 16'h6996;
    SB_LUT4 i3_2_lut (.I0(\data_in_frame[3] [4]), .I1(\data_in_frame[8] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n16_adj_5304));
    defparam i3_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i9_4_lut_adj_1325 (.I0(n48768), .I1(n53547), .I2(n53445), 
            .I3(n53183), .O(n22_adj_5305));
    defparam i9_4_lut_adj_1325.LUT_INIT = 16'h6996;
    SB_LUT4 i12992_3_lut_4_lut (.I0(n8_adj_5139), .I1(n52890), .I2(rx_data[4]), 
            .I3(\data_in_frame[16] [4]), .O(n26596));
    defparam i12992_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i12989_3_lut_4_lut (.I0(n8_adj_5139), .I1(n52890), .I2(rx_data[3]), 
            .I3(\data_in_frame[16] [3]), .O(n26593));
    defparam i12989_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i7_3_lut_adj_1326 (.I0(n53601), .I1(\data_in_frame[8] [6]), 
            .I2(n53589), .I3(GND_net), .O(n20_adj_5306));
    defparam i7_3_lut_adj_1326.LUT_INIT = 16'h9696;
    SB_LUT4 i12900_3_lut_4_lut (.I0(n8_adj_5139), .I1(n52890), .I2(rx_data[0]), 
            .I3(\data_in_frame[16] [0]), .O(n26504));
    defparam i12900_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i11_4_lut_adj_1327 (.I0(\data_in_frame[8] [3]), .I1(n22_adj_5305), 
            .I2(n16_adj_5304), .I3(n22713), .O(n24_adj_5307));
    defparam i11_4_lut_adj_1327.LUT_INIT = 16'h6996;
    SB_LUT4 i12_4_lut_adj_1328 (.I0(n53285), .I1(n24_adj_5307), .I2(n20_adj_5306), 
            .I3(Kp_23__N_915), .O(n55472));
    defparam i12_4_lut_adj_1328.LUT_INIT = 16'h6996;
    SB_LUT4 i12903_3_lut_4_lut (.I0(n8_adj_5139), .I1(n52890), .I2(rx_data[1]), 
            .I3(\data_in_frame[16] [1]), .O(n26507));
    defparam i12903_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i6_4_lut_adj_1329 (.I0(\data_in_frame[12] [0]), .I1(n55472), 
            .I2(\data_in_frame[2] [1]), .I3(\data_in_frame[8] [0]), .O(n16_adj_5308));
    defparam i6_4_lut_adj_1329.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut_adj_1330 (.I0(\data_in_frame[8] [1]), .I1(\data_in_frame[8] [7]), 
            .I2(\data_in_frame[8] [2]), .I3(n47554), .O(n17_adj_5309));
    defparam i7_4_lut_adj_1330.LUT_INIT = 16'h6996;
    SB_LUT4 i9_4_lut_adj_1331 (.I0(n17_adj_5309), .I1(\data_in_frame[9] [6]), 
            .I2(n16_adj_5308), .I3(\data_in_frame[5] [5]), .O(n53465));
    defparam i9_4_lut_adj_1331.LUT_INIT = 16'h6996;
    SB_LUT4 i12906_3_lut_4_lut (.I0(n8_adj_5139), .I1(n52890), .I2(rx_data[2]), 
            .I3(\data_in_frame[16] [2]), .O(n26510));
    defparam i12906_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 equal_288_i8_2_lut_3_lut (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(\FRAME_MATCHER.i [0]), .I3(GND_net), .O(n8_adj_5074));   // verilog/coms.v(154[7:23])
    defparam equal_288_i8_2_lut_3_lut.LUT_INIT = 16'hefef;
    SB_LUT4 i4_4_lut_adj_1332 (.I0(\data_in_frame[7] [2]), .I1(n22818), 
            .I2(n53449), .I3(n6_adj_5310), .O(n23144));
    defparam i4_4_lut_adj_1332.LUT_INIT = 16'h6996;
    SB_LUT4 equal_281_i8_2_lut_3_lut (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(\FRAME_MATCHER.i [0]), .I3(GND_net), .O(n8_adj_5139));   // verilog/coms.v(154[7:23])
    defparam equal_281_i8_2_lut_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i1_2_lut_adj_1333 (.I0(\data_in_frame[1] [0]), .I1(Kp_23__N_602), 
            .I2(GND_net), .I3(GND_net), .O(n53135));   // verilog/coms.v(78[16:27])
    defparam i1_2_lut_adj_1333.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1334 (.I0(\data_in_frame[1][3] ), .I1(\data_in_frame[1][2] ), 
            .I2(GND_net), .I3(GND_net), .O(n53050));
    defparam i1_2_lut_adj_1334.LUT_INIT = 16'h6666;
    SB_LUT4 data_in_frame_1__7__I_0_2_lut (.I0(\data_in_frame[1][7] ), .I1(\data_in_frame[1][6] ), 
            .I2(GND_net), .I3(GND_net), .O(Kp_23__N_607));   // verilog/coms.v(79[16:27])
    defparam data_in_frame_1__7__I_0_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_3_lut_adj_1335 (.I0(n48787), .I1(n21971), .I2(n47956), 
            .I3(GND_net), .O(n47851));
    defparam i1_2_lut_3_lut_adj_1335.LUT_INIT = 16'h9696;
    SB_LUT4 i3_4_lut_adj_1336 (.I0(Kp_23__N_607), .I1(Kp_23__N_679), .I2(n53050), 
            .I3(\data_in_frame[1] [1]), .O(Kp_23__N_602));   // verilog/coms.v(86[17:63])
    defparam i3_4_lut_adj_1336.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1337 (.I0(\data_in_frame[3][1] ), .I1(Kp_23__N_602), 
            .I2(\data_in_frame[0] [7]), .I3(n23046), .O(n47950));   // verilog/coms.v(72[16:69])
    defparam i3_4_lut_adj_1337.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1338 (.I0(n48787), .I1(n21971), .I2(\data_out_frame[22] [7]), 
            .I3(GND_net), .O(n53498));
    defparam i1_2_lut_3_lut_adj_1338.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1339 (.I0(\data_in_frame[7] [3]), .I1(n47950), 
            .I2(GND_net), .I3(GND_net), .O(n53318));
    defparam i1_2_lut_adj_1339.LUT_INIT = 16'h6666;
    SB_LUT4 i2_2_lut_3_lut (.I0(n55268), .I1(n48824), .I2(n53097), .I3(GND_net), 
            .O(n6_adj_5311));
    defparam i2_2_lut_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1340 (.I0(\data_in_frame[5] [1]), .I1(n53456), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_5312));
    defparam i1_2_lut_adj_1340.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1341 (.I0(\data_in_frame[5] [2]), .I1(\data_in_frame[4][7] ), 
            .I2(n53318), .I3(n6_adj_5312), .O(n53458));
    defparam i4_4_lut_adj_1341.LUT_INIT = 16'h6996;
    SB_LUT4 data_in_frame_9__7__I_0_2_lut (.I0(\data_in_frame[9] [7]), .I1(\data_in_frame[9] [6]), 
            .I2(GND_net), .I3(GND_net), .O(Kp_23__N_920));   // verilog/coms.v(86[17:28])
    defparam data_in_frame_9__7__I_0_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1342 (.I0(\data_in_frame[9] [4]), .I1(\data_in_frame[9] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n52934));
    defparam i1_2_lut_adj_1342.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1343 (.I0(\data_in_frame[9] [1]), .I1(\data_in_frame[9] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n22594));   // verilog/coms.v(73[16:41])
    defparam i1_2_lut_adj_1343.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_1344 (.I0(n22594), .I1(n52934), .I2(Kp_23__N_920), 
            .I3(\data_in_frame[9] [3]), .O(Kp_23__N_915));
    defparam i3_4_lut_adj_1344.LUT_INIT = 16'h6996;
    SB_LUT4 select_715_Select_223_i3_3_lut_4_lut (.I0(n55268), .I1(n48824), 
            .I2(n48809), .I3(\FRAME_MATCHER.state[3] ), .O(n3_adj_5151));
    defparam select_715_Select_223_i3_3_lut_4_lut.LUT_INIT = 16'h6900;
    SB_LUT4 i2_3_lut_adj_1345 (.I0(\data_in_frame[9] [3]), .I1(\data_in_frame[9] [4]), 
            .I2(n53458), .I3(GND_net), .O(n22610));   // verilog/coms.v(75[16:43])
    defparam i2_3_lut_adj_1345.LUT_INIT = 16'h6969;
    SB_LUT4 i3_4_lut_adj_1346 (.I0(\data_in_frame[12] [2]), .I1(n22610), 
            .I2(Kp_23__N_915), .I3(n23741), .O(n55482));
    defparam i3_4_lut_adj_1346.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1347 (.I0(n48777), .I1(n53498), .I2(n53207), 
            .I3(GND_net), .O(n53474));
    defparam i1_2_lut_3_lut_adj_1347.LUT_INIT = 16'h9696;
    SB_LUT4 i2_2_lut_adj_1348 (.I0(\data_in_frame[12] [1]), .I1(\data_in_frame[10] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_5313));
    defparam i2_2_lut_adj_1348.LUT_INIT = 16'h6666;
    SB_LUT4 i1_4_lut_adj_1349 (.I0(\data_in_frame[14] [3]), .I1(n53147), 
            .I2(n6_adj_5313), .I3(n55482), .O(n23039));
    defparam i1_4_lut_adj_1349.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1350 (.I0(n23039), .I1(\data_in_frame[16] [4]), 
            .I2(\data_in_frame[16] [3]), .I3(GND_net), .O(n53298));
    defparam i2_3_lut_adj_1350.LUT_INIT = 16'h9696;
    SB_LUT4 i6_4_lut_adj_1351 (.I0(\data_in_frame[13] [7]), .I1(\data_in_frame[14] [1]), 
            .I2(n53168), .I3(n22658), .O(n16_adj_5314));   // verilog/coms.v(75[16:43])
    defparam i6_4_lut_adj_1351.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut_adj_1352 (.I0(n23144), .I1(n53058), .I2(n53465), 
            .I3(n53458), .O(n17_adj_5315));   // verilog/coms.v(75[16:43])
    defparam i7_4_lut_adj_1352.LUT_INIT = 16'h9669;
    SB_LUT4 i2_3_lut_4_lut (.I0(n48777), .I1(n53498), .I2(n48824), .I3(n47851), 
            .O(n48239));
    defparam i2_3_lut_4_lut.LUT_INIT = 16'h9669;
    SB_LUT4 i9_4_lut_adj_1353 (.I0(n17_adj_5315), .I1(\data_in_frame[11] [5]), 
            .I2(n16_adj_5314), .I3(n23741), .O(n48392));   // verilog/coms.v(75[16:43])
    defparam i9_4_lut_adj_1353.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1354 (.I0(\FRAME_MATCHER.i_31__N_2322 ), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n1_adj_5245));
    defparam i1_2_lut_3_lut_adj_1354.LUT_INIT = 16'h1010;
    SB_LUT4 i1_2_lut_adj_1355 (.I0(\data_in_frame[16] [3]), .I1(n53252), 
            .I2(GND_net), .I3(GND_net), .O(n53253));
    defparam i1_2_lut_adj_1355.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1356 (.I0(\data_in_frame[18] [0]), .I1(n53598), 
            .I2(GND_net), .I3(GND_net), .O(n52995));
    defparam i1_2_lut_adj_1356.LUT_INIT = 16'h6666;
    SB_LUT4 i5_3_lut_adj_1357 (.I0(\data_in_frame[15] [7]), .I1(n22828), 
            .I2(\data_in_frame[13] [2]), .I3(GND_net), .O(n14_adj_5316));
    defparam i5_3_lut_adj_1357.LUT_INIT = 16'h9696;
    SB_LUT4 select_717_Select_7_i1_2_lut_3_lut (.I0(\FRAME_MATCHER.i_31__N_2322 ), 
            .I1(\FRAME_MATCHER.state[3] ), .I2(byte_transmit_counter_c[7]), 
            .I3(GND_net), .O(n1_adj_5157));
    defparam select_717_Select_7_i1_2_lut_3_lut.LUT_INIT = 16'h1010;
    SB_LUT4 select_717_Select_6_i1_2_lut_3_lut (.I0(\FRAME_MATCHER.i_31__N_2322 ), 
            .I1(\FRAME_MATCHER.state[3] ), .I2(byte_transmit_counter_c[6]), 
            .I3(GND_net), .O(n1_adj_5156));
    defparam select_717_Select_6_i1_2_lut_3_lut.LUT_INIT = 16'h1010;
    SB_LUT4 i8_4_lut_adj_1358 (.I0(n15_adj_5317), .I1(n22822), .I2(n14_adj_5316), 
            .I3(n53512), .O(n55195));
    defparam i8_4_lut_adj_1358.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1359 (.I0(\FRAME_MATCHER.i_31__N_2322 ), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(byte_transmit_counter_c[5]), .I3(GND_net), .O(n1_adj_5155));
    defparam i1_2_lut_3_lut_adj_1359.LUT_INIT = 16'h1010;
    SB_LUT4 i4_4_lut_adj_1360 (.I0(n55195), .I1(n52995), .I2(n53253), 
            .I3(n48794), .O(n10_adj_5318));
    defparam i4_4_lut_adj_1360.LUT_INIT = 16'h6996;
    SB_LUT4 i5_3_lut_adj_1361 (.I0(n22021), .I1(n10_adj_5318), .I2(n20730), 
            .I3(GND_net), .O(n53311));
    defparam i5_3_lut_adj_1361.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1362 (.I0(\FRAME_MATCHER.i_31__N_2322 ), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(byte_transmit_counter_c[4]), .I3(GND_net), .O(n1_adj_5154));
    defparam i1_2_lut_3_lut_adj_1362.LUT_INIT = 16'h1010;
    SB_LUT4 i1_2_lut_3_lut_adj_1363 (.I0(\FRAME_MATCHER.i_31__N_2322 ), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(byte_transmit_counter_c[3]), .I3(GND_net), .O(n1_adj_5153));
    defparam i1_2_lut_3_lut_adj_1363.LUT_INIT = 16'h1010;
    SB_LUT4 i1_2_lut_3_lut_adj_1364 (.I0(\FRAME_MATCHER.i_31__N_2322 ), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(byte_transmit_counter_c[1]), .I3(GND_net), .O(n1_c));
    defparam i1_2_lut_3_lut_adj_1364.LUT_INIT = 16'h1010;
    SB_LUT4 i2_2_lut_3_lut_4_lut (.I0(\FRAME_MATCHER.i_31__N_2322 ), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(\FRAME_MATCHER.i_31__N_2323 ), .I3(\FRAME_MATCHER.i_31__N_2325 ), 
            .O(n6_adj_5319));
    defparam i2_2_lut_3_lut_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_3_lut_adj_1365 (.I0(\FRAME_MATCHER.i_31__N_2322 ), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(\byte_transmit_counter[2] ), .I3(GND_net), .O(n1_adj_5152));
    defparam i1_2_lut_3_lut_adj_1365.LUT_INIT = 16'h1010;
    SB_LUT4 i12876_3_lut_4_lut (.I0(n35372), .I1(n52882), .I2(rx_data[0]), 
            .I3(\data_in_frame[15] [0]), .O(n26480));
    defparam i12876_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i3_4_lut_adj_1366 (.I0(\data_in_frame[17] [4]), .I1(n22898), 
            .I2(\data_in_frame[15] [3]), .I3(n47764), .O(n47876));
    defparam i3_4_lut_adj_1366.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1367 (.I0(\data_in_frame[17] [6]), .I1(n22623), 
            .I2(\data_in_frame[20] [0]), .I3(GND_net), .O(n52924));
    defparam i2_3_lut_adj_1367.LUT_INIT = 16'h9696;
    SB_LUT4 i4_4_lut_adj_1368 (.I0(n52924), .I1(n47876), .I2(\data_in_frame[20] [1]), 
            .I3(n53311), .O(n10_adj_5320));
    defparam i4_4_lut_adj_1368.LUT_INIT = 16'h6996;
    SB_LUT4 i2_2_lut_adj_1369 (.I0(\data_in_frame[22] [3]), .I1(n53276), 
            .I2(GND_net), .I3(GND_net), .O(n8_adj_5321));
    defparam i2_2_lut_adj_1369.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1370 (.I0(\data_in_frame[20] [1]), .I1(n8_adj_5321), 
            .I2(n53400), .I3(\data_in_frame[20] [2]), .O(n10_adj_5322));
    defparam i4_4_lut_adj_1370.LUT_INIT = 16'h6996;
    SB_LUT4 i5_4_lut_adj_1371 (.I0(\data_in_frame[19] [2]), .I1(n53246), 
            .I2(\data_in_frame[23] [4]), .I3(n48844), .O(n12_adj_5323));
    defparam i5_4_lut_adj_1371.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1372 (.I0(\data_in_frame[23] [6]), .I1(n53409), 
            .I2(n53015), .I3(\data_in_frame[21] [4]), .O(n54668));
    defparam i3_4_lut_adj_1372.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_1373 (.I0(\data_in_frame[21] [2]), .I1(n12_adj_5323), 
            .I2(n53329), .I3(\data_in_frame[21] [3]), .O(n54475));
    defparam i6_4_lut_adj_1373.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_1374 (.I0(\data_in_frame[22] [6]), .I1(n20730), 
            .I2(n22631), .I3(n6_adj_5324), .O(n54715));
    defparam i4_4_lut_adj_1374.LUT_INIT = 16'h6996;
    SB_LUT4 i12879_3_lut_4_lut (.I0(n35372), .I1(n52882), .I2(rx_data[1]), 
            .I3(\data_in_frame[15] [1]), .O(n26483));
    defparam i12879_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1_3_lut_adj_1375 (.I0(\data_in_frame[23] [5]), .I1(\data_in_frame[21] [4]), 
            .I2(\data_in_frame[21] [3]), .I3(GND_net), .O(n5_adj_5325));
    defparam i1_3_lut_adj_1375.LUT_INIT = 16'h9696;
    SB_LUT4 i4_4_lut_adj_1376 (.I0(\data_in_frame[20] [2]), .I1(\data_in_frame[18] [2]), 
            .I2(n20730), .I3(\data_in_frame[22] [4]), .O(n10_adj_5326));
    defparam i4_4_lut_adj_1376.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1377 (.I0(n55426), .I1(n5_adj_5325), .I2(n53489), 
            .I3(n48904), .O(n18_adj_5327));
    defparam i1_4_lut_adj_1377.LUT_INIT = 16'h1441;
    SB_LUT4 i1_rep_170_2_lut (.I0(\data_in_frame[19] [6]), .I1(\data_in_frame[21] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n63878));
    defparam i1_rep_170_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_1378 (.I0(\data_in_frame[22] [0]), .I1(n63878), 
            .I2(n53228), .I3(n47882), .O(n54852));
    defparam i3_4_lut_adj_1378.LUT_INIT = 16'h6996;
    SB_LUT4 i12882_3_lut_4_lut (.I0(n35372), .I1(n52882), .I2(rx_data[2]), 
            .I3(\data_in_frame[15] [2]), .O(n26486));
    defparam i12882_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1_4_lut_adj_1379 (.I0(\data_in_frame[21] [6]), .I1(n47876), 
            .I2(\data_in_frame[19] [5]), .I3(n23006), .O(n5_adj_5328));
    defparam i1_4_lut_adj_1379.LUT_INIT = 16'h9669;
    SB_LUT4 i12885_3_lut_4_lut (.I0(n35372), .I1(n52882), .I2(rx_data[3]), 
            .I3(\data_in_frame[15] [3]), .O(n26489));
    defparam i12885_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1_3_lut_adj_1380 (.I0(n52924), .I1(\data_in_frame[19] [7]), 
            .I2(\data_in_frame[19] [5]), .I3(GND_net), .O(n6_adj_5329));
    defparam i1_3_lut_adj_1380.LUT_INIT = 16'h9696;
    SB_LUT4 i5_3_lut_adj_1381 (.I0(\data_in_frame[19] [6]), .I1(n10_adj_5320), 
            .I2(\data_in_frame[22] [2]), .I3(GND_net), .O(n54458));
    defparam i5_3_lut_adj_1381.LUT_INIT = 16'h9696;
    SB_LUT4 i12888_3_lut_4_lut (.I0(n35372), .I1(n52882), .I2(rx_data[4]), 
            .I3(\data_in_frame[15] [4]), .O(n26492));
    defparam i12888_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i2_3_lut_adj_1382 (.I0(\data_in_frame[23] [1]), .I1(n53240), 
            .I2(n48923), .I3(GND_net), .O(n54948));
    defparam i2_3_lut_adj_1382.LUT_INIT = 16'h9696;
    SB_LUT4 i4_4_lut_adj_1383 (.I0(\data_in_frame[22] [1]), .I1(n23006), 
            .I2(n53228), .I3(n6_adj_5329), .O(n54867));
    defparam i4_4_lut_adj_1383.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1384 (.I0(\data_in_frame[22] [5]), .I1(n53400), 
            .I2(n52980), .I3(\data_in_frame[18] [3]), .O(n54619));
    defparam i3_4_lut_adj_1384.LUT_INIT = 16'h6996;
    SB_LUT4 i5_4_lut_adj_1385 (.I0(n48794), .I1(\data_in_frame[20] [6]), 
            .I2(n54876), .I3(n55195), .O(n12_adj_5330));
    defparam i5_4_lut_adj_1385.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1386 (.I0(\data_in_frame[23] [3]), .I1(n53240), 
            .I2(\data_in_frame[21] [2]), .I3(\data_in_frame[21] [1]), .O(n54950));
    defparam i3_4_lut_adj_1386.LUT_INIT = 16'h6996;
    SB_LUT4 i12891_3_lut_4_lut (.I0(n35372), .I1(n52882), .I2(rx_data[5]), 
            .I3(\data_in_frame[15] [5]), .O(n26495));
    defparam i12891_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i3_4_lut_adj_1387 (.I0(n9), .I1(\data_in_frame[23] [0]), .I2(n10_adj_5322), 
            .I3(n54876), .O(n20_adj_5331));
    defparam i3_4_lut_adj_1387.LUT_INIT = 16'h4812;
    SB_LUT4 i11_4_lut_adj_1388 (.I0(n54715), .I1(n54475), .I2(n54880), 
            .I3(n54668), .O(n28_adj_5332));
    defparam i11_4_lut_adj_1388.LUT_INIT = 16'h2000;
    SB_LUT4 i12894_3_lut_4_lut (.I0(n35372), .I1(n52882), .I2(rx_data[6]), 
            .I3(\data_in_frame[15] [6]), .O(n26498));
    defparam i12894_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i6_4_lut_adj_1389 (.I0(\data_in_frame[20] [5]), .I1(n12_adj_5330), 
            .I2(n22677), .I3(\data_in_frame[22] [7]), .O(n55002));
    defparam i6_4_lut_adj_1389.LUT_INIT = 16'h6996;
    SB_LUT4 i12897_3_lut_4_lut (.I0(n35372), .I1(n52882), .I2(rx_data[7]), 
            .I3(\data_in_frame[15] [7]), .O(n26501));
    defparam i12897_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i39056_3_lut_4_lut (.I0(n10_adj_5333), .I1(n53712), .I2(n8_adj_5220), 
            .I3(reset), .O(n7));
    defparam i39056_3_lut_4_lut.LUT_INIT = 16'hfffb;
    SB_LUT4 i9_4_lut_adj_1390 (.I0(\data_in_frame[20] [3]), .I1(n18_adj_5327), 
            .I2(n10_adj_5326), .I3(n53276), .O(n26_adj_5334));
    defparam i9_4_lut_adj_1390.LUT_INIT = 16'h4884;
    SB_LUT4 i41892_4_lut (.I0(n5_adj_5328), .I1(n54852), .I2(n53015), 
            .I3(\data_in_frame[23] [7]), .O(n56589));
    defparam i41892_4_lut.LUT_INIT = 16'hedde;
    SB_LUT4 i11554_3_lut_4_lut (.I0(n10_adj_5333), .I1(n53712), .I2(reset), 
            .I3(n8_adj_5335), .O(n25157));
    defparam i11554_3_lut_4_lut.LUT_INIT = 16'hfffb;
    SB_LUT4 i12_4_lut_adj_1391 (.I0(n54619), .I1(n54867), .I2(n54948), 
            .I3(n54458), .O(n29_adj_5336));
    defparam i12_4_lut_adj_1391.LUT_INIT = 16'h8000;
    SB_LUT4 i14_4_lut (.I0(n55002), .I1(n28_adj_5332), .I2(n20_adj_5331), 
            .I3(n54950), .O(n31_adj_5337));
    defparam i14_4_lut.LUT_INIT = 16'h0080;
    SB_LUT4 i16_4_lut_adj_1392 (.I0(n31_adj_5337), .I1(n29_adj_5336), .I2(n56589), 
            .I3(n26_adj_5334), .O(n29100));
    defparam i16_4_lut_adj_1392.LUT_INIT = 16'h0800;
    SB_LUT4 i1_2_lut_3_lut_adj_1393 (.I0(n10_adj_5333), .I1(n53712), .I2(n8), 
            .I3(GND_net), .O(n25103));
    defparam i1_2_lut_3_lut_adj_1393.LUT_INIT = 16'hfbfb;
    SB_LUT4 i11558_3_lut_4_lut (.I0(n10_adj_5333), .I1(n53712), .I2(reset), 
            .I3(n8_adj_5074), .O(n25161));
    defparam i11558_3_lut_4_lut.LUT_INIT = 16'hfffb;
    SB_LUT4 i12852_3_lut_4_lut (.I0(n8_adj_5286), .I1(n52882), .I2(rx_data[0]), 
            .I3(\data_in_frame[14] [0]), .O(n26456));
    defparam i12852_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i12855_3_lut_4_lut (.I0(n8_adj_5286), .I1(n52882), .I2(rx_data[1]), 
            .I3(\data_in_frame[14] [1]), .O(n26459));
    defparam i12855_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i41879_2_lut (.I0(n23288), .I1(n22713), .I2(GND_net), .I3(GND_net), 
            .O(n56574));
    defparam i41879_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i4_4_lut_adj_1394 (.I0(n52989), .I1(\data_in_frame[1][5] ), 
            .I2(\data_in_frame[8] [1]), .I3(n53243), .O(n10_adj_5338));
    defparam i4_4_lut_adj_1394.LUT_INIT = 16'h6996;
    SB_LUT4 i41881_4_lut (.I0(n48768), .I1(n52972), .I2(n10_adj_5338), 
            .I3(\data_in_frame[1][3] ), .O(n56576));
    defparam i41881_4_lut.LUT_INIT = 16'hebbe;
    SB_LUT4 i12858_3_lut_4_lut (.I0(n8_adj_5286), .I1(n52882), .I2(rx_data[2]), 
            .I3(\data_in_frame[14] [2]), .O(n26462));
    defparam i12858_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13_4_lut_adj_1395 (.I0(n56574), .I1(n23753), .I2(n23193), 
            .I3(n20820), .O(n30_adj_5339));
    defparam i13_4_lut_adj_1395.LUT_INIT = 16'h0100;
    SB_LUT4 i12861_3_lut_4_lut (.I0(n8_adj_5286), .I1(n52882), .I2(rx_data[3]), 
            .I3(\data_in_frame[14] [3]), .O(n26465));
    defparam i12861_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i5_3_lut_adj_1396 (.I0(n48354), .I1(n53458), .I2(\data_in_frame[7] [7]), 
            .I3(GND_net), .O(n22_adj_5340));
    defparam i5_3_lut_adj_1396.LUT_INIT = 16'h8484;
    SB_LUT4 i41883_2_lut (.I0(n23479), .I1(n55426), .I2(GND_net), .I3(GND_net), 
            .O(n56578));
    defparam i41883_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i15_4_lut_adj_1397 (.I0(n20816), .I1(n30_adj_5339), .I2(n56576), 
            .I3(n53192), .O(n32_adj_5341));
    defparam i15_4_lut_adj_1397.LUT_INIT = 16'h0800;
    SB_LUT4 i42021_4_lut (.I0(n3_adj_5274), .I1(n23152), .I2(n23144), 
            .I3(n22813), .O(n56724));
    defparam i42021_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i16_4_lut_adj_1398 (.I0(n56724), .I1(n32_adj_5341), .I2(n56578), 
            .I3(n22_adj_5340), .O(n22333));
    defparam i16_4_lut_adj_1398.LUT_INIT = 16'h0400;
    SB_LUT4 i12864_3_lut_4_lut (.I0(n8_adj_5286), .I1(n52882), .I2(rx_data[4]), 
            .I3(\data_in_frame[14] [4]), .O(n26468));
    defparam i12864_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15500_4_lut (.I0(n22333), .I1(Kp_23__N_1583), .I2(\FRAME_MATCHER.i_31__N_2324 ), 
            .I3(n29100), .O(n24563));   // verilog/coms.v(18[27:29])
    defparam i15500_4_lut.LUT_INIT = 16'hac20;
    SB_LUT4 i12867_3_lut_4_lut (.I0(n8_adj_5286), .I1(n52882), .I2(rx_data[5]), 
            .I3(\data_in_frame[14] [5]), .O(n26471));
    defparam i12867_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i12870_3_lut_4_lut (.I0(n8_adj_5286), .I1(n52882), .I2(rx_data[6]), 
            .I3(\data_in_frame[14] [6]), .O(n26474));
    defparam i12870_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i12873_3_lut_4_lut (.I0(n8_adj_5286), .I1(n52882), .I2(rx_data[7]), 
            .I3(\data_in_frame[14] [7]), .O(n26477));
    defparam i12873_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i6_4_lut_adj_1399 (.I0(\FRAME_MATCHER.i [13]), .I1(\FRAME_MATCHER.i [16]), 
            .I2(\FRAME_MATCHER.i [28]), .I3(\FRAME_MATCHER.i [20]), .O(n16_adj_5342));
    defparam i6_4_lut_adj_1399.LUT_INIT = 16'hfffe;
    SB_LUT4 i7_4_lut_adj_1400 (.I0(\FRAME_MATCHER.i [14]), .I1(\FRAME_MATCHER.i [7]), 
            .I2(\FRAME_MATCHER.i [11]), .I3(\FRAME_MATCHER.i [9]), .O(n17_adj_5343));
    defparam i7_4_lut_adj_1400.LUT_INIT = 16'hfffe;
    SB_LUT4 i3_4_lut_adj_1401 (.I0(\FRAME_MATCHER.i [15]), .I1(\FRAME_MATCHER.i [17]), 
            .I2(\FRAME_MATCHER.i [18]), .I3(\FRAME_MATCHER.i [21]), .O(n55383));
    defparam i3_4_lut_adj_1401.LUT_INIT = 16'hfffe;
    SB_LUT4 i3_4_lut_adj_1402 (.I0(\FRAME_MATCHER.i [10]), .I1(\FRAME_MATCHER.i [25]), 
            .I2(\FRAME_MATCHER.i [23]), .I3(\FRAME_MATCHER.i [19]), .O(n55141));
    defparam i3_4_lut_adj_1402.LUT_INIT = 16'hfffe;
    SB_LUT4 i9_4_lut_adj_1403 (.I0(n17_adj_5343), .I1(\FRAME_MATCHER.i [27]), 
            .I2(n16_adj_5342), .I3(\FRAME_MATCHER.i [12]), .O(n55476));
    defparam i9_4_lut_adj_1403.LUT_INIT = 16'hfffe;
    SB_LUT4 i2_3_lut_4_lut_adj_1404 (.I0(n29111), .I1(n4425), .I2(n1702), 
            .I3(n1705), .O(n54660));   // verilog/coms.v(143[4] 145[7])
    defparam i2_3_lut_4_lut_adj_1404.LUT_INIT = 16'h2000;
    SB_LUT4 i7_4_lut_adj_1405 (.I0(n55383), .I1(\FRAME_MATCHER.i [26]), 
            .I2(\FRAME_MATCHER.i [22]), .I3(\FRAME_MATCHER.i [6]), .O(n18_adj_5344));
    defparam i7_4_lut_adj_1405.LUT_INIT = 16'hfffe;
    SB_LUT4 i5_2_lut_adj_1406 (.I0(\FRAME_MATCHER.i [30]), .I1(\FRAME_MATCHER.i [5]), 
            .I2(GND_net), .I3(GND_net), .O(n16_adj_5345));
    defparam i5_2_lut_adj_1406.LUT_INIT = 16'heeee;
    SB_LUT4 i9_4_lut_adj_1407 (.I0(\FRAME_MATCHER.i [24]), .I1(n18_adj_5344), 
            .I2(n55476), .I3(n55141), .O(n20_adj_5346));
    defparam i9_4_lut_adj_1407.LUT_INIT = 16'hfffe;
    SB_LUT4 i2_3_lut_4_lut_adj_1408 (.I0(n29111), .I1(n4425), .I2(\FRAME_MATCHER.i_31__N_2325 ), 
            .I3(n4_adj_5347), .O(n54478));   // verilog/coms.v(143[4] 145[7])
    defparam i2_3_lut_4_lut_adj_1408.LUT_INIT = 16'hff20;
    SB_LUT4 i10_4_lut_adj_1409 (.I0(\FRAME_MATCHER.i [8]), .I1(n20_adj_5346), 
            .I2(n16_adj_5345), .I3(\FRAME_MATCHER.i [29]), .O(n22428));
    defparam i10_4_lut_adj_1409.LUT_INIT = 16'hfffe;
    SB_LUT4 i21944_4_lut (.I0(\FRAME_MATCHER.i [3]), .I1(\FRAME_MATCHER.i [31]), 
            .I2(n22428), .I3(\FRAME_MATCHER.i [4]), .O(n4425));   // verilog/coms.v(254[9:58])
    defparam i21944_4_lut.LUT_INIT = 16'h3230;
    SB_LUT4 i452_2_lut (.I0(n4425), .I1(\FRAME_MATCHER.i_31__N_2325 ), .I2(GND_net), 
            .I3(GND_net), .O(n1816));   // verilog/coms.v(146[4] 295[11])
    defparam i452_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i13112_3_lut_4_lut (.I0(n8_adj_5202), .I1(n52890), .I2(rx_data[1]), 
            .I3(\data_in_frame[21] [1]), .O(n26716));
    defparam i13112_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13115_3_lut_4_lut (.I0(n8_adj_5202), .I1(n52890), .I2(rx_data[2]), 
            .I3(\data_in_frame[21] [2]), .O(n26719));
    defparam i13115_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13118_3_lut_4_lut (.I0(n8_adj_5202), .I1(n52890), .I2(rx_data[3]), 
            .I3(\data_in_frame[21] [3]), .O(n26722));
    defparam i13118_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13121_3_lut_4_lut (.I0(n8_adj_5202), .I1(n52890), .I2(rx_data[4]), 
            .I3(\data_in_frame[21] [4]), .O(n26725));
    defparam i13121_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13125_3_lut_4_lut (.I0(n8_adj_5202), .I1(n52890), .I2(rx_data[5]), 
            .I3(\data_in_frame[21] [5]), .O(n26729));
    defparam i13125_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13128_3_lut_4_lut (.I0(n8_adj_5202), .I1(n52890), .I2(rx_data[6]), 
            .I3(\data_in_frame[21] [6]), .O(n26732));
    defparam i13128_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13136_3_lut_4_lut (.I0(n8_adj_5202), .I1(n52890), .I2(rx_data[7]), 
            .I3(\data_in_frame[21] [7]), .O(n26740));
    defparam i13136_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13109_3_lut_4_lut (.I0(n8_adj_5202), .I1(n52890), .I2(rx_data[0]), 
            .I3(\data_in_frame[21] [0]), .O(n26713));
    defparam i13109_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 select_715_Select_15_i2_3_lut (.I0(\data_out_frame[1][7] ), .I1(\FRAME_MATCHER.i_31__N_2320 ), 
            .I2(\FRAME_MATCHER.state_31__N_2423 [3]), .I3(GND_net), .O(n2_adj_5059));   // verilog/coms.v(146[4] 295[11])
    defparam select_715_Select_15_i2_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 select_715_Select_14_i2_3_lut (.I0(\data_out_frame[1][6] ), .I1(\FRAME_MATCHER.i_31__N_2320 ), 
            .I2(\FRAME_MATCHER.state_31__N_2423 [3]), .I3(GND_net), .O(n2_adj_5058));   // verilog/coms.v(146[4] 295[11])
    defparam select_715_Select_14_i2_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i1_3_lut_adj_1410 (.I0(\FRAME_MATCHER.i_31__N_2320 ), .I1(\FRAME_MATCHER.state_31__N_2423 [3]), 
            .I2(\data_out_frame[1][5] ), .I3(GND_net), .O(n2_adj_5057));   // verilog/coms.v(146[4] 295[11])
    defparam i1_3_lut_adj_1410.LUT_INIT = 16'ha8a8;
    SB_LUT4 select_715_Select_11_i2_3_lut (.I0(\data_out_frame[1][3] ), .I1(\FRAME_MATCHER.i_31__N_2320 ), 
            .I2(\FRAME_MATCHER.state_31__N_2423 [3]), .I3(GND_net), .O(n2_adj_5056));   // verilog/coms.v(146[4] 295[11])
    defparam select_715_Select_11_i2_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 select_715_Select_9_i2_3_lut (.I0(\data_out_frame[1][1] ), .I1(\FRAME_MATCHER.i_31__N_2320 ), 
            .I2(\FRAME_MATCHER.state_31__N_2423 [3]), .I3(GND_net), .O(n2_adj_5055));   // verilog/coms.v(146[4] 295[11])
    defparam select_715_Select_9_i2_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 select_715_Select_8_i2_3_lut (.I0(\FRAME_MATCHER.state_31__N_2423 [3]), 
            .I1(\FRAME_MATCHER.i_31__N_2320 ), .I2(\data_out_frame[1][0] ), 
            .I3(GND_net), .O(n2_adj_5054));   // verilog/coms.v(146[4] 295[11])
    defparam select_715_Select_8_i2_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i42160_4_lut (.I0(\data_out_frame[0][4] ), .I1(\data_out_frame[3][4] ), 
            .I2(byte_transmit_counter_c[1]), .I3(byte_transmit_counter[0]), 
            .O(n56872));
    defparam i42160_4_lut.LUT_INIT = 16'hc00a;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_2_i21_4_lut (.I0(\data_out_frame[21] [2]), 
            .I1(\data_out_frame[22] [2]), .I2(byte_transmit_counter_c[1]), 
            .I3(byte_transmit_counter[0]), .O(n21));   // verilog/coms.v(107[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_2_i21_4_lut.LUT_INIT = 16'h0ac0;
    SB_LUT4 i11145_3_lut (.I0(\data_out_frame[1][6] ), .I1(\data_out_frame[3][6] ), 
            .I2(byte_transmit_counter_c[1]), .I3(GND_net), .O(n24742));   // verilog/coms.v(107[34:55])
    defparam i11145_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i42215_3_lut (.I0(\data_out_frame[6] [6]), .I1(\data_out_frame[7] [6]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n56927));
    defparam i42215_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i42216_4_lut (.I0(n56927), .I1(n24742), .I2(\byte_transmit_counter[2] ), 
            .I3(byte_transmit_counter[0]), .O(n56928));
    defparam i42216_4_lut.LUT_INIT = 16'haca0;
    SB_LUT4 i42214_3_lut (.I0(\data_out_frame[4] [6]), .I1(\data_out_frame[5] [6]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n56926));
    defparam i42214_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2227687_i1_3_lut (.I0(n63320), .I1(n63386), .I2(\byte_transmit_counter[2] ), 
            .I3(GND_net), .O(n14_adj_5348));
    defparam i2227687_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_6_i16_3_lut (.I0(\data_out_frame[16] [6]), 
            .I1(\data_out_frame[17] [6]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n16_adj_5349));   // verilog/coms.v(107[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_6_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i47275_4_lut (.I0(n16_adj_5349), .I1(\data_out_frame[21] [6]), 
            .I2(\byte_transmit_counter[2] ), .I3(byte_transmit_counter[0]), 
            .O(n61988));
    defparam i47275_4_lut.LUT_INIT = 16'hca0a;
    SB_LUT4 i47276_4_lut (.I0(n61988), .I1(n59927), .I2(byte_transmit_counter_c[1]), 
            .I3(\data_out_frame[22] [6]), .O(n61989));
    defparam i47276_4_lut.LUT_INIT = 16'hca0a;
    SB_LUT4 i42121_3_lut (.I0(\data_out_frame[8] [1]), .I1(\data_out_frame[9] [1]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n56833));
    defparam i42121_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i42122_3_lut (.I0(\data_out_frame[10] [1]), .I1(\data_out_frame[11] [1]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n56834));
    defparam i42122_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i42233_3_lut (.I0(\data_out_frame[14] [1]), .I1(\data_out_frame[15] [1]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n56945));
    defparam i42233_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i42232_3_lut (.I0(\data_out_frame[12] [1]), .I1(\data_out_frame[13] [1]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n56944));
    defparam i42232_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i42229_3_lut (.I0(\data_out_frame[8] [0]), .I1(\data_out_frame[9] [0]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n56941));
    defparam i42229_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i42230_3_lut (.I0(\data_out_frame[10] [0]), .I1(\data_out_frame[11] [0]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n56942));
    defparam i42230_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i42296_3_lut (.I0(\data_out_frame[14] [0]), .I1(\data_out_frame[15] [0]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n57008));
    defparam i42296_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i42295_3_lut (.I0(\data_out_frame[12] [0]), .I1(\data_out_frame[13] [0]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n57007));
    defparam i42295_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i42211_3_lut (.I0(\data_out_frame[4] [5]), .I1(\data_out_frame[5] [5]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n56923));
    defparam i42211_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i42212_3_lut (.I0(\data_out_frame[6] [5]), .I1(\data_out_frame[7] [5]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n56924));
    defparam i42212_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i45412_2_lut (.I0(\data_out_frame[22] [5]), .I1(byte_transmit_counter[0]), 
            .I2(GND_net), .I3(GND_net), .O(n59727));   // verilog/coms.v(107[34:55])
    defparam i45412_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i45407_2_lut (.I0(\data_out_frame[21] [5]), .I1(byte_transmit_counter[0]), 
            .I2(GND_net), .I3(GND_net), .O(n59726));   // verilog/coms.v(107[34:55])
    defparam i45407_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i11119_3_lut (.I0(\data_out_frame[1][1] ), .I1(\data_out_frame[3][1] ), 
            .I2(byte_transmit_counter_c[1]), .I3(GND_net), .O(n24714));   // verilog/coms.v(107[34:55])
    defparam i11119_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i42218_3_lut (.I0(\data_out_frame[6] [1]), .I1(\data_out_frame[7] [1]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n56930));
    defparam i42218_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i42219_4_lut (.I0(n56930), .I1(n24714), .I2(\byte_transmit_counter[2] ), 
            .I3(byte_transmit_counter[0]), .O(n56931));
    defparam i42219_4_lut.LUT_INIT = 16'haca0;
    SB_LUT4 i42217_3_lut (.I0(\data_out_frame[4] [1]), .I1(\data_out_frame[5] [1]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n56929));
    defparam i42217_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_3_i1_3_lut (.I0(\data_out_frame[0][3] ), 
            .I1(\data_out_frame[1][3] ), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n1_adj_5350));   // verilog/coms.v(107[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_3_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i42151_4_lut (.I0(n1_adj_5350), .I1(\data_out_frame[3][3] ), 
            .I2(byte_transmit_counter_c[1]), .I3(byte_transmit_counter[0]), 
            .O(n56863));
    defparam i42151_4_lut.LUT_INIT = 16'hca0a;
    SB_LUT4 i45353_4_lut (.I0(\data_out_frame[26] [1]), .I1(n24840), .I2(\data_out_frame[27] [1]), 
            .I3(byte_transmit_counter[0]), .O(n59910));
    defparam i45353_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_1_i21_4_lut (.I0(\data_out_frame[21] [1]), 
            .I1(\data_out_frame[22] [1]), .I2(byte_transmit_counter_c[1]), 
            .I3(byte_transmit_counter[0]), .O(n21_adj_5351));   // verilog/coms.v(107[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_1_i21_4_lut.LUT_INIT = 16'h0ac0;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_1_i16_3_lut (.I0(\data_out_frame[16] [1]), 
            .I1(\data_out_frame[17] [1]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n16_adj_5352));   // verilog/coms.v(107[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_1_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_1_i22_4_lut (.I0(n16_adj_5352), 
            .I1(n21_adj_5351), .I2(\byte_transmit_counter[2] ), .I3(byte_transmit_counter_c[1]), 
            .O(n22_adj_5353));   // verilog/coms.v(107[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_1_i22_4_lut.LUT_INIT = 16'hc0ca;
    SB_LUT4 i42206_3_lut (.I0(\data_out_frame[6] [0]), .I1(\data_out_frame[7] [0]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n56918));
    defparam i42206_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i42207_4_lut (.I0(n56918), .I1(n24853), .I2(\byte_transmit_counter[2] ), 
            .I3(\data_out_frame[1][0] ), .O(n56919));
    defparam i42207_4_lut.LUT_INIT = 16'ha3a0;
    SB_LUT4 i42205_3_lut (.I0(\data_out_frame[4] [0]), .I1(\data_out_frame[5] [0]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n56917));
    defparam i42205_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i45555_4_lut (.I0(\data_out_frame[26] [0]), .I1(n24840), .I2(\data_out_frame[27] [0]), 
            .I3(byte_transmit_counter[0]), .O(n59912));
    defparam i45555_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_0_i21_4_lut (.I0(\data_out_frame[21] [0]), 
            .I1(\data_out_frame[22] [0]), .I2(byte_transmit_counter_c[1]), 
            .I3(byte_transmit_counter[0]), .O(n21_adj_5354));   // verilog/coms.v(107[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_0_i21_4_lut.LUT_INIT = 16'h0ac0;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_0_i16_3_lut (.I0(\data_out_frame[16] [0]), 
            .I1(\data_out_frame[17] [0]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n16_adj_5355));   // verilog/coms.v(107[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_0_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_0_i22_4_lut (.I0(n16_adj_5355), 
            .I1(n21_adj_5354), .I2(\byte_transmit_counter[2] ), .I3(byte_transmit_counter_c[1]), 
            .O(n22_adj_5356));   // verilog/coms.v(107[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_0_i22_4_lut.LUT_INIT = 16'hc0ca;
    SB_LUT4 i20257_4_lut (.I0(encoder0_position[6]), .I1(encoder1_position[6]), 
            .I2(n15_adj_3), .I3(n15), .O(n33792));
    defparam i20257_4_lut.LUT_INIT = 16'hf535;
    SB_LUT4 byte_transmit_counter_3__bdd_4_lut_48837 (.I0(byte_transmit_counter_c[3]), 
            .I1(n22_adj_5356), .I2(n59912), .I3(byte_transmit_counter_c[4]), 
            .O(n63557));
    defparam byte_transmit_counter_3__bdd_4_lut_48837.LUT_INIT = 16'he4aa;
    SB_LUT4 i1_3_lut_adj_1411 (.I0(\control_mode[1] ), .I1(n22431), .I2(\control_mode[0] ), 
            .I3(GND_net), .O(n15_adj_3));   // verilog/coms.v(128[12] 296[6])
    defparam i1_3_lut_adj_1411.LUT_INIT = 16'hfefe;
    SB_LUT4 n63557_bdd_4_lut (.I0(n63557), .I1(n63332), .I2(n7_adj_5358), 
            .I3(byte_transmit_counter_c[4]), .O(tx_data[0]));
    defparam n63557_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_2_lut_adj_1412 (.I0(control_mode_c[2]), .I1(control_mode_c[3]), 
            .I2(GND_net), .I3(GND_net), .O(n1));
    defparam i1_2_lut_adj_1412.LUT_INIT = 16'heeee;
    SB_LUT4 select_715_Select_82_i2_4_lut (.I0(\data_out_frame[10] [2]), .I1(\FRAME_MATCHER.i_31__N_2320 ), 
            .I2(encoder1_position[10]), .I3(\FRAME_MATCHER.state_31__N_2423 [3]), 
            .O(n2_adj_5279));   // verilog/coms.v(146[4] 295[11])
    defparam select_715_Select_82_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i18452_1_lut (.I0(deadband_c[2]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n32007));   // verilog/coms.v(128[12] 296[6])
    defparam i18452_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i2_3_lut_4_lut_adj_1413 (.I0(\data_out_frame[16] [7]), .I1(n53195), 
            .I2(\data_out_frame[17] [2]), .I3(n23375), .O(n53267));
    defparam i2_3_lut_4_lut_adj_1413.LUT_INIT = 16'h6996;
    SB_LUT4 i2_2_lut_3_lut_4_lut_adj_1414 (.I0(\data_out_frame[16] [7]), .I1(n53195), 
            .I2(\data_out_frame[16] [5]), .I3(\data_out_frame[16] [6]), 
            .O(n10_adj_5122));
    defparam i2_2_lut_3_lut_4_lut_adj_1414.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut (.I0(\data_out_frame[4] [3]), .I1(\data_out_frame[4] [2]), 
            .I2(\data_out_frame[6] [4]), .I3(\data_out_frame[8] [5]), .O(n53043));   // verilog/coms.v(76[16:43])
    defparam i1_2_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_adj_1415 (.I0(\data_out_frame[4] [3]), .I1(\data_out_frame[4] [2]), 
            .I2(\data_out_frame[6] [4]), .I3(\data_out_frame[8] [6]), .O(n23635));   // verilog/coms.v(76[16:43])
    defparam i1_2_lut_4_lut_adj_1415.LUT_INIT = 16'h6996;
    SB_LUT4 i17425_3_lut (.I0(\control_mode[0] ), .I1(\data_in_frame[1] [0]), 
            .I2(n19639), .I3(GND_net), .O(n26082));
    defparam i17425_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i5_3_lut_4_lut (.I0(\data_out_frame[5] [3]), .I1(\data_out_frame[8] [1]), 
            .I2(\data_out_frame[5] [7]), .I3(n10_adj_5131), .O(n52968));   // verilog/coms.v(76[16:27])
    defparam i5_3_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 select_715_Select_81_i2_4_lut (.I0(\data_out_frame[10] [1]), .I1(\FRAME_MATCHER.i_31__N_2320 ), 
            .I2(encoder1_position[9]), .I3(\FRAME_MATCHER.state_31__N_2423 [3]), 
            .O(n2_adj_5273));   // verilog/coms.v(146[4] 295[11])
    defparam select_715_Select_81_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_715_Select_80_i2_4_lut (.I0(\data_out_frame[10] [0]), .I1(\FRAME_MATCHER.i_31__N_2320 ), 
            .I2(encoder1_position[8]), .I3(\FRAME_MATCHER.state_31__N_2423 [3]), 
            .O(n2_adj_5272));   // verilog/coms.v(146[4] 295[11])
    defparam select_715_Select_80_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i2_3_lut_4_lut_adj_1416 (.I0(\data_out_frame[10] [2]), .I1(\data_out_frame[10] [3]), 
            .I2(\data_out_frame[4] [0]), .I3(\data_out_frame[6] [0]), .O(n8_adj_5130));   // verilog/coms.v(86[17:70])
    defparam i2_3_lut_4_lut_adj_1416.LUT_INIT = 16'h6996;
    SB_LUT4 select_715_Select_79_i2_4_lut (.I0(\data_out_frame[9] [7]), .I1(\FRAME_MATCHER.i_31__N_2320 ), 
            .I2(encoder1_position[23]), .I3(\FRAME_MATCHER.state_31__N_2423 [3]), 
            .O(n2_adj_5271));   // verilog/coms.v(146[4] 295[11])
    defparam select_715_Select_79_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_715_Select_78_i2_4_lut (.I0(\data_out_frame[9] [6]), .I1(\FRAME_MATCHER.i_31__N_2320 ), 
            .I2(encoder1_position[22]), .I3(\FRAME_MATCHER.state_31__N_2423 [3]), 
            .O(n2_adj_5270));   // verilog/coms.v(146[4] 295[11])
    defparam select_715_Select_78_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i4_2_lut_3_lut (.I0(\data_out_frame[10] [2]), .I1(\data_out_frame[10] [3]), 
            .I2(n53515), .I3(GND_net), .O(n18));   // verilog/coms.v(86[17:70])
    defparam i4_2_lut_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 select_715_Select_77_i2_4_lut (.I0(\data_out_frame[9] [5]), .I1(\FRAME_MATCHER.i_31__N_2320 ), 
            .I2(encoder1_position[21]), .I3(\FRAME_MATCHER.state_31__N_2423 [3]), 
            .O(n2_adj_5269));   // verilog/coms.v(146[4] 295[11])
    defparam select_715_Select_77_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_715_Select_76_i2_4_lut (.I0(\data_out_frame[9] [4]), .I1(\FRAME_MATCHER.i_31__N_2320 ), 
            .I2(encoder1_position[20]), .I3(\FRAME_MATCHER.state_31__N_2423 [3]), 
            .O(n2_adj_5268));   // verilog/coms.v(146[4] 295[11])
    defparam select_715_Select_76_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_715_Select_75_i2_4_lut (.I0(\data_out_frame[9] [3]), .I1(\FRAME_MATCHER.i_31__N_2320 ), 
            .I2(encoder1_position[19]), .I3(\FRAME_MATCHER.state_31__N_2423 [3]), 
            .O(n2_adj_5267));   // verilog/coms.v(146[4] 295[11])
    defparam select_715_Select_75_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_715_Select_74_i2_4_lut (.I0(\data_out_frame[9] [2]), .I1(\FRAME_MATCHER.i_31__N_2320 ), 
            .I2(encoder1_position[18]), .I3(\FRAME_MATCHER.state_31__N_2423 [3]), 
            .O(n2_adj_5266));   // verilog/coms.v(146[4] 295[11])
    defparam select_715_Select_74_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_715_Select_73_i2_4_lut (.I0(\data_out_frame[9] [1]), .I1(\FRAME_MATCHER.i_31__N_2320 ), 
            .I2(encoder1_position[17]), .I3(\FRAME_MATCHER.state_31__N_2423 [3]), 
            .O(n2_adj_5265));   // verilog/coms.v(146[4] 295[11])
    defparam select_715_Select_73_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_715_Select_72_i2_4_lut (.I0(\data_out_frame[9] [0]), .I1(\FRAME_MATCHER.i_31__N_2320 ), 
            .I2(encoder1_position[16]), .I3(\FRAME_MATCHER.state_31__N_2423 [3]), 
            .O(n2_adj_5264));   // verilog/coms.v(146[4] 295[11])
    defparam select_715_Select_72_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_715_Select_71_i2_4_lut (.I0(\data_out_frame[8] [7]), .I1(\FRAME_MATCHER.i_31__N_2320 ), 
            .I2(encoder0_position[7]), .I3(\FRAME_MATCHER.state_31__N_2423 [3]), 
            .O(n2_adj_5263));   // verilog/coms.v(146[4] 295[11])
    defparam select_715_Select_71_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_715_Select_70_i2_4_lut (.I0(\data_out_frame[8] [6]), .I1(\FRAME_MATCHER.i_31__N_2320 ), 
            .I2(encoder0_position[6]), .I3(\FRAME_MATCHER.state_31__N_2423 [3]), 
            .O(n2_adj_5262));   // verilog/coms.v(146[4] 295[11])
    defparam select_715_Select_70_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_715_Select_69_i2_4_lut (.I0(\data_out_frame[8] [5]), .I1(\FRAME_MATCHER.i_31__N_2320 ), 
            .I2(encoder0_position[5]), .I3(\FRAME_MATCHER.state_31__N_2423 [3]), 
            .O(n2_adj_5261));   // verilog/coms.v(146[4] 295[11])
    defparam select_715_Select_69_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_715_Select_68_i2_4_lut (.I0(\data_out_frame[8] [4]), .I1(\FRAME_MATCHER.i_31__N_2320 ), 
            .I2(encoder0_position[4]), .I3(\FRAME_MATCHER.state_31__N_2423 [3]), 
            .O(n2_adj_5260));   // verilog/coms.v(146[4] 295[11])
    defparam select_715_Select_68_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_715_Select_67_i2_4_lut (.I0(\data_out_frame[8] [3]), .I1(\FRAME_MATCHER.i_31__N_2320 ), 
            .I2(encoder0_position[3]), .I3(\FRAME_MATCHER.state_31__N_2423 [3]), 
            .O(n2_adj_5259));   // verilog/coms.v(146[4] 295[11])
    defparam select_715_Select_67_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_715_Select_66_i2_4_lut (.I0(\data_out_frame[8] [2]), .I1(\FRAME_MATCHER.i_31__N_2320 ), 
            .I2(encoder0_position[2]), .I3(\FRAME_MATCHER.state_31__N_2423 [3]), 
            .O(n2_adj_5258));   // verilog/coms.v(146[4] 295[11])
    defparam select_715_Select_66_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_4_lut_adj_1417 (.I0(\FRAME_MATCHER.i_31__N_2320 ), .I1(\data_out_frame[8] [1]), 
            .I2(encoder0_position[1]), .I3(\FRAME_MATCHER.state_31__N_2423 [3]), 
            .O(n2_adj_5257));   // verilog/coms.v(146[4] 295[11])
    defparam i1_4_lut_adj_1417.LUT_INIT = 16'ha088;
    SB_LUT4 select_715_Select_64_i2_4_lut (.I0(\data_out_frame[8] [0]), .I1(\FRAME_MATCHER.i_31__N_2320 ), 
            .I2(encoder0_position[0]), .I3(\FRAME_MATCHER.state_31__N_2423 [3]), 
            .O(n2_adj_5256));   // verilog/coms.v(146[4] 295[11])
    defparam select_715_Select_64_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_715_Select_63_i2_4_lut (.I0(\data_out_frame[7] [7]), .I1(\FRAME_MATCHER.i_31__N_2320 ), 
            .I2(encoder0_position[15]), .I3(\FRAME_MATCHER.state_31__N_2423 [3]), 
            .O(n2_adj_5255));   // verilog/coms.v(146[4] 295[11])
    defparam select_715_Select_63_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_715_Select_62_i2_4_lut (.I0(\data_out_frame[7] [6]), .I1(\FRAME_MATCHER.i_31__N_2320 ), 
            .I2(encoder0_position[14]), .I3(\FRAME_MATCHER.state_31__N_2423 [3]), 
            .O(n2_adj_5254));   // verilog/coms.v(146[4] 295[11])
    defparam select_715_Select_62_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_715_Select_61_i2_4_lut (.I0(\data_out_frame[7] [5]), .I1(\FRAME_MATCHER.i_31__N_2320 ), 
            .I2(encoder0_position[13]), .I3(\FRAME_MATCHER.state_31__N_2423 [3]), 
            .O(n2_adj_5253));   // verilog/coms.v(146[4] 295[11])
    defparam select_715_Select_61_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_715_Select_60_i2_4_lut (.I0(\data_out_frame[7] [4]), .I1(\FRAME_MATCHER.i_31__N_2320 ), 
            .I2(encoder0_position[12]), .I3(\FRAME_MATCHER.state_31__N_2423 [3]), 
            .O(n2_adj_5252));   // verilog/coms.v(146[4] 295[11])
    defparam select_715_Select_60_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_4_lut_adj_1418 (.I0(\FRAME_MATCHER.i_31__N_2320 ), .I1(\data_out_frame[7] [3]), 
            .I2(encoder0_position[11]), .I3(\FRAME_MATCHER.state_31__N_2423 [3]), 
            .O(n2_adj_5251));   // verilog/coms.v(146[4] 295[11])
    defparam i1_4_lut_adj_1418.LUT_INIT = 16'ha088;
    SB_LUT4 select_715_Select_58_i2_4_lut (.I0(\data_out_frame[7] [2]), .I1(\FRAME_MATCHER.i_31__N_2320 ), 
            .I2(encoder0_position[10]), .I3(\FRAME_MATCHER.state_31__N_2423 [3]), 
            .O(n2_adj_5250));   // verilog/coms.v(146[4] 295[11])
    defparam select_715_Select_58_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_715_Select_57_i2_4_lut (.I0(\data_out_frame[7] [1]), .I1(\FRAME_MATCHER.i_31__N_2320 ), 
            .I2(encoder0_position[9]), .I3(\FRAME_MATCHER.state_31__N_2423 [3]), 
            .O(n2_adj_5249));   // verilog/coms.v(146[4] 295[11])
    defparam select_715_Select_57_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_715_Select_56_i2_4_lut (.I0(\data_out_frame[7] [0]), .I1(\FRAME_MATCHER.i_31__N_2320 ), 
            .I2(encoder0_position[8]), .I3(\FRAME_MATCHER.state_31__N_2423 [3]), 
            .O(n2_adj_5248));   // verilog/coms.v(146[4] 295[11])
    defparam select_715_Select_56_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i6_3_lut_4_lut (.I0(n53439), .I1(n53559), .I2(n53436), .I3(n53012), 
            .O(n17_adj_5360));
    defparam i6_3_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_1419 (.I0(n53439), .I1(n53559), .I2(\data_out_frame[14] [7]), 
            .I3(n53391), .O(n48497));
    defparam i2_3_lut_4_lut_adj_1419.LUT_INIT = 16'h6996;
    SB_LUT4 i12627_3_lut_4_lut (.I0(n25103), .I1(reset), .I2(rx_data[7]), 
            .I3(\data_in_frame[2] [7]), .O(n26231));
    defparam i12627_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i12623_3_lut_4_lut (.I0(n25103), .I1(reset), .I2(rx_data[6]), 
            .I3(\data_in_frame[2] [6]), .O(n26227));
    defparam i12623_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_3_lut_4_lut (.I0(n23110), .I1(\data_out_frame[15] [4]), 
            .I2(\data_out_frame[15] [3]), .I3(n53559), .O(n47634));
    defparam i1_2_lut_3_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1420 (.I0(\data_out_frame[6] [1]), .I1(\data_out_frame[4] [0]), 
            .I2(\data_out_frame[4] [1]), .I3(\data_out_frame[6] [2]), .O(n22526));   // verilog/coms.v(74[16:42])
    defparam i1_2_lut_3_lut_4_lut_adj_1420.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1421 (.I0(n22822), .I1(n23402), .I2(n53144), 
            .I3(n54891), .O(n22623));
    defparam i1_2_lut_3_lut_4_lut_adj_1421.LUT_INIT = 16'h9669;
    SB_LUT4 i12620_3_lut_4_lut (.I0(n25103), .I1(reset), .I2(rx_data[5]), 
            .I3(\data_in_frame[2] [5]), .O(n26224));
    defparam i12620_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i6_4_lut_3_lut_4_lut (.I0(n52952), .I1(n48392), .I2(\data_in_frame[16] [1]), 
            .I3(\data_in_frame[16] [2]), .O(n15_adj_5317));
    defparam i6_4_lut_3_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1422 (.I0(\data_in_frame[15] [6]), .I1(\data_in_frame[13] [4]), 
            .I2(\data_in_frame[13] [5]), .I3(\data_in_frame[13] [6]), .O(n6_adj_5246));   // verilog/coms.v(77[16:43])
    defparam i1_2_lut_3_lut_4_lut_adj_1422.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1423 (.I0(n47766), .I1(n53394), .I2(\data_out_frame[14] [5]), 
            .I3(n52968), .O(n53436));
    defparam i1_2_lut_3_lut_4_lut_adj_1423.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1424 (.I0(\data_in_frame[13] [1]), .I1(\data_in_frame[13] [3]), 
            .I2(\data_in_frame[13] [4]), .I3(\data_in_frame[13] [2]), .O(n53529));   // verilog/coms.v(86[17:63])
    defparam i1_2_lut_3_lut_4_lut_adj_1424.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1425 (.I0(\data_in_frame[13] [1]), .I1(\data_in_frame[13] [3]), 
            .I2(\data_in_frame[13] [4]), .I3(\data_in_frame[13] [7]), .O(n53512));   // verilog/coms.v(86[17:63])
    defparam i1_2_lut_3_lut_4_lut_adj_1425.LUT_INIT = 16'h6996;
    SB_LUT4 i12617_3_lut_4_lut (.I0(n25103), .I1(reset), .I2(rx_data[4]), 
            .I3(\data_in_frame[2] [4]), .O(n26221));
    defparam i12617_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_3_lut_adj_1426 (.I0(n10_adj_5280), .I1(n53712), .I2(n8_adj_5335), 
            .I3(GND_net), .O(n25071));
    defparam i1_2_lut_3_lut_adj_1426.LUT_INIT = 16'hfbfb;
    SB_LUT4 i11_4_lut_4_lut_adj_1427 (.I0(n25103), .I1(reset), .I2(rx_data[3]), 
            .I3(\data_in_frame[2] [3]), .O(n52143));
    defparam i11_4_lut_4_lut_adj_1427.LUT_INIT = 16'hfe10;
    SB_LUT4 i12611_3_lut_4_lut (.I0(n25103), .I1(reset), .I2(rx_data[2]), 
            .I3(\data_in_frame[2] [2]), .O(n26215));
    defparam i12611_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i12608_3_lut_4_lut (.I0(n25103), .I1(reset), .I2(rx_data[1]), 
            .I3(\data_in_frame[2] [1]), .O(n26212));
    defparam i12608_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i12604_3_lut_4_lut (.I0(n25103), .I1(reset), .I2(rx_data[0]), 
            .I3(\data_in_frame[2] [0]), .O(n26208));
    defparam i12604_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_4_lut_adj_1428 (.I0(DE_c), .I1(\FRAME_MATCHER.i_31__N_2320 ), 
            .I2(n6_adj_5319), .I3(n29098), .O(n23764));   // verilog/coms.v(146[4] 295[11])
    defparam i1_4_lut_adj_1428.LUT_INIT = 16'haaa8;
    SB_LUT4 select_1656_Select_0_i1_2_lut (.I0(tx_transmit_N_3189), .I1(\FRAME_MATCHER.i_31__N_2322 ), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5244));   // verilog/coms.v(146[4] 295[11])
    defparam select_1656_Select_0_i1_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 equal_295_i8_2_lut_3_lut (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(\FRAME_MATCHER.i [0]), .I3(GND_net), .O(n8));   // verilog/coms.v(154[7:23])
    defparam equal_295_i8_2_lut_3_lut.LUT_INIT = 16'hfdfd;
    SB_LUT4 select_715_Select_183_i2_4_lut (.I0(\data_out_frame[22] [7]), 
            .I1(\FRAME_MATCHER.i_31__N_2320 ), .I2(\current[7] ), .I3(\FRAME_MATCHER.state_31__N_2423 [3]), 
            .O(n2_adj_5243));   // verilog/coms.v(146[4] 295[11])
    defparam select_715_Select_183_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_4_lut_adj_1429 (.I0(\FRAME_MATCHER.i_31__N_2320 ), .I1(\data_out_frame[22] [6]), 
            .I2(\current[6] ), .I3(\FRAME_MATCHER.state_31__N_2423 [3]), 
            .O(n2_adj_5242));   // verilog/coms.v(146[4] 295[11])
    defparam i1_4_lut_adj_1429.LUT_INIT = 16'ha088;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1430 (.I0(\data_in_frame[7] [6]), .I1(n23666), 
            .I2(\data_in_frame[10] [2]), .I3(n48354), .O(n6_adj_5283));
    defparam i1_2_lut_3_lut_4_lut_adj_1430.LUT_INIT = 16'h6996;
    SB_LUT4 select_715_Select_181_i2_4_lut (.I0(\data_out_frame[22] [5]), 
            .I1(\FRAME_MATCHER.i_31__N_2320 ), .I2(\current[5] ), .I3(\FRAME_MATCHER.state_31__N_2423 [3]), 
            .O(n2_adj_5241));   // verilog/coms.v(146[4] 295[11])
    defparam select_715_Select_181_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_715_Select_180_i2_4_lut (.I0(\data_out_frame[22] [4]), 
            .I1(\FRAME_MATCHER.i_31__N_2320 ), .I2(\current[4] ), .I3(\FRAME_MATCHER.state_31__N_2423 [3]), 
            .O(n2_adj_5240));   // verilog/coms.v(146[4] 295[11])
    defparam select_715_Select_180_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i11524_3_lut_4_lut (.I0(n10_adj_5280), .I1(n53712), .I2(reset), 
            .I3(n8), .O(n25127));
    defparam i11524_3_lut_4_lut.LUT_INIT = 16'hfffb;
    SB_LUT4 select_715_Select_179_i2_4_lut (.I0(\data_out_frame[22] [3]), 
            .I1(\FRAME_MATCHER.i_31__N_2320 ), .I2(\current[3] ), .I3(\FRAME_MATCHER.state_31__N_2423 [3]), 
            .O(n2_adj_5239));   // verilog/coms.v(146[4] 295[11])
    defparam select_715_Select_179_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_715_Select_178_i2_4_lut (.I0(\data_out_frame[22] [2]), 
            .I1(\FRAME_MATCHER.i_31__N_2320 ), .I2(\current[2] ), .I3(\FRAME_MATCHER.state_31__N_2423 [3]), 
            .O(n2_adj_5238));   // verilog/coms.v(146[4] 295[11])
    defparam select_715_Select_178_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_715_Select_177_i2_4_lut (.I0(\data_out_frame[22] [1]), 
            .I1(\FRAME_MATCHER.i_31__N_2320 ), .I2(\current[1] ), .I3(\FRAME_MATCHER.state_31__N_2423 [3]), 
            .O(n2_adj_5237));   // verilog/coms.v(146[4] 295[11])
    defparam select_715_Select_177_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_715_Select_176_i2_4_lut (.I0(\data_out_frame[22] [0]), 
            .I1(\FRAME_MATCHER.i_31__N_2320 ), .I2(\current[0] ), .I3(\FRAME_MATCHER.state_31__N_2423 [3]), 
            .O(n2_adj_5236));   // verilog/coms.v(146[4] 295[11])
    defparam select_715_Select_176_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_715_Select_175_i2_4_lut (.I0(\data_out_frame[21] [7]), 
            .I1(\FRAME_MATCHER.i_31__N_2320 ), .I2(\current[15] ), .I3(\FRAME_MATCHER.state_31__N_2423 [3]), 
            .O(n2_adj_5235));   // verilog/coms.v(146[4] 295[11])
    defparam select_715_Select_175_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_715_Select_174_i2_4_lut (.I0(\data_out_frame[21] [6]), 
            .I1(\FRAME_MATCHER.i_31__N_2320 ), .I2(\current[15] ), .I3(\FRAME_MATCHER.state_31__N_2423 [3]), 
            .O(n2_adj_5234));   // verilog/coms.v(146[4] 295[11])
    defparam select_715_Select_174_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_715_Select_173_i2_4_lut (.I0(\data_out_frame[21] [5]), 
            .I1(\FRAME_MATCHER.i_31__N_2320 ), .I2(\current[15] ), .I3(\FRAME_MATCHER.state_31__N_2423 [3]), 
            .O(n2_adj_5233));   // verilog/coms.v(146[4] 295[11])
    defparam select_715_Select_173_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_715_Select_172_i2_4_lut (.I0(\data_out_frame[21] [4]), 
            .I1(\FRAME_MATCHER.i_31__N_2320 ), .I2(\current[15] ), .I3(\FRAME_MATCHER.state_31__N_2423 [3]), 
            .O(n2_adj_5232));   // verilog/coms.v(146[4] 295[11])
    defparam select_715_Select_172_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_715_Select_171_i2_4_lut (.I0(\data_out_frame[21] [3]), 
            .I1(\FRAME_MATCHER.i_31__N_2320 ), .I2(\current[11] ), .I3(\FRAME_MATCHER.state_31__N_2423 [3]), 
            .O(n2_adj_5231));   // verilog/coms.v(146[4] 295[11])
    defparam select_715_Select_171_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_3_lut_4_lut_4_lut (.I0(\data_in_frame[0] [5]), .I1(\data_in_frame[0] [4]), 
            .I2(\data_in_frame[2] [5]), .I3(\data_in_frame[0] [3]), .O(n22818));   // verilog/coms.v(77[16:27])
    defparam i1_2_lut_3_lut_4_lut_4_lut.LUT_INIT = 16'ha55a;
    SB_LUT4 select_715_Select_170_i2_4_lut (.I0(\data_out_frame[21] [2]), 
            .I1(\FRAME_MATCHER.i_31__N_2320 ), .I2(\current[10] ), .I3(\FRAME_MATCHER.state_31__N_2423 [3]), 
            .O(n2_adj_5230));   // verilog/coms.v(146[4] 295[11])
    defparam select_715_Select_170_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_715_Select_169_i2_4_lut (.I0(\data_out_frame[21] [1]), 
            .I1(\FRAME_MATCHER.i_31__N_2320 ), .I2(\current[9] ), .I3(\FRAME_MATCHER.state_31__N_2423 [3]), 
            .O(n2_adj_5229));   // verilog/coms.v(146[4] 295[11])
    defparam select_715_Select_169_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_715_Select_168_i2_4_lut (.I0(\data_out_frame[21] [0]), 
            .I1(\FRAME_MATCHER.i_31__N_2320 ), .I2(\current[8] ), .I3(\FRAME_MATCHER.state_31__N_2423 [3]), 
            .O(n2_adj_5228));   // verilog/coms.v(146[4] 295[11])
    defparam select_715_Select_168_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1431 (.I0(\data_in_frame[5] [4]), .I1(\data_in_frame[3][3] ), 
            .I2(\data_in_frame[0] [7]), .I3(\data_in_frame[1] [1]), .O(n53427));
    defparam i1_2_lut_3_lut_4_lut_adj_1431.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1432 (.I0(\data_in_frame[5] [6]), .I1(\data_in_frame[6] [0]), 
            .I2(\data_in_frame[1][5] ), .I3(\data_in_frame[1][4] ), .O(n6_adj_5290));   // verilog/coms.v(77[16:43])
    defparam i1_2_lut_3_lut_4_lut_adj_1432.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1433 (.I0(\data_in_frame[1][6] ), .I1(\data_in_frame[3][7] ), 
            .I2(\data_in_frame[1][4] ), .I3(\data_in_frame[1][3] ), .O(n6_adj_5294));   // verilog/coms.v(76[16:27])
    defparam i1_2_lut_3_lut_4_lut_adj_1433.LUT_INIT = 16'h6996;
    SB_LUT4 byte_transmit_counter_2__bdd_4_lut (.I0(\byte_transmit_counter[2] ), 
            .I1(n63302), .I2(n56844), .I3(byte_transmit_counter_c[3]), 
            .O(n63371));
    defparam byte_transmit_counter_2__bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_LUT4 equal_286_i8_2_lut_3_lut (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(\FRAME_MATCHER.i [0]), .I3(GND_net), .O(n8_adj_5335));   // verilog/coms.v(154[7:23])
    defparam equal_286_i8_2_lut_3_lut.LUT_INIT = 16'hdfdf;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1434 (.I0(\data_in_frame[3] [4]), .I1(\data_in_frame[3][3] ), 
            .I2(\data_in_frame[0] [7]), .I3(\data_in_frame[1] [1]), .O(n53424));
    defparam i1_2_lut_3_lut_4_lut_adj_1434.LUT_INIT = 16'h6996;
    SB_LUT4 select_715_Select_143_i2_4_lut (.I0(\data_out_frame[17] [7]), 
            .I1(\FRAME_MATCHER.i_31__N_2320 ), .I2(pwm_setpoint[7]), .I3(\FRAME_MATCHER.state_31__N_2423 [3]), 
            .O(n2_adj_5227));   // verilog/coms.v(146[4] 295[11])
    defparam select_715_Select_143_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1435 (.I0(n23083), .I1(\data_out_frame[5] [3]), 
            .I2(\data_out_frame[5] [5]), .I3(\data_out_frame[5] [0]), .O(n52912));   // verilog/coms.v(72[16:62])
    defparam i1_2_lut_3_lut_4_lut_adj_1435.LUT_INIT = 16'h6996;
    SB_LUT4 select_715_Select_142_i2_4_lut (.I0(\data_out_frame[17] [6]), 
            .I1(\FRAME_MATCHER.i_31__N_2320 ), .I2(pwm_setpoint[6]), .I3(\FRAME_MATCHER.state_31__N_2423 [3]), 
            .O(n2_adj_5226));   // verilog/coms.v(146[4] 295[11])
    defparam select_715_Select_142_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_4_lut_adj_1436 (.I0(n54765), .I1(n47634), .I2(\data_out_frame[17] [5]), 
            .I3(n47851), .O(n48790));
    defparam i1_2_lut_4_lut_adj_1436.LUT_INIT = 16'h9669;
    SB_LUT4 i1_4_lut_adj_1437 (.I0(\FRAME_MATCHER.i_31__N_2320 ), .I1(\data_out_frame[17] [5]), 
            .I2(pwm_setpoint[5]), .I3(\FRAME_MATCHER.state_31__N_2423 [3]), 
            .O(n2_adj_5225));   // verilog/coms.v(146[4] 295[11])
    defparam i1_4_lut_adj_1437.LUT_INIT = 16'ha088;
    SB_LUT4 i5_3_lut_4_lut_adj_1438 (.I0(n47766), .I1(n33_c), .I2(\data_out_frame[17] [2]), 
            .I3(\data_out_frame[17] [3]), .O(n14_adj_5361));   // verilog/coms.v(98[12:26])
    defparam i5_3_lut_4_lut_adj_1438.LUT_INIT = 16'h6996;
    SB_LUT4 select_715_Select_140_i2_4_lut (.I0(\data_out_frame[17] [4]), 
            .I1(\FRAME_MATCHER.i_31__N_2320 ), .I2(pwm_setpoint[4]), .I3(\FRAME_MATCHER.state_31__N_2423 [3]), 
            .O(n2_adj_5224));   // verilog/coms.v(146[4] 295[11])
    defparam select_715_Select_140_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i2_3_lut_4_lut_adj_1439 (.I0(\data_out_frame[16] [4]), .I1(n47766), 
            .I2(n53574), .I3(n47853), .O(n55349));
    defparam i2_3_lut_4_lut_adj_1439.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1440 (.I0(\data_out_frame[16] [6]), .I1(\data_out_frame[16] [5]), 
            .I2(\data_out_frame[16] [7]), .I3(GND_net), .O(n4_adj_5124));
    defparam i1_2_lut_3_lut_adj_1440.LUT_INIT = 16'h9696;
    SB_LUT4 select_715_Select_139_i2_4_lut (.I0(\data_out_frame[17] [3]), 
            .I1(\FRAME_MATCHER.i_31__N_2320 ), .I2(pwm_setpoint[3]), .I3(\FRAME_MATCHER.state_31__N_2423 [3]), 
            .O(n2_adj_5223));   // verilog/coms.v(146[4] 295[11])
    defparam select_715_Select_139_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_715_Select_221_i3_2_lut_3_lut (.I0(n48239), .I1(n48259), 
            .I2(\FRAME_MATCHER.state[3] ), .I3(GND_net), .O(n3_adj_5149));   // verilog/coms.v(146[4] 295[11])
    defparam select_715_Select_221_i3_2_lut_3_lut.LUT_INIT = 16'h9090;
    SB_LUT4 select_715_Select_138_i2_4_lut (.I0(\data_out_frame[17] [2]), 
            .I1(\FRAME_MATCHER.i_31__N_2320 ), .I2(pwm_setpoint[2]), .I3(\FRAME_MATCHER.state_31__N_2423 [3]), 
            .O(n2_adj_5222));   // verilog/coms.v(146[4] 295[11])
    defparam select_715_Select_138_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1441 (.I0(\data_out_frame[16] [3]), .I1(n47750), 
            .I2(n33_c), .I3(\data_out_frame[16] [4]), .O(n47956));
    defparam i1_2_lut_3_lut_4_lut_adj_1441.LUT_INIT = 16'h6996;
    SB_LUT4 i2_2_lut_3_lut_4_lut_adj_1442 (.I0(\data_out_frame[16] [3]), .I1(n47750), 
            .I2(n47956), .I3(\data_out_frame[16] [4]), .O(n15_adj_5362));
    defparam i2_2_lut_3_lut_4_lut_adj_1442.LUT_INIT = 16'h6996;
    SB_LUT4 select_715_Select_137_i2_4_lut (.I0(\data_out_frame[17] [1]), 
            .I1(\FRAME_MATCHER.i_31__N_2320 ), .I2(pwm_setpoint[1]), .I3(\FRAME_MATCHER.state_31__N_2423 [3]), 
            .O(n2_adj_5209));   // verilog/coms.v(146[4] 295[11])
    defparam select_715_Select_137_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_3_lut_adj_1443 (.I0(\data_out_frame[16] [3]), .I1(n47750), 
            .I2(n54719), .I3(GND_net), .O(n53291));
    defparam i1_2_lut_3_lut_adj_1443.LUT_INIT = 16'h6969;
    SB_LUT4 i2_3_lut_4_lut_adj_1444 (.I0(\data_out_frame[4] [6]), .I1(\data_out_frame[5] [0]), 
            .I2(\data_out_frame[7] [2]), .I3(n52976), .O(n53397));   // verilog/coms.v(86[17:28])
    defparam i2_3_lut_4_lut_adj_1444.LUT_INIT = 16'h6996;
    SB_LUT4 select_715_Select_136_i2_4_lut (.I0(\data_out_frame[17] [0]), 
            .I1(\FRAME_MATCHER.i_31__N_2320 ), .I2(pwm_setpoint[0]), .I3(\FRAME_MATCHER.state_31__N_2423 [3]), 
            .O(n2_adj_5208));   // verilog/coms.v(146[4] 295[11])
    defparam select_715_Select_136_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 byte_transmit_counter_3__bdd_4_lut_48792 (.I0(byte_transmit_counter_c[3]), 
            .I1(n22_adj_5353), .I2(n59910), .I3(byte_transmit_counter_c[4]), 
            .O(n63533));
    defparam byte_transmit_counter_3__bdd_4_lut_48792.LUT_INIT = 16'he4aa;
    SB_LUT4 n63371_bdd_4_lut (.I0(n63371), .I1(n56864), .I2(n56863), .I3(byte_transmit_counter_c[3]), 
            .O(n63374));
    defparam n63371_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n63533_bdd_4_lut (.I0(n63533), .I1(n63326), .I2(n7_adj_5363), 
            .I3(byte_transmit_counter_c[4]), .O(tx_data[1]));
    defparam n63533_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 select_715_Select_135_i2_4_lut (.I0(\data_out_frame[16] [7]), 
            .I1(\FRAME_MATCHER.i_31__N_2320 ), .I2(pwm_setpoint[15]), .I3(\FRAME_MATCHER.state_31__N_2423 [3]), 
            .O(n2_adj_5207));   // verilog/coms.v(146[4] 295[11])
    defparam select_715_Select_135_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i2_3_lut_4_lut_adj_1445 (.I0(\data_out_frame[4] [6]), .I1(\data_out_frame[5] [0]), 
            .I2(\data_out_frame[7] [2]), .I3(\data_out_frame[5] [1]), .O(n23720));   // verilog/coms.v(86[17:28])
    defparam i2_3_lut_4_lut_adj_1445.LUT_INIT = 16'h6996;
    SB_LUT4 select_715_Select_134_i2_4_lut (.I0(\data_out_frame[16] [6]), 
            .I1(\FRAME_MATCHER.i_31__N_2320 ), .I2(pwm_setpoint[14]), .I3(\FRAME_MATCHER.state_31__N_2423 [3]), 
            .O(n2_adj_5206));   // verilog/coms.v(146[4] 295[11])
    defparam select_715_Select_134_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_4_lut_adj_1446 (.I0(n22545), .I1(n52968), .I2(\data_out_frame[14] [4]), 
            .I3(\data_out_frame[16] [6]), .O(n53094));   // verilog/coms.v(76[16:43])
    defparam i1_2_lut_4_lut_adj_1446.LUT_INIT = 16'h6996;
    SB_LUT4 select_715_Select_133_i2_4_lut (.I0(\data_out_frame[16] [5]), 
            .I1(\FRAME_MATCHER.i_31__N_2320 ), .I2(pwm_setpoint[13]), .I3(\FRAME_MATCHER.state_31__N_2423 [3]), 
            .O(n2_adj_5205));   // verilog/coms.v(146[4] 295[11])
    defparam select_715_Select_133_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_715_Select_132_i2_4_lut (.I0(\data_out_frame[16] [4]), 
            .I1(\FRAME_MATCHER.i_31__N_2320 ), .I2(pwm_setpoint[12]), .I3(\FRAME_MATCHER.state_31__N_2423 [3]), 
            .O(n2_adj_5204));   // verilog/coms.v(146[4] 295[11])
    defparam select_715_Select_132_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_4_lut_adj_1447 (.I0(\FRAME_MATCHER.i_31__N_2322 ), .I1(r_SM_Main_2__N_3318[0]), 
            .I2(tx_active), .I3(n44_adj_5364), .O(n22342));   // verilog/coms.v(146[4] 295[11])
    defparam i1_2_lut_4_lut_adj_1447.LUT_INIT = 16'ha8aa;
    SB_LUT4 i45642_2_lut (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i_31__N_2318 ), 
            .I2(GND_net), .I3(GND_net), .O(n59871));   // verilog/coms.v(155[12:15])
    defparam i45642_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i45641_2_lut (.I0(\FRAME_MATCHER.i [2]), .I1(\FRAME_MATCHER.i_31__N_2318 ), 
            .I2(GND_net), .I3(GND_net), .O(n59870));   // verilog/coms.v(155[12:15])
    defparam i45641_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i1_3_lut_4_lut (.I0(\FRAME_MATCHER.i [0]), .I1(\FRAME_MATCHER.i [4]), 
            .I2(n22428), .I3(\FRAME_MATCHER.i [1]), .O(n5_adj_5365));
    defparam i1_3_lut_4_lut.LUT_INIT = 16'hfefc;
    SB_LUT4 i45634_2_lut (.I0(\FRAME_MATCHER.i [3]), .I1(\FRAME_MATCHER.i_31__N_2318 ), 
            .I2(GND_net), .I3(GND_net), .O(n59869));   // verilog/coms.v(155[12:15])
    defparam i45634_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i46198_2_lut (.I0(\FRAME_MATCHER.i [4]), .I1(\FRAME_MATCHER.i_31__N_2318 ), 
            .I2(GND_net), .I3(GND_net), .O(n59862));   // verilog/coms.v(155[12:15])
    defparam i46198_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i45600_2_lut (.I0(\FRAME_MATCHER.i [5]), .I1(\FRAME_MATCHER.i_31__N_2318 ), 
            .I2(GND_net), .I3(GND_net), .O(n59857));   // verilog/coms.v(155[12:15])
    defparam i45600_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i45599_2_lut (.I0(\FRAME_MATCHER.i [6]), .I1(\FRAME_MATCHER.i_31__N_2318 ), 
            .I2(GND_net), .I3(GND_net), .O(n59856));   // verilog/coms.v(155[12:15])
    defparam i45599_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i1_4_lut_4_lut (.I0(n29111), .I1(\FRAME_MATCHER.i_31__N_2323 ), 
            .I2(n52615), .I3(n3302), .O(n4_adj_5347));   // verilog/coms.v(146[4] 295[11])
    defparam i1_4_lut_4_lut.LUT_INIT = 16'ha0a8;
    SB_LUT4 select_715_Select_131_i2_4_lut (.I0(\data_out_frame[16] [3]), 
            .I1(\FRAME_MATCHER.i_31__N_2320 ), .I2(pwm_setpoint[11]), .I3(\FRAME_MATCHER.state_31__N_2423 [3]), 
            .O(n2_adj_5200));   // verilog/coms.v(146[4] 295[11])
    defparam select_715_Select_131_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i45592_2_lut (.I0(\FRAME_MATCHER.i [7]), .I1(\FRAME_MATCHER.i_31__N_2318 ), 
            .I2(GND_net), .I3(GND_net), .O(n59855));   // verilog/coms.v(155[12:15])
    defparam i45592_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i1_2_lut_4_lut_adj_1448 (.I0(\FRAME_MATCHER.i_31__N_2319 ), .I1(n771), 
            .I2(\FRAME_MATCHER.i_31__N_2318 ), .I3(n22342), .O(n52615));   // verilog/coms.v(146[4] 295[11])
    defparam i1_2_lut_4_lut_adj_1448.LUT_INIT = 16'hfff2;
    SB_LUT4 i45590_2_lut (.I0(\FRAME_MATCHER.i [8]), .I1(\FRAME_MATCHER.i_31__N_2318 ), 
            .I2(GND_net), .I3(GND_net), .O(n59853));   // verilog/coms.v(155[12:15])
    defparam i45590_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_48832 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[6] [3]), .I2(\data_out_frame[7] [3]), .I3(byte_transmit_counter_c[1]), 
            .O(n63527));
    defparam byte_transmit_counter_0__bdd_4_lut_48832.LUT_INIT = 16'he4aa;
    SB_LUT4 i1_2_lut_4_lut_adj_1449 (.I0(n22545), .I1(n52968), .I2(\data_out_frame[14] [4]), 
            .I3(\data_out_frame[16] [5]), .O(n53574));   // verilog/coms.v(76[16:43])
    defparam i1_2_lut_4_lut_adj_1449.LUT_INIT = 16'h6996;
    SB_LUT4 n63527_bdd_4_lut (.I0(n63527), .I1(\data_out_frame[5] [3]), 
            .I2(\data_out_frame[4] [3]), .I3(byte_transmit_counter_c[1]), 
            .O(n56864));
    defparam n63527_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i41900_3_lut_4_lut (.I0(n23252), .I1(\data_in_frame[2] [7]), 
            .I2(\data_in_frame[0] [6]), .I3(\data_in_frame[0] [5]), .O(n56597));
    defparam i41900_3_lut_4_lut.LUT_INIT = 16'hebbe;
    SB_LUT4 i7_3_lut_4_lut (.I0(Kp_23__N_583), .I1(n23201), .I2(\data_in_frame[0] [0]), 
            .I3(\data_in_frame[1][7] ), .O(n24_adj_5366));
    defparam i7_3_lut_4_lut.LUT_INIT = 16'h2112;
    SB_LUT4 select_715_Select_130_i2_4_lut (.I0(\data_out_frame[16] [2]), 
            .I1(\FRAME_MATCHER.i_31__N_2320 ), .I2(pwm_setpoint[10]), .I3(\FRAME_MATCHER.state_31__N_2423 [3]), 
            .O(n2_adj_5199));   // verilog/coms.v(146[4] 295[11])
    defparam select_715_Select_130_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i45582_2_lut (.I0(\FRAME_MATCHER.i [9]), .I1(\FRAME_MATCHER.i_31__N_2318 ), 
            .I2(GND_net), .I3(GND_net), .O(n59850));   // verilog/coms.v(155[12:15])
    defparam i45582_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i1_2_lut_3_lut_adj_1450 (.I0(\data_in_frame[2] [5]), .I1(\data_in_frame[0] [4]), 
            .I2(\data_in_frame[0] [3]), .I3(GND_net), .O(n23201));   // verilog/coms.v(75[16:43])
    defparam i1_2_lut_3_lut_adj_1450.LUT_INIT = 16'h9696;
    SB_LUT4 select_715_Select_129_i2_4_lut (.I0(\data_out_frame[16] [1]), 
            .I1(\FRAME_MATCHER.i_31__N_2320 ), .I2(pwm_setpoint[9]), .I3(\FRAME_MATCHER.state_31__N_2423 [3]), 
            .O(n2_adj_5198));   // verilog/coms.v(146[4] 295[11])
    defparam select_715_Select_129_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_715_Select_128_i2_4_lut (.I0(\data_out_frame[16] [0]), 
            .I1(\FRAME_MATCHER.i_31__N_2320 ), .I2(pwm_setpoint[8]), .I3(\FRAME_MATCHER.state_31__N_2423 [3]), 
            .O(n2_adj_5197));   // verilog/coms.v(146[4] 295[11])
    defparam select_715_Select_128_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_715_Select_127_i2_4_lut (.I0(\data_out_frame[15] [7]), 
            .I1(\FRAME_MATCHER.i_31__N_2320 ), .I2(pwm_setpoint[23]), .I3(\FRAME_MATCHER.state_31__N_2423 [3]), 
            .O(n2_adj_5196));   // verilog/coms.v(146[4] 295[11])
    defparam select_715_Select_127_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_715_Select_126_i2_4_lut (.I0(\data_out_frame[15] [6]), 
            .I1(\FRAME_MATCHER.i_31__N_2320 ), .I2(pwm_setpoint[22]), .I3(\FRAME_MATCHER.state_31__N_2423 [3]), 
            .O(n2_adj_5195));   // verilog/coms.v(146[4] 295[11])
    defparam select_715_Select_126_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_715_Select_125_i2_4_lut (.I0(\data_out_frame[15] [5]), 
            .I1(\FRAME_MATCHER.i_31__N_2320 ), .I2(pwm_setpoint[21]), .I3(\FRAME_MATCHER.state_31__N_2423 [3]), 
            .O(n2_adj_5194));   // verilog/coms.v(146[4] 295[11])
    defparam select_715_Select_125_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_715_Select_124_i2_4_lut (.I0(\data_out_frame[15] [4]), 
            .I1(\FRAME_MATCHER.i_31__N_2320 ), .I2(pwm_setpoint[20]), .I3(\FRAME_MATCHER.state_31__N_2423 [3]), 
            .O(n2_adj_5193));   // verilog/coms.v(146[4] 295[11])
    defparam select_715_Select_124_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_715_Select_123_i2_4_lut (.I0(\data_out_frame[15] [3]), 
            .I1(\FRAME_MATCHER.i_31__N_2320 ), .I2(pwm_setpoint[19]), .I3(\FRAME_MATCHER.state_31__N_2423 [3]), 
            .O(n2_adj_5192));   // verilog/coms.v(146[4] 295[11])
    defparam select_715_Select_123_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_715_Select_122_i2_4_lut (.I0(\data_out_frame[15] [2]), 
            .I1(\FRAME_MATCHER.i_31__N_2320 ), .I2(pwm_setpoint[18]), .I3(\FRAME_MATCHER.state_31__N_2423 [3]), 
            .O(n2_adj_5191));   // verilog/coms.v(146[4] 295[11])
    defparam select_715_Select_122_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_715_Select_121_i2_4_lut (.I0(\data_out_frame[15] [1]), 
            .I1(\FRAME_MATCHER.i_31__N_2320 ), .I2(pwm_setpoint[17]), .I3(\FRAME_MATCHER.state_31__N_2423 [3]), 
            .O(n2_adj_5190));   // verilog/coms.v(146[4] 295[11])
    defparam select_715_Select_121_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_715_Select_120_i2_4_lut (.I0(\data_out_frame[15] [0]), 
            .I1(\FRAME_MATCHER.i_31__N_2320 ), .I2(pwm_setpoint[16]), .I3(\FRAME_MATCHER.state_31__N_2423 [3]), 
            .O(n2_adj_5189));   // verilog/coms.v(146[4] 295[11])
    defparam select_715_Select_120_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_715_Select_119_i2_4_lut (.I0(\data_out_frame[14] [7]), 
            .I1(\FRAME_MATCHER.i_31__N_2320 ), .I2(setpoint[7]), .I3(\FRAME_MATCHER.state_31__N_2423 [3]), 
            .O(n2_adj_5188));   // verilog/coms.v(146[4] 295[11])
    defparam select_715_Select_119_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_715_Select_118_i2_4_lut (.I0(\data_out_frame[14] [6]), 
            .I1(\FRAME_MATCHER.i_31__N_2320 ), .I2(setpoint[6]), .I3(\FRAME_MATCHER.state_31__N_2423 [3]), 
            .O(n2_adj_5187));   // verilog/coms.v(146[4] 295[11])
    defparam select_715_Select_118_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_3_lut_adj_1451 (.I0(\data_in_frame[2] [3]), .I1(\data_in_frame[0] [1]), 
            .I2(\data_in_frame[0] [2]), .I3(GND_net), .O(n23252));   // verilog/coms.v(166[9:87])
    defparam i1_2_lut_3_lut_adj_1451.LUT_INIT = 16'h9696;
    SB_LUT4 select_715_Select_117_i2_4_lut (.I0(\data_out_frame[14] [5]), 
            .I1(\FRAME_MATCHER.i_31__N_2320 ), .I2(setpoint[5]), .I3(\FRAME_MATCHER.state_31__N_2423 [3]), 
            .O(n2_adj_5186));   // verilog/coms.v(146[4] 295[11])
    defparam select_715_Select_117_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_715_Select_116_i2_4_lut (.I0(\data_out_frame[14] [4]), 
            .I1(\FRAME_MATCHER.i_31__N_2320 ), .I2(setpoint[4]), .I3(\FRAME_MATCHER.state_31__N_2423 [3]), 
            .O(n2_adj_5185));   // verilog/coms.v(146[4] 295[11])
    defparam select_715_Select_116_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_715_Select_115_i2_4_lut (.I0(\data_out_frame[14] [3]), 
            .I1(\FRAME_MATCHER.i_31__N_2320 ), .I2(setpoint[3]), .I3(\FRAME_MATCHER.state_31__N_2423 [3]), 
            .O(n2_adj_5184));   // verilog/coms.v(146[4] 295[11])
    defparam select_715_Select_115_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i45581_2_lut (.I0(\FRAME_MATCHER.i [10]), .I1(\FRAME_MATCHER.i_31__N_2318 ), 
            .I2(GND_net), .I3(GND_net), .O(n59849));   // verilog/coms.v(155[12:15])
    defparam i45581_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 select_715_Select_114_i2_4_lut (.I0(\data_out_frame[14] [2]), 
            .I1(\FRAME_MATCHER.i_31__N_2320 ), .I2(setpoint[2]), .I3(\FRAME_MATCHER.state_31__N_2423 [3]), 
            .O(n2_adj_5183));   // verilog/coms.v(146[4] 295[11])
    defparam select_715_Select_114_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_4_lut_adj_1452 (.I0(\FRAME_MATCHER.i_31__N_2320 ), .I1(\data_out_frame[14] [1]), 
            .I2(setpoint[1]), .I3(\FRAME_MATCHER.state_31__N_2423 [3]), 
            .O(n2_adj_5182));   // verilog/coms.v(146[4] 295[11])
    defparam i1_4_lut_adj_1452.LUT_INIT = 16'ha088;
    SB_LUT4 select_715_Select_112_i2_4_lut (.I0(\data_out_frame[14] [0]), 
            .I1(\FRAME_MATCHER.i_31__N_2320 ), .I2(setpoint[0]), .I3(\FRAME_MATCHER.state_31__N_2423 [3]), 
            .O(n2_adj_5181));   // verilog/coms.v(146[4] 295[11])
    defparam select_715_Select_112_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_715_Select_111_i2_4_lut (.I0(\data_out_frame[13] [7]), 
            .I1(\FRAME_MATCHER.i_31__N_2320 ), .I2(setpoint[15]), .I3(\FRAME_MATCHER.state_31__N_2423 [3]), 
            .O(n2_adj_5180));   // verilog/coms.v(146[4] 295[11])
    defparam select_715_Select_111_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_715_Select_110_i2_4_lut (.I0(\data_out_frame[13] [6]), 
            .I1(\FRAME_MATCHER.i_31__N_2320 ), .I2(setpoint[14]), .I3(\FRAME_MATCHER.state_31__N_2423 [3]), 
            .O(n2_adj_5179));   // verilog/coms.v(146[4] 295[11])
    defparam select_715_Select_110_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_715_Select_109_i2_4_lut (.I0(\data_out_frame[13] [5]), 
            .I1(\FRAME_MATCHER.i_31__N_2320 ), .I2(setpoint[13]), .I3(\FRAME_MATCHER.state_31__N_2423 [3]), 
            .O(n2_adj_5178));   // verilog/coms.v(146[4] 295[11])
    defparam select_715_Select_109_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_715_Select_108_i2_4_lut (.I0(\data_out_frame[13] [4]), 
            .I1(\FRAME_MATCHER.i_31__N_2320 ), .I2(setpoint[12]), .I3(\FRAME_MATCHER.state_31__N_2423 [3]), 
            .O(n2_adj_5177));   // verilog/coms.v(146[4] 295[11])
    defparam select_715_Select_108_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i45580_2_lut (.I0(\FRAME_MATCHER.i [11]), .I1(\FRAME_MATCHER.i_31__N_2318 ), 
            .I2(GND_net), .I3(GND_net), .O(n59848));   // verilog/coms.v(155[12:15])
    defparam i45580_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i45579_2_lut (.I0(\FRAME_MATCHER.i [12]), .I1(\FRAME_MATCHER.i_31__N_2318 ), 
            .I2(GND_net), .I3(GND_net), .O(n59847));   // verilog/coms.v(155[12:15])
    defparam i45579_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i45578_2_lut (.I0(\FRAME_MATCHER.i [13]), .I1(\FRAME_MATCHER.i_31__N_2318 ), 
            .I2(GND_net), .I3(GND_net), .O(n59846));   // verilog/coms.v(155[12:15])
    defparam i45578_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i45552_2_lut (.I0(\FRAME_MATCHER.i [14]), .I1(\FRAME_MATCHER.i_31__N_2318 ), 
            .I2(GND_net), .I3(GND_net), .O(n59845));   // verilog/coms.v(155[12:15])
    defparam i45552_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i45573_2_lut (.I0(\FRAME_MATCHER.i [15]), .I1(\FRAME_MATCHER.i_31__N_2318 ), 
            .I2(GND_net), .I3(GND_net), .O(n59844));   // verilog/coms.v(155[12:15])
    defparam i45573_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i45543_2_lut (.I0(\FRAME_MATCHER.i [16]), .I1(\FRAME_MATCHER.i_31__N_2318 ), 
            .I2(GND_net), .I3(GND_net), .O(n59841));   // verilog/coms.v(155[12:15])
    defparam i45543_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i45542_2_lut (.I0(\FRAME_MATCHER.i [17]), .I1(\FRAME_MATCHER.i_31__N_2318 ), 
            .I2(GND_net), .I3(GND_net), .O(n59840));   // verilog/coms.v(155[12:15])
    defparam i45542_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i45594_2_lut (.I0(\FRAME_MATCHER.i [18]), .I1(\FRAME_MATCHER.i_31__N_2318 ), 
            .I2(GND_net), .I3(GND_net), .O(n59838));   // verilog/coms.v(155[12:15])
    defparam i45594_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i45534_2_lut (.I0(\FRAME_MATCHER.i [19]), .I1(\FRAME_MATCHER.i_31__N_2318 ), 
            .I2(GND_net), .I3(GND_net), .O(n59829));   // verilog/coms.v(155[12:15])
    defparam i45534_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 select_715_Select_107_i2_4_lut (.I0(\data_out_frame[13] [3]), 
            .I1(\FRAME_MATCHER.i_31__N_2320 ), .I2(setpoint[11]), .I3(\FRAME_MATCHER.state_31__N_2423 [3]), 
            .O(n2_adj_5176));   // verilog/coms.v(146[4] 295[11])
    defparam select_715_Select_107_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_715_Select_106_i2_4_lut (.I0(\data_out_frame[13] [2]), 
            .I1(\FRAME_MATCHER.i_31__N_2320 ), .I2(setpoint[10]), .I3(\FRAME_MATCHER.state_31__N_2423 [3]), 
            .O(n2_adj_5175));   // verilog/coms.v(146[4] 295[11])
    defparam select_715_Select_106_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i45514_2_lut (.I0(\FRAME_MATCHER.i [20]), .I1(\FRAME_MATCHER.i_31__N_2318 ), 
            .I2(GND_net), .I3(GND_net), .O(n59816));   // verilog/coms.v(155[12:15])
    defparam i45514_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 select_715_Select_4_i2_3_lut (.I0(\data_out_frame[0][4] ), .I1(\FRAME_MATCHER.i_31__N_2320 ), 
            .I2(\FRAME_MATCHER.state_31__N_2423 [3]), .I3(GND_net), .O(n2_adj_5053));   // verilog/coms.v(146[4] 295[11])
    defparam select_715_Select_4_i2_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i1_4_lut_adj_1453 (.I0(\FRAME_MATCHER.i_31__N_2320 ), .I1(\data_out_frame[13] [1]), 
            .I2(setpoint[9]), .I3(\FRAME_MATCHER.state_31__N_2423 [3]), 
            .O(n2_adj_5174));   // verilog/coms.v(146[4] 295[11])
    defparam i1_4_lut_adj_1453.LUT_INIT = 16'ha088;
    SB_LUT4 select_715_Select_104_i2_4_lut (.I0(\data_out_frame[13] [0]), 
            .I1(\FRAME_MATCHER.i_31__N_2320 ), .I2(setpoint[8]), .I3(\FRAME_MATCHER.state_31__N_2423 [3]), 
            .O(n2_adj_5173));   // verilog/coms.v(146[4] 295[11])
    defparam select_715_Select_104_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_715_Select_103_i2_4_lut (.I0(\data_out_frame[12] [7]), 
            .I1(\FRAME_MATCHER.i_31__N_2320 ), .I2(setpoint[23]), .I3(\FRAME_MATCHER.state_31__N_2423 [3]), 
            .O(n2_adj_5172));   // verilog/coms.v(146[4] 295[11])
    defparam select_715_Select_103_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_715_Select_102_i2_4_lut (.I0(\data_out_frame[12] [6]), 
            .I1(\FRAME_MATCHER.i_31__N_2320 ), .I2(setpoint[22]), .I3(\FRAME_MATCHER.state_31__N_2423 [3]), 
            .O(n2_adj_5171));   // verilog/coms.v(146[4] 295[11])
    defparam select_715_Select_102_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_715_Select_101_i2_4_lut (.I0(\data_out_frame[12] [5]), 
            .I1(\FRAME_MATCHER.i_31__N_2320 ), .I2(setpoint[21]), .I3(\FRAME_MATCHER.state_31__N_2423 [3]), 
            .O(n2_adj_5170));   // verilog/coms.v(146[4] 295[11])
    defparam select_715_Select_101_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_715_Select_100_i2_4_lut (.I0(\data_out_frame[12] [4]), 
            .I1(\FRAME_MATCHER.i_31__N_2320 ), .I2(setpoint[20]), .I3(\FRAME_MATCHER.state_31__N_2423 [3]), 
            .O(n2_adj_5169));   // verilog/coms.v(146[4] 295[11])
    defparam select_715_Select_100_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i45513_2_lut (.I0(\FRAME_MATCHER.i [21]), .I1(\FRAME_MATCHER.i_31__N_2318 ), 
            .I2(GND_net), .I3(GND_net), .O(n59815));   // verilog/coms.v(155[12:15])
    defparam i45513_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i45508_2_lut (.I0(\FRAME_MATCHER.i [22]), .I1(\FRAME_MATCHER.i_31__N_2318 ), 
            .I2(GND_net), .I3(GND_net), .O(n59814));   // verilog/coms.v(155[12:15])
    defparam i45508_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i45502_2_lut (.I0(\FRAME_MATCHER.i [23]), .I1(\FRAME_MATCHER.i_31__N_2318 ), 
            .I2(GND_net), .I3(GND_net), .O(n59813));   // verilog/coms.v(155[12:15])
    defparam i45502_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 select_715_Select_3_i2_3_lut (.I0(\data_out_frame[0][3] ), .I1(\FRAME_MATCHER.i_31__N_2320 ), 
            .I2(\FRAME_MATCHER.state_31__N_2423 [3]), .I3(GND_net), .O(n2_adj_5052));   // verilog/coms.v(146[4] 295[11])
    defparam select_715_Select_3_i2_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i1_2_lut_adj_1454 (.I0(\data_in_frame[0] [6]), .I1(\data_in_frame[0] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n52983));   // verilog/coms.v(78[16:27])
    defparam i1_2_lut_adj_1454.LUT_INIT = 16'h6666;
    SB_LUT4 i11147_3_lut (.I0(\data_out_frame[1][7] ), .I1(\data_out_frame[3][7] ), 
            .I2(byte_transmit_counter_c[1]), .I3(GND_net), .O(n24745));   // verilog/coms.v(107[34:55])
    defparam i11147_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i42221_3_lut (.I0(\data_out_frame[6] [7]), .I1(\data_out_frame[7] [7]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n56933));
    defparam i42221_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i42222_4_lut (.I0(n56933), .I1(n24745), .I2(\byte_transmit_counter[2] ), 
            .I3(byte_transmit_counter[0]), .O(n56934));
    defparam i42222_4_lut.LUT_INIT = 16'haca0;
    SB_LUT4 i42220_3_lut (.I0(\data_out_frame[4] [7]), .I1(\data_out_frame[5] [7]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n56932));
    defparam i42220_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2227084_i1_3_lut (.I0(n63338), .I1(n63284), .I2(\byte_transmit_counter[2] ), 
            .I3(GND_net), .O(n14_adj_5167));
    defparam i2227084_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i46177_4_lut (.I0(\data_out_frame[26] [7]), .I1(n24840), .I2(\data_out_frame[27] [7]), 
            .I3(byte_transmit_counter[0]), .O(n59919));
    defparam i46177_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_adj_1455 (.I0(\data_in_frame[0] [1]), .I1(\data_in_frame[0] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n53122));   // verilog/coms.v(166[9:87])
    defparam i1_2_lut_adj_1455.LUT_INIT = 16'h6666;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_7_i21_4_lut (.I0(\data_out_frame[21] [7]), 
            .I1(\data_out_frame[22] [7]), .I2(byte_transmit_counter_c[1]), 
            .I3(byte_transmit_counter[0]), .O(n21_adj_5367));   // verilog/coms.v(107[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_7_i21_4_lut.LUT_INIT = 16'h0ac0;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_7_i16_3_lut (.I0(\data_out_frame[16] [7]), 
            .I1(\data_out_frame[17] [7]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n16_adj_5368));   // verilog/coms.v(107[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_7_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_7_i22_4_lut (.I0(n16_adj_5368), 
            .I1(n21_adj_5367), .I2(\byte_transmit_counter[2] ), .I3(byte_transmit_counter_c[1]), 
            .O(n22_adj_5166));   // verilog/coms.v(107[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_7_i22_4_lut.LUT_INIT = 16'hc0ca;
    SB_LUT4 select_715_Select_55_i2_4_lut (.I0(\data_out_frame[6] [7]), .I1(\FRAME_MATCHER.i_31__N_2320 ), 
            .I2(encoder0_position[23]), .I3(\FRAME_MATCHER.state_31__N_2423 [3]), 
            .O(n2_adj_5165));   // verilog/coms.v(146[4] 295[11])
    defparam select_715_Select_55_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_715_Select_54_i2_4_lut (.I0(\data_out_frame[6] [6]), .I1(\FRAME_MATCHER.i_31__N_2320 ), 
            .I2(encoder0_position[22]), .I3(\FRAME_MATCHER.state_31__N_2423 [3]), 
            .O(n2_adj_5164));   // verilog/coms.v(146[4] 295[11])
    defparam select_715_Select_54_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_715_Select_53_i2_4_lut (.I0(\data_out_frame[6] [5]), .I1(\FRAME_MATCHER.i_31__N_2320 ), 
            .I2(encoder0_position[21]), .I3(\FRAME_MATCHER.state_31__N_2423 [3]), 
            .O(n2_adj_5163));   // verilog/coms.v(146[4] 295[11])
    defparam select_715_Select_53_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_715_Select_52_i2_4_lut (.I0(\data_out_frame[6] [4]), .I1(\FRAME_MATCHER.i_31__N_2320 ), 
            .I2(encoder0_position[20]), .I3(\FRAME_MATCHER.state_31__N_2423 [3]), 
            .O(n2_adj_5162));   // verilog/coms.v(146[4] 295[11])
    defparam select_715_Select_52_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_adj_1456 (.I0(\data_in_frame[0] [6]), .I1(\data_in_frame[1] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n53201));   // verilog/coms.v(71[16:27])
    defparam i1_2_lut_adj_1456.LUT_INIT = 16'h6666;
    SB_LUT4 i1_4_lut_adj_1457 (.I0(n24840), .I1(\data_out_frame[26] [2]), 
            .I2(\data_out_frame[27] [2]), .I3(byte_transmit_counter[0]), 
            .O(n33004));   // verilog/coms.v(107[34:55])
    defparam i1_4_lut_adj_1457.LUT_INIT = 16'ha088;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_2_i16_3_lut (.I0(\data_out_frame[16] [2]), 
            .I1(\data_out_frame[17] [2]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n16_adj_5369));   // verilog/coms.v(107[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_2_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i42238_4_lut (.I0(\data_out_frame[0][2] ), .I1(n16_adj_5369), 
            .I2(byte_transmit_counter_c[4]), .I3(byte_transmit_counter[0]), 
            .O(n61082));
    defparam i42238_4_lut.LUT_INIT = 16'hc0ca;
    SB_LUT4 i42202_3_lut (.I0(\data_out_frame[8] [2]), .I1(\data_out_frame[9] [2]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n56914));
    defparam i42202_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2_3_lut_adj_1458 (.I0(\data_in_frame[2] [2]), .I1(\data_in_frame[0] [0]), 
            .I2(\data_in_frame[0] [1]), .I3(GND_net), .O(n23221));   // verilog/coms.v(166[9:87])
    defparam i2_3_lut_adj_1458.LUT_INIT = 16'h9696;
    SB_LUT4 i4_4_lut_adj_1459 (.I0(\data_in_frame[0] [4]), .I1(\data_in_frame[0] [6]), 
            .I2(ID[4]), .I3(ID[6]), .O(n12_adj_5370));   // verilog/coms.v(237[12:32])
    defparam i4_4_lut_adj_1459.LUT_INIT = 16'h7bde;
    SB_LUT4 i2_4_lut_adj_1460 (.I0(\data_in_frame[0] [1]), .I1(\data_in_frame[0] [2]), 
            .I2(ID[1]), .I3(ID[2]), .O(n10_adj_5371));   // verilog/coms.v(237[12:32])
    defparam i2_4_lut_adj_1460.LUT_INIT = 16'h7bde;
    SB_LUT4 i42203_3_lut (.I0(\data_out_frame[10] [2]), .I1(\data_out_frame[11] [2]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n56915));
    defparam i42203_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i42239_4_lut (.I0(n56914), .I1(byte_transmit_counter_c[1]), 
            .I2(byte_transmit_counter_c[3]), .I3(n61082), .O(n56951));
    defparam i42239_4_lut.LUT_INIT = 16'ha3a0;
    SB_LUT4 i2_3_lut_4_lut_adj_1461 (.I0(\data_in_frame[0] [5]), .I1(\data_in_frame[0] [4]), 
            .I2(\data_in_frame[7] [4]), .I3(n23046), .O(n53571));   // verilog/coms.v(77[16:27])
    defparam i2_3_lut_4_lut_adj_1461.LUT_INIT = 16'h6996;
    SB_LUT4 i42204_3_lut (.I0(n56915), .I1(n33004), .I2(byte_transmit_counter_c[4]), 
            .I3(GND_net), .O(n56916));
    defparam i42204_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i42240_3_lut (.I0(n56916), .I1(n56951), .I2(n57324), .I3(GND_net), 
            .O(n56952));
    defparam i42240_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i22306102_i1_3_lut (.I0(n56952), .I1(n63296), .I2(\byte_transmit_counter[2] ), 
            .I3(GND_net), .O(tx_data[2]));
    defparam i22306102_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3_4_lut_adj_1462 (.I0(\data_in_frame[0] [7]), .I1(\data_in_frame[0] [5]), 
            .I2(ID[7]), .I3(ID[5]), .O(n11));   // verilog/coms.v(237[12:32])
    defparam i3_4_lut_adj_1462.LUT_INIT = 16'h7bde;
    SB_LUT4 equal_1931_i7_2_lut_3_lut (.I0(\data_in_frame[0] [5]), .I1(\data_in_frame[0] [4]), 
            .I2(\data_in_frame[2] [6]), .I3(GND_net), .O(n7_adj_5277));   // verilog/coms.v(77[16:27])
    defparam equal_1931_i7_2_lut_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_3_i21_4_lut (.I0(\data_out_frame[21] [3]), 
            .I1(\data_out_frame[22] [3]), .I2(byte_transmit_counter_c[1]), 
            .I3(byte_transmit_counter[0]), .O(n21_adj_5372));   // verilog/coms.v(107[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_3_i21_4_lut.LUT_INIT = 16'h0ac0;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_3_i16_3_lut (.I0(\data_out_frame[16] [3]), 
            .I1(\data_out_frame[17] [3]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n16_adj_5373));   // verilog/coms.v(107[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_3_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_3_i24_3_lut (.I0(\data_out_frame[26] [3]), 
            .I1(\data_out_frame[27] [3]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n24_adj_5374));   // verilog/coms.v(107[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_3_i24_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_3_i22_4_lut (.I0(n16_adj_5373), 
            .I1(n21_adj_5372), .I2(\byte_transmit_counter[2] ), .I3(byte_transmit_counter_c[1]), 
            .O(n22_adj_5375));   // verilog/coms.v(107[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_3_i22_4_lut.LUT_INIT = 16'hc0ca;
    SB_LUT4 i42368_4_lut (.I0(n22_adj_5375), .I1(n24_adj_5374), .I2(byte_transmit_counter_c[3]), 
            .I3(n24840), .O(n57080));
    defparam i42368_4_lut.LUT_INIT = 16'hca0a;
    SB_LUT4 i42369_3_lut (.I0(n63374), .I1(n57080), .I2(byte_transmit_counter_c[4]), 
            .I3(GND_net), .O(tx_data[3]));
    defparam i42369_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_6_i7_3_lut_4_lut (.I0(\byte_transmit_counter[2] ), 
            .I1(byte_transmit_counter_c[1]), .I2(n56928), .I3(n56926), 
            .O(n7_adj_5376));   // verilog/coms.v(107[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_6_i7_3_lut_4_lut.LUT_INIT = 16'hf2d0;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_1_i7_3_lut_4_lut (.I0(\byte_transmit_counter[2] ), 
            .I1(byte_transmit_counter_c[1]), .I2(n56931), .I3(n56929), 
            .O(n7_adj_5363));   // verilog/coms.v(107[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_1_i7_3_lut_4_lut.LUT_INIT = 16'hf2d0;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_4_i21_4_lut (.I0(\data_out_frame[21] [4]), 
            .I1(\data_out_frame[22] [4]), .I2(byte_transmit_counter_c[1]), 
            .I3(byte_transmit_counter[0]), .O(n21_adj_5377));   // verilog/coms.v(107[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_4_i21_4_lut.LUT_INIT = 16'h0ac0;
    SB_LUT4 i1_4_lut_adj_1463 (.I0(\data_in_frame[0] [0]), .I1(\data_in_frame[0] [3]), 
            .I2(ID[0]), .I3(ID[3]), .O(n9_adj_5378));   // verilog/coms.v(237[12:32])
    defparam i1_4_lut_adj_1463.LUT_INIT = 16'h7bde;
    SB_LUT4 i7_4_lut_adj_1464 (.I0(n9_adj_5378), .I1(n11), .I2(n10_adj_5371), 
            .I3(n12_adj_5370), .O(n55426));   // verilog/coms.v(237[12:32])
    defparam i7_4_lut_adj_1464.LUT_INIT = 16'hfffe;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_4_i16_3_lut (.I0(\data_out_frame[16] [4]), 
            .I1(\data_out_frame[17] [4]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n16_adj_5379));   // verilog/coms.v(107[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_4_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_4_i24_3_lut (.I0(\data_out_frame[26] [4]), 
            .I1(\data_out_frame[27] [4]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n24_adj_5380));   // verilog/coms.v(107[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_4_i24_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_4_i22_4_lut (.I0(n16_adj_5379), 
            .I1(n21_adj_5377), .I2(\byte_transmit_counter[2] ), .I3(byte_transmit_counter_c[1]), 
            .O(n22_adj_5381));   // verilog/coms.v(107[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_4_i22_4_lut.LUT_INIT = 16'hc0ca;
    SB_LUT4 i1_2_lut_adj_1465 (.I0(\data_in_frame[2] [0]), .I1(Kp_23__N_583), 
            .I2(GND_net), .I3(GND_net), .O(n53141));   // verilog/coms.v(71[16:69])
    defparam i1_2_lut_adj_1465.LUT_INIT = 16'h6666;
    SB_LUT4 i42134_4_lut (.I0(n22_adj_5381), .I1(n24_adj_5380), .I2(byte_transmit_counter_c[3]), 
            .I3(n24840), .O(n56846));
    defparam i42134_4_lut.LUT_INIT = 16'hca0a;
    SB_LUT4 i42135_3_lut (.I0(n63290), .I1(n56846), .I2(byte_transmit_counter_c[4]), 
            .I3(GND_net), .O(tx_data[4]));
    defparam i42135_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 equal_1931_i10_2_lut (.I0(\data_in_frame[0] [7]), .I1(\data_in_frame[1] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n10_adj_5382));   // verilog/coms.v(166[9:87])
    defparam equal_1931_i10_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i10_3_lut_4_lut (.I0(\byte_transmit_counter[2] ), .I1(byte_transmit_counter_c[1]), 
            .I2(n56919), .I3(n56917), .O(n7_adj_5358));   // verilog/coms.v(107[34:55])
    defparam i10_3_lut_4_lut.LUT_INIT = 16'hf2d0;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_7_i7_3_lut_4_lut (.I0(\byte_transmit_counter[2] ), 
            .I1(byte_transmit_counter_c[1]), .I2(n56934), .I3(n56932), 
            .O(n7_adj_5168));   // verilog/coms.v(107[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_7_i7_3_lut_4_lut.LUT_INIT = 16'hf2d0;
    SB_LUT4 i2_3_lut_adj_1466 (.I0(\data_in_frame[0] [3]), .I1(\data_in_frame[0] [2]), 
            .I2(\data_in_frame[2] [4]), .I3(GND_net), .O(n23536));   // verilog/coms.v(75[16:43])
    defparam i2_3_lut_adj_1466.LUT_INIT = 16'h9696;
    SB_LUT4 i42612_3_lut (.I0(byte_transmit_counter_c[3]), .I1(byte_transmit_counter_c[4]), 
            .I2(byte_transmit_counter_c[1]), .I3(GND_net), .O(n57324));
    defparam i42612_3_lut.LUT_INIT = 16'ha8a8;
    SB_LUT4 i1_2_lut_adj_1467 (.I0(\data_in_frame[0] [4]), .I1(\data_in_frame[0] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n52956));   // verilog/coms.v(75[16:43])
    defparam i1_2_lut_adj_1467.LUT_INIT = 16'h6666;
    SB_LUT4 i11160_2_lut (.I0(byte_transmit_counter_c[1]), .I1(\byte_transmit_counter[2] ), 
            .I2(GND_net), .I3(GND_net), .O(n24840));   // verilog/coms.v(107[34:55])
    defparam i11160_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i1_4_lut_adj_1468 (.I0(n24840), .I1(\data_out_frame[26] [5]), 
            .I2(\data_out_frame[27] [5]), .I3(byte_transmit_counter[0]), 
            .O(n33453));   // verilog/coms.v(107[34:55])
    defparam i1_4_lut_adj_1468.LUT_INIT = 16'ha088;
    SB_LUT4 i1_2_lut_adj_1469 (.I0(byte_transmit_counter[0]), .I1(byte_transmit_counter_c[1]), 
            .I2(GND_net), .I3(GND_net), .O(n24853));   // verilog/coms.v(128[12] 296[6])
    defparam i1_2_lut_adj_1469.LUT_INIT = 16'hdddd;
    SB_LUT4 i1_2_lut_adj_1470 (.I0(\data_in_frame[0] [0]), .I1(\data_in_frame[1][7] ), 
            .I2(GND_net), .I3(GND_net), .O(n53186));   // verilog/coms.v(71[16:69])
    defparam i1_2_lut_adj_1470.LUT_INIT = 16'h6666;
    SB_LUT4 i42208_3_lut (.I0(\data_out_frame[8] [5]), .I1(\data_out_frame[9] [5]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n56920));
    defparam i42208_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3_4_lut_adj_1471 (.I0(\data_in_frame[0] [7]), .I1(n53122), 
            .I2(n52983), .I3(n52956), .O(Kp_23__N_583));   // verilog/coms.v(71[16:27])
    defparam i3_4_lut_adj_1471.LUT_INIT = 16'h6996;
    SB_LUT4 i42209_3_lut (.I0(\data_out_frame[10] [5]), .I1(\data_out_frame[11] [5]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n56921));
    defparam i42209_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i42210_3_lut (.I0(n56921), .I1(n33453), .I2(byte_transmit_counter_c[4]), 
            .I3(GND_net), .O(n56922));
    defparam i42210_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i5_3_lut_adj_1472 (.I0(n23536), .I1(Kp_23__N_583), .I2(\data_in_frame[2] [1]), 
            .I3(GND_net), .O(n22_adj_5383));
    defparam i5_3_lut_adj_1472.LUT_INIT = 16'h1414;
    SB_LUT4 i10_4_lut_adj_1473 (.I0(\data_in_frame[1][4] ), .I1(\data_in_frame[1][3] ), 
            .I2(\data_in_frame[1][2] ), .I3(\data_in_frame[1][6] ), .O(n27_adj_5384));
    defparam i10_4_lut_adj_1473.LUT_INIT = 16'h8000;
    SB_LUT4 i9_4_lut_adj_1474 (.I0(\data_in_frame[0] [0]), .I1(n10_adj_5382), 
            .I2(n53141), .I3(\data_in_frame[1][5] ), .O(n26_adj_5385));
    defparam i9_4_lut_adj_1474.LUT_INIT = 16'h2100;
    SB_LUT4 select_715_Select_51_i2_4_lut (.I0(\data_out_frame[6] [3]), .I1(\FRAME_MATCHER.i_31__N_2320 ), 
            .I2(encoder0_position[19]), .I3(\FRAME_MATCHER.state_31__N_2423 [3]), 
            .O(n2_adj_5161));   // verilog/coms.v(146[4] 295[11])
    defparam select_715_Select_51_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i11164_4_lut (.I0(\FRAME_MATCHER.i [0]), .I1(n133[0]), .I2(n3133), 
            .I3(\FRAME_MATCHER.i_31__N_2318 ), .O(n24764));   // verilog/coms.v(155[12:15])
    defparam i11164_4_lut.LUT_INIT = 16'hc0ca;
    SB_LUT4 i12_4_lut_adj_1475 (.I0(n7_adj_5277), .I1(n24_adj_5366), .I2(\data_in_frame[0] [7]), 
            .I3(n53201), .O(n29_adj_5386));
    defparam i12_4_lut_adj_1475.LUT_INIT = 16'h0440;
    SB_LUT4 i14_4_lut_adj_1476 (.I0(n27_adj_5384), .I1(n55426), .I2(n22_adj_5383), 
            .I3(n23221), .O(n31_adj_5387));
    defparam i14_4_lut_adj_1476.LUT_INIT = 16'h0020;
    SB_LUT4 i16_4_lut_adj_1477 (.I0(n31_adj_5387), .I1(n29_adj_5386), .I2(n56597), 
            .I3(n26_adj_5385), .O(\FRAME_MATCHER.state_31__N_2423 [3]));
    defparam i16_4_lut_adj_1477.LUT_INIT = 16'h0800;
    SB_LUT4 i11973_2_lut_2_lut (.I0(reset), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(GND_net), .I3(GND_net), .O(n25577));   // verilog/coms.v(128[12] 296[6])
    defparam i11973_2_lut_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i11972_2_lut_2_lut (.I0(reset), .I1(\FRAME_MATCHER.i_31__N_2319 ), 
            .I2(GND_net), .I3(GND_net), .O(n25576));   // verilog/coms.v(128[12] 296[6])
    defparam i11972_2_lut_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i4910_4_lut (.I0(\FRAME_MATCHER.i_31__N_2325 ), .I1(n29111), 
            .I2(n54660), .I3(n4425), .O(n18187));   // verilog/coms.v(146[4] 295[11])
    defparam i4910_4_lut.LUT_INIT = 16'ha0a2;
    SB_LUT4 i1_4_lut_adj_1478 (.I0(n18187), .I1(n29111), .I2(n52615), 
            .I3(n19648), .O(n23848));   // verilog/coms.v(146[4] 295[11])
    defparam i1_4_lut_adj_1478.LUT_INIT = 16'hbbba;
    SB_LUT4 select_715_Select_50_i2_4_lut (.I0(\data_out_frame[6] [2]), .I1(\FRAME_MATCHER.i_31__N_2320 ), 
            .I2(encoder0_position[18]), .I3(\FRAME_MATCHER.state_31__N_2423 [3]), 
            .O(n2_adj_5160));   // verilog/coms.v(146[4] 295[11])
    defparam select_715_Select_50_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i444_2_lut (.I0(n3302), .I1(\FRAME_MATCHER.i_31__N_2323 ), .I2(GND_net), 
            .I3(GND_net), .O(n1808));   // verilog/coms.v(146[4] 295[11])
    defparam i444_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_1479 (.I0(n3302), .I1(n29111), .I2(GND_net), 
            .I3(GND_net), .O(n29112));   // verilog/coms.v(226[9:54])
    defparam i1_2_lut_adj_1479.LUT_INIT = 16'h4444;
    SB_LUT4 i1_2_lut_adj_1480 (.I0(\FRAME_MATCHER.i_31__N_2323 ), .I1(n1705), 
            .I2(GND_net), .I3(GND_net), .O(n5_adj_5388));   // verilog/coms.v(140[7:80])
    defparam i1_2_lut_adj_1480.LUT_INIT = 16'h8888;
    SB_LUT4 i1_4_lut_adj_1481 (.I0(n5_adj_5388), .I1(n1702), .I2(n29112), 
            .I3(n54478), .O(n51969));   // verilog/coms.v(146[4] 295[11])
    defparam i1_4_lut_adj_1481.LUT_INIT = 16'hb380;
    SB_LUT4 i4915_4_lut (.I0(n1703), .I1(\FRAME_MATCHER.state[3] ), .I2(n1705), 
            .I3(n22342), .O(n18192));   // verilog/coms.v(146[4] 295[11])
    defparam i4915_4_lut.LUT_INIT = 16'heccc;
    SB_LUT4 i433_2_lut (.I0(\FRAME_MATCHER.state_31__N_2423 [3]), .I1(\FRAME_MATCHER.i_31__N_2320 ), 
            .I2(GND_net), .I3(GND_net), .O(n1797));   // verilog/coms.v(146[4] 295[11])
    defparam i433_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1_3_lut_adj_1482 (.I0(\FRAME_MATCHER.i_31__N_2320 ), .I1(\FRAME_MATCHER.state_31__N_2423 [3]), 
            .I2(\data_out_frame[0][2] ), .I3(GND_net), .O(n2));   // verilog/coms.v(146[4] 295[11])
    defparam i1_3_lut_adj_1482.LUT_INIT = 16'ha8a8;
    SB_LUT4 i1_2_lut_adj_1483 (.I0(\FRAME_MATCHER.i_31__N_2319 ), .I1(n771), 
            .I2(GND_net), .I3(GND_net), .O(n1796));   // verilog/coms.v(146[4] 295[11])
    defparam i1_2_lut_adj_1483.LUT_INIT = 16'h8888;
    SB_LUT4 i21942_4_lut (.I0(n8_adj_5139), .I1(\FRAME_MATCHER.i [31]), 
            .I2(n22258), .I3(\FRAME_MATCHER.i [3]), .O(n3302));   // verilog/coms.v(226[9:54])
    defparam i21942_4_lut.LUT_INIT = 16'h3230;
    SB_LUT4 i1_2_lut_adj_1484 (.I0(\FRAME_MATCHER.i [4]), .I1(n22428), .I2(GND_net), 
            .I3(GND_net), .O(n22258));   // verilog/coms.v(154[7:23])
    defparam i1_2_lut_adj_1484.LUT_INIT = 16'heeee;
    SB_LUT4 i21939_4_lut (.I0(n5_adj_5365), .I1(\FRAME_MATCHER.i [31]), 
            .I2(\FRAME_MATCHER.i [3]), .I3(\FRAME_MATCHER.i [2]), .O(n771));   // verilog/coms.v(157[9:60])
    defparam i21939_4_lut.LUT_INIT = 16'h3332;
    SB_LUT4 i1_2_lut_adj_1485 (.I0(\FRAME_MATCHER.i_31__N_2319 ), .I1(n771), 
            .I2(GND_net), .I3(GND_net), .O(n30_adj_5389));   // verilog/coms.v(146[4] 295[11])
    defparam i1_2_lut_adj_1485.LUT_INIT = 16'h2222;
    SB_LUT4 i1_2_lut_adj_1486 (.I0(\FRAME_MATCHER.i_31__N_2318 ), .I1(n22342), 
            .I2(GND_net), .I3(GND_net), .O(n52879));   // verilog/coms.v(146[4] 295[11])
    defparam i1_2_lut_adj_1486.LUT_INIT = 16'heeee;
    SB_LUT4 i2_2_lut_adj_1487 (.I0(n3302), .I1(\FRAME_MATCHER.i_31__N_2323 ), 
            .I2(GND_net), .I3(GND_net), .O(n19648));   // verilog/coms.v(146[4] 295[11])
    defparam i2_2_lut_adj_1487.LUT_INIT = 16'h4444;
    SB_LUT4 i2_4_lut_adj_1488 (.I0(n4425), .I1(n19648), .I2(\FRAME_MATCHER.i_31__N_2325 ), 
            .I3(n52879), .O(n54832));   // verilog/coms.v(146[4] 295[11])
    defparam i2_4_lut_adj_1488.LUT_INIT = 16'hffdc;
    SB_LUT4 i41906_4_lut (.I0(n1703), .I1(n30_adj_5389), .I2(n1705), .I3(n54832), 
            .O(n56605));   // verilog/coms.v(146[4] 295[11])
    defparam i41906_4_lut.LUT_INIT = 16'h8a88;
    SB_LUT4 i1_2_lut_adj_1489 (.I0(Kp_23__N_1583), .I1(\FRAME_MATCHER.i_31__N_2324 ), 
            .I2(GND_net), .I3(GND_net), .O(n29098));   // verilog/coms.v(146[4] 295[11])
    defparam i1_2_lut_adj_1489.LUT_INIT = 16'heeee;
    SB_LUT4 i2_2_lut_adj_1490 (.I0(\data_in[2] [3]), .I1(\data_in[3] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n10_adj_5390));
    defparam i2_2_lut_adj_1490.LUT_INIT = 16'heeee;
    SB_LUT4 i6_4_lut_adj_1491 (.I0(\data_in[0] [2]), .I1(\data_in[3] [3]), 
            .I2(\data_in[3] [1]), .I3(\data_in[0] [7]), .O(n14_adj_5391));
    defparam i6_4_lut_adj_1491.LUT_INIT = 16'hfeff;
    SB_LUT4 i7_4_lut_adj_1492 (.I0(\data_in[3] [6]), .I1(n14_adj_5391), 
            .I2(n10_adj_5390), .I3(\data_in[2] [1]), .O(n22352));
    defparam i7_4_lut_adj_1492.LUT_INIT = 16'hfffd;
    SB_LUT4 i8_4_lut_adj_1493 (.I0(\data_in[2] [6]), .I1(\data_in[1] [3]), 
            .I2(\data_in[1] [6]), .I3(\data_in[1] [2]), .O(n20_adj_5392));
    defparam i8_4_lut_adj_1493.LUT_INIT = 16'hfbff;
    SB_LUT4 i7_4_lut_adj_1494 (.I0(n22352), .I1(n22277), .I2(\data_in[3] [7]), 
            .I3(\data_in[0] [1]), .O(n19));
    defparam i7_4_lut_adj_1494.LUT_INIT = 16'hfeff;
    SB_LUT4 i42025_4_lut (.I0(\data_in[2] [5]), .I1(\data_in[2] [0]), .I2(\data_in[3] [2]), 
            .I3(\data_in[0] [5]), .O(n56728));
    defparam i42025_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i11_3_lut_adj_1495 (.I0(n56728), .I1(n19), .I2(n20_adj_5392), 
            .I3(GND_net), .O(n29111));
    defparam i11_3_lut_adj_1495.LUT_INIT = 16'hfdfd;
    SB_LUT4 i7_4_lut_adj_1496 (.I0(\data_in[2] [4]), .I1(n22352), .I2(\data_in[1] [5]), 
            .I3(n22425), .O(n18_adj_5393));
    defparam i7_4_lut_adj_1496.LUT_INIT = 16'hfffd;
    SB_LUT4 i9_4_lut_adj_1497 (.I0(\data_in[0] [6]), .I1(n18_adj_5393), 
            .I2(\data_in[3] [0]), .I3(n22419), .O(n20_adj_5394));
    defparam i9_4_lut_adj_1497.LUT_INIT = 16'hfffd;
    SB_LUT4 i4_2_lut_adj_1498 (.I0(\data_in[1] [0]), .I1(\data_in[0] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n15_adj_5395));
    defparam i4_2_lut_adj_1498.LUT_INIT = 16'heeee;
    SB_LUT4 i10_4_lut_adj_1499 (.I0(n15_adj_5395), .I1(n20_adj_5394), .I2(\data_in[2] [2]), 
            .I3(\data_in[1] [4]), .O(n1702));
    defparam i10_4_lut_adj_1499.LUT_INIT = 16'hfeff;
    SB_LUT4 i1_2_lut_adj_1500 (.I0(n1702), .I1(n29111), .I2(GND_net), 
            .I3(GND_net), .O(n1703));   // verilog/coms.v(146[4] 295[11])
    defparam i1_2_lut_adj_1500.LUT_INIT = 16'h8888;
    SB_LUT4 i4_4_lut_adj_1501 (.I0(\data_in[1] [7]), .I1(\data_in[0] [0]), 
            .I2(\data_in[1] [1]), .I3(\data_in[0] [4]), .O(n10_adj_5396));
    defparam i4_4_lut_adj_1501.LUT_INIT = 16'hfdff;
    SB_LUT4 i5_3_lut_adj_1502 (.I0(\data_in[3] [4]), .I1(n10_adj_5396), 
            .I2(\data_in[2] [7]), .I3(GND_net), .O(n22419));
    defparam i5_3_lut_adj_1502.LUT_INIT = 16'hdfdf;
    SB_LUT4 i42027_3_lut (.I0(\data_in[3] [0]), .I1(\data_in[2] [2]), .I2(\data_in[1] [5]), 
            .I3(GND_net), .O(n56730));
    defparam i42027_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 i6_4_lut_adj_1503 (.I0(\data_in[1] [0]), .I1(\data_in[0] [6]), 
            .I2(\data_in[2] [4]), .I3(\data_in[0] [3]), .O(n15_adj_5397));
    defparam i6_4_lut_adj_1503.LUT_INIT = 16'hfdff;
    SB_LUT4 i8_4_lut_adj_1504 (.I0(n15_adj_5397), .I1(\data_in[1] [4]), 
            .I2(n56730), .I3(n22419), .O(n22277));
    defparam i8_4_lut_adj_1504.LUT_INIT = 16'hffef;
    SB_LUT4 i6_4_lut_adj_1505 (.I0(\data_in[0] [1]), .I1(\data_in[1] [2]), 
            .I2(\data_in[3] [2]), .I3(\data_in[0] [5]), .O(n16_adj_5398));
    defparam i6_4_lut_adj_1505.LUT_INIT = 16'hfffe;
    SB_LUT4 i7_4_lut_adj_1506 (.I0(\data_in[1] [6]), .I1(\data_in[2] [5]), 
            .I2(\data_in[2] [0]), .I3(\data_in[1] [3]), .O(n17_adj_5399));
    defparam i7_4_lut_adj_1506.LUT_INIT = 16'hfffd;
    SB_LUT4 i9_4_lut_adj_1507 (.I0(n17_adj_5399), .I1(\data_in[3] [7]), 
            .I2(n16_adj_5398), .I3(\data_in[2] [6]), .O(n22425));
    defparam i9_4_lut_adj_1507.LUT_INIT = 16'hfbff;
    SB_LUT4 i6_4_lut_adj_1508 (.I0(\data_in[3] [6]), .I1(\data_in[0] [7]), 
            .I2(\data_in[2] [1]), .I3(n22277), .O(n16_adj_5400));
    defparam i6_4_lut_adj_1508.LUT_INIT = 16'hffef;
    SB_LUT4 i7_4_lut_adj_1509 (.I0(n22425), .I1(\data_in[2] [3]), .I2(\data_in[0] [2]), 
            .I3(\data_in[3] [5]), .O(n17_adj_5401));
    defparam i7_4_lut_adj_1509.LUT_INIT = 16'hbfff;
    SB_LUT4 i9_4_lut_adj_1510 (.I0(n17_adj_5401), .I1(\data_in[3] [3]), 
            .I2(n16_adj_5400), .I3(\data_in[3] [1]), .O(n1705));
    defparam i9_4_lut_adj_1510.LUT_INIT = 16'hfbff;
    SB_LUT4 i1_2_lut_adj_1511 (.I0(n1705), .I1(\FRAME_MATCHER.i_31__N_2318 ), 
            .I2(GND_net), .I3(GND_net), .O(n4_adj_5402));   // verilog/coms.v(146[4] 295[11])
    defparam i1_2_lut_adj_1511.LUT_INIT = 16'h8888;
    SB_LUT4 i2_4_lut_adj_1512 (.I0(\FRAME_MATCHER.state_31__N_2423 [3]), .I1(n1703), 
            .I2(\FRAME_MATCHER.i_31__N_2320 ), .I3(n4_adj_5402), .O(n6_adj_5403));   // verilog/coms.v(146[4] 295[11])
    defparam i2_4_lut_adj_1512.LUT_INIT = 16'hdc50;
    SB_LUT4 i3_4_lut_adj_1513 (.I0(n29098), .I1(n6_adj_5403), .I2(\FRAME_MATCHER.i_31__N_2322 ), 
            .I3(n36757), .O(n63712));   // verilog/coms.v(146[4] 295[11])
    defparam i3_4_lut_adj_1513.LUT_INIT = 16'heefe;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1514 (.I0(\data_out_frame[5] [3]), .I1(\data_out_frame[8] [1]), 
            .I2(\data_out_frame[5] [4]), .I3(\data_out_frame[8] [2]), .O(n6_adj_5066));   // verilog/coms.v(76[16:27])
    defparam i1_2_lut_3_lut_4_lut_adj_1514.LUT_INIT = 16'h6996;
    SB_LUT4 select_715_Select_99_i2_4_lut (.I0(\data_out_frame[12] [3]), .I1(\FRAME_MATCHER.i_31__N_2320 ), 
            .I2(setpoint[19]), .I3(\FRAME_MATCHER.state_31__N_2423 [3]), 
            .O(n2_adj_5159));   // verilog/coms.v(146[4] 295[11])
    defparam select_715_Select_99_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_715_Select_98_i2_4_lut (.I0(\data_out_frame[12] [2]), .I1(\FRAME_MATCHER.i_31__N_2320 ), 
            .I2(setpoint[18]), .I3(\FRAME_MATCHER.state_31__N_2423 [3]), 
            .O(n2_adj_5158));   // verilog/coms.v(146[4] 295[11])
    defparam select_715_Select_98_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_4_lut_4_lut (.I0(reset), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(\FRAME_MATCHER.i_31__N_2320 ), .I3(\data_out_frame[26] [0]), 
            .O(n52841));   // verilog/coms.v(128[12] 296[6])
    defparam i1_2_lut_4_lut_4_lut.LUT_INIT = 16'h5100;
    SB_LUT4 i45501_2_lut (.I0(\FRAME_MATCHER.i [24]), .I1(\FRAME_MATCHER.i_31__N_2318 ), 
            .I2(GND_net), .I3(GND_net), .O(n59812));   // verilog/coms.v(155[12:15])
    defparam i45501_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1515 (.I0(reset), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(\FRAME_MATCHER.i_31__N_2320 ), .I3(\data_out_frame[26] [1]), 
            .O(n52840));   // verilog/coms.v(128[12] 296[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1515.LUT_INIT = 16'h5100;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1516 (.I0(reset), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(\FRAME_MATCHER.i_31__N_2320 ), .I3(\data_out_frame[26] [2]), 
            .O(n52839));   // verilog/coms.v(128[12] 296[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1516.LUT_INIT = 16'h5100;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1517 (.I0(reset), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(\FRAME_MATCHER.i_31__N_2320 ), .I3(\data_out_frame[26] [3]), 
            .O(n52838));   // verilog/coms.v(128[12] 296[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1517.LUT_INIT = 16'h5100;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1518 (.I0(reset), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(\FRAME_MATCHER.i_31__N_2320 ), .I3(\data_out_frame[26] [4]), 
            .O(n52837));   // verilog/coms.v(128[12] 296[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1518.LUT_INIT = 16'h5100;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1519 (.I0(reset), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(\FRAME_MATCHER.i_31__N_2320 ), .I3(\data_out_frame[26] [5]), 
            .O(n52836));   // verilog/coms.v(128[12] 296[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1519.LUT_INIT = 16'h5100;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1520 (.I0(reset), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(\FRAME_MATCHER.i_31__N_2320 ), .I3(\data_out_frame[26][6] ), 
            .O(n52835));   // verilog/coms.v(128[12] 296[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1520.LUT_INIT = 16'h5100;
    SB_LUT4 select_715_Select_222_i3_4_lut (.I0(n48259), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(n48764), .I3(n48824), .O(n3_adj_5150));   // verilog/coms.v(146[4] 295[11])
    defparam select_715_Select_222_i3_4_lut.LUT_INIT = 16'h4884;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1521 (.I0(reset), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(\FRAME_MATCHER.i_31__N_2320 ), .I3(\data_out_frame[26] [7]), 
            .O(n52834));   // verilog/coms.v(128[12] 296[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1521.LUT_INIT = 16'h5100;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1522 (.I0(reset), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(\FRAME_MATCHER.i_31__N_2320 ), .I3(\data_out_frame[27] [0]), 
            .O(n52833));   // verilog/coms.v(128[12] 296[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1522.LUT_INIT = 16'h5100;
    SB_LUT4 select_715_Select_220_i3_4_lut (.I0(n48239), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(n53474), .I3(n48758), .O(n3_adj_5148));   // verilog/coms.v(146[4] 295[11])
    defparam select_715_Select_220_i3_4_lut.LUT_INIT = 16'h8448;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1523 (.I0(reset), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(\FRAME_MATCHER.i_31__N_2320 ), .I3(\data_out_frame[27] [1]), 
            .O(n52832));   // verilog/coms.v(128[12] 296[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1523.LUT_INIT = 16'h5100;
    SB_LUT4 select_715_Select_219_i3_3_lut (.I0(n53097), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(n53335), .I3(GND_net), .O(n3_adj_5147));   // verilog/coms.v(146[4] 295[11])
    defparam select_715_Select_219_i3_3_lut.LUT_INIT = 16'h8484;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1524 (.I0(reset), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(\FRAME_MATCHER.i_31__N_2320 ), .I3(\data_out_frame[27] [2]), 
            .O(n52831));   // verilog/coms.v(128[12] 296[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1524.LUT_INIT = 16'h5100;
    SB_LUT4 i9_4_lut_adj_1525 (.I0(n53477), .I1(\data_out_frame[17] [6]), 
            .I2(\data_out_frame[22] [7]), .I3(\data_out_frame[17] [2]), 
            .O(n22_adj_5404));
    defparam i9_4_lut_adj_1525.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1526 (.I0(reset), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(\FRAME_MATCHER.i_31__N_2320 ), .I3(\data_out_frame[27] [3]), 
            .O(n52830));   // verilog/coms.v(128[12] 296[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1526.LUT_INIT = 16'h5100;
    SB_LUT4 i11_4_lut_adj_1527 (.I0(n15_adj_5362), .I1(n22_adj_5404), .I2(n48497), 
            .I3(n55349), .O(n24_adj_5405));
    defparam i11_4_lut_adj_1527.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1528 (.I0(reset), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(\FRAME_MATCHER.i_31__N_2320 ), .I3(\data_out_frame[27] [4]), 
            .O(n52829));   // verilog/coms.v(128[12] 296[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1528.LUT_INIT = 16'h5100;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1529 (.I0(reset), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(\FRAME_MATCHER.i_31__N_2320 ), .I3(\data_out_frame[27] [5]), 
            .O(n52828));   // verilog/coms.v(128[12] 296[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1529.LUT_INIT = 16'h5100;
    SB_LUT4 i12_4_lut_adj_1530 (.I0(\data_out_frame[22] [6]), .I1(n24_adj_5405), 
            .I2(n20_adj_5406), .I3(n47634), .O(n48758));
    defparam i12_4_lut_adj_1530.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1531 (.I0(reset), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(\FRAME_MATCHER.i_31__N_2320 ), .I3(\data_out_frame[27][6] ), 
            .O(n52827));   // verilog/coms.v(128[12] 296[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1531.LUT_INIT = 16'h5100;
    SB_LUT4 select_715_Select_218_i3_4_lut (.I0(n53335), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(n48758), .I3(n52908), .O(n3_adj_5146));   // verilog/coms.v(146[4] 295[11])
    defparam select_715_Select_218_i3_4_lut.LUT_INIT = 16'h8448;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1532 (.I0(reset), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(\FRAME_MATCHER.i_31__N_2320 ), .I3(\data_out_frame[27] [7]), 
            .O(n52826));   // verilog/coms.v(128[12] 296[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1532.LUT_INIT = 16'h5100;
    SB_LUT4 i12497_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(\data_in[1] [0]), 
            .I3(\data_in[0] [0]), .O(n26101));   // verilog/coms.v(128[12] 296[6])
    defparam i12497_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i2_3_lut_adj_1533 (.I0(n55349), .I1(n55268), .I2(\data_out_frame[21] [0]), 
            .I3(GND_net), .O(n48259));
    defparam i2_3_lut_adj_1533.LUT_INIT = 16'h9696;
    SB_LUT4 i12787_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(\data_in[1] [2]), 
            .I3(\data_in[0] [2]), .O(n26391));   // verilog/coms.v(128[12] 296[6])
    defparam i12787_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1_2_lut_adj_1534 (.I0(n48239), .I1(n48259), .I2(GND_net), 
            .I3(GND_net), .O(n23272));
    defparam i1_2_lut_adj_1534.LUT_INIT = 16'h6666;
    SB_LUT4 i12786_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(\data_in[1] [3]), 
            .I3(\data_in[0] [3]), .O(n26390));   // verilog/coms.v(128[12] 296[6])
    defparam i12786_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i12785_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(\data_in[1] [4]), 
            .I3(\data_in[0] [4]), .O(n26389));   // verilog/coms.v(128[12] 296[6])
    defparam i12785_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i12784_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(\data_in[1] [5]), 
            .I3(\data_in[0] [5]), .O(n26388));   // verilog/coms.v(128[12] 296[6])
    defparam i12784_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 select_715_Select_217_i3_4_lut (.I0(n23272), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(n6_adj_5311), .I3(n48935), .O(n3_adj_5145));   // verilog/coms.v(146[4] 295[11])
    defparam select_715_Select_217_i3_4_lut.LUT_INIT = 16'h8448;
    SB_LUT4 select_715_Select_216_i3_3_lut (.I0(n48935), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(n52908), .I3(GND_net), .O(n3_adj_5144));   // verilog/coms.v(146[4] 295[11])
    defparam select_715_Select_216_i3_3_lut.LUT_INIT = 16'h4848;
    SB_LUT4 i12783_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(\data_in[1] [6]), 
            .I3(\data_in[0] [6]), .O(n26387));   // verilog/coms.v(128[12] 296[6])
    defparam i12783_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1_2_lut_adj_1535 (.I0(n47766), .I1(n53574), .I2(GND_net), 
            .I3(GND_net), .O(n53282));
    defparam i1_2_lut_adj_1535.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_1536 (.I0(\data_out_frame[21] [1]), .I1(n53291), 
            .I2(n53282), .I3(n33_c), .O(n48824));
    defparam i3_4_lut_adj_1536.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1537 (.I0(n55349), .I1(\data_out_frame[21] [0]), 
            .I2(n47851), .I3(GND_net), .O(n53207));
    defparam i2_3_lut_adj_1537.LUT_INIT = 16'h6969;
    SB_LUT4 i2_3_lut_adj_1538 (.I0(n54590), .I1(\data_out_frame[22] [5]), 
            .I2(n54765), .I3(GND_net), .O(n53335));
    defparam i2_3_lut_adj_1538.LUT_INIT = 16'h9696;
    SB_LUT4 i11_4_lut_adj_1539 (.I0(n55477), .I1(n53207), .I2(n53506), 
            .I3(n55268), .O(n26_adj_5407));
    defparam i11_4_lut_adj_1539.LUT_INIT = 16'h6996;
    SB_LUT4 i9_4_lut_adj_1540 (.I0(n53302), .I1(n53498), .I2(n48764), 
            .I3(n52931), .O(n24_adj_5408));
    defparam i9_4_lut_adj_1540.LUT_INIT = 16'h6996;
    SB_LUT4 i10_4_lut_adj_1541 (.I0(\data_out_frame[22] [6]), .I1(n48777), 
            .I2(n48858), .I3(n53219), .O(n25_adj_5409));
    defparam i10_4_lut_adj_1541.LUT_INIT = 16'h9669;
    SB_LUT4 i8_3_lut (.I0(n48824), .I1(n48885), .I2(n23712), .I3(GND_net), 
            .O(n23_adj_5410));
    defparam i8_3_lut.LUT_INIT = 16'h6969;
    SB_LUT4 i14_4_lut_adj_1542 (.I0(n23_adj_5410), .I1(n25_adj_5409), .I2(n24_adj_5408), 
            .I3(n26_adj_5407), .O(n48935));
    defparam i14_4_lut_adj_1542.LUT_INIT = 16'h6996;
    SB_LUT4 select_715_Select_215_i3_4_lut (.I0(n48935), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(n53335), .I3(n52932), .O(n3_adj_5143));   // verilog/coms.v(146[4] 295[11])
    defparam select_715_Select_215_i3_4_lut.LUT_INIT = 16'h4884;
    SB_LUT4 i12782_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(\data_in[1] [7]), 
            .I3(\data_in[0] [7]), .O(n26386));   // verilog/coms.v(128[12] 296[6])
    defparam i12782_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 select_715_Select_214_i3_3_lut (.I0(n52932), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(n47815), .I3(GND_net), .O(n3_adj_5142));   // verilog/coms.v(146[4] 295[11])
    defparam select_715_Select_214_i3_3_lut.LUT_INIT = 16'h4848;
    SB_LUT4 select_715_Select_213_i3_2_lut_3_lut (.I0(n47815), .I1(n55276), 
            .I2(\FRAME_MATCHER.state[3] ), .I3(GND_net), .O(n3_adj_5141));
    defparam select_715_Select_213_i3_2_lut_3_lut.LUT_INIT = 16'h9090;
    SB_LUT4 i3_3_lut_4_lut (.I0(n47815), .I1(n55276), .I2(n52908), .I3(n54489), 
            .O(n8_adj_5102));
    defparam i3_3_lut_4_lut.LUT_INIT = 16'h9669;
    SB_LUT4 i12781_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(\data_in[2] [0]), 
            .I3(\data_in[1] [0]), .O(n26385));   // verilog/coms.v(128[12] 296[6])
    defparam i12781_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i12780_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(\data_in[2] [1]), 
            .I3(\data_in[1] [1]), .O(n26384));   // verilog/coms.v(128[12] 296[6])
    defparam i12780_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i12779_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(\data_in[2] [2]), 
            .I3(\data_in[1] [2]), .O(n26383));   // verilog/coms.v(128[12] 296[6])
    defparam i12779_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i12778_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(\data_in[2] [3]), 
            .I3(\data_in[1] [3]), .O(n26382));   // verilog/coms.v(128[12] 296[6])
    defparam i12778_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1_2_lut_3_lut_adj_1543 (.I0(n10_adj_5280), .I1(n53712), .I2(n8_adj_5074), 
            .I3(GND_net), .O(n25077));
    defparam i1_2_lut_3_lut_adj_1543.LUT_INIT = 16'hfbfb;
    SB_LUT4 i12777_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(\data_in[2] [4]), 
            .I3(\data_in[1] [4]), .O(n26381));   // verilog/coms.v(128[12] 296[6])
    defparam i12777_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i12776_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(\data_in[2] [5]), 
            .I3(\data_in[1] [5]), .O(n26380));   // verilog/coms.v(128[12] 296[6])
    defparam i12776_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i7_4_lut_adj_1544 (.I0(\data_out_frame[14] [4]), .I1(\data_out_frame[13] [0]), 
            .I2(n53342), .I3(n53501), .O(n18_adj_5411));
    defparam i7_4_lut_adj_1544.LUT_INIT = 16'h6996;
    SB_LUT4 i12775_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(\data_in[2] [6]), 
            .I3(\data_in[1] [6]), .O(n26379));   // verilog/coms.v(128[12] 296[6])
    defparam i12775_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i8_4_lut_adj_1545 (.I0(n53360), .I1(n21993), .I2(n53273), 
            .I3(\data_out_frame[14] [1]), .O(n19_adj_5412));
    defparam i8_4_lut_adj_1545.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_1546 (.I0(n19_adj_5412), .I1(\data_out_frame[15] [7]), 
            .I2(n17_adj_5360), .I3(n18_adj_5411), .O(n12_adj_5413));
    defparam i4_4_lut_adj_1546.LUT_INIT = 16'h9669;
    SB_LUT4 i5_4_lut_adj_1547 (.I0(\data_out_frame[15] [0]), .I1(n53305), 
            .I2(n23432), .I3(n23361), .O(n13_adj_5414));
    defparam i5_4_lut_adj_1547.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut_adj_1548 (.I0(n13_adj_5414), .I1(n53391), .I2(n12_adj_5413), 
            .I3(n22958), .O(n54606));
    defparam i7_4_lut_adj_1548.LUT_INIT = 16'h6996;
    SB_LUT4 i5_4_lut_adj_1549 (.I0(\data_out_frame[16] [0]), .I1(n54606), 
            .I2(\data_out_frame[17] [1]), .I3(\data_out_frame[16] [7]), 
            .O(n12_adj_5415));
    defparam i5_4_lut_adj_1549.LUT_INIT = 16'h9669;
    SB_LUT4 i6_4_lut_adj_1550 (.I0(\data_out_frame[17] [7]), .I1(n12_adj_5415), 
            .I2(n53524), .I3(n54719), .O(n53477));
    defparam i6_4_lut_adj_1550.LUT_INIT = 16'h9669;
    SB_LUT4 i6_4_lut_adj_1551 (.I0(n53477), .I1(n53574), .I2(\data_out_frame[17] [5]), 
            .I3(n53237), .O(n15_adj_5416));   // verilog/coms.v(98[12:26])
    defparam i6_4_lut_adj_1551.LUT_INIT = 16'h6996;
    SB_LUT4 i8_4_lut_adj_1552 (.I0(n15_adj_5416), .I1(\data_out_frame[17] [0]), 
            .I2(n14_adj_5361), .I3(\data_out_frame[16] [4]), .O(n21971));   // verilog/coms.v(98[12:26])
    defparam i8_4_lut_adj_1552.LUT_INIT = 16'h6996;
    SB_LUT4 i12774_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(\data_in[2] [7]), 
            .I3(\data_in[1] [7]), .O(n26378));   // verilog/coms.v(128[12] 296[6])
    defparam i12774_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i12773_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(\data_in[3] [0]), 
            .I3(\data_in[2] [0]), .O(n26377));   // verilog/coms.v(128[12] 296[6])
    defparam i12773_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i12772_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(\data_in[3] [1]), 
            .I3(\data_in[2] [1]), .O(n26376));   // verilog/coms.v(128[12] 296[6])
    defparam i12772_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i12771_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(\data_in[3] [2]), 
            .I3(\data_in[2] [2]), .O(n26375));   // verilog/coms.v(128[12] 296[6])
    defparam i12771_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i2_3_lut_adj_1553 (.I0(\FRAME_MATCHER.i [3]), .I1(\FRAME_MATCHER.i [4]), 
            .I2(\FRAME_MATCHER.i [5]), .I3(GND_net), .O(n10_adj_5280));   // verilog/coms.v(154[7:23])
    defparam i2_3_lut_adj_1553.LUT_INIT = 16'hfbfb;
    SB_LUT4 i12770_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(\data_in[3] [3]), 
            .I3(\data_in[2] [3]), .O(n26374));   // verilog/coms.v(128[12] 296[6])
    defparam i12770_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1_2_lut_adj_1554 (.I0(n53339), .I1(n48790), .I2(GND_net), 
            .I3(GND_net), .O(n8_adj_5417));
    defparam i1_2_lut_adj_1554.LUT_INIT = 16'h6666;
    SB_LUT4 i5_4_lut_adj_1555 (.I0(n21971), .I1(\data_out_frame[21] [6]), 
            .I2(n55276), .I3(n48833), .O(n12_adj_5418));
    defparam i5_4_lut_adj_1555.LUT_INIT = 16'h9669;
    SB_LUT4 select_715_Select_212_i3_4_lut (.I0(n23712), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(n12_adj_5418), .I3(n8_adj_5417), .O(n3_adj_5140));   // verilog/coms.v(146[4] 295[11])
    defparam select_715_Select_212_i3_4_lut.LUT_INIT = 16'h4884;
    SB_LUT4 i45500_2_lut (.I0(\FRAME_MATCHER.i [25]), .I1(\FRAME_MATCHER.i_31__N_2318 ), 
            .I2(GND_net), .I3(GND_net), .O(n59811));   // verilog/coms.v(155[12:15])
    defparam i45500_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i45499_2_lut (.I0(\FRAME_MATCHER.i [26]), .I1(\FRAME_MATCHER.i_31__N_2318 ), 
            .I2(GND_net), .I3(GND_net), .O(n59810));   // verilog/coms.v(155[12:15])
    defparam i45499_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i12769_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(\data_in[3] [4]), 
            .I3(\data_in[2] [4]), .O(n26373));   // verilog/coms.v(128[12] 296[6])
    defparam i12769_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i12768_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(\data_in[3] [5]), 
            .I3(\data_in[2] [5]), .O(n26372));   // verilog/coms.v(128[12] 296[6])
    defparam i12768_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i12767_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(\data_in[3] [6]), 
            .I3(\data_in[2] [6]), .O(n26371));   // verilog/coms.v(128[12] 296[6])
    defparam i12767_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i12766_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(\data_in[3] [7]), 
            .I3(\data_in[2] [7]), .O(n26370));   // verilog/coms.v(128[12] 296[6])
    defparam i12766_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i12765_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(rx_data[0]), 
            .I3(\data_in[3] [0]), .O(n26369));   // verilog/coms.v(128[12] 296[6])
    defparam i12765_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i12764_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(rx_data[1]), 
            .I3(\data_in[3] [1]), .O(n26368));   // verilog/coms.v(128[12] 296[6])
    defparam i12764_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i12763_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(rx_data[2]), 
            .I3(\data_in[3] [2]), .O(n26367));   // verilog/coms.v(128[12] 296[6])
    defparam i12763_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i7_3_lut_4_lut_adj_1556 (.I0(n22564), .I1(n53068), .I2(n48790), 
            .I3(\data_out_frame[17] [0]), .O(n20_adj_5406));
    defparam i7_3_lut_4_lut_adj_1556.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_3_lut_adj_1557 (.I0(n22564), .I1(n53068), .I2(\data_out_frame[17] [4]), 
            .I3(GND_net), .O(n53088));
    defparam i1_2_lut_3_lut_adj_1557.LUT_INIT = 16'h9696;
    SB_LUT4 i12762_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(rx_data[3]), 
            .I3(\data_in[3] [3]), .O(n26366));   // verilog/coms.v(128[12] 296[6])
    defparam i12762_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i12761_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(rx_data[4]), 
            .I3(\data_in[3] [4]), .O(n26365));   // verilog/coms.v(128[12] 296[6])
    defparam i12761_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i12760_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(rx_data[5]), 
            .I3(\data_in[3] [5]), .O(n26364));   // verilog/coms.v(128[12] 296[6])
    defparam i12760_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i12759_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(rx_data[6]), 
            .I3(\data_in[3] [6]), .O(n26363));   // verilog/coms.v(128[12] 296[6])
    defparam i12759_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i12758_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(rx_data[7]), 
            .I3(\data_in[3] [7]), .O(n26362));   // verilog/coms.v(128[12] 296[6])
    defparam i12758_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 select_715_Select_211_i3_2_lut (.I0(n54489), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_5138));   // verilog/coms.v(146[4] 295[11])
    defparam select_715_Select_211_i3_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i12788_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(\data_in[1] [1]), 
            .I3(\data_in[0] [1]), .O(n26392));   // verilog/coms.v(128[12] 296[6])
    defparam i12788_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i2_3_lut_4_lut_adj_1558 (.I0(\data_in_frame[21] [1]), .I1(n53521), 
            .I2(n53495), .I3(\data_in_frame[23] [2]), .O(n54880));
    defparam i2_3_lut_4_lut_adj_1558.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_adj_1559 (.I0(\data_in_frame[20] [4]), .I1(\data_in_frame[20] [5]), 
            .I2(\data_in_frame[16] [3]), .I3(n53252), .O(n6_adj_5324));
    defparam i1_2_lut_4_lut_adj_1559.LUT_INIT = 16'h9669;
    SB_LUT4 i3_2_lut_4_lut (.I0(\data_in_frame[19] [7]), .I1(n22021), .I2(n10_adj_5318), 
            .I3(n20730), .O(n9));
    defparam i3_2_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_adj_1560 (.I0(n48392), .I1(n23039), .I2(\data_in_frame[16] [4]), 
            .I3(\data_in_frame[16] [3]), .O(n48794));
    defparam i1_2_lut_4_lut_adj_1560.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1561 (.I0(\data_in_frame[9] [1]), .I1(\data_in_frame[9] [2]), 
            .I2(\data_in_frame[11] [7]), .I3(GND_net), .O(n23741));
    defparam i1_2_lut_3_lut_adj_1561.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_4_lut_adj_1562 (.I0(\data_in_frame[2] [6]), .I1(\data_in_frame[0] [5]), 
            .I2(\data_in_frame[0] [4]), .I3(n23201), .O(n53456));
    defparam i1_2_lut_4_lut_adj_1562.LUT_INIT = 16'h6996;
    SB_LUT4 i1_3_lut_4_lut_adj_1563 (.I0(\data_in_frame[2] [7]), .I1(\data_in_frame[0] [5]), 
            .I2(\data_in_frame[1] [0]), .I3(Kp_23__N_602), .O(n23046));
    defparam i1_3_lut_4_lut_adj_1563.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_adj_1564 (.I0(\data_in_frame[5] [0]), .I1(n53471), 
            .I2(\data_in_frame[5] [1]), .I3(n23046), .O(n6_adj_5310));
    defparam i1_2_lut_4_lut_adj_1564.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1565 (.I0(\data_in_frame[3][3] ), .I1(\data_in_frame[0] [7]), 
            .I2(\data_in_frame[1] [1]), .I3(GND_net), .O(n53058));   // verilog/coms.v(75[16:43])
    defparam i1_2_lut_3_lut_adj_1565.LUT_INIT = 16'h9696;
    SB_LUT4 i45494_2_lut (.I0(\FRAME_MATCHER.i [27]), .I1(\FRAME_MATCHER.i_31__N_2318 ), 
            .I2(GND_net), .I3(GND_net), .O(n59809));   // verilog/coms.v(155[12:15])
    defparam i45494_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i1_2_lut_3_lut_adj_1566 (.I0(\data_in_frame[3][7] ), .I1(\data_in_frame[1][4] ), 
            .I2(\data_in_frame[1][3] ), .I3(GND_net), .O(n53445));   // verilog/coms.v(76[16:27])
    defparam i1_2_lut_3_lut_adj_1566.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1567 (.I0(\data_in_frame[6] [0]), .I1(\data_in_frame[1][5] ), 
            .I2(\data_in_frame[1][4] ), .I3(GND_net), .O(n53183));   // verilog/coms.v(77[16:43])
    defparam i1_2_lut_3_lut_adj_1567.LUT_INIT = 16'h9696;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_48648 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[10] [7]), .I2(\data_out_frame[11] [7]), 
            .I3(byte_transmit_counter_c[1]), .O(n63335));
    defparam byte_transmit_counter_0__bdd_4_lut_48648.LUT_INIT = 16'he4aa;
    SB_LUT4 i2_3_lut_4_lut_adj_1568 (.I0(\data_in_frame[3][6] ), .I1(\data_in_frame[3] [5]), 
            .I2(\data_in_frame[5] [7]), .I3(n23252), .O(n52989));   // verilog/coms.v(79[16:27])
    defparam i2_3_lut_4_lut_adj_1568.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1569 (.I0(n47634), .I1(\data_out_frame[17] [5]), 
            .I2(n47851), .I3(GND_net), .O(n53302));
    defparam i1_2_lut_3_lut_adj_1569.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1570 (.I0(n47634), .I1(\data_out_frame[17] [5]), 
            .I2(n23712), .I3(GND_net), .O(n5));
    defparam i1_2_lut_3_lut_adj_1570.LUT_INIT = 16'h9696;
    SB_LUT4 i13178_3_lut_4_lut (.I0(n8_adj_5286), .I1(n52895), .I2(rx_data[2]), 
            .I3(\data_in_frame[6] [2]), .O(n26782));
    defparam i13178_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13388_3_lut_4_lut (.I0(n8_adj_5074), .I1(n52882), .I2(rx_data[0]), 
            .I3(\data_in_frame[9] [0]), .O(n26992));
    defparam i13388_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13313_3_lut_4_lut (.I0(n8_adj_5286), .I1(n52895), .I2(rx_data[3]), 
            .I3(\data_in_frame[6] [3]), .O(n26917));
    defparam i13313_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_3_lut_4_lut_adj_1571 (.I0(\data_in_frame[8] [0]), .I1(n48415), 
            .I2(n53550), .I3(n53050), .O(n53541));
    defparam i2_3_lut_4_lut_adj_1571.LUT_INIT = 16'h6996;
    SB_LUT4 i13327_3_lut_4_lut (.I0(n8_adj_5286), .I1(n52895), .I2(rx_data[4]), 
            .I3(\data_in_frame[6] [4]), .O(n26931));
    defparam i13327_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_3_lut_adj_1572 (.I0(\data_in_frame[4] [2]), .I1(\data_in_frame[1][7] ), 
            .I2(\data_in_frame[1][6] ), .I3(GND_net), .O(n53418));   // verilog/coms.v(74[16:42])
    defparam i1_2_lut_3_lut_adj_1572.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1573 (.I0(\data_in_frame[3] [4]), .I1(\data_in_frame[1][3] ), 
            .I2(\data_in_frame[1][2] ), .I3(GND_net), .O(n22652));
    defparam i1_2_lut_3_lut_adj_1573.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_4_lut_adj_1574 (.I0(\data_in_frame[9] [7]), .I1(\data_in_frame[9] [6]), 
            .I2(n20816), .I3(n20820), .O(n47554));
    defparam i2_3_lut_4_lut_adj_1574.LUT_INIT = 16'h6996;
    SB_LUT4 i45493_2_lut (.I0(\FRAME_MATCHER.i [28]), .I1(\FRAME_MATCHER.i_31__N_2318 ), 
            .I2(GND_net), .I3(GND_net), .O(n59808));   // verilog/coms.v(155[12:15])
    defparam i45493_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i45285_2_lut (.I0(\FRAME_MATCHER.i [29]), .I1(\FRAME_MATCHER.i_31__N_2318 ), 
            .I2(GND_net), .I3(GND_net), .O(n59807));   // verilog/coms.v(155[12:15])
    defparam i45285_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i1_2_lut_4_lut_adj_1575 (.I0(\data_in_frame[1] [1]), .I1(\data_in_frame[3][2] ), 
            .I2(\data_in_frame[0] [6]), .I3(\data_in_frame[1] [0]), .O(n23666));   // verilog/coms.v(71[16:27])
    defparam i1_2_lut_4_lut_adj_1575.LUT_INIT = 16'h6996;
    SB_LUT4 i13330_3_lut_4_lut (.I0(n8_adj_5286), .I1(n52895), .I2(rx_data[5]), 
            .I3(\data_in_frame[6] [5]), .O(n26934));
    defparam i13330_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i46079_2_lut (.I0(\FRAME_MATCHER.i [30]), .I1(\FRAME_MATCHER.i_31__N_2318 ), 
            .I2(GND_net), .I3(GND_net), .O(n59793));   // verilog/coms.v(155[12:15])
    defparam i46079_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i1_2_lut_3_lut_adj_1576 (.I0(\data_in_frame[4]_c [4]), .I1(n23536), 
            .I2(\data_in_frame[4]_c [5]), .I3(GND_net), .O(n22688));   // verilog/coms.v(97[12:25])
    defparam i1_2_lut_3_lut_adj_1576.LUT_INIT = 16'h9696;
    SB_LUT4 i5_3_lut_4_lut_adj_1577 (.I0(\data_in_frame[6] [6]), .I1(n10_adj_5287), 
            .I2(\data_in_frame[2] [5]), .I3(n52956), .O(n23753));   // verilog/coms.v(75[16:43])
    defparam i5_3_lut_4_lut_adj_1577.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_1578 (.I0(\data_in_frame[4]_c [4]), .I1(\data_in_frame[6] [7]), 
            .I2(\data_in_frame[2] [3]), .I3(n53122), .O(n53168));   // verilog/coms.v(75[16:43])
    defparam i2_3_lut_4_lut_adj_1578.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1579 (.I0(\data_in_frame[12] [2]), .I1(n47554), 
            .I2(\data_in_frame[10] [0]), .I3(GND_net), .O(n53288));
    defparam i1_2_lut_3_lut_adj_1579.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_4_lut_adj_1580 (.I0(\data_in_frame[1][3] ), .I1(n53424), 
            .I2(n53073), .I3(\data_in_frame[5] [5]), .O(n48354));   // verilog/coms.v(86[17:70])
    defparam i2_3_lut_4_lut_adj_1580.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_1581 (.I0(\data_in_frame[6] [4]), .I1(\data_in_frame[8] [6]), 
            .I2(n53345), .I3(Kp_23__N_710), .O(n23193));   // verilog/coms.v(77[16:43])
    defparam i2_3_lut_4_lut_adj_1581.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_1582 (.I0(\data_in_frame[13] [0]), .I1(n52940), 
            .I2(n48942), .I3(n22898), .O(n53580));
    defparam i2_3_lut_4_lut_adj_1582.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_3_lut_adj_1583 (.I0(\data_in_frame[9] [1]), .I1(\data_in_frame[9] [2]), 
            .I2(\data_in_frame[11] [3]), .I3(GND_net), .O(n53430));   // verilog/coms.v(73[16:41])
    defparam i1_2_lut_3_lut_adj_1583.LUT_INIT = 16'h9696;
    SB_LUT4 i5_3_lut_4_lut_adj_1584 (.I0(\data_in_frame[15] [7]), .I1(\data_in_frame[16] [0]), 
            .I2(n10_adj_5247), .I3(\data_in_frame[17] [7]), .O(n22021));   // verilog/coms.v(86[17:28])
    defparam i5_3_lut_4_lut_adj_1584.LUT_INIT = 16'h6996;
    SB_LUT4 i13333_3_lut_4_lut (.I0(n8_adj_5286), .I1(n52895), .I2(rx_data[6]), 
            .I3(\data_in_frame[6] [6]), .O(n26937));
    defparam i13333_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_4_lut_adj_1585 (.I0(n22610), .I1(n23152), .I2(\data_in_frame[11] [5]), 
            .I3(n23002), .O(n53509));   // verilog/coms.v(86[17:28])
    defparam i1_2_lut_4_lut_adj_1585.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_1586 (.I0(n23152), .I1(n22594), .I2(\data_in_frame[11] [3]), 
            .I3(n23479), .O(n22822));   // verilog/coms.v(73[16:41])
    defparam i2_3_lut_4_lut_adj_1586.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_4_lut (.I0(n22843), .I1(\data_in_frame[13] [5]), .I2(n23402), 
            .I3(GND_net), .O(n53079));   // verilog/coms.v(77[16:43])
    defparam i3_4_lut_4_lut.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_4_lut_adj_1587 (.I0(\data_in_frame[18] [1]), .I1(n53321), 
            .I2(n10_adj_5247), .I3(\data_in_frame[17] [7]), .O(n53400));
    defparam i1_2_lut_4_lut_adj_1587.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1588 (.I0(n55031), .I1(n53085), .I2(\data_in_frame[18]_c [6]), 
            .I3(GND_net), .O(n53348));
    defparam i1_2_lut_3_lut_adj_1588.LUT_INIT = 16'h6969;
    SB_LUT4 select_715_Select_49_i2_4_lut (.I0(\data_out_frame[6] [1]), .I1(\FRAME_MATCHER.i_31__N_2320 ), 
            .I2(encoder0_position[17]), .I3(\FRAME_MATCHER.state_31__N_2423 [3]), 
            .O(n2_adj_5136));   // verilog/coms.v(146[4] 295[11])
    defparam select_715_Select_49_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_3_lut_adj_1589 (.I0(\data_in_frame[20] [5]), .I1(\data_in_frame[16] [3]), 
            .I2(n53252), .I3(GND_net), .O(n53234));
    defparam i1_2_lut_3_lut_adj_1589.LUT_INIT = 16'h6969;
    SB_LUT4 n63335_bdd_4_lut (.I0(n63335), .I1(\data_out_frame[9] [7]), 
            .I2(\data_out_frame[8] [7]), .I3(byte_transmit_counter_c[1]), 
            .O(n63338));
    defparam n63335_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_2_lut_4_lut_adj_1590 (.I0(\data_in_frame[15] [0]), .I1(n22813), 
            .I2(n23288), .I3(\data_in_frame[10] [5]), .O(n53375));   // verilog/coms.v(72[16:27])
    defparam i1_2_lut_4_lut_adj_1590.LUT_INIT = 16'h6996;
    SB_LUT4 i13336_3_lut_4_lut (.I0(n8_adj_5286), .I1(n52895), .I2(rx_data[7]), 
            .I3(\data_in_frame[6] [7]), .O(n26940));
    defparam i13336_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_4_lut_adj_1591 (.I0(\data_in_frame[17] [1]), .I1(n54710), 
            .I2(n10_adj_5218), .I3(\data_in_frame[14] [5]), .O(n53329));
    defparam i1_2_lut_4_lut_adj_1591.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_3_lut_adj_1592 (.I0(\data_in_frame[19] [4]), .I1(n23006), 
            .I2(n48781), .I3(GND_net), .O(n47882));
    defparam i1_2_lut_3_lut_adj_1592.LUT_INIT = 16'h9696;
    SB_LUT4 i12980_3_lut_4_lut (.I0(n8_adj_5286), .I1(n52895), .I2(rx_data[1]), 
            .I3(\data_in_frame[6] [1]), .O(n26584));
    defparam i12980_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_4_lut_adj_1593 (.I0(\data_in_frame[17] [0]), .I1(\data_in_frame[19] [1]), 
            .I2(n55031), .I3(n47932), .O(n53489));
    defparam i1_2_lut_4_lut_adj_1593.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_4_lut_adj_1594 (.I0(n47876), .I1(n54891), .I2(n47756), 
            .I3(\data_in_frame[17] [5]), .O(n48785));
    defparam i1_2_lut_4_lut_adj_1594.LUT_INIT = 16'h9669;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_48767 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[6] [4]), .I2(\data_out_frame[7] [4]), .I3(byte_transmit_counter_c[1]), 
            .O(n63497));
    defparam byte_transmit_counter_0__bdd_4_lut_48767.LUT_INIT = 16'he4aa;
    SB_LUT4 i1_2_lut_3_lut_adj_1595 (.I0(\data_in_frame[15] [5]), .I1(\data_in_frame[13] [4]), 
            .I2(n53091), .I3(GND_net), .O(n53144));
    defparam i1_2_lut_3_lut_adj_1595.LUT_INIT = 16'h9696;
    SB_LUT4 i12923_3_lut_4_lut (.I0(n8_adj_5286), .I1(n52895), .I2(rx_data[0]), 
            .I3(\data_in_frame[6] [0]), .O(n26527));
    defparam i12923_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_3_lut_adj_1596 (.I0(\data_in_frame[2] [0]), .I1(\data_in_frame[4]_c [3]), 
            .I2(\data_in_frame[7] [7]), .I3(GND_net), .O(n53589));   // verilog/coms.v(74[16:42])
    defparam i1_2_lut_3_lut_adj_1596.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_4_lut_adj_1597 (.I0(\data_in_frame[2] [0]), .I1(\data_in_frame[4]_c [3]), 
            .I2(n23221), .I3(n53418), .O(Kp_23__N_710));   // verilog/coms.v(74[16:42])
    defparam i2_3_lut_4_lut_adj_1597.LUT_INIT = 16'h6996;
    SB_LUT4 n63497_bdd_4_lut (.I0(n63497), .I1(\data_out_frame[5] [4]), 
            .I2(\data_out_frame[4] [4]), .I3(byte_transmit_counter_c[1]), 
            .O(n56873));
    defparam n63497_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i2_3_lut_4_lut_adj_1598 (.I0(n23252), .I1(n52972), .I2(\data_in_frame[7] [1]), 
            .I3(\data_in_frame[6] [7]), .O(n53607));
    defparam i2_3_lut_4_lut_adj_1598.LUT_INIT = 16'h6996;
    SB_LUT4 i1_3_lut_4_lut_adj_1599 (.I0(n23252), .I1(n52972), .I2(n53243), 
            .I3(\data_in_frame[6] [0]), .O(n53073));
    defparam i1_3_lut_4_lut_adj_1599.LUT_INIT = 16'h9669;
    SB_LUT4 i2_3_lut_4_lut_adj_1600 (.I0(\data_in_frame[7] [6]), .I1(n23666), 
            .I2(n22652), .I3(n53213), .O(n20820));
    defparam i2_3_lut_4_lut_adj_1600.LUT_INIT = 16'h6996;
    SB_LUT4 i21862_2_lut_3_lut (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(\FRAME_MATCHER.i [0]), .I3(GND_net), .O(n35372));
    defparam i21862_2_lut_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 i13391_3_lut_4_lut (.I0(n8_adj_5074), .I1(n52882), .I2(rx_data[1]), 
            .I3(\data_in_frame[9] [1]), .O(n26995));
    defparam i13391_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_3_lut_4_lut_adj_1601 (.I0(\data_in_frame[13] [5]), .I1(n53529), 
            .I2(\data_in_frame[13] [7]), .I3(\data_in_frame[13] [6]), .O(n52952));
    defparam i2_3_lut_4_lut_adj_1601.LUT_INIT = 16'h6996;
    SB_LUT4 equal_291_i8_2_lut_3_lut (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(\FRAME_MATCHER.i [0]), .I3(GND_net), .O(n8_adj_5286));
    defparam equal_291_i8_2_lut_3_lut.LUT_INIT = 16'hf7f7;
    SB_LUT4 i1_2_lut_3_lut_adj_1602 (.I0(reset), .I1(n53712), .I2(n10_adj_5280), 
            .I3(GND_net), .O(n52890));
    defparam i1_2_lut_3_lut_adj_1602.LUT_INIT = 16'hfbfb;
    SB_LUT4 i2_3_lut_4_lut_adj_1603 (.I0(\data_in_frame[16] [4]), .I1(n48798), 
            .I2(n23039), .I3(n53348), .O(n22056));
    defparam i2_3_lut_4_lut_adj_1603.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1604 (.I0(\data_in_frame[16] [4]), .I1(n48798), 
            .I2(n47898), .I3(GND_net), .O(n6_adj_5284));
    defparam i1_2_lut_3_lut_adj_1604.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1605 (.I0(reset), .I1(n53712), .I2(n10_adj_5419), 
            .I3(GND_net), .O(n52882));
    defparam i1_2_lut_3_lut_adj_1605.LUT_INIT = 16'hfbfb;
    SB_LUT4 i2_3_lut_4_lut_adj_1606 (.I0(\data_in_frame[13] [2]), .I1(\data_in_frame[13] [1]), 
            .I2(\data_in_frame[15] [3]), .I3(n53532), .O(n47756));
    defparam i2_3_lut_4_lut_adj_1606.LUT_INIT = 16'h6996;
    SB_LUT4 i5_3_lut_4_lut_adj_1607 (.I0(\data_in_frame[13] [2]), .I1(\data_in_frame[13] [1]), 
            .I2(\data_in_frame[21] [3]), .I3(\data_in_frame[21] [4]), .O(n26_adj_5211));
    defparam i5_3_lut_4_lut_adj_1607.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1608 (.I0(reset), .I1(n53712), .I2(n10_adj_5333), 
            .I3(GND_net), .O(n52895));
    defparam i1_2_lut_3_lut_adj_1608.LUT_INIT = 16'hfbfb;
    SB_LUT4 i1_2_lut_3_lut_adj_1609 (.I0(n22713), .I1(n53352), .I2(\data_in_frame[10] [7]), 
            .I3(GND_net), .O(n23002));
    defparam i1_2_lut_3_lut_adj_1609.LUT_INIT = 16'h9696;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_48619 (.I0(byte_transmit_counter_c[1]), 
            .I1(n57007), .I2(n57008), .I3(\byte_transmit_counter[2] ), 
            .O(n63329));
    defparam byte_transmit_counter_1__bdd_4_lut_48619.LUT_INIT = 16'he4aa;
    SB_LUT4 i5_3_lut_4_lut_adj_1610 (.I0(n22713), .I1(n53352), .I2(n10_adj_5282), 
            .I3(n23509), .O(n54891));
    defparam i5_3_lut_4_lut_adj_1610.LUT_INIT = 16'h6996;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_48743 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[6] [2]), .I2(\data_out_frame[7] [2]), .I3(byte_transmit_counter_c[1]), 
            .O(n63491));
    defparam byte_transmit_counter_0__bdd_4_lut_48743.LUT_INIT = 16'he4aa;
    SB_LUT4 i1_2_lut_3_lut_adj_1611 (.I0(n52952), .I1(n53580), .I2(n22822), 
            .I3(GND_net), .O(n48511));
    defparam i1_2_lut_3_lut_adj_1611.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_4_lut_adj_1612 (.I0(n20672), .I1(n53157), .I2(\data_in_frame[10] [3]), 
            .I3(\data_in_frame[12] [4]), .O(n52937));
    defparam i1_2_lut_4_lut_adj_1612.LUT_INIT = 16'h6996;
    SB_LUT4 equal_290_i10_2_lut_3_lut (.I0(\FRAME_MATCHER.i [4]), .I1(\FRAME_MATCHER.i [5]), 
            .I2(\FRAME_MATCHER.i [3]), .I3(GND_net), .O(n10_adj_5419));   // verilog/coms.v(154[7:23])
    defparam equal_290_i10_2_lut_3_lut.LUT_INIT = 16'hefef;
    SB_LUT4 i1_2_lut_4_lut_adj_1613 (.I0(n20672), .I1(n53157), .I2(\data_in_frame[10] [3]), 
            .I3(\data_in_frame[12] [5]), .O(n52940));
    defparam i1_2_lut_4_lut_adj_1613.LUT_INIT = 16'h6996;
    SB_LUT4 equal_298_i10_2_lut_3_lut (.I0(\FRAME_MATCHER.i [4]), .I1(\FRAME_MATCHER.i [5]), 
            .I2(\FRAME_MATCHER.i [3]), .I3(GND_net), .O(n10_adj_5333));   // verilog/coms.v(154[7:23])
    defparam equal_298_i10_2_lut_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i1_2_lut_2_lut (.I0(reset), .I1(\FRAME_MATCHER.i_31__N_2322 ), 
            .I2(GND_net), .I3(GND_net), .O(n52664));   // verilog/coms.v(128[12] 296[6])
    defparam i1_2_lut_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i2_2_lut_3_lut_3_lut (.I0(Kp_23__N_1583), .I1(n29100), .I2(reset), 
            .I3(GND_net), .O(n19639));
    defparam i2_2_lut_3_lut_3_lut.LUT_INIT = 16'h0808;
    SB_LUT4 i1_2_lut_4_lut_adj_1614 (.I0(n48497), .I1(n10_adj_5135), .I2(n4), 
            .I3(n53314), .O(n53315));
    defparam i1_2_lut_4_lut_adj_1614.LUT_INIT = 16'h6996;
    SB_LUT4 i2_2_lut_3_lut_adj_1615 (.I0(\data_out_frame[10] [4]), .I1(\data_out_frame[10] [6]), 
            .I2(\data_out_frame[6] [0]), .I3(GND_net), .O(n10_adj_5133));   // verilog/coms.v(86[17:70])
    defparam i2_2_lut_3_lut_adj_1615.LUT_INIT = 16'h9696;
    SB_LUT4 n63329_bdd_4_lut (.I0(n63329), .I1(n56942), .I2(n56941), .I3(\byte_transmit_counter[2] ), 
            .O(n63332));
    defparam n63329_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i13394_3_lut_4_lut (.I0(n8_adj_5074), .I1(n52882), .I2(rx_data[2]), 
            .I3(\data_in_frame[9] [2]), .O(n26998));
    defparam i13394_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_4_lut_adj_1616 (.I0(\data_out_frame[10] [1]), .I1(\data_out_frame[9] [7]), 
            .I2(\data_out_frame[7] [5]), .I3(\data_out_frame[7] [6]), .O(n53518));
    defparam i1_2_lut_4_lut_adj_1616.LUT_INIT = 16'h6996;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_48604 (.I0(byte_transmit_counter_c[1]), 
            .I1(n56944), .I2(n56945), .I3(\byte_transmit_counter[2] ), 
            .O(n63323));
    defparam byte_transmit_counter_1__bdd_4_lut_48604.LUT_INIT = 16'he4aa;
    SB_LUT4 i13412_3_lut_4_lut (.I0(n8), .I1(n52882), .I2(rx_data[0]), 
            .I3(\data_in_frame[10] [0]), .O(n27016));
    defparam i13412_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 n63323_bdd_4_lut (.I0(n63323), .I1(n56834), .I2(n56833), .I3(\byte_transmit_counter[2] ), 
            .O(n63326));
    defparam n63323_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i2_2_lut_3_lut_adj_1617 (.I0(\data_in_frame[15] [6]), .I1(\data_in_frame[13] [4]), 
            .I2(\data_in_frame[18] [0]), .I3(GND_net), .O(n7_adj_5221));   // verilog/coms.v(77[16:43])
    defparam i2_2_lut_3_lut_adj_1617.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1618 (.I0(\data_out_frame[9] [7]), .I1(\data_out_frame[7] [5]), 
            .I2(\data_out_frame[7] [6]), .I3(GND_net), .O(n23123));   // verilog/coms.v(76[16:27])
    defparam i1_2_lut_3_lut_adj_1618.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_4_lut_adj_1619 (.I0(\data_out_frame[14] [6]), .I1(n53535), 
            .I2(n10_adj_5129), .I3(\data_out_frame[10] [3]), .O(n4));   // verilog/coms.v(86[17:63])
    defparam i1_2_lut_4_lut_adj_1619.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1620 (.I0(\data_out_frame[4] [1]), .I1(\data_out_frame[4] [2]), 
            .I2(\data_out_frame[6] [3]), .I3(GND_net), .O(n22533));   // verilog/coms.v(76[16:43])
    defparam i1_2_lut_3_lut_adj_1620.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1621 (.I0(\data_out_frame[5] [6]), .I1(\data_out_frame[10] [4]), 
            .I2(\data_out_frame[6] [1]), .I3(GND_net), .O(n53332));   // verilog/coms.v(86[17:70])
    defparam i1_2_lut_3_lut_adj_1621.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1622 (.I0(\data_out_frame[5] [5]), .I1(\data_out_frame[7] [7]), 
            .I2(\data_out_frame[6] [0]), .I3(GND_net), .O(n53535));   // verilog/coms.v(76[16:27])
    defparam i1_2_lut_3_lut_adj_1622.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_4_lut_adj_1623 (.I0(\data_out_frame[17] [0]), .I1(n53094), 
            .I2(n53267), .I3(\data_out_frame[21] [4]), .O(n55477));
    defparam i2_3_lut_4_lut_adj_1623.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_1624 (.I0(\data_out_frame[12] [1]), .I1(\data_out_frame[14] [3]), 
            .I2(n22545), .I3(n21977), .O(n47750));
    defparam i2_3_lut_4_lut_adj_1624.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1625 (.I0(\data_out_frame[5] [6]), .I1(\data_out_frame[5] [2]), 
            .I2(\data_out_frame[7] [4]), .I3(GND_net), .O(n6_adj_5120));
    defparam i1_2_lut_3_lut_adj_1625.LUT_INIT = 16'h9696;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_48609 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[10] [6]), .I2(\data_out_frame[11] [6]), 
            .I3(byte_transmit_counter_c[1]), .O(n63317));
    defparam byte_transmit_counter_0__bdd_4_lut_48609.LUT_INIT = 16'he4aa;
    SB_LUT4 n63317_bdd_4_lut (.I0(n63317), .I1(\data_out_frame[9] [6]), 
            .I2(\data_out_frame[8] [6]), .I3(byte_transmit_counter_c[1]), 
            .O(n63320));
    defparam n63317_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_3__bdd_4_lut_48772 (.I0(byte_transmit_counter_c[3]), 
            .I1(n61989), .I2(n59928), .I3(byte_transmit_counter_c[4]), 
            .O(n63311));
    defparam byte_transmit_counter_3__bdd_4_lut_48772.LUT_INIT = 16'he4aa;
    SB_LUT4 n63311_bdd_4_lut (.I0(n63311), .I1(n14_adj_5348), .I2(n7_adj_5376), 
            .I3(byte_transmit_counter_c[4]), .O(tx_data[6]));
    defparam n63311_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i13415_3_lut_4_lut (.I0(n8), .I1(n52882), .I2(rx_data[1]), 
            .I3(\data_in_frame[10] [1]), .O(n27019));
    defparam i13415_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i45286_2_lut (.I0(\FRAME_MATCHER.i [31]), .I1(\FRAME_MATCHER.i_31__N_2318 ), 
            .I2(GND_net), .I3(GND_net), .O(n59781));   // verilog/coms.v(155[12:15])
    defparam i45286_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i48560_1_lut (.I0(n3133), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n63273));   // verilog/coms.v(146[4] 295[11])
    defparam i48560_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i13397_3_lut_4_lut (.I0(n8_adj_5074), .I1(n52882), .I2(rx_data[3]), 
            .I3(\data_in_frame[9] [3]), .O(n27001));
    defparam i13397_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_48595 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[10] [4]), .I2(\data_out_frame[11] [4]), 
            .I3(byte_transmit_counter_c[1]), .O(n63305));
    defparam byte_transmit_counter_0__bdd_4_lut_48595.LUT_INIT = 16'he4aa;
    SB_LUT4 n63305_bdd_4_lut (.I0(n63305), .I1(\data_out_frame[9] [4]), 
            .I2(\data_out_frame[8] [4]), .I3(byte_transmit_counter_c[1]), 
            .O(n56961));
    defparam n63305_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i20308_3_lut (.I0(\control_mode[4] ), .I1(\data_in_frame[1][4] ), 
            .I2(n19639), .I3(GND_net), .O(n26912));
    defparam i20308_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i20307_3_lut (.I0(control_mode_c[3]), .I1(\data_in_frame[1][3] ), 
            .I2(n19639), .I3(GND_net), .O(n26913));
    defparam i20307_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i20306_3_lut (.I0(control_mode_c[2]), .I1(\data_in_frame[1][2] ), 
            .I2(n19639), .I3(GND_net), .O(n26914));
    defparam i20306_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_48586 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[10] [3]), .I2(\data_out_frame[11] [3]), 
            .I3(byte_transmit_counter_c[1]), .O(n63299));
    defparam byte_transmit_counter_0__bdd_4_lut_48586.LUT_INIT = 16'he4aa;
    SB_LUT4 i17375_3_lut (.I0(\control_mode[1] ), .I1(\data_in_frame[1] [1]), 
            .I2(n19639), .I3(GND_net), .O(n26915));
    defparam i17375_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11538_4_lut (.I0(n10_adj_5419), .I1(reset), .I2(n53712), 
            .I3(n8_adj_5335), .O(n25141));
    defparam i11538_4_lut.LUT_INIT = 16'hffef;
    SB_LUT4 n63491_bdd_4_lut (.I0(n63491), .I1(\data_out_frame[5] [2]), 
            .I2(\data_out_frame[4] [2]), .I3(byte_transmit_counter_c[1]), 
            .O(n56877));
    defparam n63491_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i13400_3_lut_4_lut (.I0(n8_adj_5074), .I1(n52882), .I2(rx_data[4]), 
            .I3(\data_in_frame[9] [4]), .O(n27004));
    defparam i13400_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13418_3_lut_4_lut (.I0(n8), .I1(n52882), .I2(rx_data[2]), 
            .I3(\data_in_frame[10] [2]), .O(n27022));
    defparam i13418_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13421_3_lut_4_lut (.I0(n8), .I1(n52882), .I2(rx_data[3]), 
            .I3(\data_in_frame[10] [3]), .O(n27025));
    defparam i13421_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 n63299_bdd_4_lut (.I0(n63299), .I1(\data_out_frame[9] [3]), 
            .I2(\data_out_frame[8] [3]), .I3(byte_transmit_counter_c[1]), 
            .O(n63302));
    defparam n63299_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_4__bdd_4_lut (.I0(byte_transmit_counter_c[4]), 
            .I1(n56886), .I2(n33004), .I3(byte_transmit_counter_c[3]), 
            .O(n63293));
    defparam byte_transmit_counter_4__bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_LUT4 i13424_3_lut_4_lut (.I0(n8), .I1(n52882), .I2(rx_data[4]), 
            .I3(\data_in_frame[10] [4]), .O(n27028));
    defparam i13424_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 n63293_bdd_4_lut (.I0(n63293), .I1(n21), .I2(n56877), .I3(byte_transmit_counter_c[3]), 
            .O(n63296));
    defparam n63293_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_2__bdd_4_lut_48638 (.I0(\byte_transmit_counter[2] ), 
            .I1(n56961), .I2(n56853), .I3(byte_transmit_counter_c[3]), 
            .O(n63287));
    defparam byte_transmit_counter_2__bdd_4_lut_48638.LUT_INIT = 16'he4aa;
    SB_LUT4 i12_4_lut_3_lut_4_lut (.I0(n22822), .I1(n23402), .I2(\data_in_frame[21] [5]), 
            .I3(n53509), .O(n33_adj_5212));   // verilog/coms.v(75[16:43])
    defparam i12_4_lut_3_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 n63287_bdd_4_lut (.I0(n63287), .I1(n56873), .I2(n56872), .I3(byte_transmit_counter_c[3]), 
            .O(n63290));
    defparam n63287_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_2_lut_3_lut_adj_1626 (.I0(n53394), .I1(\data_out_frame[14] [5]), 
            .I2(n52968), .I3(GND_net), .O(n23432));   // verilog/coms.v(76[16:43])
    defparam i1_2_lut_3_lut_adj_1626.LUT_INIT = 16'h9696;
    SB_LUT4 i12460_3_lut_4_lut (.I0(Kp_23__N_1583), .I1(n29100), .I2(\data_in_frame[16] [0]), 
            .I3(\deadband[0] ), .O(n26064));
    defparam i12460_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_48581 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[14] [7]), .I2(\data_out_frame[15] [7]), 
            .I3(byte_transmit_counter_c[1]), .O(n63281));
    defparam byte_transmit_counter_0__bdd_4_lut_48581.LUT_INIT = 16'he4aa;
    SB_LUT4 i12461_3_lut_4_lut (.I0(Kp_23__N_1583), .I1(n29100), .I2(\data_in_frame[13] [0]), 
            .I3(IntegralLimit[0]), .O(n26065));
    defparam i12461_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 n63281_bdd_4_lut (.I0(n63281), .I1(\data_out_frame[13] [7]), 
            .I2(\data_out_frame[12] [7]), .I3(byte_transmit_counter_c[1]), 
            .O(n63284));
    defparam n63281_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i13427_3_lut_4_lut (.I0(n8), .I1(n52882), .I2(rx_data[5]), 
            .I3(\data_in_frame[10] [5]), .O(n27031));
    defparam i13427_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i12468_3_lut_4_lut (.I0(Kp_23__N_1583), .I1(n29100), .I2(\data_in_frame[3] [0]), 
            .I3(\Kp[0] ), .O(n26072));
    defparam i12468_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i12979_3_lut_4_lut (.I0(Kp_23__N_1583), .I1(n29100), .I2(\data_in_frame[12] [4]), 
            .I3(IntegralLimit[12]), .O(n26583));
    defparam i12979_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i11_3_lut_4_lut_adj_1627 (.I0(n8), .I1(n52882), .I2(\data_in_frame[10] [7]), 
            .I3(rx_data[7]), .O(n52311));
    defparam i11_3_lut_4_lut_adj_1627.LUT_INIT = 16'hf1e0;
    SB_LUT4 i12985_3_lut_4_lut (.I0(Kp_23__N_1583), .I1(n29100), .I2(\data_in_frame[12] [3]), 
            .I3(IntegralLimit[11]), .O(n26589));
    defparam i12985_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i12988_3_lut_4_lut (.I0(Kp_23__N_1583), .I1(n29100), .I2(\data_in_frame[12] [2]), 
            .I3(IntegralLimit[10]), .O(n26592));
    defparam i12988_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i13004_3_lut_4_lut (.I0(Kp_23__N_1583), .I1(n29100), .I2(\data_in_frame[12] [1]), 
            .I3(IntegralLimit[9]), .O(n26608));
    defparam i13004_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i17129_3_lut_4_lut (.I0(Kp_23__N_1583), .I1(n29100), .I2(\data_in_frame[5] [0]), 
            .I3(\Ki[0] ), .O(n26081));
    defparam i17129_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i12480_3_lut_4_lut (.I0(Kp_23__N_1583), .I1(n29100), .I2(\data_in_frame[10] [0]), 
            .I3(PWMLimit[0]), .O(n26084));
    defparam i12480_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i12482_3_lut_4_lut (.I0(Kp_23__N_1583), .I1(n29100), .I2(\data_in_frame[3][6] ), 
            .I3(\Kp[6] ), .O(n26086));
    defparam i12482_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i13048_3_lut (.I0(\data_in_frame[18]_c [6]), .I1(rx_data[6]), 
            .I2(n25127), .I3(GND_net), .O(n26652));   // verilog/coms.v(128[12] 296[6])
    defparam i13048_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_4_lut_adj_1628 (.I0(n54590), .I1(n47956), .I2(n48787), 
            .I3(\data_out_frame[21] [7]), .O(n6_adj_5099));
    defparam i1_2_lut_4_lut_adj_1628.LUT_INIT = 16'h9669;
    SB_LUT4 i13057_3_lut_4_lut (.I0(Kp_23__N_1583), .I1(n29100), .I2(\data_in_frame[12] [0]), 
            .I3(IntegralLimit[8]), .O(n26661));
    defparam i13057_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1_2_lut_3_lut_adj_1629 (.I0(\data_out_frame[4] [0]), .I1(\data_out_frame[4] [1]), 
            .I2(\data_out_frame[6] [2]), .I3(GND_net), .O(n22529));   // verilog/coms.v(75[16:43])
    defparam i1_2_lut_3_lut_adj_1629.LUT_INIT = 16'h9696;
    SB_LUT4 i13076_3_lut_4_lut (.I0(Kp_23__N_1583), .I1(n29100), .I2(\data_in_frame[13] [7]), 
            .I3(IntegralLimit[7]), .O(n26680));
    defparam i13076_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2_2_lut_4_lut (.I0(n23083), .I1(n22519), .I2(\data_out_frame[4] [7]), 
            .I3(n53131), .O(n6_adj_5093));
    defparam i2_2_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i13101_3_lut_4_lut (.I0(Kp_23__N_1583), .I1(n29100), .I2(\data_in_frame[13] [6]), 
            .I3(IntegralLimit[6]), .O(n26705));
    defparam i13101_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1_2_lut_3_lut_adj_1630 (.I0(\data_out_frame[7] [1]), .I1(\data_out_frame[9] [3]), 
            .I2(n23720), .I3(GND_net), .O(n53459));
    defparam i1_2_lut_3_lut_adj_1630.LUT_INIT = 16'h9696;
    SB_LUT4 i13124_3_lut_4_lut (.I0(Kp_23__N_1583), .I1(n29100), .I2(\data_in_frame[2] [7]), 
            .I3(\Kp[15] ), .O(n26728));
    defparam i13124_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2_2_lut_3_lut_adj_1631 (.I0(\data_out_frame[5] [5]), .I1(\data_out_frame[5] [4]), 
            .I2(n53308), .I3(GND_net), .O(n6_adj_5078));   // verilog/coms.v(86[17:70])
    defparam i2_2_lut_3_lut_adj_1631.LUT_INIT = 16'h9696;
    SB_LUT4 i3_2_lut_4_lut_adj_1632 (.I0(n22533), .I1(n53043), .I2(\data_out_frame[9] [4]), 
            .I3(\data_out_frame[9] [7]), .O(n12_adj_5072));
    defparam i3_2_lut_4_lut_adj_1632.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1633 (.I0(n22533), .I1(n53043), .I2(\data_out_frame[11] [2]), 
            .I3(GND_net), .O(n53453));
    defparam i1_2_lut_3_lut_adj_1633.LUT_INIT = 16'h9696;
    SB_LUT4 i13132_3_lut_4_lut (.I0(Kp_23__N_1583), .I1(n29100), .I2(\data_in_frame[13] [5]), 
            .I3(IntegralLimit[5]), .O(n26736));
    defparam i13132_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i13133_3_lut_4_lut (.I0(Kp_23__N_1583), .I1(n29100), .I2(\data_in_frame[13] [4]), 
            .I3(IntegralLimit[4]), .O(n26737));
    defparam i13133_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1_2_lut_3_lut_adj_1634 (.I0(n54765), .I1(n47853), .I2(n48777), 
            .I3(GND_net), .O(n47777));
    defparam i1_2_lut_3_lut_adj_1634.LUT_INIT = 16'h6969;
    SB_LUT4 i1_2_lut_4_lut_adj_1635 (.I0(\data_out_frame[22] [1]), .I1(n47853), 
            .I2(n47956), .I3(n48773), .O(n48885));
    defparam i1_2_lut_4_lut_adj_1635.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1636 (.I0(n53068), .I1(\data_out_frame[17] [6]), 
            .I2(\data_out_frame[17] [4]), .I3(GND_net), .O(n6_adj_5063));
    defparam i1_2_lut_3_lut_adj_1636.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_4_lut_adj_1637 (.I0(\data_out_frame[11] [3]), .I1(n23083), 
            .I2(n22519), .I3(\data_out_frame[4] [7]), .O(n53462));
    defparam i1_2_lut_4_lut_adj_1637.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_adj_1638 (.I0(\data_out_frame[15] [7]), .I1(n23256), 
            .I2(n47860), .I3(\data_out_frame[13] [6]), .O(n53357));
    defparam i1_2_lut_4_lut_adj_1638.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1639 (.I0(\data_out_frame[9] [1]), .I1(\data_out_frame[8] [7]), 
            .I2(n23417), .I3(GND_net), .O(n52998));
    defparam i1_2_lut_3_lut_adj_1639.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_4_lut_adj_1640 (.I0(n54590), .I1(n2142), .I2(\data_out_frame[22] [3]), 
            .I3(\data_out_frame[22] [4]), .O(n52932));
    defparam i1_2_lut_4_lut_adj_1640.LUT_INIT = 16'h9669;
    SB_LUT4 i13134_3_lut_4_lut (.I0(Kp_23__N_1583), .I1(n29100), .I2(\data_in_frame[2] [6]), 
            .I3(\Kp[14] ), .O(n26738));
    defparam i13134_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i13135_3_lut_4_lut (.I0(Kp_23__N_1583), .I1(n29100), .I2(\data_in_frame[13] [3]), 
            .I3(IntegralLimit[3]), .O(n26739));
    defparam i13135_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1_2_lut_3_lut_adj_1641 (.I0(\data_out_frame[15] [4]), .I1(\data_out_frame[15] [3]), 
            .I2(n53559), .I3(GND_net), .O(n53082));
    defparam i1_2_lut_3_lut_adj_1641.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1642 (.I0(\data_out_frame[21] [7]), .I1(\data_out_frame[21] [6]), 
            .I2(n53314), .I3(GND_net), .O(n53279));
    defparam i1_2_lut_3_lut_adj_1642.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_4_lut_adj_1643 (.I0(\data_out_frame[22] [0]), .I1(n22564), 
            .I2(n53068), .I3(\data_out_frame[17] [4]), .O(n23712));
    defparam i1_2_lut_4_lut_adj_1643.LUT_INIT = 16'h6996;
    SB_LUT4 i13150_3_lut_4_lut (.I0(Kp_23__N_1583), .I1(n29100), .I2(\data_in_frame[2] [5]), 
            .I3(\Kp[13] ), .O(n26754));
    defparam i13150_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i13151_3_lut_4_lut (.I0(Kp_23__N_1583), .I1(n29100), .I2(\data_in_frame[13] [2]), 
            .I3(IntegralLimit[2]), .O(n26755));
    defparam i13151_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i39052_2_lut_3_lut (.I0(n3133), .I1(rx_data_ready), .I2(\FRAME_MATCHER.rx_data_ready_prev ), 
            .I3(GND_net), .O(n53712));
    defparam i39052_2_lut_3_lut.LUT_INIT = 16'h0808;
    uart_tx tx (.r_Clock_Count({r_Clock_Count}), .clk16MHz(clk16MHz), .n24612(n24612), 
            .n36763(n36763), .GND_net(GND_net), .VCC_net(VCC_net), .tx_o(tx_o), 
            .tx_data({tx_data[7:6], Open_24, Open_25, Open_26, Open_27, 
            Open_28, tx_data[0]}), .byte_transmit_counter({byte_transmit_counter_c[7:3], 
            \byte_transmit_counter[2] , byte_transmit_counter_c[1], byte_transmit_counter[0]}), 
            .n44(n44_adj_5364), .n26829(n26829), .\r_Bit_Index[0] (\r_Bit_Index[0] ), 
            .\data_out_frame[14][5] (\data_out_frame[14] [5]), .\data_out_frame[15][5] (\data_out_frame[15] [5]), 
            .\data_out_frame[13][5] (\data_out_frame[13] [5]), .\data_out_frame[12][5] (\data_out_frame[12] [5]), 
            .\tx_data[4] (tx_data[4]), .\tx_data[3] (tx_data[3]), .\tx_data[2] (tx_data[2]), 
            .\tx_data[1] (tx_data[1]), .tx_active(tx_active), .\o_Rx_DV_N_3261[12] (\o_Rx_DV_N_3261[12] ), 
            .n4837(n4837), .\o_Rx_DV_N_3261[24] (\o_Rx_DV_N_3261[24] ), 
            .n29(n29), .n23(n23), .\r_SM_Main_2__N_3318[0] (r_SM_Main_2__N_3318[0]), 
            .n27(n27), .n36757(n36757), .n47(n47), .tx_transmit_N_3189(tx_transmit_N_3189), 
            .\data_out_frame[16][5] (\data_out_frame[16] [5]), .\data_out_frame[17][5] (\data_out_frame[17] [5]), 
            .n24853(n24853), .\data_out_frame[1][5] (\data_out_frame[1][5] ), 
            .n33453(n33453), .n56920(n56920), .n56922(n56922), .n57324(n57324), 
            .n59726(n59726), .n59727(n59727), .n56924(n56924), .n56923(n56923), 
            .tx_enable(tx_enable)) /* synthesis syn_module_defined=1 */ ;   // verilog/coms.v(108[25:94])
    uart_rx rx (.baudrate({baudrate}), .n24621(n24621), .clk16MHz(clk16MHz), 
            .n53789(n53789), .GND_net(GND_net), .r_Clock_Count({r_Clock_Count_adj_13}), 
            .VCC_net(VCC_net), .n26516(n26516), .rx_data({rx_data}), .\r_SM_Main[2] (\r_SM_Main[2] ), 
            .r_Rx_Data(r_Rx_Data), .RX_N_42(RX_N_42), .\o_Rx_DV_N_3261[24] (\o_Rx_DV_N_3261[24] ), 
            .n27(n27), .n29(n29), .\r_Bit_Index[0] (\r_Bit_Index[0]_adj_12 ), 
            .n55980(n55980), .n23(n23), .n55948(n55948), .\o_Rx_DV_N_3261[12] (\o_Rx_DV_N_3261[12] ), 
            .n26445(n26445), .\o_Rx_DV_N_3261[8] (\o_Rx_DV_N_3261[8] ), 
            .n26443(n26443), .\o_Rx_DV_N_3261[7] (\o_Rx_DV_N_3261[7] ), 
            .\o_Rx_DV_N_3261[6] (\o_Rx_DV_N_3261[6] ), .\o_Rx_DV_N_3261[5] (\o_Rx_DV_N_3261[5] ), 
            .n33(n33), .\o_Rx_DV_N_3261[4] (\o_Rx_DV_N_3261[4] ), .\o_Rx_DV_N_3261[3] (\o_Rx_DV_N_3261[3] ), 
            .\o_Rx_DV_N_3261[2] (\o_Rx_DV_N_3261[2] ), .\o_Rx_DV_N_3261[1] (\o_Rx_DV_N_3261[1] ), 
            .\o_Rx_DV_N_3261[0] (\o_Rx_DV_N_3261[0] ), .n27051(n27051), 
            .n26970(n26970), .n4834(n4834), .n52823(n52823), .n26836(n26836), 
            .n48959(n48959), .rx_data_ready(rx_data_ready), .n26832(n26832), 
            .n55964(n55964), .n55996(n55996), .\r_SM_Main[1] (\r_SM_Main[1] ), 
            .\r_SM_Main_2__N_3219[1] (\r_SM_Main_2__N_3219[1] ), .n55461(n55461), 
            .n26587(n26587), .n26062(n26062), .n55884(n55884), .n55900(n55900), 
            .n55916(n55916), .n55932(n55932), .n55814(n55814), .n24535(n24535), 
            .n34(n34)) /* synthesis syn_module_defined=1 */ ;   // verilog/coms.v(94[25:68])
    
endmodule
//
// Verilog Description of module uart_tx
//

module uart_tx (r_Clock_Count, clk16MHz, n24612, n36763, GND_net, 
            VCC_net, tx_o, tx_data, byte_transmit_counter, n44, n26829, 
            \r_Bit_Index[0] , \data_out_frame[14][5] , \data_out_frame[15][5] , 
            \data_out_frame[13][5] , \data_out_frame[12][5] , \tx_data[4] , 
            \tx_data[3] , \tx_data[2] , \tx_data[1] , tx_active, \o_Rx_DV_N_3261[12] , 
            n4837, \o_Rx_DV_N_3261[24] , n29, n23, \r_SM_Main_2__N_3318[0] , 
            n27, n36757, n47, tx_transmit_N_3189, \data_out_frame[16][5] , 
            \data_out_frame[17][5] , n24853, \data_out_frame[1][5] , n33453, 
            n56920, n56922, n57324, n59726, n59727, n56924, n56923, 
            tx_enable) /* synthesis syn_module_defined=1 */ ;
    output [8:0]r_Clock_Count;
    input clk16MHz;
    output n24612;
    input n36763;
    input GND_net;
    input VCC_net;
    output tx_o;
    input [7:0]tx_data;
    input [7:0]byte_transmit_counter;
    output n44;
    input n26829;
    output \r_Bit_Index[0] ;
    input \data_out_frame[14][5] ;
    input \data_out_frame[15][5] ;
    input \data_out_frame[13][5] ;
    input \data_out_frame[12][5] ;
    input \tx_data[4] ;
    input \tx_data[3] ;
    input \tx_data[2] ;
    input \tx_data[1] ;
    output tx_active;
    input \o_Rx_DV_N_3261[12] ;
    input n4837;
    input \o_Rx_DV_N_3261[24] ;
    input n29;
    input n23;
    input \r_SM_Main_2__N_3318[0] ;
    input n27;
    output n36757;
    output n47;
    output tx_transmit_N_3189;
    input \data_out_frame[16][5] ;
    input \data_out_frame[17][5] ;
    input n24853;
    input \data_out_frame[1][5] ;
    input n33453;
    input n56920;
    input n56922;
    input n57324;
    input n59726;
    input n59727;
    input n56924;
    input n56923;
    output tx_enable;
    
    wire clk16MHz /* synthesis SET_AS_NETWORK=clk16MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(31[6:14])
    wire [8:0]n41;
    
    wire n1, n25952;
    wire [2:0]n460;
    wire [2:0]r_Bit_Index;   // verilog/uart_tx.v(34[16:27])
    
    wire n36762;
    wire [2:0]r_SM_Main;   // verilog/uart_tx.v(32[16:25])
    
    wire n46684, n46683, n46682, n46681, n46680, n46679, n46678, 
        n46677, n3, n21898;
    wire [7:0]r_Tx_Data;   // verilog/uart_tx.v(35[16:25])
    
    wire n19213, n109, n55301, n63413, n63416, n3_adj_5049;
    wire [7:0]tx_data_c;   // verilog/coms.v(106[13:20])
    
    wire n48965, n63731, n38, n59798, n59795, n3_adj_5050, n63362, 
        n56836, n56837, n56840, n56839, n14, n15, n55736, n36774, 
        n53849, n63359, n59753, n57004, n57002, n57005, n63350, 
        n57003, n57006, n55742, n63347;
    
    SB_DFFESR r_Clock_Count_1951__i0 (.Q(r_Clock_Count[0]), .C(clk16MHz), 
            .E(n1), .D(n41[0]), .R(n25952));   // verilog/uart_tx.v(119[34:51])
    SB_DFFESR r_Bit_Index_i1 (.Q(r_Bit_Index[1]), .C(clk16MHz), .E(n24612), 
            .D(n460[1]), .R(n36762));   // verilog/uart_tx.v(41[10] 144[8])
    SB_DFFESR r_Bit_Index_i2 (.Q(r_Bit_Index[2]), .C(clk16MHz), .E(n24612), 
            .D(n460[2]), .R(n36762));   // verilog/uart_tx.v(41[10] 144[8])
    SB_LUT4 i48314_4_lut (.I0(r_SM_Main[2]), .I1(n36763), .I2(r_SM_Main[1]), 
            .I3(r_SM_Main[0]), .O(n25952));
    defparam i48314_4_lut.LUT_INIT = 16'h1115;
    SB_DFFESR r_Clock_Count_1951__i8 (.Q(r_Clock_Count[8]), .C(clk16MHz), 
            .E(n1), .D(n41[8]), .R(n25952));   // verilog/uart_tx.v(119[34:51])
    SB_DFFESR r_Clock_Count_1951__i7 (.Q(r_Clock_Count[7]), .C(clk16MHz), 
            .E(n1), .D(n41[7]), .R(n25952));   // verilog/uart_tx.v(119[34:51])
    SB_DFFESR r_Clock_Count_1951__i6 (.Q(r_Clock_Count[6]), .C(clk16MHz), 
            .E(n1), .D(n41[6]), .R(n25952));   // verilog/uart_tx.v(119[34:51])
    SB_DFFESR r_Clock_Count_1951__i5 (.Q(r_Clock_Count[5]), .C(clk16MHz), 
            .E(n1), .D(n41[5]), .R(n25952));   // verilog/uart_tx.v(119[34:51])
    SB_DFFESR r_Clock_Count_1951__i4 (.Q(r_Clock_Count[4]), .C(clk16MHz), 
            .E(n1), .D(n41[4]), .R(n25952));   // verilog/uart_tx.v(119[34:51])
    SB_DFFESR r_Clock_Count_1951__i3 (.Q(r_Clock_Count[3]), .C(clk16MHz), 
            .E(n1), .D(n41[3]), .R(n25952));   // verilog/uart_tx.v(119[34:51])
    SB_DFFESR r_Clock_Count_1951__i2 (.Q(r_Clock_Count[2]), .C(clk16MHz), 
            .E(n1), .D(n41[2]), .R(n25952));   // verilog/uart_tx.v(119[34:51])
    SB_DFFESR r_Clock_Count_1951__i1 (.Q(r_Clock_Count[1]), .C(clk16MHz), 
            .E(n1), .D(n41[1]), .R(n25952));   // verilog/uart_tx.v(119[34:51])
    SB_LUT4 i1_1_lut (.I0(r_SM_Main[2]), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n1));
    defparam i1_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 r_Clock_Count_1951_add_4_10_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[8]), .I3(n46684), .O(n41[8])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1951_add_4_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 r_Clock_Count_1951_add_4_9_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[7]), .I3(n46683), .O(n41[7])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1951_add_4_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_1951_add_4_9 (.CI(n46683), .I0(GND_net), .I1(r_Clock_Count[7]), 
            .CO(n46684));
    SB_LUT4 r_Clock_Count_1951_add_4_8_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[6]), .I3(n46682), .O(n41[6])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1951_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_1951_add_4_8 (.CI(n46682), .I0(GND_net), .I1(r_Clock_Count[6]), 
            .CO(n46683));
    SB_LUT4 r_Clock_Count_1951_add_4_7_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[5]), .I3(n46681), .O(n41[5])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1951_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_1951_add_4_7 (.CI(n46681), .I0(GND_net), .I1(r_Clock_Count[5]), 
            .CO(n46682));
    SB_LUT4 r_Clock_Count_1951_add_4_6_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[4]), .I3(n46680), .O(n41[4])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1951_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_1951_add_4_6 (.CI(n46680), .I0(GND_net), .I1(r_Clock_Count[4]), 
            .CO(n46681));
    SB_LUT4 r_Clock_Count_1951_add_4_5_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[3]), .I3(n46679), .O(n41[3])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1951_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_1951_add_4_5 (.CI(n46679), .I0(GND_net), .I1(r_Clock_Count[3]), 
            .CO(n46680));
    SB_LUT4 r_Clock_Count_1951_add_4_4_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[2]), .I3(n46678), .O(n41[2])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1951_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_1951_add_4_4 (.CI(n46678), .I0(GND_net), .I1(r_Clock_Count[2]), 
            .CO(n46679));
    SB_LUT4 r_Clock_Count_1951_add_4_3_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[1]), .I3(n46677), .O(n41[1])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1951_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_1951_add_4_3 (.CI(n46677), .I0(GND_net), .I1(r_Clock_Count[1]), 
            .CO(n46678));
    SB_LUT4 r_Clock_Count_1951_add_4_2_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[0]), .I3(VCC_net), .O(n41[0])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1951_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_1951_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(r_Clock_Count[0]), 
            .CO(n46677));
    SB_DFFE o_Tx_Serial_51 (.Q(tx_o), .C(clk16MHz), .E(n1), .D(n3));   // verilog/uart_tx.v(41[10] 144[8])
    SB_DFFE r_Tx_Data_i0 (.Q(r_Tx_Data[0]), .C(clk16MHz), .E(n21898), 
            .D(tx_data[0]));   // verilog/uart_tx.v(41[10] 144[8])
    SB_DFFSR r_SM_Main_i0 (.Q(r_SM_Main[0]), .C(clk16MHz), .D(n19213), 
            .R(r_SM_Main[2]));   // verilog/uart_tx.v(41[10] 144[8])
    SB_LUT4 i1_2_lut (.I0(byte_transmit_counter[0]), .I1(byte_transmit_counter[1]), 
            .I2(GND_net), .I3(GND_net), .O(n109));   // verilog/coms.v(103[12:33])
    defparam i1_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i2_4_lut (.I0(byte_transmit_counter[3]), .I1(n109), .I2(byte_transmit_counter[4]), 
            .I3(byte_transmit_counter[2]), .O(n55301));   // verilog/coms.v(103[12:33])
    defparam i2_4_lut.LUT_INIT = 16'ha080;
    SB_LUT4 i3_4_lut (.I0(byte_transmit_counter[5]), .I1(byte_transmit_counter[6]), 
            .I2(byte_transmit_counter[7]), .I3(n55301), .O(n44));
    defparam i3_4_lut.LUT_INIT = 16'hfffe;
    SB_DFFE r_Bit_Index_i0 (.Q(\r_Bit_Index[0] ), .C(clk16MHz), .E(VCC_net), 
            .D(n26829));   // verilog/uart_tx.v(41[10] 144[8])
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_48723 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[14][5] ), .I2(\data_out_frame[15][5] ), 
            .I3(byte_transmit_counter[1]), .O(n63413));
    defparam byte_transmit_counter_0__bdd_4_lut_48723.LUT_INIT = 16'he4aa;
    SB_LUT4 n63413_bdd_4_lut (.I0(n63413), .I1(\data_out_frame[13][5] ), 
            .I2(\data_out_frame[12][5] ), .I3(byte_transmit_counter[1]), 
            .O(n63416));
    defparam n63413_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFFSR r_SM_Main_i1 (.Q(r_SM_Main[1]), .C(clk16MHz), .D(n3_adj_5049), 
            .R(r_SM_Main[2]));   // verilog/uart_tx.v(41[10] 144[8])
    SB_DFFE r_Tx_Data_i7 (.Q(r_Tx_Data[7]), .C(clk16MHz), .E(n21898), 
            .D(tx_data[7]));   // verilog/uart_tx.v(41[10] 144[8])
    SB_DFFE r_Tx_Data_i6 (.Q(r_Tx_Data[6]), .C(clk16MHz), .E(n21898), 
            .D(tx_data[6]));   // verilog/uart_tx.v(41[10] 144[8])
    SB_DFFE r_Tx_Data_i5 (.Q(r_Tx_Data[5]), .C(clk16MHz), .E(n21898), 
            .D(tx_data_c[5]));   // verilog/uart_tx.v(41[10] 144[8])
    SB_DFFE r_Tx_Data_i4 (.Q(r_Tx_Data[4]), .C(clk16MHz), .E(n21898), 
            .D(\tx_data[4] ));   // verilog/uart_tx.v(41[10] 144[8])
    SB_DFFE r_Tx_Data_i3 (.Q(r_Tx_Data[3]), .C(clk16MHz), .E(n21898), 
            .D(\tx_data[3] ));   // verilog/uart_tx.v(41[10] 144[8])
    SB_DFFE r_Tx_Data_i2 (.Q(r_Tx_Data[2]), .C(clk16MHz), .E(n21898), 
            .D(\tx_data[2] ));   // verilog/uart_tx.v(41[10] 144[8])
    SB_DFFE r_Tx_Data_i1 (.Q(r_Tx_Data[1]), .C(clk16MHz), .E(n21898), 
            .D(\tx_data[1] ));   // verilog/uart_tx.v(41[10] 144[8])
    SB_DFF r_Tx_Active_53 (.Q(tx_active), .C(clk16MHz), .D(n48965));   // verilog/uart_tx.v(41[10] 144[8])
    SB_DFF r_SM_Main_i2 (.Q(r_SM_Main[2]), .C(clk16MHz), .D(n63731));   // verilog/uart_tx.v(41[10] 144[8])
    SB_LUT4 i46163_3_lut (.I0(n38), .I1(\o_Rx_DV_N_3261[12] ), .I2(n4837), 
            .I3(GND_net), .O(n59798));   // verilog/uart_tx.v(32[16:25])
    defparam i46163_3_lut.LUT_INIT = 16'h0202;
    SB_LUT4 i46158_4_lut (.I0(n59798), .I1(\o_Rx_DV_N_3261[24] ), .I2(n29), 
            .I3(n23), .O(n59795));   // verilog/uart_tx.v(32[16:25])
    defparam i46158_4_lut.LUT_INIT = 16'h0002;
    SB_LUT4 i7_4_lut (.I0(\r_SM_Main_2__N_3318[0] ), .I1(n59795), .I2(r_SM_Main[1]), 
            .I3(n27), .O(n3_adj_5050));   // verilog/uart_tx.v(32[16:25])
    defparam i7_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i8_3_lut (.I0(n3_adj_5050), .I1(n36763), .I2(r_SM_Main[0]), 
            .I3(GND_net), .O(n19213));   // verilog/uart_tx.v(32[16:25])
    defparam i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i23278_3_lut (.I0(r_SM_Main[0]), .I1(n63362), .I2(r_SM_Main[1]), 
            .I3(GND_net), .O(n3));   // verilog/uart_tx.v(32[16:25])
    defparam i23278_3_lut.LUT_INIT = 16'he5e5;
    SB_LUT4 i42124_3_lut (.I0(r_Tx_Data[0]), .I1(r_Tx_Data[1]), .I2(\r_Bit_Index[0] ), 
            .I3(GND_net), .O(n56836));
    defparam i42124_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i42125_3_lut (.I0(r_Tx_Data[2]), .I1(r_Tx_Data[3]), .I2(\r_Bit_Index[0] ), 
            .I3(GND_net), .O(n56837));
    defparam i42125_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i42128_3_lut (.I0(r_Tx_Data[6]), .I1(r_Tx_Data[7]), .I2(\r_Bit_Index[0] ), 
            .I3(GND_net), .O(n56840));
    defparam i42128_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i42127_3_lut (.I0(r_Tx_Data[4]), .I1(r_Tx_Data[5]), .I2(\r_Bit_Index[0] ), 
            .I3(GND_net), .O(n56839));
    defparam i42127_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i5_3_lut (.I0(r_SM_Main[0]), .I1(\o_Rx_DV_N_3261[24] ), .I2(n27), 
            .I3(GND_net), .O(n14));
    defparam i5_3_lut.LUT_INIT = 16'h0202;
    SB_LUT4 i6_4_lut (.I0(n29), .I1(\o_Rx_DV_N_3261[12] ), .I2(n23), .I3(n4837), 
            .O(n15));
    defparam i6_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 i8_4_lut (.I0(n15), .I1(n1), .I2(n14), .I3(r_SM_Main[1]), 
            .O(n63731));
    defparam i8_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i12_4_lut (.I0(tx_active), .I1(r_SM_Main[1]), .I2(n55736), 
            .I3(n36774), .O(n48965));   // verilog/uart_tx.v(32[16:25])
    defparam i12_4_lut.LUT_INIT = 16'h3aba;
    SB_LUT4 i46058_3_lut (.I0(r_Bit_Index[2]), .I1(r_Bit_Index[1]), .I2(\r_Bit_Index[0] ), 
            .I3(GND_net), .O(n460[2]));
    defparam i46058_3_lut.LUT_INIT = 16'h6a6a;
    SB_LUT4 i1_3_lut_4_lut_4_lut (.I0(r_SM_Main[0]), .I1(\r_SM_Main_2__N_3318[0] ), 
            .I2(r_SM_Main[1]), .I3(r_SM_Main[2]), .O(n55736));   // verilog/uart_tx.v(41[10] 144[8])
    defparam i1_3_lut_4_lut_4_lut.LUT_INIT = 16'h00f4;
    SB_LUT4 i2_3_lut_4_lut_4_lut (.I0(r_SM_Main[0]), .I1(\r_SM_Main_2__N_3318[0] ), 
            .I2(r_SM_Main[1]), .I3(r_SM_Main[2]), .O(n21898));   // verilog/uart_tx.v(41[10] 144[8])
    defparam i2_3_lut_4_lut_4_lut.LUT_INIT = 16'h0004;
    SB_LUT4 i1_2_lut_3_lut (.I0(\r_SM_Main_2__N_3318[0] ), .I1(tx_active), 
            .I2(n44), .I3(GND_net), .O(n36757));
    defparam i1_2_lut_3_lut.LUT_INIT = 16'hefef;
    SB_LUT4 i48558_2_lut_3_lut_4_lut (.I0(r_SM_Main[2]), .I1(r_SM_Main[0]), 
            .I2(n36763), .I3(r_SM_Main[1]), .O(n24612));
    defparam i48558_2_lut_3_lut_4_lut.LUT_INIT = 16'h0111;
    SB_LUT4 i67_2_lut_4_lut (.I0(r_SM_Main[1]), .I1(\r_Bit_Index[0] ), .I2(r_Bit_Index[1]), 
            .I3(r_Bit_Index[2]), .O(n47));   // verilog/uart_tx.v(32[16:25])
    defparam i67_2_lut_4_lut.LUT_INIT = 16'hd555;
    SB_LUT4 i48419_2_lut_3_lut (.I0(\r_SM_Main_2__N_3318[0] ), .I1(tx_active), 
            .I2(n44), .I3(GND_net), .O(tx_transmit_N_3189));
    defparam i48419_2_lut_3_lut.LUT_INIT = 16'h0101;
    SB_LUT4 i2_3_lut (.I0(\r_Bit_Index[0] ), .I1(r_Bit_Index[1]), .I2(r_Bit_Index[2]), 
            .I3(GND_net), .O(n38));   // verilog/uart_tx.v(41[10] 144[8])
    defparam i2_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 i38969_rep_5_2_lut (.I0(n36763), .I1(r_SM_Main[1]), .I2(GND_net), 
            .I3(GND_net), .O(n53849));
    defparam i38969_rep_5_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 r_Bit_Index_1__bdd_4_lut (.I0(r_Bit_Index[1]), .I1(n56839), 
            .I2(n56840), .I3(r_Bit_Index[2]), .O(n63359));
    defparam r_Bit_Index_1__bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_LUT4 n63359_bdd_4_lut (.I0(n63359), .I1(n56837), .I2(n56836), .I3(r_Bit_Index[2]), 
            .O(n63362));
    defparam n63359_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i45676_4_lut (.I0(\data_out_frame[16][5] ), .I1(byte_transmit_counter[1]), 
            .I2(\data_out_frame[17][5] ), .I3(byte_transmit_counter[0]), 
            .O(n59753));
    defparam i45676_4_lut.LUT_INIT = 16'h3022;
    SB_LUT4 i42292_4_lut (.I0(n24853), .I1(n59753), .I2(byte_transmit_counter[4]), 
            .I3(\data_out_frame[1][5] ), .O(n57004));
    defparam i42292_4_lut.LUT_INIT = 16'hc5c0;
    SB_LUT4 i42290_3_lut (.I0(n63416), .I1(n33453), .I2(byte_transmit_counter[4]), 
            .I3(GND_net), .O(n57002));
    defparam i42290_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i42293_3_lut (.I0(n56920), .I1(n57004), .I2(byte_transmit_counter[3]), 
            .I3(GND_net), .O(n57005));
    defparam i42293_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i42291_3_lut (.I0(n63350), .I1(n57002), .I2(byte_transmit_counter[3]), 
            .I3(GND_net), .O(n57003));
    defparam i42291_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i42294_3_lut (.I0(n56922), .I1(n57005), .I2(n57324), .I3(GND_net), 
            .O(n57006));
    defparam i42294_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i2230099_i1_3_lut (.I0(n57006), .I1(n57003), .I2(byte_transmit_counter[2]), 
            .I3(GND_net), .O(tx_data_c[5]));
    defparam i2230099_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_3_lut_4_lut (.I0(r_SM_Main[2]), .I1(r_SM_Main[0]), .I2(n53849), 
            .I3(n47), .O(n36762));
    defparam i1_3_lut_4_lut.LUT_INIT = 16'h0100;
    SB_LUT4 i1_4_lut (.I0(n23), .I1(\o_Rx_DV_N_3261[12] ), .I2(n4837), 
            .I3(r_SM_Main[0]), .O(n55742));
    defparam i1_4_lut.LUT_INIT = 16'h0100;
    SB_LUT4 i1_4_lut_adj_1043 (.I0(\o_Rx_DV_N_3261[24] ), .I1(n27), .I2(n29), 
            .I3(n55742), .O(n36774));
    defparam i1_4_lut_adj_1043.LUT_INIT = 16'h0100;
    SB_LUT4 i17_2_lut (.I0(n36774), .I1(r_SM_Main[1]), .I2(GND_net), .I3(GND_net), 
            .O(n3_adj_5049));   // verilog/uart_tx.v(32[16:25])
    defparam i17_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i20_2_lut (.I0(r_Bit_Index[1]), .I1(\r_Bit_Index[0] ), .I2(GND_net), 
            .I3(GND_net), .O(n460[1]));   // verilog/uart_tx.v(34[16:27])
    defparam i20_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut (.I0(byte_transmit_counter[1]), 
            .I1(n59726), .I2(n59727), .I3(byte_transmit_counter[4]), .O(n63347));
    defparam byte_transmit_counter_1__bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_LUT4 n63347_bdd_4_lut (.I0(n63347), .I1(n56924), .I2(n56923), .I3(byte_transmit_counter[4]), 
            .O(n63350));
    defparam n63347_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 o_Tx_Serial_I_0_1_lut (.I0(tx_o), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(tx_enable));   // verilog/uart_tx.v(39[24:36])
    defparam o_Tx_Serial_I_0_1_lut.LUT_INIT = 16'h5555;
    
endmodule
//
// Verilog Description of module uart_rx
//

module uart_rx (baudrate, n24621, clk16MHz, n53789, GND_net, r_Clock_Count, 
            VCC_net, n26516, rx_data, \r_SM_Main[2] , r_Rx_Data, RX_N_42, 
            \o_Rx_DV_N_3261[24] , n27, n29, \r_Bit_Index[0] , n55980, 
            n23, n55948, \o_Rx_DV_N_3261[12] , n26445, \o_Rx_DV_N_3261[8] , 
            n26443, \o_Rx_DV_N_3261[7] , \o_Rx_DV_N_3261[6] , \o_Rx_DV_N_3261[5] , 
            n33, \o_Rx_DV_N_3261[4] , \o_Rx_DV_N_3261[3] , \o_Rx_DV_N_3261[2] , 
            \o_Rx_DV_N_3261[1] , \o_Rx_DV_N_3261[0] , n27051, n26970, 
            n4834, n52823, n26836, n48959, rx_data_ready, n26832, 
            n55964, n55996, \r_SM_Main[1] , \r_SM_Main_2__N_3219[1] , 
            n55461, n26587, n26062, n55884, n55900, n55916, n55932, 
            n55814, n24535, n34) /* synthesis syn_module_defined=1 */ ;
    input [31:0]baudrate;
    output n24621;
    input clk16MHz;
    output n53789;
    input GND_net;
    output [7:0]r_Clock_Count;
    input VCC_net;
    input n26516;
    output [7:0]rx_data;
    output \r_SM_Main[2] ;
    output r_Rx_Data;
    input RX_N_42;
    output \o_Rx_DV_N_3261[24] ;
    output n27;
    output n29;
    output \r_Bit_Index[0] ;
    output n55980;
    output n23;
    output n55948;
    output \o_Rx_DV_N_3261[12] ;
    input n26445;
    output \o_Rx_DV_N_3261[8] ;
    input n26443;
    output \o_Rx_DV_N_3261[7] ;
    output \o_Rx_DV_N_3261[6] ;
    output \o_Rx_DV_N_3261[5] ;
    output n33;
    output \o_Rx_DV_N_3261[4] ;
    output \o_Rx_DV_N_3261[3] ;
    output \o_Rx_DV_N_3261[2] ;
    output \o_Rx_DV_N_3261[1] ;
    output \o_Rx_DV_N_3261[0] ;
    input n27051;
    input n26970;
    input n4834;
    input n52823;
    input n26836;
    input n48959;
    output rx_data_ready;
    input n26832;
    output n55964;
    output n55996;
    output \r_SM_Main[1] ;
    input \r_SM_Main_2__N_3219[1] ;
    output n55461;
    input n26587;
    input n26062;
    output n55884;
    output n55900;
    output n55916;
    output n55932;
    input n55814;
    output n24535;
    output n34;
    
    wire clk16MHz /* synthesis SET_AS_NETWORK=clk16MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(31[6:14])
    
    wire n3169;
    wire [23:0]n7806;
    wire [23:0]n294;
    
    wire n11;
    wire [2:0]n479;
    wire [2:0]r_Bit_Index;   // verilog/uart_rx.v(34[17:28])
    
    wire n46444, n2832, n2519, n46445, n2599;
    wire [23:0]n7676;
    
    wire n2716, n3168, n13, n3167, n15, n1412;
    wire [23:0]n7442;
    
    wire n1556;
    wire [7:0]n1;
    
    wire n24619, n25950;
    wire [23:0]n7468;
    
    wire n1697, n3161, n27_c, n60335, n33_c, n12;
    wire [23:0]n7494;
    
    wire n1835, n60313;
    wire [23:0]n7728;
    
    wire n2833, n2397, n46443, n10, n35, n30, n21, n19, n17, 
        n9, n60359, n43, n16, n60218, n2834, n2272, n46442, 
        n8, n2835, n2144, n46441, n2836, n2013, n46440, n2837, 
        n1879, n46439, n45_adj_4766, n24, n3172, n3274, n2838, 
        n1742, n46438, n2839, n1602, n46437, n7, n60425, n2840, 
        n1459, n46436, n61377, n2841, n1460, n46435, n2842, n1011, 
        n46434, n2843, n856, n46433, n2844, n698, n46432, n2845, 
        n858, n46431, n55690, n538, n53871;
    wire [23:0]n7702;
    
    wire n2713, n2977, n46430, n2714, n2867, n46429, n61359, n2715, 
        n2754, n46428, n25, n23_c, n62621, n2638, n46427, n31, 
        n29_c, n61927, n2717, n46426, n37, n62792, n2718, n46425, 
        n2719, n46424, n6, n62629, n2720, n46423, n62630, n2721, 
        n46422, n2722, n46421, n2723, n46420, n2724, n46419, n55696, 
        n48, n4, n2725, n46418, n2726, n46417, n62396, n2727, 
        n46416, n2728, n46415, n2729, n46414, n2730, n46413, n55688, 
        n53875, n2596, n46412, n62397, n60321, n2597, n46411, 
        n2598, n46410, n46409, n2600, n46408;
    wire [23:0]n7520;
    
    wire n1970, n2601, n46407, n2602, n46406, n2603, n46405, n2604, 
        n46404, n2605, n46403, n2606, n46402, n2607, n46401, n62851, 
        n804, n42, n960, n62351, n62991, n62992;
    wire [23:0]n7546;
    
    wire n2102, n39, n62970;
    wire [23:0]n7572;
    
    wire n2231, n60230, n61948, n2608, n46400, n62349, n41, n60256, 
        n2609, n46399, n62635, n40, n2610, n46398, n3151, n3253, 
        n62637, n56554, n56484, n56430, n56356, n55652, n54733, 
        n2611, n46397;
    wire [23:0]n7598;
    
    wire n2357, n2612, n46396;
    wire [23:0]n7624;
    
    wire n2480, n55686, n53879;
    wire [23:0]n7650;
    
    wire n2476, n46395, n2477, n46394, n3046;
    wire [23:0]n7780;
    
    wire n3049, n3154, n3047, n3152, n3048, n3153, n3050, n3155, 
        n3053, n3158, n33_adj_4768, n3051, n3156, n37_adj_4769, 
        n3052, n3157, n35_adj_4770, n3054, n3159, n31_adj_4771, 
        n3056, n3057, n3162, n25_adj_4772, n27_adj_4773, n3058, 
        n3163, n3059, n3164, n2478, n46393, n22504, n48_adj_4774, 
        n35471, n54412, n21_adj_4775, n23_adj_4776, n3065, n3170, 
        n3066, n3171, n9_adj_4777, n3060, n3165, n3064, n11_adj_4778, 
        n19_adj_4779, n3062, n3055, n3160, n3061, n3166, n3063, 
        n13_adj_4781, n15_adj_4782, n17_adj_4783, n29_adj_4784, n56556, 
        n56558, n644, n44, n46, n42_adj_4787, n1113, n53644, n53646;
    wire [23:0]n7390;
    
    wire n1263, n56560, n22434, n1264, n41_adj_4790, n60473, n61469, 
        n62008, n62002, n60481, n6_adj_4791, n62178, n14, n32, 
        n62179, n60467, n12_adj_4792, n60463, n62721, n61334, n8_adj_4793, 
        n62180, n2479, n46392, n62181, n60503, n61447, n10_adj_4794, 
        n61944, n61332, n62386, n62916, n62398, n62997, n62998, 
        n62850, n62761, n62762, n2938;
    wire [23:0]n7754;
    
    wire n2946, n2941, n2939, n2940, n2944, n35_adj_4795, n2942, 
        n39_adj_4796, n2945, n33_adj_4797, n2943, n37_adj_4798, n2947, 
        n2948, n46391, n27_adj_4799, n29_adj_4800, n2949, n39_adj_4801, 
        n2950, n2481, n46390, n2482, n46389, n2483, n46388, n23_adj_4802, 
        n25_adj_4803, n803, n9112, n18960, n46_adj_4804, n2956, 
        n2484, n46387, n2957, n11_adj_4805, n2951, n2955, n2485, 
        n46386, n13_adj_4806, n21_adj_4807, n3;
    wire [2:0]r_SM_Main;   // verilog/uart_rx.v(37[17:26])
    
    wire n2952, n2953, n2486, n46385, n2487, n46384, n2954, r_Rx_Data_R, 
        n41_adj_4808, n43_adj_4809, n15_adj_4810, n17_adj_4811, n19_adj_4812, 
        n31_adj_4813, n60563, n2488, n46383, n2489, n46382, n61543, 
        n62038, n62034, n60567, n8_adj_4814, n1409, n1553, n62186, 
        n62187, n2490, n46381, n16_adj_4815, n34_c, n60547, n46149, 
        n46148, n55658, n14_adj_4817, n60539, n62697, n1267, n36, 
        n61322, n10_adj_4818, n62188, n2491, n46380, n62189, n60579, 
        n61521, n12_adj_4819, n20, n61320, n55684, n53883, n2353, 
        n46379, n1694, n62428, n62914, n61942, n62993, n1832, 
        n53648, n1967, n62994, n2099, n2228, n62400, n56822, n46147, 
        n55708, n62401, n4_adj_4821, n2354, n46378, n38_adj_4822, 
        n40_adj_4823, n46146;
    wire [24:0]o_Rx_DV_N_3261;
    
    wire n2355, n46377, n2356, n46376, n2827, n46375, n46145, 
        n55706, n2358, n46374, n959, n9283, n19010, n46_adj_4825, 
        n1111, n1261, n2359, n46373, n2828;
    wire [23:0]n7416;
    
    wire n1408, n2829, n2360, n46372, n37_adj_4826, n1552, n2830, 
        n2361, n46371, n41_adj_4827, n60459, n62591, n46144, n55704, 
        n1693, n35_adj_4828, n22501, n2362, n46370, n2831, n39_adj_4829, 
        n29_adj_4830, n31_adj_4831, n23_adj_4832, n25_adj_4833, n27_adj_4834, 
        n13_adj_4835, n15_adj_4836, n17_adj_4837, n2363, n46369, n46143, 
        n2364, n46368, n19_adj_4838, n2365, n46367, n21_adj_4839, 
        n33_adj_4840, n46142, n55702, n2366, n46366, n46141, n55700, 
        n2367, n46365, n55682, n53887, n2227, n46364, n56428, 
        n46140, n55656, n46363, n2229, n46362, n56488, n2230, 
        n46361, n56486, n56490, n56354, n22476, n46139, n55698, 
        n60640, n61635, n62084, n62080, n60646, n10_adj_4841, n62192, 
        n62193, n18, n36_adj_4842, n1831, n46360, n2232, n46359, 
        n60626, n16_adj_4843, n60618, n62659, n2233, n46358, n2234, 
        n46357, n62592, n61308, n1966, n2235, n46356, n2236, n46355, 
        n14_adj_4844, n22, n12_adj_4845, n60675, n62655, n46138, 
        n62656, n2237, n46354, n62528, n62461, n62910, n2238, 
        n46353, n2239, n46352, n61306, n2240, n46351, n63011, 
        n63012, n55680, n53891, n63004, n37_adj_4846, n43_adj_4847, 
        n1262, n62568, n41_adj_4848, n2098, n39_adj_4849, n39_adj_4850, 
        n37_adj_4851, n43_adj_4852, n31_adj_4853, n41_adj_4854, n33_adj_4855, 
        n31_adj_4856, n35_adj_4857, n45_adj_4858, n33_adj_4859, n46137, 
        n25_adj_4860, n27_adj_4861, n29_adj_4862, n27_adj_4863, n25_adj_4864, 
        n46350, n29_adj_4865, n15_adj_4866, n46349, n2100, n46348, 
        n21_adj_4867, n27_adj_4868, n25_adj_4869, n23_adj_4870, n60116, 
        n2101, n46347, n19_adj_4871, n46346, n46136, n33_adj_4872, 
        n31_adj_4873, n29_adj_4874, n60091, n2103, n46345, n1415, 
        n1559, n46645, n1700, n46135, n2104, n46344, n46644, n17_adj_4875, 
        n21_adj_4876, n19_adj_4877, n21_adj_4878, n23_adj_4879, n2105, 
        n46343, n46134, n46643, n35_adj_4880, n60730, n61711, n1838, 
        n62120, n46642, n2106, n46342, n23_adj_4881, n2107, n46341, 
        n46641, n62116, n46133, n63689, n60736, n962, n40_adj_4882, 
        n12_adj_4883, n62198, n17_adj_4884, n20_adj_4885, n59971, 
        n59959, n20_adj_4886, n38_adj_4887, n62199, n60714, n62164, 
        n18_adj_4888, n60712, n62763, n46640, n46132, n61300, n46639, 
        n2108, n46340, n1973, n16_adj_4889, n16_adj_4890, n24_adj_4891, 
        n2109, n46339, n2110, n26, n28, n14_adj_4892, n60755, 
        n62651, n62652, n62532, n62477, n24_adj_4893, n35_adj_4894, 
        n32_adj_4895, n22_adj_4896, n60085, n62842, n46338, n46337, 
        n1968, n46336, n46131, n1969, n46335, n62888, n46334, 
        n46130, n1971, n46333, n37_adj_4897, n62843, n39_adj_4898, 
        n62774, n62194, n61298, n62999, n63000, n60109, n62844, 
        n961, n1114, n805, n22_adj_4899, n23_adj_4900, n56292, n56264, 
        n56274, n56376, n56456, n24_adj_4901, n59864, n46_adj_4903, 
        n48_adj_4904, n31_adj_4905, n56416, n22484, n35469, n62224, 
        n62225, n59963, n61785, n22_adj_4906, n62334, n61282, n20_adj_4907, 
        n28_adj_4908, n18_adj_4909, n59955, n62848, n62849, n62766, 
        n60931, n62541, n36_adj_4910, n62743, n62744, n39_adj_4911, 
        n45_adj_4912, n43_adj_4913, n41_adj_4914, n33_adj_4915, n35_adj_4916, 
        n37_adj_4917, n27_adj_4918, n29_adj_4919, n31_adj_4920, n21_adj_4921, 
        n1972, n46332, n46331, n46129, n1974, n46330, n1975, n46329, 
        n46128, n1976, n46328, n1977, n46327, n46127, n46326, 
        n46325, n1833, n46324, n19008, n23_adj_4922, n46126, n1834, 
        n46323, n46322, n1836, n46321, n1837, n46320, n46319, 
        n1839, n46318, n1840, n46317, n25_adj_4923, n1841, n46316, 
        n55678, n53900, n46315, n46314, n1695, n46313, n1696, 
        n46312, n41_adj_4924, n62612, n46311, n1698, n46310, n1699, 
        n46309, n46308, n19_adj_4925, n62904, n60028, n60012, n62174, 
        n1701, n46307, n18_adj_4926, n1702, n62406, n62407, n60021, 
        n60979, n46306, n33_adj_4927, n24_adj_4928, n26_adj_4929, 
        n56818, n54397, n42_adj_4930, n46305, n1554, n46304, n1555, 
        n46303, n14_adj_4931, n15_adj_4932, n56176, n56710, n56184, 
        n46302, n22_adj_4933, n30_adj_4934, n1557, n46301, n20_adj_4935, 
        n60008, n62846, n1558, n46300, n56792, n46299, n1560, 
        n46298, n62847, n46297, n62768, n60983, n46296, n61935, 
        n62620, n61937, n1410, n46295, n1411, n46294, n62905, 
        n62868, n56182, n22498, n56180, n17_adj_4936, n19_adj_4937, 
        n27_adj_4938, n56470, n56156, n56308, n37_adj_4939, n25_adj_4940, 
        n23_adj_4941, n21_adj_4942, n60817, n61767, n62148, n46293, 
        n31_adj_4943, n29_adj_4944, n62144, n35_adj_4945, n60819, 
        n60180, n14_adj_4946, n62204, n62205, n42_adj_4947, n62254, 
        n62255, n56786, n1413, n46292, n1414, n46291, n46290, 
        n55676, n53909, n48_adj_4948, n56814, n1115, n1265, n3_adj_4949, 
        n43_adj_4950, n41_adj_4951, n46289, n46288, n46287, n46286, 
        n39_adj_4952, n37_adj_4953, n33_adj_4954, n46285, n35_adj_4955, 
        n56208, n56206, n56464, n22385, n25_adj_4956, n27_adj_4957, 
        n29_adj_4958, n1266, n46284, n31_adj_4959, n23_adj_4960, n60195, 
        n60172, n46283, n22_adj_4961, n28_adj_4962, n30_adj_4963, 
        n55674, n53913, n46282, n1112, n46281, n26_adj_4964, n34_adj_4965, 
        n24_adj_4966, n60166, n62808, n62809, n62778, n62244, n60187, 
        n62414, n42_adj_4967, n56458, n62675, n56474, n56472, n22473, 
        n62676, n46280, n46279, n46278, n37_adj_4968, n35_adj_4969, 
        n1116, n46277, n41_adj_4970, n39_adj_4971, n29_adj_4972, n55672, 
        n53917, n31_adj_4973, n43_adj_4974, n33_adj_4975, n27_adj_4976, 
        n60262, n56346, n56762, n38_adj_4977, n40_adj_4978, n42_adj_4979, 
        n30_adj_4980, n38_adj_4981, n53894, n60469, n62785, n62786, 
        n26_adj_4982, n62420, n62421, n60233, n28_adj_4983, n60227, 
        n62806, n62313, n62971, n62972, n62891, n48_adj_4984, n56410, 
        n56418, n22464, n6_adj_4985, n56242, n56344, n56118, n48_adj_4986, 
        n56382, n3186, n46513, n3082, n46512, n3188, n46511, n3084, 
        n46510, n46509, n46508, n46507, n46506, n25_adj_4987, n46505, 
        n46504, n46503, n46502, n46501, n46500, n46499, n46498, 
        n46497, n46496, n46495, n46494, n46493, n46492, n46491, 
        n53859, n46490, n46489, n46488, n46487, n46486, n46485, 
        n46484, n46483, n46482, n46481, n46480, n46479, n46478, 
        n46477, n46476, n46475, n46474, n46473, n46472, n46471, 
        n46470, n55694, n53863, n46469, n56358, n46468, n46467, 
        n46466, n46465, n46464, n56452, n56772, n46463, n46462, 
        n46461, n46460, n46459, n46458, n46457, n56774, n46456, 
        n46455, n46454, n46453, n48_adj_4988, n46452, n46451, n46450, 
        n55692, n53867, n46449, n46448, n46447, n46446, n37_adj_4989, 
        n35_adj_4990, n41_adj_4991, n43_adj_4992, n29_adj_4993, n39_adj_4994, 
        n31_adj_4995, n33_adj_4996, n39_adj_4997, n56388, n27_adj_4998, 
        n60328, n30_adj_4999, n38_adj_5000, n26_adj_5001, n62424, 
        n62425, n56318, n22481, n53920, n60317, n42_adj_5002, n28_adj_5003, 
        n60315, n62869, n62309, n22444, n62292, n22_adj_5004, n40_adj_5005, 
        n62293, n48_adj_5006, n60805, n62967, n22507, n62968, n62895, 
        n37_adj_5007, n48_adj_5008, n22470, n20_adj_5009, n60792, 
        n62338, n41_adj_5010, n60170, n53903, n32_adj_5011, n62228, 
        n62229, n61292, n60410, n61373, n34_adj_5012, n62304, n39_adj_5013, 
        n61271, n43_adj_5014, n37_adj_5015, n62545, n31_adj_5016, 
        n35_adj_5017, n62546, n52650, n56700, n33_adj_5018, n41_adj_5019, 
        n56780, n2, n9473, n29_adj_5020, n60364, n41_adj_5021, n43_adj_5022, 
        n39_adj_5023, n41_adj_5024, n37_adj_5025, n43_adj_5026, n56160, 
        n18896, n48_adj_5027, n32_adj_5028, n40_adj_5029, n56386, 
        n28_adj_5030, n62226, n62227, n60349, n30_adj_5031, n60347, 
        n62426, n61274, n62804, n44_adj_5032, n62805, n22492, n44_adj_5033, 
        n9276, n35725, n56804, n45_adj_5034, n39_adj_5035, n56800, 
        n56802, n34_adj_5036, n16_adj_5037, n18_adj_5038, n26_adj_5039, 
        n62250, n60840, n62649, n62251, n62650, n60449, n61405, 
        n36_adj_5040, n38_adj_5041, n62534, n61264, n62491, n62298, 
        n59759, n59765, n59756, n59762, n62799, n62797, n61290, 
        n32_adj_5042, n62248, n56246, n3_adj_5043, n56250, n5, n62249, 
        n56254, n8_adj_5044, n59788, n59785, n60433, n61391, n59782, 
        n34_adj_5045, n62302, n55766, n61268, n62549, n55772, n62550, 
        n56738, n28_adj_5046, n59876, n59873, n56448, n56174, n56748, 
        n56080, n56768, n56766, n56764, n56098, n54439;
    
    SB_LUT4 div_37_LessThan_2210_i11_4_lut (.I0(n3169), .I1(baudrate[5]), 
            .I2(n7806[5]), .I3(n294[1]), .O(n11));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i11_4_lut.LUT_INIT = 16'h3c66;
    SB_DFFESR r_Bit_Index_i1 (.Q(r_Bit_Index[1]), .C(clk16MHz), .E(n24621), 
            .D(n479[1]), .R(n53789));   // verilog/uart_rx.v(50[10] 145[8])
    SB_DFFESR r_Bit_Index_i2 (.Q(r_Bit_Index[2]), .C(clk16MHz), .E(n24621), 
            .D(n479[2]), .R(n53789));   // verilog/uart_rx.v(50[10] 145[8])
    SB_CARRY add_2551_16 (.CI(n46444), .I0(n2832), .I1(n2519), .CO(n46445));
    SB_LUT4 div_37_i1825_3_lut (.I0(n2599), .I1(n7676[20]), .I2(n294[6]), 
            .I3(GND_net), .O(n2716));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1825_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_2210_i13_4_lut (.I0(n3168), .I1(baudrate[6]), 
            .I2(n7806[6]), .I3(n294[1]), .O(n13));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i13_4_lut.LUT_INIT = 16'h3c66;
    SB_LUT4 div_37_LessThan_2210_i15_4_lut (.I0(n3167), .I1(baudrate[7]), 
            .I2(n7806[7]), .I3(n294[1]), .O(n15));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i15_4_lut.LUT_INIT = 16'h3c66;
    SB_LUT4 div_37_i1043_3_lut (.I0(n1412), .I1(n7442[19]), .I2(n294[15]), 
            .I3(GND_net), .O(n1556));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1043_3_lut.LUT_INIT = 16'hcaca;
    SB_DFFESR r_Clock_Count_1948__i0 (.Q(r_Clock_Count[0]), .C(clk16MHz), 
            .E(n24619), .D(n1[0]), .R(n25950));   // verilog/uart_rx.v(121[34:51])
    SB_LUT4 div_37_i1138_3_lut (.I0(n1556), .I1(n7468[19]), .I2(n294[14]), 
            .I3(GND_net), .O(n1697));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1138_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_2210_i27_4_lut (.I0(n3161), .I1(baudrate[13]), 
            .I2(n7806[13]), .I3(n294[1]), .O(n27_c));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i27_4_lut.LUT_INIT = 16'h3c66;
    SB_LUT4 i45623_4_lut (.I0(n27_c), .I1(n15), .I2(n13), .I3(n11), 
            .O(n60335));
    defparam i45623_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 div_37_LessThan_2210_i12_3_lut (.I0(baudrate[7]), .I1(baudrate[16]), 
            .I2(n33_c), .I3(GND_net), .O(n12));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1231_3_lut (.I0(n1697), .I1(n7494[19]), .I2(n294[13]), 
            .I3(GND_net), .O(n1835));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1231_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i45601_2_lut (.I0(n33_c), .I1(n15), .I2(GND_net), .I3(GND_net), 
            .O(n60313));
    defparam i45601_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 add_2551_15_lut (.I0(GND_net), .I1(n2833), .I2(n2397), .I3(n46443), 
            .O(n7728[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2551_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_LessThan_2210_i10_3_lut (.I0(baudrate[5]), .I1(baudrate[6]), 
            .I2(n13), .I3(GND_net), .O(n10));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i10_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_2210_i30_3_lut (.I0(n12), .I1(baudrate[17]), 
            .I2(n35), .I3(GND_net), .O(n30));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i30_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_2551_15 (.CI(n46443), .I0(n2833), .I1(n2397), .CO(n46444));
    SB_LUT4 i45647_4_lut (.I0(n21), .I1(n19), .I2(n17), .I3(n9), .O(n60359));
    defparam i45647_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 div_37_LessThan_2210_i16_3_lut (.I0(baudrate[9]), .I1(baudrate[21]), 
            .I2(n43), .I3(GND_net), .O(n16));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i45506_2_lut (.I0(n43), .I1(n19), .I2(GND_net), .I3(GND_net), 
            .O(n60218));
    defparam i45506_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 add_2551_14_lut (.I0(GND_net), .I1(n2834), .I2(n2272), .I3(n46442), 
            .O(n7728[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2551_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2551_14 (.CI(n46442), .I0(n2834), .I1(n2272), .CO(n46443));
    SB_LUT4 div_37_LessThan_2210_i8_3_lut (.I0(baudrate[4]), .I1(baudrate[8]), 
            .I2(n17), .I3(GND_net), .O(n8));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_2551_13_lut (.I0(GND_net), .I1(n2835), .I2(n2144), .I3(n46441), 
            .O(n7728[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2551_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2551_13 (.CI(n46441), .I0(n2835), .I1(n2144), .CO(n46442));
    SB_LUT4 add_2551_12_lut (.I0(GND_net), .I1(n2836), .I2(n2013), .I3(n46440), 
            .O(n7728[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2551_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2551_12 (.CI(n46440), .I0(n2836), .I1(n2013), .CO(n46441));
    SB_LUT4 add_2551_11_lut (.I0(GND_net), .I1(n2837), .I2(n1879), .I3(n46439), 
            .O(n7728[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2551_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2551_11 (.CI(n46439), .I0(n2837), .I1(n1879), .CO(n46440));
    SB_LUT4 div_37_LessThan_2210_i24_3_lut (.I0(n16), .I1(baudrate[22]), 
            .I2(n45_adj_4766), .I3(GND_net), .O(n24));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i24_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2208_3_lut (.I0(n3172), .I1(n7806[2]), .I2(n294[1]), 
            .I3(GND_net), .O(n3274));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2208_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_2551_10_lut (.I0(GND_net), .I1(n2838), .I2(n1742), .I3(n46438), 
            .O(n7728[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2551_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2551_10 (.CI(n46438), .I0(n2838), .I1(n1742), .CO(n46439));
    SB_LUT4 add_2551_9_lut (.I0(GND_net), .I1(n2839), .I2(n1602), .I3(n46437), 
            .O(n7728[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2551_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2551_9 (.CI(n46437), .I0(n2839), .I1(n1602), .CO(n46438));
    SB_LUT4 i45713_3_lut (.I0(n7), .I1(n3274), .I2(baudrate[2]), .I3(GND_net), 
            .O(n60425));
    defparam i45713_3_lut.LUT_INIT = 16'hbebe;
    SB_LUT4 add_2551_8_lut (.I0(GND_net), .I1(n2840), .I2(n1459), .I3(n46436), 
            .O(n7728[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2551_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2551_8 (.CI(n46436), .I0(n2840), .I1(n1459), .CO(n46437));
    SB_LUT4 i46664_4_lut (.I0(n13), .I1(n11), .I2(n9), .I3(n60425), 
            .O(n61377));
    defparam i46664_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 add_2551_7_lut (.I0(GND_net), .I1(n2841), .I2(n1460), .I3(n46435), 
            .O(n7728[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2551_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2551_7 (.CI(n46435), .I0(n2841), .I1(n1460), .CO(n46436));
    SB_LUT4 add_2551_6_lut (.I0(GND_net), .I1(n2842), .I2(n1011), .I3(n46434), 
            .O(n7728[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2551_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2551_6 (.CI(n46434), .I0(n2842), .I1(n1011), .CO(n46435));
    SB_LUT4 add_2551_5_lut (.I0(GND_net), .I1(n2843), .I2(n856), .I3(n46433), 
            .O(n7728[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2551_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2551_5 (.CI(n46433), .I0(n2843), .I1(n856), .CO(n46434));
    SB_LUT4 add_2551_4_lut (.I0(GND_net), .I1(n2844), .I2(n698), .I3(n46432), 
            .O(n7728[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2551_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2551_4 (.CI(n46432), .I0(n2844), .I1(n698), .CO(n46433));
    SB_LUT4 add_2551_3_lut (.I0(GND_net), .I1(n2845), .I2(n858), .I3(n46431), 
            .O(n7728[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2551_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2551_3 (.CI(n46431), .I0(n2845), .I1(n858), .CO(n46432));
    SB_LUT4 add_2551_2_lut (.I0(n53871), .I1(GND_net), .I2(n538), .I3(VCC_net), 
            .O(n55690)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2551_2_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_2551_2 (.CI(VCC_net), .I0(GND_net), .I1(n538), .CO(n46431));
    SB_LUT4 add_2550_20_lut (.I0(GND_net), .I1(n2713), .I2(n2977), .I3(n46430), 
            .O(n7702[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2550_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2550_19_lut (.I0(GND_net), .I1(n2714), .I2(n2867), .I3(n46429), 
            .O(n7702[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2550_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2550_19 (.CI(n46429), .I0(n2714), .I1(n2867), .CO(n46430));
    SB_LUT4 i46646_4_lut (.I0(n19), .I1(n17), .I2(n15), .I3(n61377), 
            .O(n61359));
    defparam i46646_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 add_2550_18_lut (.I0(GND_net), .I1(n2715), .I2(n2754), .I3(n46428), 
            .O(n7702[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2550_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2550_18 (.CI(n46428), .I0(n2715), .I1(n2754), .CO(n46429));
    SB_LUT4 i47908_4_lut (.I0(n25), .I1(n23_c), .I2(n21), .I3(n61359), 
            .O(n62621));
    defparam i47908_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 add_2550_17_lut (.I0(GND_net), .I1(n2716), .I2(n2638), .I3(n46427), 
            .O(n7702[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2550_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2550_17 (.CI(n46427), .I0(n2716), .I1(n2638), .CO(n46428));
    SB_LUT4 i47214_4_lut (.I0(n31), .I1(n29_c), .I2(n27_c), .I3(n62621), 
            .O(n61927));
    defparam i47214_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 add_2550_16_lut (.I0(GND_net), .I1(n2717), .I2(n2519), .I3(n46426), 
            .O(n7702[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2550_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2550_16 (.CI(n46426), .I0(n2717), .I1(n2519), .CO(n46427));
    SB_LUT4 i48079_4_lut (.I0(n37), .I1(n35), .I2(n33_c), .I3(n61927), 
            .O(n62792));
    defparam i48079_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 add_2550_15_lut (.I0(GND_net), .I1(n2718), .I2(n2397), .I3(n46425), 
            .O(n7702[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2550_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2550_15 (.CI(n46425), .I0(n2718), .I1(n2397), .CO(n46426));
    SB_LUT4 add_2550_14_lut (.I0(GND_net), .I1(n2719), .I2(n2272), .I3(n46424), 
            .O(n7702[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2550_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2550_14 (.CI(n46424), .I0(n2719), .I1(n2272), .CO(n46425));
    SB_LUT4 div_37_LessThan_2210_i6_3_lut (.I0(baudrate[2]), .I1(baudrate[3]), 
            .I2(n7), .I3(GND_net), .O(n6));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i6_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i47916_3_lut (.I0(n6), .I1(baudrate[10]), .I2(n21), .I3(GND_net), 
            .O(n62629));   // verilog/uart_rx.v(119[33:55])
    defparam i47916_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_2550_13_lut (.I0(GND_net), .I1(n2720), .I2(n2144), .I3(n46423), 
            .O(n7702[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2550_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2550_13 (.CI(n46423), .I0(n2720), .I1(n2144), .CO(n46424));
    SB_LUT4 i47917_3_lut (.I0(n62629), .I1(baudrate[11]), .I2(n23_c), 
            .I3(GND_net), .O(n62630));   // verilog/uart_rx.v(119[33:55])
    defparam i47917_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_2550_12_lut (.I0(GND_net), .I1(n2721), .I2(n2013), .I3(n46422), 
            .O(n7702[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2550_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2550_12 (.CI(n46422), .I0(n2721), .I1(n2013), .CO(n46423));
    SB_LUT4 add_2550_11_lut (.I0(GND_net), .I1(n2722), .I2(n1879), .I3(n46421), 
            .O(n7702[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2550_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2550_11 (.CI(n46421), .I0(n2722), .I1(n1879), .CO(n46422));
    SB_LUT4 add_2550_10_lut (.I0(GND_net), .I1(n2723), .I2(n1742), .I3(n46420), 
            .O(n7702[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2550_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2550_10 (.CI(n46420), .I0(n2723), .I1(n1742), .CO(n46421));
    SB_LUT4 add_2550_9_lut (.I0(GND_net), .I1(n2724), .I2(n1602), .I3(n46419), 
            .O(n7702[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2550_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_LessThan_2210_i4_4_lut (.I0(baudrate[0]), .I1(baudrate[1]), 
            .I2(n55696), .I3(n48), .O(n4));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i4_4_lut.LUT_INIT = 16'hee8e;
    SB_CARRY add_2550_9 (.CI(n46419), .I0(n2724), .I1(n1602), .CO(n46420));
    SB_LUT4 add_2550_8_lut (.I0(GND_net), .I1(n2725), .I2(n1459), .I3(n46418), 
            .O(n7702[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2550_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2550_8 (.CI(n46418), .I0(n2725), .I1(n1459), .CO(n46419));
    SB_LUT4 add_2550_7_lut (.I0(GND_net), .I1(n2726), .I2(n1460), .I3(n46417), 
            .O(n7702[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2550_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i47683_3_lut (.I0(n4), .I1(baudrate[13]), .I2(n27_c), .I3(GND_net), 
            .O(n62396));   // verilog/uart_rx.v(119[33:55])
    defparam i47683_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_2550_7 (.CI(n46417), .I0(n2726), .I1(n1460), .CO(n46418));
    SB_LUT4 add_2550_6_lut (.I0(GND_net), .I1(n2727), .I2(n1011), .I3(n46416), 
            .O(n7702[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2550_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2550_6 (.CI(n46416), .I0(n2727), .I1(n1011), .CO(n46417));
    SB_LUT4 add_2550_5_lut (.I0(GND_net), .I1(n2728), .I2(n856), .I3(n46415), 
            .O(n7702[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2550_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2550_5 (.CI(n46415), .I0(n2728), .I1(n856), .CO(n46416));
    SB_LUT4 add_2550_4_lut (.I0(GND_net), .I1(n2729), .I2(n698), .I3(n46414), 
            .O(n7702[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2550_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2550_4 (.CI(n46414), .I0(n2729), .I1(n698), .CO(n46415));
    SB_LUT4 add_2550_3_lut (.I0(GND_net), .I1(n2730), .I2(n858), .I3(n46413), 
            .O(n7702[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2550_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2550_3 (.CI(n46413), .I0(n2730), .I1(n858), .CO(n46414));
    SB_LUT4 add_2550_2_lut (.I0(n53875), .I1(GND_net), .I2(n538), .I3(VCC_net), 
            .O(n55688)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2550_2_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_2550_2 (.CI(VCC_net), .I0(GND_net), .I1(n538), .CO(n46413));
    SB_LUT4 add_2549_19_lut (.I0(GND_net), .I1(n2596), .I2(n2867), .I3(n46412), 
            .O(n7676[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2549_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i47684_3_lut (.I0(n62396), .I1(baudrate[14]), .I2(n29_c), 
            .I3(GND_net), .O(n62397));   // verilog/uart_rx.v(119[33:55])
    defparam i47684_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i45609_4_lut (.I0(n33_c), .I1(n31), .I2(n29_c), .I3(n60335), 
            .O(n60321));
    defparam i45609_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 add_2549_18_lut (.I0(GND_net), .I1(n2597), .I2(n2754), .I3(n46411), 
            .O(n7676[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2549_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2549_18 (.CI(n46411), .I0(n2597), .I1(n2754), .CO(n46412));
    SB_LUT4 add_2549_17_lut (.I0(GND_net), .I1(n2598), .I2(n2638), .I3(n46410), 
            .O(n7676[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2549_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2549_17 (.CI(n46410), .I0(n2598), .I1(n2638), .CO(n46411));
    SB_LUT4 add_2549_16_lut (.I0(GND_net), .I1(n2599), .I2(n2519), .I3(n46409), 
            .O(n7676[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2549_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2549_16 (.CI(n46409), .I0(n2599), .I1(n2519), .CO(n46410));
    SB_LUT4 add_2549_15_lut (.I0(GND_net), .I1(n2600), .I2(n2397), .I3(n46408), 
            .O(n7676[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2549_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2549_15 (.CI(n46408), .I0(n2600), .I1(n2397), .CO(n46409));
    SB_LUT4 div_37_i1322_3_lut (.I0(n1835), .I1(n7520[19]), .I2(n294[12]), 
            .I3(GND_net), .O(n1970));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1322_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_2549_14_lut (.I0(GND_net), .I1(n2601), .I2(n2272), .I3(n46407), 
            .O(n7676[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2549_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2549_14 (.CI(n46407), .I0(n2601), .I1(n2272), .CO(n46408));
    SB_LUT4 add_2549_13_lut (.I0(GND_net), .I1(n2602), .I2(n2144), .I3(n46406), 
            .O(n7676[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2549_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2549_13 (.CI(n46406), .I0(n2602), .I1(n2144), .CO(n46407));
    SB_LUT4 add_2549_12_lut (.I0(GND_net), .I1(n2603), .I2(n2013), .I3(n46405), 
            .O(n7676[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2549_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2549_12 (.CI(n46405), .I0(n2603), .I1(n2013), .CO(n46406));
    SB_LUT4 add_2549_11_lut (.I0(GND_net), .I1(n2604), .I2(n1879), .I3(n46404), 
            .O(n7676[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2549_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2549_11 (.CI(n46404), .I0(n2604), .I1(n1879), .CO(n46405));
    SB_LUT4 add_2549_10_lut (.I0(GND_net), .I1(n2605), .I2(n1742), .I3(n46403), 
            .O(n7676[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2549_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2549_10 (.CI(n46403), .I0(n2605), .I1(n1742), .CO(n46404));
    SB_LUT4 add_2549_9_lut (.I0(GND_net), .I1(n2606), .I2(n1602), .I3(n46402), 
            .O(n7676[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2549_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2549_9 (.CI(n46402), .I0(n2606), .I1(n1602), .CO(n46403));
    SB_LUT4 add_2549_8_lut (.I0(GND_net), .I1(n2607), .I2(n1459), .I3(n46401), 
            .O(n7676[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2549_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2549_8 (.CI(n46401), .I0(n2607), .I1(n1459), .CO(n46402));
    SB_LUT4 i48138_4_lut (.I0(n30), .I1(n10), .I2(n35), .I3(n60313), 
            .O(n62851));   // verilog/uart_rx.v(119[33:55])
    defparam i48138_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 div_37_i641_4_lut (.I0(n804), .I1(n42), .I2(n294[19]), .I3(baudrate[2]), 
            .O(n960));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i641_4_lut.LUT_INIT = 16'h6a9a;
    SB_LUT4 i47638_3_lut (.I0(n62397), .I1(baudrate[15]), .I2(n31), .I3(GND_net), 
            .O(n62351));   // verilog/uart_rx.v(119[33:55])
    defparam i47638_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i48278_4_lut (.I0(n62351), .I1(n62851), .I2(n35), .I3(n60321), 
            .O(n62991));   // verilog/uart_rx.v(119[33:55])
    defparam i48278_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i48279_3_lut (.I0(n62991), .I1(baudrate[18]), .I2(n37), .I3(GND_net), 
            .O(n62992));   // verilog/uart_rx.v(119[33:55])
    defparam i48279_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1411_3_lut (.I0(n1970), .I1(n7546[19]), .I2(n294[11]), 
            .I3(GND_net), .O(n2102));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1411_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i48257_3_lut (.I0(n62992), .I1(baudrate[19]), .I2(n39), .I3(GND_net), 
            .O(n62970));   // verilog/uart_rx.v(119[33:55])
    defparam i48257_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1498_3_lut (.I0(n2102), .I1(n7572[19]), .I2(n294[10]), 
            .I3(GND_net), .O(n2231));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1498_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i45518_4_lut (.I0(n43), .I1(n25), .I2(n23_c), .I3(n60359), 
            .O(n60230));
    defparam i45518_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i47235_4_lut (.I0(n24), .I1(n8), .I2(n45_adj_4766), .I3(n60218), 
            .O(n61948));   // verilog/uart_rx.v(119[33:55])
    defparam i47235_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 add_2549_7_lut (.I0(GND_net), .I1(n2608), .I2(n1460), .I3(n46400), 
            .O(n7676[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2549_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i47636_3_lut (.I0(n62630), .I1(baudrate[12]), .I2(n25), .I3(GND_net), 
            .O(n62349));   // verilog/uart_rx.v(119[33:55])
    defparam i47636_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i45544_4_lut (.I0(n43), .I1(n41), .I2(n39), .I3(n62792), 
            .O(n60256));
    defparam i45544_4_lut.LUT_INIT = 16'haaab;
    SB_CARRY add_2549_7 (.CI(n46400), .I0(n2608), .I1(n1460), .CO(n46401));
    SB_LUT4 add_2549_6_lut (.I0(GND_net), .I1(n2609), .I2(n1011), .I3(n46399), 
            .O(n7676[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2549_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i47922_4_lut (.I0(n62349), .I1(n61948), .I2(n45_adj_4766), 
            .I3(n60230), .O(n62635));   // verilog/uart_rx.v(119[33:55])
    defparam i47922_4_lut.LUT_INIT = 16'hccca;
    SB_CARRY add_2549_6 (.CI(n46399), .I0(n2609), .I1(n1011), .CO(n46400));
    SB_LUT4 i48180_3_lut (.I0(n62970), .I1(baudrate[20]), .I2(n41), .I3(GND_net), 
            .O(n40));   // verilog/uart_rx.v(119[33:55])
    defparam i48180_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF r_Rx_Byte_i3 (.Q(rx_data[3]), .C(clk16MHz), .D(n26516));   // verilog/uart_rx.v(50[10] 145[8])
    SB_LUT4 add_2549_5_lut (.I0(GND_net), .I1(n2610), .I2(n856), .I3(n46398), 
            .O(n7676[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2549_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2549_5 (.CI(n46398), .I0(n2610), .I1(n856), .CO(n46399));
    SB_LUT4 div_37_i2187_3_lut (.I0(n3151), .I1(n7806[23]), .I2(n294[1]), 
            .I3(GND_net), .O(n3253));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2187_3_lut.LUT_INIT = 16'hcaca;
    SB_DFFESR r_Clock_Count_1948__i7 (.Q(r_Clock_Count[7]), .C(clk16MHz), 
            .E(n24619), .D(n1[7]), .R(n25950));   // verilog/uart_rx.v(121[34:51])
    SB_LUT4 i47924_4_lut (.I0(n40), .I1(n62635), .I2(n45_adj_4766), .I3(n60256), 
            .O(n62637));   // verilog/uart_rx.v(119[33:55])
    defparam i47924_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i1_4_lut (.I0(n56554), .I1(n56484), .I2(n56430), .I3(n56356), 
            .O(n55652));
    defparam i1_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i48434_4_lut (.I0(n55652), .I1(n62637), .I2(baudrate[23]), 
            .I3(n3253), .O(n54733));   // verilog/uart_rx.v(119[33:55])
    defparam i48434_4_lut.LUT_INIT = 16'h1501;
    SB_LUT4 add_2549_4_lut (.I0(GND_net), .I1(n2611), .I2(n698), .I3(n46397), 
            .O(n7676[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2549_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2549_4 (.CI(n46397), .I0(n2611), .I1(n698), .CO(n46398));
    SB_LUT4 div_37_i1583_3_lut (.I0(n2231), .I1(n7598[19]), .I2(n294[9]), 
            .I3(GND_net), .O(n2357));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1583_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_2549_3_lut (.I0(GND_net), .I1(n2612), .I2(n858), .I3(n46396), 
            .O(n7676[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2549_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_i1666_3_lut (.I0(n2357), .I1(n7624[19]), .I2(n294[8]), 
            .I3(GND_net), .O(n2480));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1666_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_2549_3 (.CI(n46396), .I0(n2612), .I1(n858), .CO(n46397));
    SB_LUT4 add_2549_2_lut (.I0(n53879), .I1(GND_net), .I2(n538), .I3(VCC_net), 
            .O(n55686)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2549_2_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_2549_2 (.CI(VCC_net), .I0(GND_net), .I1(n538), .CO(n46396));
    SB_LUT4 add_2548_18_lut (.I0(GND_net), .I1(n2476), .I2(n2754), .I3(n46395), 
            .O(n7650[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2548_18_lut.LUT_INIT = 16'hC33C;
    SB_DFFESR r_Clock_Count_1948__i6 (.Q(r_Clock_Count[6]), .C(clk16MHz), 
            .E(n24619), .D(n1[6]), .R(n25950));   // verilog/uart_rx.v(121[34:51])
    SB_LUT4 add_2548_17_lut (.I0(GND_net), .I1(n2477), .I2(n2638), .I3(n46394), 
            .O(n7650[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2548_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_i2118_3_lut (.I0(n3046), .I1(n7780[23]), .I2(n294[2]), 
            .I3(GND_net), .O(n3151));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2118_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2121_3_lut (.I0(n3049), .I1(n7780[20]), .I2(n294[2]), 
            .I3(GND_net), .O(n3154));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2121_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2119_3_lut (.I0(n3047), .I1(n7780[22]), .I2(n294[2]), 
            .I3(GND_net), .O(n3152));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2119_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2120_3_lut (.I0(n3048), .I1(n7780[21]), .I2(n294[2]), 
            .I3(GND_net), .O(n3153));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2120_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2122_3_lut (.I0(n3050), .I1(n7780[19]), .I2(n294[2]), 
            .I3(GND_net), .O(n3155));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2122_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2125_3_lut (.I0(n3053), .I1(n7780[16]), .I2(n294[2]), 
            .I3(GND_net), .O(n3158));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2125_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_2141_i33_2_lut (.I0(n3158), .I1(baudrate[15]), 
            .I2(GND_net), .I3(GND_net), .O(n33_adj_4768));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2141_i33_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i2123_3_lut (.I0(n3051), .I1(n7780[18]), .I2(n294[2]), 
            .I3(GND_net), .O(n3156));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2123_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_2141_i37_2_lut (.I0(n3156), .I1(baudrate[17]), 
            .I2(GND_net), .I3(GND_net), .O(n37_adj_4769));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2141_i37_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i2124_3_lut (.I0(n3052), .I1(n7780[17]), .I2(n294[2]), 
            .I3(GND_net), .O(n3157));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2124_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_2141_i35_2_lut (.I0(n3157), .I1(baudrate[16]), 
            .I2(GND_net), .I3(GND_net), .O(n35_adj_4770));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2141_i35_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i2126_3_lut (.I0(n3054), .I1(n7780[15]), .I2(n294[2]), 
            .I3(GND_net), .O(n3159));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2126_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_2141_i31_2_lut (.I0(n3159), .I1(baudrate[14]), 
            .I2(GND_net), .I3(GND_net), .O(n31_adj_4771));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2141_i31_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i2128_3_lut (.I0(n3056), .I1(n7780[13]), .I2(n294[2]), 
            .I3(GND_net), .O(n3161));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2128_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1747_3_lut (.I0(n2480), .I1(n7650[19]), .I2(n294[7]), 
            .I3(GND_net), .O(n2600));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1747_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2129_3_lut (.I0(n3057), .I1(n7780[12]), .I2(n294[2]), 
            .I3(GND_net), .O(n3162));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2129_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_2141_i25_2_lut (.I0(n3162), .I1(baudrate[11]), 
            .I2(GND_net), .I3(GND_net), .O(n25_adj_4772));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2141_i25_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_2141_i27_2_lut (.I0(n3161), .I1(baudrate[12]), 
            .I2(GND_net), .I3(GND_net), .O(n27_adj_4773));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2141_i27_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_2548_17 (.CI(n46394), .I0(n2477), .I1(n2638), .CO(n46395));
    SB_LUT4 div_37_i2130_3_lut (.I0(n3058), .I1(n7780[11]), .I2(n294[2]), 
            .I3(GND_net), .O(n3163));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2130_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2131_3_lut (.I0(n3059), .I1(n7780[10]), .I2(n294[2]), 
            .I3(GND_net), .O(n3164));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2131_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_2548_16_lut (.I0(GND_net), .I1(n2478), .I2(n2519), .I3(n46393), 
            .O(n7650[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2548_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_4_lut_adj_948 (.I0(n22504), .I1(n48_adj_4774), .I2(n35471), 
            .I3(baudrate[2]), .O(n54412));
    defparam i1_4_lut_adj_948.LUT_INIT = 16'hefff;
    SB_LUT4 div_37_LessThan_2141_i21_2_lut (.I0(n3164), .I1(baudrate[9]), 
            .I2(GND_net), .I3(GND_net), .O(n21_adj_4775));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2141_i21_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_2141_i23_2_lut (.I0(n3163), .I1(baudrate[10]), 
            .I2(GND_net), .I3(GND_net), .O(n23_adj_4776));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2141_i23_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i2137_3_lut (.I0(n3065), .I1(n7780[4]), .I2(n294[2]), 
            .I3(GND_net), .O(n3170));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2137_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2138_3_lut (.I0(n3066), .I1(n7780[3]), .I2(n294[2]), 
            .I3(GND_net), .O(n3171));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2138_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_2141_i9_2_lut (.I0(n3170), .I1(baudrate[3]), 
            .I2(GND_net), .I3(GND_net), .O(n9_adj_4777));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2141_i9_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i2132_3_lut (.I0(n3060), .I1(n7780[9]), .I2(n294[2]), 
            .I3(GND_net), .O(n3165));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2132_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1826_3_lut (.I0(n2600), .I1(n7676[19]), .I2(n294[6]), 
            .I3(GND_net), .O(n2717));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1826_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2136_3_lut (.I0(n3064), .I1(n7780[5]), .I2(n294[2]), 
            .I3(GND_net), .O(n3169));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2136_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_2141_i11_2_lut (.I0(n3169), .I1(baudrate[4]), 
            .I2(GND_net), .I3(GND_net), .O(n11_adj_4778));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2141_i11_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_2141_i19_2_lut (.I0(n3165), .I1(baudrate[8]), 
            .I2(GND_net), .I3(GND_net), .O(n19_adj_4779));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2141_i19_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i2134_3_lut (.I0(n3062), .I1(n7780[7]), .I2(n294[2]), 
            .I3(GND_net), .O(n3167));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2134_3_lut.LUT_INIT = 16'hcaca;
    SB_DFFESR r_Clock_Count_1948__i5 (.Q(r_Clock_Count[5]), .C(clk16MHz), 
            .E(n24619), .D(n1[5]), .R(n25950));   // verilog/uart_rx.v(121[34:51])
    SB_LUT4 div_37_i2127_3_lut (.I0(n3055), .I1(n7780[14]), .I2(n294[2]), 
            .I3(GND_net), .O(n3160));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2127_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2133_3_lut (.I0(n3061), .I1(n7780[8]), .I2(n294[2]), 
            .I3(GND_net), .O(n3166));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2133_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2135_3_lut (.I0(n3063), .I1(n7780[6]), .I2(n294[2]), 
            .I3(GND_net), .O(n3168));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2135_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_2141_i13_2_lut (.I0(n3168), .I1(baudrate[5]), 
            .I2(GND_net), .I3(GND_net), .O(n13_adj_4781));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2141_i13_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_2141_i15_2_lut (.I0(n3167), .I1(baudrate[6]), 
            .I2(GND_net), .I3(GND_net), .O(n15_adj_4782));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2141_i15_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_2141_i17_2_lut (.I0(n3166), .I1(baudrate[7]), 
            .I2(GND_net), .I3(GND_net), .O(n17_adj_4783));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2141_i17_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_2141_i29_2_lut (.I0(n3160), .I1(baudrate[13]), 
            .I2(GND_net), .I3(GND_net), .O(n29_adj_4784));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2141_i29_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut (.I0(baudrate[25]), .I1(baudrate[29]), .I2(GND_net), 
            .I3(GND_net), .O(n56556));
    defparam i1_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i1_2_lut_adj_949 (.I0(baudrate[24]), .I1(baudrate[31]), .I2(GND_net), 
            .I3(GND_net), .O(n56558));
    defparam i1_2_lut_adj_949.LUT_INIT = 16'heeee;
    SB_DFFESR r_Clock_Count_1948__i4 (.Q(r_Clock_Count[4]), .C(clk16MHz), 
            .E(n24619), .D(n1[4]), .R(n25950));   // verilog/uart_rx.v(121[34:51])
    SB_DFFESR r_Clock_Count_1948__i3 (.Q(r_Clock_Count[3]), .C(clk16MHz), 
            .E(n24619), .D(n1[3]), .R(n25950));   // verilog/uart_rx.v(121[34:51])
    SB_LUT4 i3672_4_lut (.I0(n644), .I1(baudrate[2]), .I2(n54412), .I3(n44), 
            .O(n46));   // verilog/uart_rx.v(119[33:55])
    defparam i3672_4_lut.LUT_INIT = 16'hb3a0;
    SB_LUT4 div_37_i744_4_lut (.I0(n960), .I1(baudrate[3]), .I2(n294[18]), 
            .I3(n42_adj_4787), .O(n1113));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i744_4_lut.LUT_INIT = 16'h6a9a;
    SB_DFFESR r_Clock_Count_1948__i2 (.Q(r_Clock_Count[2]), .C(clk16MHz), 
            .E(n24619), .D(n1[2]), .R(n25950));   // verilog/uart_rx.v(121[34:51])
    SB_LUT4 div_37_i534_4_lut (.I0(n53644), .I1(n294[20]), .I2(n46), .I3(baudrate[3]), 
            .O(n53646));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i534_4_lut.LUT_INIT = 16'h6aa6;
    SB_DFFESR r_Clock_Count_1948__i1 (.Q(r_Clock_Count[1]), .C(clk16MHz), 
            .E(n24619), .D(n1[1]), .R(n25950));   // verilog/uart_rx.v(121[34:51])
    SB_LUT4 div_37_i845_3_lut (.I0(n1113), .I1(n7390[21]), .I2(n294[17]), 
            .I3(GND_net), .O(n1263));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i845_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_adj_950 (.I0(baudrate[26]), .I1(baudrate[30]), .I2(GND_net), 
            .I3(GND_net), .O(n56554));
    defparam i1_2_lut_adj_950.LUT_INIT = 16'heeee;
    SB_LUT4 i1_4_lut_adj_951 (.I0(n56558), .I1(n56560), .I2(n56356), .I3(n56556), 
            .O(n22434));
    defparam i1_4_lut_adj_951.LUT_INIT = 16'hfffe;
    SB_LUT4 div_37_LessThan_866_i41_2_lut (.I0(n1264), .I1(baudrate[4]), 
            .I2(GND_net), .I3(GND_net), .O(n41_adj_4790));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_866_i41_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i45761_4_lut (.I0(n29_adj_4784), .I1(n17_adj_4783), .I2(n15_adj_4782), 
            .I3(n13_adj_4781), .O(n60473));
    defparam i45761_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i46756_4_lut (.I0(n11_adj_4778), .I1(n9_adj_4777), .I2(n3171), 
            .I3(baudrate[2]), .O(n61469));
    defparam i46756_4_lut.LUT_INIT = 16'heffe;
    SB_LUT4 i47295_4_lut (.I0(n17_adj_4783), .I1(n15_adj_4782), .I2(n13_adj_4781), 
            .I3(n61469), .O(n62008));
    defparam i47295_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i47289_4_lut (.I0(n23_adj_4776), .I1(n21_adj_4775), .I2(n19_adj_4779), 
            .I3(n62008), .O(n62002));
    defparam i47289_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i45769_4_lut (.I0(n29_adj_4784), .I1(n27_adj_4773), .I2(n25_adj_4772), 
            .I3(n62002), .O(n60481));
    defparam i45769_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 div_37_LessThan_2141_i6_3_lut (.I0(baudrate[0]), .I1(baudrate[1]), 
            .I2(n3172), .I3(GND_net), .O(n6_adj_4791));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2141_i6_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i47465_3_lut (.I0(n6_adj_4791), .I1(baudrate[13]), .I2(n29_adj_4784), 
            .I3(GND_net), .O(n62178));   // verilog/uart_rx.v(119[33:55])
    defparam i47465_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_2141_i32_3_lut (.I0(n14), .I1(baudrate[17]), 
            .I2(n37_adj_4769), .I3(GND_net), .O(n32));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2141_i32_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i47466_3_lut (.I0(n62178), .I1(baudrate[14]), .I2(n31_adj_4771), 
            .I3(GND_net), .O(n62179));   // verilog/uart_rx.v(119[33:55])
    defparam i47466_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i45755_4_lut (.I0(n35_adj_4770), .I1(n33_adj_4768), .I2(n31_adj_4771), 
            .I3(n60473), .O(n60467));
    defparam i45755_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i48008_4_lut (.I0(n32), .I1(n12_adj_4792), .I2(n37_adj_4769), 
            .I3(n60463), .O(n62721));   // verilog/uart_rx.v(119[33:55])
    defparam i48008_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i46621_3_lut (.I0(n62179), .I1(baudrate[15]), .I2(n33_adj_4768), 
            .I3(GND_net), .O(n61334));   // verilog/uart_rx.v(119[33:55])
    defparam i46621_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i47467_3_lut (.I0(n8_adj_4793), .I1(baudrate[10]), .I2(n23_adj_4776), 
            .I3(GND_net), .O(n62180));   // verilog/uart_rx.v(119[33:55])
    defparam i47467_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_2548_16 (.CI(n46393), .I0(n2478), .I1(n2519), .CO(n46394));
    SB_LUT4 add_2548_15_lut (.I0(GND_net), .I1(n2479), .I2(n2397), .I3(n46392), 
            .O(n7650[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2548_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i47468_3_lut (.I0(n62180), .I1(baudrate[11]), .I2(n25_adj_4772), 
            .I3(GND_net), .O(n62181));   // verilog/uart_rx.v(119[33:55])
    defparam i47468_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i46734_4_lut (.I0(n25_adj_4772), .I1(n23_adj_4776), .I2(n21_adj_4775), 
            .I3(n60503), .O(n61447));
    defparam i46734_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i47231_3_lut (.I0(n10_adj_4794), .I1(baudrate[9]), .I2(n21_adj_4775), 
            .I3(GND_net), .O(n61944));   // verilog/uart_rx.v(119[33:55])
    defparam i47231_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i46619_3_lut (.I0(n62181), .I1(baudrate[12]), .I2(n27_adj_4773), 
            .I3(GND_net), .O(n61332));   // verilog/uart_rx.v(119[33:55])
    defparam i46619_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i47673_4_lut (.I0(n35_adj_4770), .I1(n33_adj_4768), .I2(n31_adj_4771), 
            .I3(n60481), .O(n62386));
    defparam i47673_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 div_37_i1824_3_lut (.I0(n2598), .I1(n7676[21]), .I2(n294[6]), 
            .I3(GND_net), .O(n2715));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1824_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i48203_4_lut (.I0(n61334), .I1(n62721), .I2(n37_adj_4769), 
            .I3(n60467), .O(n62916));   // verilog/uart_rx.v(119[33:55])
    defparam i48203_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i47685_4_lut (.I0(n61332), .I1(n61944), .I2(n27_adj_4773), 
            .I3(n61447), .O(n62398));   // verilog/uart_rx.v(119[33:55])
    defparam i47685_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i48284_4_lut (.I0(n62398), .I1(n62916), .I2(n37_adj_4769), 
            .I3(n62386), .O(n62997));   // verilog/uart_rx.v(119[33:55])
    defparam i48284_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i48285_3_lut (.I0(n62997), .I1(baudrate[18]), .I2(n3155), 
            .I3(GND_net), .O(n62998));   // verilog/uart_rx.v(119[33:55])
    defparam i48285_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i48137_3_lut (.I0(n62998), .I1(baudrate[19]), .I2(n3154), 
            .I3(GND_net), .O(n62850));   // verilog/uart_rx.v(119[33:55])
    defparam i48137_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i48048_3_lut (.I0(n62850), .I1(baudrate[20]), .I2(n3153), 
            .I3(GND_net), .O(n62761));   // verilog/uart_rx.v(119[33:55])
    defparam i48048_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i48049_3_lut (.I0(n62761), .I1(baudrate[21]), .I2(n3152), 
            .I3(GND_net), .O(n62762));   // verilog/uart_rx.v(119[33:55])
    defparam i48049_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i47915_3_lut (.I0(n62762), .I1(baudrate[22]), .I2(n3151), 
            .I3(GND_net), .O(n48));   // verilog/uart_rx.v(119[33:55])
    defparam i47915_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_i2047_3_lut (.I0(n2938), .I1(n7754[23]), .I2(n294[3]), 
            .I3(GND_net), .O(n3046));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2047_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2055_3_lut (.I0(n2946), .I1(n7754[15]), .I2(n294[3]), 
            .I3(GND_net), .O(n3054));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2055_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2050_3_lut (.I0(n2941), .I1(n7754[20]), .I2(n294[3]), 
            .I3(GND_net), .O(n3049));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2050_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2048_3_lut (.I0(n2939), .I1(n7754[22]), .I2(n294[3]), 
            .I3(GND_net), .O(n3047));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2048_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2049_3_lut (.I0(n2940), .I1(n7754[21]), .I2(n294[3]), 
            .I3(GND_net), .O(n3048));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2049_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2053_3_lut (.I0(n2944), .I1(n7754[17]), .I2(n294[3]), 
            .I3(GND_net), .O(n3052));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2053_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_2070_i35_2_lut (.I0(n3052), .I1(baudrate[15]), 
            .I2(GND_net), .I3(GND_net), .O(n35_adj_4795));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2070_i35_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i2051_3_lut (.I0(n2942), .I1(n7754[19]), .I2(n294[3]), 
            .I3(GND_net), .O(n3050));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2051_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_2070_i39_2_lut (.I0(n3050), .I1(baudrate[17]), 
            .I2(GND_net), .I3(GND_net), .O(n39_adj_4796));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2070_i39_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i2054_3_lut (.I0(n2945), .I1(n7754[16]), .I2(n294[3]), 
            .I3(GND_net), .O(n3053));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2054_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_2070_i33_2_lut (.I0(n3053), .I1(baudrate[14]), 
            .I2(GND_net), .I3(GND_net), .O(n33_adj_4797));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2070_i33_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i2052_3_lut (.I0(n2943), .I1(n7754[18]), .I2(n294[3]), 
            .I3(GND_net), .O(n3051));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2052_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_2070_i37_2_lut (.I0(n3051), .I1(baudrate[16]), 
            .I2(GND_net), .I3(GND_net), .O(n37_adj_4798));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2070_i37_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i2056_3_lut (.I0(n2947), .I1(n7754[14]), .I2(n294[3]), 
            .I3(GND_net), .O(n3055));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2056_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2057_3_lut (.I0(n2948), .I1(n7754[13]), .I2(n294[3]), 
            .I3(GND_net), .O(n3056));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2057_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_2548_15 (.CI(n46392), .I0(n2479), .I1(n2397), .CO(n46393));
    SB_LUT4 add_2548_14_lut (.I0(GND_net), .I1(n2480), .I2(n2272), .I3(n46391), 
            .O(n7650[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2548_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_LessThan_2070_i27_2_lut (.I0(n3056), .I1(baudrate[11]), 
            .I2(GND_net), .I3(GND_net), .O(n27_adj_4799));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2070_i27_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_2070_i29_2_lut (.I0(n3055), .I1(baudrate[12]), 
            .I2(GND_net), .I3(GND_net), .O(n29_adj_4800));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2070_i29_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_2548_14 (.CI(n46391), .I0(n2480), .I1(n2272), .CO(n46392));
    SB_LUT4 div_37_i2058_3_lut (.I0(n2949), .I1(n7754[12]), .I2(n294[3]), 
            .I3(GND_net), .O(n3057));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2058_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1845_i39_2_lut (.I0(n2717), .I1(baudrate[14]), 
            .I2(GND_net), .I3(GND_net), .O(n39_adj_4801));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1845_i39_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i2059_3_lut (.I0(n2950), .I1(n7754[11]), .I2(n294[3]), 
            .I3(GND_net), .O(n3058));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2059_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_2548_13_lut (.I0(GND_net), .I1(n2481), .I2(n2144), .I3(n46390), 
            .O(n7650[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2548_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2548_13 (.CI(n46390), .I0(n2481), .I1(n2144), .CO(n46391));
    SB_LUT4 add_2548_12_lut (.I0(GND_net), .I1(n2482), .I2(n2013), .I3(n46389), 
            .O(n7650[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2548_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2548_12 (.CI(n46389), .I0(n2482), .I1(n2013), .CO(n46390));
    SB_LUT4 add_2548_11_lut (.I0(GND_net), .I1(n2483), .I2(n1879), .I3(n46388), 
            .O(n7650[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2548_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_LessThan_2070_i23_2_lut (.I0(n3058), .I1(baudrate[9]), 
            .I2(GND_net), .I3(GND_net), .O(n23_adj_4802));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2070_i23_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_2070_i25_2_lut (.I0(n3057), .I1(baudrate[10]), 
            .I2(GND_net), .I3(GND_net), .O(n25_adj_4803));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2070_i25_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i3841_4_lut (.I0(n803), .I1(baudrate[3]), .I2(n9112), .I3(n18960), 
            .O(n46_adj_4804));   // verilog/uart_rx.v(119[33:55])
    defparam i3841_4_lut.LUT_INIT = 16'hbbb2;
    SB_LUT4 div_37_i2065_3_lut (.I0(n2956), .I1(n7754[5]), .I2(n294[3]), 
            .I3(GND_net), .O(n3064));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2065_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_2548_11 (.CI(n46388), .I0(n2483), .I1(n1879), .CO(n46389));
    SB_LUT4 add_2548_10_lut (.I0(GND_net), .I1(n2484), .I2(n1742), .I3(n46387), 
            .O(n7650[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2548_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_i2066_3_lut (.I0(n2957), .I1(n7754[4]), .I2(n294[3]), 
            .I3(GND_net), .O(n3065));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2066_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_2548_10 (.CI(n46387), .I0(n2484), .I1(n1742), .CO(n46388));
    SB_LUT4 div_37_LessThan_2070_i11_2_lut (.I0(n3064), .I1(baudrate[3]), 
            .I2(GND_net), .I3(GND_net), .O(n11_adj_4805));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2070_i11_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i2060_3_lut (.I0(n2951), .I1(n7754[10]), .I2(n294[3]), 
            .I3(GND_net), .O(n3059));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2060_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2064_3_lut (.I0(n2955), .I1(n7754[6]), .I2(n294[3]), 
            .I3(GND_net), .O(n3063));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2064_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_2548_9_lut (.I0(GND_net), .I1(n2485), .I2(n1602), .I3(n46386), 
            .O(n7650[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2548_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_LessThan_2070_i13_2_lut (.I0(n3063), .I1(baudrate[4]), 
            .I2(GND_net), .I3(GND_net), .O(n13_adj_4806));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2070_i13_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_2070_i21_2_lut (.I0(n3059), .I1(baudrate[8]), 
            .I2(GND_net), .I3(GND_net), .O(n21_adj_4807));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2070_i21_2_lut.LUT_INIT = 16'h6666;
    SB_DFFSR r_SM_Main_i0 (.Q(r_SM_Main[0]), .C(clk16MHz), .D(n3), .R(\r_SM_Main[2] ));   // verilog/uart_rx.v(50[10] 145[8])
    SB_CARRY add_2548_9 (.CI(n46386), .I0(n2485), .I1(n1602), .CO(n46387));
    SB_LUT4 div_37_i2061_3_lut (.I0(n2952), .I1(n7754[9]), .I2(n294[3]), 
            .I3(GND_net), .O(n3060));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2061_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2062_3_lut (.I0(n2953), .I1(n7754[8]), .I2(n294[3]), 
            .I3(GND_net), .O(n3061));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2062_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_2548_8_lut (.I0(GND_net), .I1(n2486), .I2(n1459), .I3(n46385), 
            .O(n7650[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2548_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2548_8 (.CI(n46385), .I0(n2486), .I1(n1459), .CO(n46386));
    SB_LUT4 add_2548_7_lut (.I0(GND_net), .I1(n2487), .I2(n1460), .I3(n46384), 
            .O(n7650[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2548_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_i2063_3_lut (.I0(n2954), .I1(n7754[7]), .I2(n294[3]), 
            .I3(GND_net), .O(n3062));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2063_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF r_Rx_Data_56 (.Q(r_Rx_Data), .C(clk16MHz), .D(r_Rx_Data_R));   // verilog/uart_rx.v(42[10] 46[8])
    SB_LUT4 div_37_LessThan_1845_i41_2_lut (.I0(n2716), .I1(baudrate[15]), 
            .I2(GND_net), .I3(GND_net), .O(n41_adj_4808));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1845_i41_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1845_i43_2_lut (.I0(n2715), .I1(baudrate[16]), 
            .I2(GND_net), .I3(GND_net), .O(n43_adj_4809));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1845_i43_2_lut.LUT_INIT = 16'h6666;
    SB_DFF r_Rx_Data_R_55 (.Q(r_Rx_Data_R), .C(clk16MHz), .D(RX_N_42));   // verilog/uart_rx.v(42[10] 46[8])
    SB_LUT4 div_37_LessThan_2070_i15_2_lut (.I0(n3062), .I1(baudrate[5]), 
            .I2(GND_net), .I3(GND_net), .O(n15_adj_4810));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2070_i15_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_2070_i17_2_lut (.I0(n3061), .I1(baudrate[6]), 
            .I2(GND_net), .I3(GND_net), .O(n17_adj_4811));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2070_i17_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_2070_i19_2_lut (.I0(n3060), .I1(baudrate[7]), 
            .I2(GND_net), .I3(GND_net), .O(n19_adj_4812));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2070_i19_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_2070_i31_2_lut (.I0(n3054), .I1(baudrate[13]), 
            .I2(GND_net), .I3(GND_net), .O(n31_adj_4813));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2070_i31_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_2548_7 (.CI(n46384), .I0(n2487), .I1(n1460), .CO(n46385));
    SB_LUT4 i45851_4_lut (.I0(n31_adj_4813), .I1(n19_adj_4812), .I2(n17_adj_4811), 
            .I3(n15_adj_4810), .O(n60563));
    defparam i45851_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 add_2548_6_lut (.I0(GND_net), .I1(n2488), .I2(n1011), .I3(n46383), 
            .O(n7650[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2548_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2548_6 (.CI(n46383), .I0(n2488), .I1(n1011), .CO(n46384));
    SB_LUT4 add_2548_5_lut (.I0(GND_net), .I1(n2489), .I2(n856), .I3(n46382), 
            .O(n7650[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2548_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i46830_4_lut (.I0(n13_adj_4806), .I1(n11_adj_4805), .I2(n3065), 
            .I3(baudrate[2]), .O(n61543));
    defparam i46830_4_lut.LUT_INIT = 16'heffe;
    SB_LUT4 i47325_4_lut (.I0(n19_adj_4812), .I1(n17_adj_4811), .I2(n15_adj_4810), 
            .I3(n61543), .O(n62038));
    defparam i47325_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i47321_4_lut (.I0(n25_adj_4803), .I1(n23_adj_4802), .I2(n21_adj_4807), 
            .I3(n62038), .O(n62034));
    defparam i47321_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i45855_4_lut (.I0(n31_adj_4813), .I1(n29_adj_4800), .I2(n27_adj_4799), 
            .I3(n62034), .O(n60567));
    defparam i45855_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 div_37_LessThan_2070_i8_3_lut (.I0(baudrate[0]), .I1(baudrate[1]), 
            .I2(n3066), .I3(GND_net), .O(n8_adj_4814));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2070_i8_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_i1040_3_lut (.I0(n1409), .I1(n7442[22]), .I2(n294[15]), 
            .I3(GND_net), .O(n1553));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1040_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i47473_3_lut (.I0(n8_adj_4814), .I1(baudrate[13]), .I2(n31_adj_4813), 
            .I3(GND_net), .O(n62186));   // verilog/uart_rx.v(119[33:55])
    defparam i47473_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i47474_3_lut (.I0(n62186), .I1(baudrate[14]), .I2(n33_adj_4797), 
            .I3(GND_net), .O(n62187));   // verilog/uart_rx.v(119[33:55])
    defparam i47474_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_2548_5 (.CI(n46382), .I0(n2489), .I1(n856), .CO(n46383));
    SB_LUT4 add_2548_4_lut (.I0(GND_net), .I1(n2490), .I2(n698), .I3(n46381), 
            .O(n7650[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2548_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_LessThan_2070_i34_3_lut (.I0(n16_adj_4815), .I1(baudrate[17]), 
            .I2(n39_adj_4796), .I3(GND_net), .O(n34_c));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2070_i34_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i45835_4_lut (.I0(n37_adj_4798), .I1(n35_adj_4795), .I2(n33_adj_4797), 
            .I3(n60563), .O(n60547));
    defparam i45835_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 sub_38_add_2_26_lut (.I0(GND_net), .I1(GND_net), .I2(VCC_net), 
            .I3(n46149), .O(\o_Rx_DV_N_3261[24] )) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_26_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_38_add_2_25_lut (.I0(n55658), .I1(n294[23]), .I2(VCC_net), 
            .I3(n46148), .O(n27)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_25_lut.LUT_INIT = 16'hebbe;
    SB_LUT4 i47984_4_lut (.I0(n34_c), .I1(n14_adj_4817), .I2(n39_adj_4796), 
            .I3(n60539), .O(n62697));   // verilog/uart_rx.v(119[33:55])
    defparam i47984_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 div_37_LessThan_866_i36_3_lut (.I0(baudrate[0]), .I1(baudrate[1]), 
            .I2(n1267), .I3(GND_net), .O(n36));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_866_i36_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i46609_3_lut (.I0(n62187), .I1(baudrate[15]), .I2(n35_adj_4795), 
            .I3(GND_net), .O(n61322));   // verilog/uart_rx.v(119[33:55])
    defparam i46609_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i47475_3_lut (.I0(n10_adj_4818), .I1(baudrate[10]), .I2(n25_adj_4803), 
            .I3(GND_net), .O(n62188));   // verilog/uart_rx.v(119[33:55])
    defparam i47475_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_2548_4 (.CI(n46381), .I0(n2490), .I1(n698), .CO(n46382));
    SB_CARRY sub_38_add_2_25 (.CI(n46148), .I0(n294[23]), .I1(VCC_net), 
            .CO(n46149));
    SB_LUT4 add_2548_3_lut (.I0(GND_net), .I1(n2491), .I2(n858), .I3(n46380), 
            .O(n7650[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2548_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i47476_3_lut (.I0(n62188), .I1(baudrate[11]), .I2(n27_adj_4799), 
            .I3(GND_net), .O(n62189));   // verilog/uart_rx.v(119[33:55])
    defparam i47476_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i46808_4_lut (.I0(n27_adj_4799), .I1(n25_adj_4803), .I2(n23_adj_4802), 
            .I3(n60579), .O(n61521));
    defparam i46808_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 div_37_LessThan_2070_i20_3_lut (.I0(n12_adj_4819), .I1(baudrate[9]), 
            .I2(n23_adj_4802), .I3(GND_net), .O(n20));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2070_i20_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2160_1_lut (.I0(baudrate[15]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n2638));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2160_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i46607_3_lut (.I0(n62189), .I1(baudrate[12]), .I2(n29_adj_4800), 
            .I3(GND_net), .O(n61320));   // verilog/uart_rx.v(119[33:55])
    defparam i46607_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_2548_3 (.CI(n46380), .I0(n2491), .I1(n858), .CO(n46381));
    SB_LUT4 add_2548_2_lut (.I0(n53883), .I1(GND_net), .I2(n538), .I3(VCC_net), 
            .O(n55684)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2548_2_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_2548_2 (.CI(VCC_net), .I0(GND_net), .I1(n538), .CO(n46380));
    SB_LUT4 add_2547_17_lut (.I0(GND_net), .I1(n2353), .I2(n2638), .I3(n46379), 
            .O(n7624[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2547_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_i1135_3_lut (.I0(n1553), .I1(n7468[22]), .I2(n294[14]), 
            .I3(GND_net), .O(n1694));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1135_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i47715_4_lut (.I0(n37_adj_4798), .I1(n35_adj_4795), .I2(n33_adj_4797), 
            .I3(n60567), .O(n62428));
    defparam i47715_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i48201_4_lut (.I0(n61322), .I1(n62697), .I2(n39_adj_4796), 
            .I3(n60547), .O(n62914));   // verilog/uart_rx.v(119[33:55])
    defparam i48201_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i47229_4_lut (.I0(n61320), .I1(n20), .I2(n29_adj_4800), .I3(n61521), 
            .O(n61942));   // verilog/uart_rx.v(119[33:55])
    defparam i47229_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i48280_4_lut (.I0(n61942), .I1(n62914), .I2(n39_adj_4796), 
            .I3(n62428), .O(n62993));   // verilog/uart_rx.v(119[33:55])
    defparam i48280_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 div_37_i1228_3_lut (.I0(n1694), .I1(n7494[22]), .I2(n294[13]), 
            .I3(GND_net), .O(n1832));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1228_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i639_4_lut (.I0(n53646), .I1(n294[19]), .I2(n46_adj_4804), 
            .I3(baudrate[4]), .O(n53648));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i639_4_lut.LUT_INIT = 16'h6aa6;
    SB_LUT4 div_37_i1319_3_lut (.I0(n1832), .I1(n7520[22]), .I2(n294[12]), 
            .I3(GND_net), .O(n1967));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1319_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i48281_3_lut (.I0(n62993), .I1(baudrate[18]), .I2(n3049), 
            .I3(GND_net), .O(n62994));   // verilog/uart_rx.v(119[33:55])
    defparam i48281_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_i1408_3_lut (.I0(n1967), .I1(n7546[22]), .I2(n294[11]), 
            .I3(GND_net), .O(n2099));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1408_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1495_3_lut (.I0(n2099), .I1(n7572[22]), .I2(n294[10]), 
            .I3(GND_net), .O(n2228));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1495_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i47687_3_lut (.I0(n62994), .I1(baudrate[19]), .I2(n3048), 
            .I3(GND_net), .O(n62400));   // verilog/uart_rx.v(119[33:55])
    defparam i47687_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 sub_38_add_2_24_lut (.I0(n55708), .I1(n56822), .I2(VCC_net), 
            .I3(n46147), .O(n29)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_24_lut.LUT_INIT = 16'hebbe;
    SB_LUT4 i47688_3_lut (.I0(n62400), .I1(baudrate[20]), .I2(n3047), 
            .I3(GND_net), .O(n62401));   // verilog/uart_rx.v(119[33:55])
    defparam i47688_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_i2159_1_lut (.I0(baudrate[16]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n2754));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2159_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY sub_38_add_2_24 (.CI(n46147), .I0(n56822), .I1(VCC_net), 
            .CO(n46148));
    SB_LUT4 i1_3_lut_4_lut (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[2]), .I2(\r_Bit_Index[0] ), 
            .I3(n4_adj_4821), .O(n55980));
    defparam i1_3_lut_4_lut.LUT_INIT = 16'hff7f;
    SB_LUT4 add_2547_16_lut (.I0(GND_net), .I1(n2354), .I2(n2519), .I3(n46378), 
            .O(n7624[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2547_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_i1580_3_lut (.I0(n2228), .I1(n7598[22]), .I2(n294[9]), 
            .I3(GND_net), .O(n2354));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1580_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_866_i40_3_lut (.I0(n38_adj_4822), .I1(baudrate[4]), 
            .I2(n41_adj_4790), .I3(GND_net), .O(n40_adj_4823));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_866_i40_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_2547_16 (.CI(n46378), .I0(n2354), .I1(n2519), .CO(n46379));
    SB_LUT4 sub_38_add_2_23_lut (.I0(o_Rx_DV_N_3261[18]), .I1(n294[21]), 
            .I2(VCC_net), .I3(n46146), .O(n23)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_23_lut.LUT_INIT = 16'hebbe;
    SB_LUT4 add_2547_15_lut (.I0(GND_net), .I1(n2355), .I2(n2397), .I3(n46377), 
            .O(n7624[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2547_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2547_15 (.CI(n46377), .I0(n2355), .I1(n2397), .CO(n46378));
    SB_LUT4 add_2547_14_lut (.I0(GND_net), .I1(n2356), .I2(n2272), .I3(n46376), 
            .O(n7624[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2547_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_i1663_3_lut (.I0(n2354), .I1(n7624[22]), .I2(n294[8]), 
            .I3(GND_net), .O(n2477));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1663_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY sub_38_add_2_23 (.CI(n46146), .I0(n294[21]), .I1(VCC_net), 
            .CO(n46147));
    SB_CARRY add_2547_14 (.CI(n46376), .I0(n2356), .I1(n2272), .CO(n46377));
    SB_LUT4 div_37_i1974_3_lut (.I0(n2827), .I1(n7728[23]), .I2(n294[4]), 
            .I3(GND_net), .O(n2938));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1974_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_2547_13_lut (.I0(GND_net), .I1(n2357), .I2(n2144), .I3(n46375), 
            .O(n7624[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2547_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2547_13 (.CI(n46375), .I0(n2357), .I1(n2144), .CO(n46376));
    SB_LUT4 sub_38_add_2_22_lut (.I0(n55706), .I1(n294[20]), .I2(VCC_net), 
            .I3(n46145), .O(n55708)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_22_lut.LUT_INIT = 16'hebbe;
    SB_LUT4 add_2547_12_lut (.I0(GND_net), .I1(n2358), .I2(n2013), .I3(n46374), 
            .O(n7624[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2547_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2547_12 (.CI(n46374), .I0(n2358), .I1(n2013), .CO(n46375));
    SB_CARRY sub_38_add_2_22 (.CI(n46145), .I0(n294[20]), .I1(VCC_net), 
            .CO(n46146));
    SB_LUT4 div_37_i1989_3_lut (.I0(n2842), .I1(n7728[8]), .I2(n294[4]), 
            .I3(GND_net), .O(n2953));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1989_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4012_4_lut (.I0(n959), .I1(baudrate[4]), .I2(n9283), .I3(n19010), 
            .O(n46_adj_4825));   // verilog/uart_rx.v(119[33:55])
    defparam i4012_4_lut.LUT_INIT = 16'hbbb2;
    SB_LUT4 div_37_i742_4_lut (.I0(n53648), .I1(n294[18]), .I2(n46_adj_4825), 
            .I3(baudrate[5]), .O(n1111));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i742_4_lut.LUT_INIT = 16'h9559;
    SB_LUT4 div_37_i2158_1_lut (.I0(baudrate[17]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n2867));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2158_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1_3_lut_4_lut_adj_952 (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[2]), 
            .I2(\r_Bit_Index[0] ), .I3(n4_adj_4821), .O(n55948));
    defparam i1_3_lut_4_lut_adj_952.LUT_INIT = 16'hfff7;
    SB_LUT4 div_37_i843_3_lut (.I0(n1111), .I1(n7390[23]), .I2(n294[17]), 
            .I3(GND_net), .O(n1261));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i843_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_2547_11_lut (.I0(GND_net), .I1(n2359), .I2(n1879), .I3(n46373), 
            .O(n7624[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2547_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_i1975_3_lut (.I0(n2828), .I1(n7728[22]), .I2(n294[4]), 
            .I3(GND_net), .O(n2939));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1975_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i942_3_lut (.I0(n1261), .I1(n7416[23]), .I2(n294[16]), 
            .I3(GND_net), .O(n1408));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i942_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1976_3_lut (.I0(n2829), .I1(n7728[21]), .I2(n294[4]), 
            .I3(GND_net), .O(n2940));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1976_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_2547_11 (.CI(n46373), .I0(n2359), .I1(n1879), .CO(n46374));
    SB_LUT4 add_2547_10_lut (.I0(GND_net), .I1(n2360), .I2(n1742), .I3(n46372), 
            .O(n7624[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2547_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_i1979_3_lut (.I0(n2832), .I1(n7728[18]), .I2(n294[4]), 
            .I3(GND_net), .O(n2943));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1979_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1997_i37_2_lut (.I0(n2943), .I1(baudrate[15]), 
            .I2(GND_net), .I3(GND_net), .O(n37_adj_4826));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1997_i37_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1039_3_lut (.I0(n1408), .I1(n7442[23]), .I2(n294[15]), 
            .I3(GND_net), .O(n1552));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1039_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2157_1_lut (.I0(baudrate[18]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n2977));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2157_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_37_i1977_3_lut (.I0(n2830), .I1(n7728[20]), .I2(n294[4]), 
            .I3(GND_net), .O(n2941));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1977_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_2547_10 (.CI(n46372), .I0(n2360), .I1(n1742), .CO(n46373));
    SB_LUT4 add_2547_9_lut (.I0(GND_net), .I1(n2361), .I2(n1602), .I3(n46371), 
            .O(n7624[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2547_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_LessThan_1997_i41_2_lut (.I0(n2941), .I1(baudrate[17]), 
            .I2(GND_net), .I3(GND_net), .O(n41_adj_4827));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1997_i41_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i47878_4_lut (.I0(n40_adj_4823), .I1(n36), .I2(n41_adj_4790), 
            .I3(n60459), .O(n62591));   // verilog/uart_rx.v(119[33:55])
    defparam i47878_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 sub_38_add_2_21_lut (.I0(n55704), .I1(n294[19]), .I2(VCC_net), 
            .I3(n46144), .O(n55706)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_21_lut.LUT_INIT = 16'hebbe;
    SB_LUT4 div_37_i1980_3_lut (.I0(n2833), .I1(n7728[17]), .I2(n294[4]), 
            .I3(GND_net), .O(n2944));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1980_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1134_3_lut (.I0(n1552), .I1(n7468[23]), .I2(n294[14]), 
            .I3(GND_net), .O(n1693));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1134_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1997_i35_2_lut (.I0(n2944), .I1(baudrate[14]), 
            .I2(GND_net), .I3(GND_net), .O(n35_adj_4828));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1997_i35_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY sub_38_add_2_21 (.CI(n46144), .I0(n294[19]), .I1(VCC_net), 
            .CO(n46145));
    SB_LUT4 i39206_1_lut (.I0(n22501), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n53871));
    defparam i39206_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_2547_9 (.CI(n46371), .I0(n2361), .I1(n1602), .CO(n46372));
    SB_LUT4 add_2547_8_lut (.I0(GND_net), .I1(n2362), .I2(n1459), .I3(n46370), 
            .O(n7624[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2547_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_i1978_3_lut (.I0(n2831), .I1(n7728[19]), .I2(n294[4]), 
            .I3(GND_net), .O(n2942));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1978_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1744_3_lut (.I0(n2477), .I1(n7650[22]), .I2(n294[7]), 
            .I3(GND_net), .O(n2597));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1744_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_2547_8 (.CI(n46370), .I0(n2362), .I1(n1459), .CO(n46371));
    SB_LUT4 div_37_LessThan_1997_i39_2_lut (.I0(n2942), .I1(baudrate[16]), 
            .I2(GND_net), .I3(GND_net), .O(n39_adj_4829));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1997_i39_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i2175_1_lut (.I0(baudrate[0]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n538));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2175_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_37_i1982_3_lut (.I0(n2835), .I1(n7728[15]), .I2(n294[4]), 
            .I3(GND_net), .O(n2946));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1982_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1983_3_lut (.I0(n2836), .I1(n7728[14]), .I2(n294[4]), 
            .I3(GND_net), .O(n2947));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1983_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1997_i29_2_lut (.I0(n2947), .I1(baudrate[11]), 
            .I2(GND_net), .I3(GND_net), .O(n29_adj_4830));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1997_i29_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1997_i31_2_lut (.I0(n2946), .I1(baudrate[12]), 
            .I2(GND_net), .I3(GND_net), .O(n31_adj_4831));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1997_i31_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1984_3_lut (.I0(n2837), .I1(n7728[13]), .I2(n294[4]), 
            .I3(GND_net), .O(n2948));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1984_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1985_3_lut (.I0(n2838), .I1(n7728[12]), .I2(n294[4]), 
            .I3(GND_net), .O(n2949));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1985_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1986_3_lut (.I0(n2839), .I1(n7728[11]), .I2(n294[4]), 
            .I3(GND_net), .O(n2950));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1986_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1997_i23_2_lut (.I0(n2950), .I1(baudrate[8]), 
            .I2(GND_net), .I3(GND_net), .O(n23_adj_4832));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1997_i23_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1997_i25_2_lut (.I0(n2949), .I1(baudrate[9]), 
            .I2(GND_net), .I3(GND_net), .O(n25_adj_4833));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1997_i25_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1997_i27_2_lut (.I0(n2948), .I1(baudrate[10]), 
            .I2(GND_net), .I3(GND_net), .O(n27_adj_4834));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1997_i27_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1990_3_lut (.I0(n2843), .I1(n7728[7]), .I2(n294[4]), 
            .I3(GND_net), .O(n2954));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1990_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1991_3_lut (.I0(n2844), .I1(n7728[6]), .I2(n294[4]), 
            .I3(GND_net), .O(n2955));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1991_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1992_3_lut (.I0(n2845), .I1(n7728[5]), .I2(n294[4]), 
            .I3(GND_net), .O(n2956));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1992_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1997_i13_2_lut (.I0(n2955), .I1(baudrate[3]), 
            .I2(GND_net), .I3(GND_net), .O(n13_adj_4835));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1997_i13_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1997_i15_2_lut (.I0(n2954), .I1(baudrate[4]), 
            .I2(GND_net), .I3(GND_net), .O(n15_adj_4836));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1997_i15_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1981_3_lut (.I0(n2834), .I1(n7728[16]), .I2(n294[4]), 
            .I3(GND_net), .O(n2945));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1981_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1988_3_lut (.I0(n2841), .I1(n7728[9]), .I2(n294[4]), 
            .I3(GND_net), .O(n2952));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1988_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1987_3_lut (.I0(n2840), .I1(n7728[10]), .I2(n294[4]), 
            .I3(GND_net), .O(n2951));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1987_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1997_i17_2_lut (.I0(n2953), .I1(baudrate[5]), 
            .I2(GND_net), .I3(GND_net), .O(n17_adj_4837));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1997_i17_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_2547_7_lut (.I0(GND_net), .I1(n2363), .I2(n1460), .I3(n46369), 
            .O(n7624[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2547_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2547_7 (.CI(n46369), .I0(n2363), .I1(n1460), .CO(n46370));
    SB_LUT4 sub_38_add_2_20_lut (.I0(GND_net), .I1(n294[18]), .I2(VCC_net), 
            .I3(n46143), .O(o_Rx_DV_N_3261[18])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2547_6_lut (.I0(GND_net), .I1(n2364), .I2(n1011), .I3(n46368), 
            .O(n7624[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2547_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2547_6 (.CI(n46368), .I0(n2364), .I1(n1011), .CO(n46369));
    SB_LUT4 div_37_LessThan_1997_i19_2_lut (.I0(n2952), .I1(baudrate[6]), 
            .I2(GND_net), .I3(GND_net), .O(n19_adj_4838));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1997_i19_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY sub_38_add_2_20 (.CI(n46143), .I0(n294[18]), .I1(VCC_net), 
            .CO(n46144));
    SB_LUT4 add_2547_5_lut (.I0(GND_net), .I1(n2365), .I2(n856), .I3(n46367), 
            .O(n7624[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2547_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_LessThan_1997_i21_2_lut (.I0(n2951), .I1(baudrate[7]), 
            .I2(GND_net), .I3(GND_net), .O(n21_adj_4839));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1997_i21_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_2547_5 (.CI(n46367), .I0(n2365), .I1(n856), .CO(n46368));
    SB_LUT4 div_37_LessThan_1997_i33_2_lut (.I0(n2945), .I1(baudrate[13]), 
            .I2(GND_net), .I3(GND_net), .O(n33_adj_4840));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1997_i33_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 sub_38_add_2_19_lut (.I0(n55702), .I1(n294[17]), .I2(VCC_net), 
            .I3(n46142), .O(n55704)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_19_lut.LUT_INIT = 16'hebbe;
    SB_LUT4 add_2547_4_lut (.I0(GND_net), .I1(n2366), .I2(n698), .I3(n46366), 
            .O(n7624[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2547_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_38_add_2_19 (.CI(n46142), .I0(n294[17]), .I1(VCC_net), 
            .CO(n46143));
    SB_CARRY add_2547_4 (.CI(n46366), .I0(n2366), .I1(n698), .CO(n46367));
    SB_LUT4 sub_38_add_2_18_lut (.I0(n55700), .I1(n294[16]), .I2(VCC_net), 
            .I3(n46141), .O(n55702)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_18_lut.LUT_INIT = 16'hebbe;
    SB_LUT4 add_2547_3_lut (.I0(GND_net), .I1(n2367), .I2(n858), .I3(n46365), 
            .O(n7624[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2547_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2547_3 (.CI(n46365), .I0(n2367), .I1(n858), .CO(n46366));
    SB_LUT4 add_2547_2_lut (.I0(n53887), .I1(GND_net), .I2(n538), .I3(VCC_net), 
            .O(n55682)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2547_2_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_2547_2 (.CI(VCC_net), .I0(GND_net), .I1(n538), .CO(n46365));
    SB_LUT4 add_2546_16_lut (.I0(GND_net), .I1(n2227), .I2(n2519), .I3(n46364), 
            .O(n7598[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2546_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_38_add_2_18 (.CI(n46141), .I0(n294[16]), .I1(VCC_net), 
            .CO(n46142));
    SB_LUT4 div_37_i1823_3_lut (.I0(n2597), .I1(n7676[22]), .I2(n294[6]), 
            .I3(GND_net), .O(n2714));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1823_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_adj_953 (.I0(baudrate[28]), .I1(baudrate[26]), .I2(GND_net), 
            .I3(GND_net), .O(n56428));
    defparam i1_2_lut_adj_953.LUT_INIT = 16'heeee;
    SB_LUT4 sub_38_add_2_17_lut (.I0(n55656), .I1(n294[15]), .I2(VCC_net), 
            .I3(n46140), .O(n55658)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_17_lut.LUT_INIT = 16'hebbe;
    SB_LUT4 add_2546_15_lut (.I0(GND_net), .I1(n2228), .I2(n2397), .I3(n46363), 
            .O(n7598[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2546_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2546_15 (.CI(n46363), .I0(n2228), .I1(n2397), .CO(n46364));
    SB_LUT4 add_2546_14_lut (.I0(GND_net), .I1(n2229), .I2(n2272), .I3(n46362), 
            .O(n7598[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2546_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2546_14 (.CI(n46362), .I0(n2229), .I1(n2272), .CO(n46363));
    SB_CARRY sub_38_add_2_17 (.CI(n46140), .I0(n294[15]), .I1(VCC_net), 
            .CO(n46141));
    SB_LUT4 i1_3_lut (.I0(baudrate[31]), .I1(baudrate[21]), .I2(baudrate[27]), 
            .I3(GND_net), .O(n56488));
    defparam i1_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 add_2546_13_lut (.I0(GND_net), .I1(n2230), .I2(n2144), .I3(n46361), 
            .O(n7598[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2546_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_4_lut_adj_954 (.I0(n56488), .I1(n56486), .I2(n56490), .I3(n56354), 
            .O(n22476));
    defparam i1_4_lut_adj_954.LUT_INIT = 16'hfffe;
    SB_LUT4 sub_38_add_2_16_lut (.I0(n55698), .I1(n294[14]), .I2(VCC_net), 
            .I3(n46139), .O(n55700)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_16_lut.LUT_INIT = 16'hebbe;
    SB_LUT4 i45928_4_lut (.I0(n33_adj_4840), .I1(n21_adj_4839), .I2(n19_adj_4838), 
            .I3(n17_adj_4837), .O(n60640));
    defparam i45928_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i46922_4_lut (.I0(n15_adj_4836), .I1(n13_adj_4835), .I2(n2956), 
            .I3(baudrate[2]), .O(n61635));
    defparam i46922_4_lut.LUT_INIT = 16'heffe;
    SB_LUT4 div_37_i2174_1_lut (.I0(baudrate[1]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n858));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2174_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i47371_4_lut (.I0(n21_adj_4839), .I1(n19_adj_4838), .I2(n17_adj_4837), 
            .I3(n61635), .O(n62084));
    defparam i47371_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i47367_4_lut (.I0(n27_adj_4834), .I1(n25_adj_4833), .I2(n23_adj_4832), 
            .I3(n62084), .O(n62080));
    defparam i47367_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i45934_4_lut (.I0(n33_adj_4840), .I1(n31_adj_4831), .I2(n29_adj_4830), 
            .I3(n62080), .O(n60646));
    defparam i45934_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 div_37_LessThan_1997_i10_3_lut (.I0(baudrate[0]), .I1(baudrate[1]), 
            .I2(n2957), .I3(GND_net), .O(n10_adj_4841));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1997_i10_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i47479_3_lut (.I0(n10_adj_4841), .I1(baudrate[13]), .I2(n33_adj_4840), 
            .I3(GND_net), .O(n62192));   // verilog/uart_rx.v(119[33:55])
    defparam i47479_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i47480_3_lut (.I0(n62192), .I1(baudrate[14]), .I2(n35_adj_4828), 
            .I3(GND_net), .O(n62193));   // verilog/uart_rx.v(119[33:55])
    defparam i47480_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1997_i36_3_lut (.I0(n18), .I1(baudrate[17]), 
            .I2(n41_adj_4827), .I3(GND_net), .O(n36_adj_4842));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1997_i36_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_2546_13 (.CI(n46361), .I0(n2230), .I1(n2144), .CO(n46362));
    SB_LUT4 div_37_i1227_3_lut (.I0(n1693), .I1(n7494[23]), .I2(n294[13]), 
            .I3(GND_net), .O(n1831));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1227_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_2546_12_lut (.I0(GND_net), .I1(n2231), .I2(n2013), .I3(n46360), 
            .O(n7598[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2546_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2546_12 (.CI(n46360), .I0(n2231), .I1(n2013), .CO(n46361));
    SB_LUT4 add_2546_11_lut (.I0(GND_net), .I1(n2232), .I2(n1879), .I3(n46359), 
            .O(n7598[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2546_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2546_11 (.CI(n46359), .I0(n2232), .I1(n1879), .CO(n46360));
    SB_LUT4 i45914_4_lut (.I0(n39_adj_4829), .I1(n37_adj_4826), .I2(n35_adj_4828), 
            .I3(n60640), .O(n60626));
    defparam i45914_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i47946_4_lut (.I0(n36_adj_4842), .I1(n16_adj_4843), .I2(n41_adj_4827), 
            .I3(n60618), .O(n62659));   // verilog/uart_rx.v(119[33:55])
    defparam i47946_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 add_2546_10_lut (.I0(GND_net), .I1(n2233), .I2(n1742), .I3(n46358), 
            .O(n7598[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2546_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2546_10 (.CI(n46358), .I0(n2233), .I1(n1742), .CO(n46359));
    SB_LUT4 add_2546_9_lut (.I0(GND_net), .I1(n2234), .I2(n1602), .I3(n46357), 
            .O(n7598[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2546_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2546_9 (.CI(n46357), .I0(n2234), .I1(n1602), .CO(n46358));
    SB_LUT4 i47879_3_lut (.I0(n62591), .I1(baudrate[5]), .I2(n1263), .I3(GND_net), 
            .O(n62592));   // verilog/uart_rx.v(119[33:55])
    defparam i47879_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i46595_3_lut (.I0(n62193), .I1(baudrate[15]), .I2(n37_adj_4826), 
            .I3(GND_net), .O(n61308));   // verilog/uart_rx.v(119[33:55])
    defparam i46595_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1318_3_lut (.I0(n1831), .I1(n7520[23]), .I2(n294[12]), 
            .I3(GND_net), .O(n1966));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1318_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY sub_38_add_2_16 (.CI(n46139), .I0(n294[14]), .I1(VCC_net), 
            .CO(n46140));
    SB_LUT4 add_2546_8_lut (.I0(GND_net), .I1(n2235), .I2(n1459), .I3(n46356), 
            .O(n7598[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2546_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2546_8 (.CI(n46356), .I0(n2235), .I1(n1459), .CO(n46357));
    SB_LUT4 add_2546_7_lut (.I0(GND_net), .I1(n2236), .I2(n1460), .I3(n46355), 
            .O(n7598[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2546_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_LessThan_1997_i22_3_lut (.I0(n14_adj_4844), .I1(baudrate[9]), 
            .I2(n25_adj_4833), .I3(GND_net), .O(n22));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1997_i22_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i47942_4_lut (.I0(n22), .I1(n12_adj_4845), .I2(n25_adj_4833), 
            .I3(n60675), .O(n62655));   // verilog/uart_rx.v(119[33:55])
    defparam i47942_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 sub_38_add_2_15_lut (.I0(o_Rx_DV_N_3261[10]), .I1(n294[13]), 
            .I2(VCC_net), .I3(n46138), .O(n55698)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_15_lut.LUT_INIT = 16'hebbe;
    SB_LUT4 i47943_3_lut (.I0(n62655), .I1(baudrate[10]), .I2(n27_adj_4834), 
            .I3(GND_net), .O(n62656));   // verilog/uart_rx.v(119[33:55])
    defparam i47943_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_2546_7 (.CI(n46355), .I0(n2236), .I1(n1460), .CO(n46356));
    SB_LUT4 add_2546_6_lut (.I0(GND_net), .I1(n2237), .I2(n1011), .I3(n46354), 
            .O(n7598[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2546_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_38_add_2_15 (.CI(n46138), .I0(n294[13]), .I1(VCC_net), 
            .CO(n46139));
    SB_LUT4 i47815_3_lut (.I0(n62656), .I1(baudrate[11]), .I2(n29_adj_4830), 
            .I3(GND_net), .O(n62528));   // verilog/uart_rx.v(119[33:55])
    defparam i47815_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i47748_4_lut (.I0(n39_adj_4829), .I1(n37_adj_4826), .I2(n35_adj_4828), 
            .I3(n60646), .O(n62461));
    defparam i47748_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i48197_4_lut (.I0(n61308), .I1(n62659), .I2(n41_adj_4827), 
            .I3(n60626), .O(n62910));   // verilog/uart_rx.v(119[33:55])
    defparam i48197_4_lut.LUT_INIT = 16'hccca;
    SB_CARRY add_2546_6 (.CI(n46354), .I0(n2237), .I1(n1011), .CO(n46355));
    SB_LUT4 add_2546_5_lut (.I0(GND_net), .I1(n2238), .I2(n856), .I3(n46353), 
            .O(n7598[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2546_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2546_5 (.CI(n46353), .I0(n2238), .I1(n856), .CO(n46354));
    SB_LUT4 add_2546_4_lut (.I0(GND_net), .I1(n2239), .I2(n698), .I3(n46352), 
            .O(n7598[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2546_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i46593_3_lut (.I0(n62528), .I1(baudrate[12]), .I2(n31_adj_4831), 
            .I3(GND_net), .O(n61306));   // verilog/uart_rx.v(119[33:55])
    defparam i46593_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_2546_4 (.CI(n46352), .I0(n2239), .I1(n698), .CO(n46353));
    SB_LUT4 add_2546_3_lut (.I0(GND_net), .I1(n2240), .I2(n858), .I3(n46351), 
            .O(n7598[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2546_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i48298_4_lut (.I0(n61306), .I1(n62910), .I2(n41_adj_4827), 
            .I3(n62461), .O(n63011));   // verilog/uart_rx.v(119[33:55])
    defparam i48298_4_lut.LUT_INIT = 16'hccca;
    SB_CARRY add_2546_3 (.CI(n46351), .I0(n2240), .I1(n858), .CO(n46352));
    SB_LUT4 i48299_3_lut (.I0(n63011), .I1(baudrate[18]), .I2(n2940), 
            .I3(GND_net), .O(n63012));   // verilog/uart_rx.v(119[33:55])
    defparam i48299_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 add_2546_2_lut (.I0(n53891), .I1(GND_net), .I2(n538), .I3(VCC_net), 
            .O(n55680)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2546_2_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i48291_3_lut (.I0(n63012), .I1(baudrate[19]), .I2(n2939), 
            .I3(GND_net), .O(n63004));   // verilog/uart_rx.v(119[33:55])
    defparam i48291_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_LessThan_1766_i37_2_lut (.I0(n2601), .I1(baudrate[12]), 
            .I2(GND_net), .I3(GND_net), .O(n37_adj_4846));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1766_i37_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1766_i43_2_lut (.I0(n2598), .I1(baudrate[15]), 
            .I2(GND_net), .I3(GND_net), .O(n43_adj_4847));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1766_i43_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i47855_3_lut (.I0(n62592), .I1(baudrate[6]), .I2(n1262), .I3(GND_net), 
            .O(n62568));   // verilog/uart_rx.v(119[33:55])
    defparam i47855_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_i1899_3_lut (.I0(n2713), .I1(n7702[23]), .I2(n294[5]), 
            .I3(GND_net), .O(n2827));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1899_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1766_i41_2_lut (.I0(n2599), .I1(baudrate[14]), 
            .I2(GND_net), .I3(GND_net), .O(n41_adj_4848));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1766_i41_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1407_3_lut (.I0(n1966), .I1(n7546[23]), .I2(n294[11]), 
            .I3(GND_net), .O(n2098));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1407_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1900_3_lut (.I0(n2714), .I1(n7702[22]), .I2(n294[5]), 
            .I3(GND_net), .O(n2828));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1900_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1903_3_lut (.I0(n2717), .I1(n7702[19]), .I2(n294[5]), 
            .I3(GND_net), .O(n2831));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1903_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1766_i39_2_lut (.I0(n2600), .I1(baudrate[13]), 
            .I2(GND_net), .I3(GND_net), .O(n39_adj_4849));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1766_i39_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1922_i39_2_lut (.I0(n2831), .I1(baudrate[15]), 
            .I2(GND_net), .I3(GND_net), .O(n39_adj_4850));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1922_i39_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1922_i37_2_lut (.I0(n2832), .I1(baudrate[14]), 
            .I2(GND_net), .I3(GND_net), .O(n37_adj_4851));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1922_i37_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1901_3_lut (.I0(n2715), .I1(n7702[21]), .I2(n294[5]), 
            .I3(GND_net), .O(n2829));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1901_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1922_i43_2_lut (.I0(n2829), .I1(baudrate[17]), 
            .I2(GND_net), .I3(GND_net), .O(n43_adj_4852));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1922_i43_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1766_i31_2_lut (.I0(n2604), .I1(baudrate[9]), 
            .I2(GND_net), .I3(GND_net), .O(n31_adj_4853));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1766_i31_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1902_3_lut (.I0(n2716), .I1(n7702[20]), .I2(n294[5]), 
            .I3(GND_net), .O(n2830));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1902_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1922_i41_2_lut (.I0(n2830), .I1(baudrate[16]), 
            .I2(GND_net), .I3(GND_net), .O(n41_adj_4854));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1922_i41_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1766_i33_2_lut (.I0(n2603), .I1(baudrate[10]), 
            .I2(GND_net), .I3(GND_net), .O(n33_adj_4855));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1766_i33_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1922_i31_2_lut (.I0(n2835), .I1(baudrate[11]), 
            .I2(GND_net), .I3(GND_net), .O(n31_adj_4856));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1922_i31_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1766_i35_2_lut (.I0(n2602), .I1(baudrate[11]), 
            .I2(GND_net), .I3(GND_net), .O(n35_adj_4857));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1766_i35_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1494_3_lut (.I0(n2098), .I1(n7572[23]), .I2(n294[10]), 
            .I3(GND_net), .O(n2227));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1494_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1845_i45_2_lut (.I0(n2714), .I1(baudrate[17]), 
            .I2(GND_net), .I3(GND_net), .O(n45_adj_4858));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1845_i45_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1922_i33_2_lut (.I0(n2834), .I1(baudrate[12]), 
            .I2(GND_net), .I3(GND_net), .O(n33_adj_4859));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1922_i33_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 sub_38_add_2_14_lut (.I0(GND_net), .I1(n294[12]), .I2(VCC_net), 
            .I3(n46137), .O(\o_Rx_DV_N_3261[12] )) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_LessThan_1922_i25_2_lut (.I0(n2838), .I1(baudrate[8]), 
            .I2(GND_net), .I3(GND_net), .O(n25_adj_4860));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1922_i25_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1766_i27_2_lut (.I0(n2606), .I1(baudrate[7]), 
            .I2(GND_net), .I3(GND_net), .O(n27_adj_4861));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1766_i27_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1766_i29_2_lut (.I0(n2605), .I1(baudrate[8]), 
            .I2(GND_net), .I3(GND_net), .O(n29_adj_4862));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1766_i29_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1922_i27_2_lut (.I0(n2837), .I1(baudrate[9]), 
            .I2(GND_net), .I3(GND_net), .O(n27_adj_4863));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1922_i27_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1766_i25_2_lut (.I0(n2607), .I1(baudrate[6]), 
            .I2(GND_net), .I3(GND_net), .O(n25_adj_4864));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1766_i25_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_2546_2 (.CI(VCC_net), .I0(GND_net), .I1(n538), .CO(n46351));
    SB_LUT4 add_2545_14_lut (.I0(GND_net), .I1(n2098), .I2(n2397), .I3(n46350), 
            .O(n7572[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2545_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_LessThan_1922_i29_2_lut (.I0(n2836), .I1(baudrate[10]), 
            .I2(GND_net), .I3(GND_net), .O(n29_adj_4865));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1922_i29_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1922_i15_2_lut (.I0(n2843), .I1(baudrate[3]), 
            .I2(GND_net), .I3(GND_net), .O(n15_adj_4866));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1922_i15_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_2545_13_lut (.I0(GND_net), .I1(n2099), .I2(n2272), .I3(n46349), 
            .O(n7572[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2545_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2545_13 (.CI(n46349), .I0(n2099), .I1(n2272), .CO(n46350));
    SB_LUT4 add_2545_12_lut (.I0(GND_net), .I1(n2100), .I2(n2144), .I3(n46348), 
            .O(n7572[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2545_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_i1579_3_lut (.I0(n2227), .I1(n7598[23]), .I2(n294[9]), 
            .I3(GND_net), .O(n2353));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1579_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY sub_38_add_2_14 (.CI(n46137), .I0(n294[12]), .I1(VCC_net), 
            .CO(n46138));
    SB_LUT4 div_37_LessThan_1602_i21_2_lut (.I0(n2366), .I1(baudrate[2]), 
            .I2(GND_net), .I3(GND_net), .O(n21_adj_4867));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1602_i21_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_2545_12 (.CI(n46348), .I0(n2100), .I1(n2144), .CO(n46349));
    SB_LUT4 i45404_4_lut (.I0(n27_adj_4868), .I1(n25_adj_4869), .I2(n23_adj_4870), 
            .I3(n21_adj_4867), .O(n60116));
    defparam i45404_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 add_2545_11_lut (.I0(GND_net), .I1(n2101), .I2(n2013), .I3(n46347), 
            .O(n7572[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2545_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_LessThan_1766_i19_2_lut (.I0(n2610), .I1(baudrate[3]), 
            .I2(GND_net), .I3(GND_net), .O(n19_adj_4871));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1766_i19_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_2545_11 (.CI(n46347), .I0(n2101), .I1(n2013), .CO(n46348));
    SB_LUT4 add_2545_10_lut (.I0(GND_net), .I1(n2102), .I2(n1879), .I3(n46346), 
            .O(n7572[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2545_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_38_add_2_13_lut (.I0(o_Rx_DV_N_3261[9]), .I1(n294[11]), 
            .I2(VCC_net), .I3(n46136), .O(n55656)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_13_lut.LUT_INIT = 16'hebbe;
    SB_LUT4 i45379_4_lut (.I0(n33_adj_4872), .I1(n31_adj_4873), .I2(n29_adj_4874), 
            .I3(n60116), .O(n60091));
    defparam i45379_4_lut.LUT_INIT = 16'haaab;
    SB_CARRY add_2545_10 (.CI(n46346), .I0(n2102), .I1(n1879), .CO(n46347));
    SB_LUT4 add_2545_9_lut (.I0(GND_net), .I1(n2103), .I2(n1742), .I3(n46345), 
            .O(n7572[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2545_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_i1046_3_lut (.I0(n1415), .I1(n7442[16]), .I2(n294[15]), 
            .I3(GND_net), .O(n1559));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1046_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_2545_9 (.CI(n46345), .I0(n2103), .I1(n1742), .CO(n46346));
    SB_LUT4 r_Clock_Count_1948_add_4_9_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[7]), .I3(n46645), .O(n1[7])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1948_add_4_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_38_add_2_13 (.CI(n46136), .I0(n294[11]), .I1(VCC_net), 
            .CO(n46137));
    SB_LUT4 div_37_i1141_3_lut (.I0(n1559), .I1(n7468[16]), .I2(n294[14]), 
            .I3(GND_net), .O(n1700));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1141_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 sub_38_add_2_12_lut (.I0(GND_net), .I1(n294[10]), .I2(VCC_net), 
            .I3(n46135), .O(o_Rx_DV_N_3261[10])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2545_8_lut (.I0(GND_net), .I1(n2104), .I2(n1602), .I3(n46344), 
            .O(n7572[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2545_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_38_add_2_12 (.CI(n46135), .I0(n294[10]), .I1(VCC_net), 
            .CO(n46136));
    SB_LUT4 r_Clock_Count_1948_add_4_8_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[6]), .I3(n46644), .O(n1[6])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1948_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_LessThan_1922_i17_2_lut (.I0(n2842), .I1(baudrate[4]), 
            .I2(GND_net), .I3(GND_net), .O(n17_adj_4875));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1922_i17_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1766_i21_2_lut (.I0(n2609), .I1(baudrate[4]), 
            .I2(GND_net), .I3(GND_net), .O(n21_adj_4876));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1766_i21_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1922_i19_2_lut (.I0(n2841), .I1(baudrate[5]), 
            .I2(GND_net), .I3(GND_net), .O(n19_adj_4877));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1922_i19_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1922_i21_2_lut (.I0(n2840), .I1(baudrate[6]), 
            .I2(GND_net), .I3(GND_net), .O(n21_adj_4878));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1922_i21_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1922_i23_2_lut (.I0(n2839), .I1(baudrate[7]), 
            .I2(GND_net), .I3(GND_net), .O(n23_adj_4879));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1922_i23_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_2545_8 (.CI(n46344), .I0(n2104), .I1(n1602), .CO(n46345));
    SB_LUT4 add_2545_7_lut (.I0(GND_net), .I1(n2105), .I2(n1459), .I3(n46343), 
            .O(n7572[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2545_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2545_7 (.CI(n46343), .I0(n2105), .I1(n1459), .CO(n46344));
    SB_CARRY r_Clock_Count_1948_add_4_8 (.CI(n46644), .I0(GND_net), .I1(r_Clock_Count[6]), 
            .CO(n46645));
    SB_LUT4 sub_38_add_2_11_lut (.I0(GND_net), .I1(n294[9]), .I2(VCC_net), 
            .I3(n46134), .O(o_Rx_DV_N_3261[9])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 r_Clock_Count_1948_add_4_7_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[5]), .I3(n46643), .O(n1[5])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1948_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_LessThan_1922_i35_2_lut (.I0(n2833), .I1(baudrate[13]), 
            .I2(GND_net), .I3(GND_net), .O(n35_adj_4880));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1922_i35_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i46018_4_lut (.I0(n35_adj_4880), .I1(n23_adj_4879), .I2(n21_adj_4878), 
            .I3(n19_adj_4877), .O(n60730));
    defparam i46018_4_lut.LUT_INIT = 16'haaab;
    SB_CARRY r_Clock_Count_1948_add_4_7 (.CI(n46643), .I0(GND_net), .I1(r_Clock_Count[5]), 
            .CO(n46644));
    SB_LUT4 i46998_4_lut (.I0(n17_adj_4875), .I1(n15_adj_4866), .I2(n2844), 
            .I3(baudrate[2]), .O(n61711));
    defparam i46998_4_lut.LUT_INIT = 16'heffe;
    SB_LUT4 div_37_i1234_3_lut (.I0(n1700), .I1(n7494[16]), .I2(n294[13]), 
            .I3(GND_net), .O(n1838));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1234_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i47407_4_lut (.I0(n23_adj_4879), .I1(n21_adj_4878), .I2(n19_adj_4877), 
            .I3(n61711), .O(n62120));
    defparam i47407_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 r_Clock_Count_1948_add_4_6_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[4]), .I3(n46642), .O(n1[4])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1948_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2545_6_lut (.I0(GND_net), .I1(n2106), .I2(n1460), .I3(n46342), 
            .O(n7572[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2545_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_1948_add_4_6 (.CI(n46642), .I0(GND_net), .I1(r_Clock_Count[4]), 
            .CO(n46643));
    SB_CARRY add_2545_6 (.CI(n46342), .I0(n2106), .I1(n1460), .CO(n46343));
    SB_LUT4 div_37_LessThan_1766_i23_2_lut (.I0(n2608), .I1(baudrate[5]), 
            .I2(GND_net), .I3(GND_net), .O(n23_adj_4881));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1766_i23_2_lut.LUT_INIT = 16'h6666;
    SB_DFF r_Rx_Byte_i2 (.Q(rx_data[2]), .C(clk16MHz), .D(n26445));   // verilog/uart_rx.v(50[10] 145[8])
    SB_LUT4 add_2545_5_lut (.I0(GND_net), .I1(n2107), .I2(n1011), .I3(n46341), 
            .O(n7572[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2545_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_38_add_2_11 (.CI(n46134), .I0(n294[9]), .I1(VCC_net), 
            .CO(n46135));
    SB_LUT4 r_Clock_Count_1948_add_4_5_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[3]), .I3(n46641), .O(n1[3])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1948_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i47403_4_lut (.I0(n29_adj_4865), .I1(n27_adj_4863), .I2(n25_adj_4860), 
            .I3(n62120), .O(n62116));
    defparam i47403_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 sub_38_add_2_10_lut (.I0(GND_net), .I1(n294[8]), .I2(VCC_net), 
            .I3(n46133), .O(\o_Rx_DV_N_3261[8] )) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_10_lut.LUT_INIT = 16'hC33C;
    SB_DFF r_Rx_Byte_i1 (.Q(rx_data[1]), .C(clk16MHz), .D(n26443));   // verilog/uart_rx.v(50[10] 145[8])
    SB_DFF r_SM_Main_i2 (.Q(\r_SM_Main[2] ), .C(clk16MHz), .D(n63689));   // verilog/uart_rx.v(50[10] 145[8])
    SB_LUT4 i46024_4_lut (.I0(n35_adj_4880), .I1(n33_adj_4859), .I2(n31_adj_4856), 
            .I3(n62116), .O(n60736));
    defparam i46024_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i3990_2_lut (.I0(n962), .I1(baudrate[1]), .I2(GND_net), .I3(GND_net), 
            .O(n40_adj_4882));   // verilog/uart_rx.v(119[33:55])
    defparam i3990_2_lut.LUT_INIT = 16'hbbbb;
    SB_CARRY sub_38_add_2_10 (.CI(n46133), .I0(n294[8]), .I1(VCC_net), 
            .CO(n46134));
    SB_LUT4 div_37_LessThan_1922_i12_3_lut (.I0(baudrate[0]), .I1(baudrate[1]), 
            .I2(n2845), .I3(GND_net), .O(n12_adj_4883));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1922_i12_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i47485_3_lut (.I0(n12_adj_4883), .I1(baudrate[13]), .I2(n35_adj_4880), 
            .I3(GND_net), .O(n62198));   // verilog/uart_rx.v(119[33:55])
    defparam i47485_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1766_i17_2_lut (.I0(n2611), .I1(baudrate[2]), 
            .I2(GND_net), .I3(GND_net), .O(n17_adj_4884));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1766_i17_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1602_i20_3_lut (.I0(baudrate[0]), .I1(baudrate[1]), 
            .I2(n2367), .I3(GND_net), .O(n20_adj_4885));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1602_i20_3_lut.LUT_INIT = 16'h8e8e;
    SB_CARRY r_Clock_Count_1948_add_4_5 (.CI(n46641), .I0(GND_net), .I1(r_Clock_Count[3]), 
            .CO(n46642));
    SB_LUT4 i45259_4_lut (.I0(n23_adj_4881), .I1(n21_adj_4876), .I2(n19_adj_4871), 
            .I3(n17_adj_4884), .O(n59971));
    defparam i45259_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i45247_4_lut (.I0(n29_adj_4862), .I1(n27_adj_4861), .I2(n25_adj_4864), 
            .I3(n59971), .O(n59959));
    defparam i45247_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 div_37_LessThan_1922_i38_3_lut (.I0(n20_adj_4886), .I1(baudrate[17]), 
            .I2(n43_adj_4852), .I3(GND_net), .O(n38_adj_4887));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1922_i38_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i47486_3_lut (.I0(n62198), .I1(baudrate[14]), .I2(n37_adj_4851), 
            .I3(GND_net), .O(n62199));   // verilog/uart_rx.v(119[33:55])
    defparam i47486_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i46002_4_lut (.I0(n41_adj_4854), .I1(n39_adj_4850), .I2(n37_adj_4851), 
            .I3(n60730), .O(n60714));
    defparam i46002_4_lut.LUT_INIT = 16'haaab;
    SB_CARRY add_2545_5 (.CI(n46341), .I0(n2107), .I1(n1011), .CO(n46342));
    SB_LUT4 i47451_4_lut (.I0(n35_adj_4857), .I1(n33_adj_4855), .I2(n31_adj_4853), 
            .I3(n59959), .O(n62164));
    defparam i47451_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i48050_4_lut (.I0(n38_adj_4887), .I1(n18_adj_4888), .I2(n43_adj_4852), 
            .I3(n60712), .O(n62763));   // verilog/uart_rx.v(119[33:55])
    defparam i48050_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 r_Clock_Count_1948_add_4_4_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[2]), .I3(n46640), .O(n1[2])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1948_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_1948_add_4_4 (.CI(n46640), .I0(GND_net), .I1(r_Clock_Count[2]), 
            .CO(n46641));
    SB_LUT4 sub_38_add_2_9_lut (.I0(GND_net), .I1(n294[7]), .I2(VCC_net), 
            .I3(n46132), .O(\o_Rx_DV_N_3261[7] )) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i46587_3_lut (.I0(n62199), .I1(baudrate[15]), .I2(n39_adj_4850), 
            .I3(GND_net), .O(n61300));   // verilog/uart_rx.v(119[33:55])
    defparam i46587_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 r_Clock_Count_1948_add_4_3_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[1]), .I3(n46639), .O(n1[1])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1948_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2545_4_lut (.I0(GND_net), .I1(n2108), .I2(n856), .I3(n46340), 
            .O(n7572[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2545_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_i1325_3_lut (.I0(n1838), .I1(n7520[16]), .I2(n294[12]), 
            .I3(GND_net), .O(n1973));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1325_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1766_i16_3_lut (.I0(baudrate[0]), .I1(baudrate[1]), 
            .I2(n2612), .I3(GND_net), .O(n16_adj_4889));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1766_i16_3_lut.LUT_INIT = 16'h8e8e;
    SB_CARRY r_Clock_Count_1948_add_4_3 (.CI(n46639), .I0(GND_net), .I1(r_Clock_Count[1]), 
            .CO(n46640));
    SB_LUT4 div_37_LessThan_1922_i24_3_lut (.I0(n16_adj_4890), .I1(baudrate[9]), 
            .I2(n27_adj_4863), .I3(GND_net), .O(n24_adj_4891));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1922_i24_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 r_Clock_Count_1948_add_4_2_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[0]), .I3(VCC_net), .O(n1[0])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1948_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2545_4 (.CI(n46340), .I0(n2108), .I1(n856), .CO(n46341));
    SB_LUT4 add_2545_3_lut (.I0(GND_net), .I1(n2109), .I2(n698), .I3(n46339), 
            .O(n7572[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2545_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2545_3 (.CI(n46339), .I0(n2109), .I1(n698), .CO(n46340));
    SB_LUT4 add_2545_2_lut (.I0(GND_net), .I1(n2110), .I2(n858), .I3(VCC_net), 
            .O(n7572[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2545_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_LessThan_1602_i28_3_lut (.I0(n26), .I1(baudrate[7]), 
            .I2(n31_adj_4873), .I3(GND_net), .O(n28));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1602_i28_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i47938_4_lut (.I0(n24_adj_4891), .I1(n14_adj_4892), .I2(n27_adj_4863), 
            .I3(n60755), .O(n62651));   // verilog/uart_rx.v(119[33:55])
    defparam i47938_4_lut.LUT_INIT = 16'haaac;
    SB_CARRY sub_38_add_2_9 (.CI(n46132), .I0(n294[7]), .I1(VCC_net), 
            .CO(n46133));
    SB_CARRY r_Clock_Count_1948_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(r_Clock_Count[0]), 
            .CO(n46639));
    SB_LUT4 i47939_3_lut (.I0(n62651), .I1(baudrate[10]), .I2(n29_adj_4865), 
            .I3(GND_net), .O(n62652));   // verilog/uart_rx.v(119[33:55])
    defparam i47939_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i47819_3_lut (.I0(n62652), .I1(baudrate[11]), .I2(n31_adj_4856), 
            .I3(GND_net), .O(n62532));   // verilog/uart_rx.v(119[33:55])
    defparam i47819_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_2545_2 (.CI(VCC_net), .I0(n2110), .I1(n858), .CO(n46339));
    SB_LUT4 i47764_4_lut (.I0(n41_adj_4854), .I1(n39_adj_4850), .I2(n37_adj_4851), 
            .I3(n60736), .O(n62477));
    defparam i47764_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 div_37_LessThan_1602_i32_3_lut (.I0(n24_adj_4893), .I1(baudrate[9]), 
            .I2(n35_adj_4894), .I3(GND_net), .O(n32_adj_4895));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1602_i32_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i48129_4_lut (.I0(n32_adj_4895), .I1(n22_adj_4896), .I2(n35_adj_4894), 
            .I3(n60085), .O(n62842));   // verilog/uart_rx.v(119[33:55])
    defparam i48129_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 add_2544_14_lut (.I0(GND_net), .I1(n1966), .I2(n2272), .I3(n46338), 
            .O(n7546[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2544_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2544_13_lut (.I0(GND_net), .I1(n1967), .I2(n2144), .I3(n46337), 
            .O(n7546[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2544_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2544_13 (.CI(n46337), .I0(n1967), .I1(n2144), .CO(n46338));
    SB_LUT4 add_2544_12_lut (.I0(GND_net), .I1(n1968), .I2(n2013), .I3(n46336), 
            .O(n7546[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2544_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_38_add_2_8_lut (.I0(GND_net), .I1(n294[6]), .I2(VCC_net), 
            .I3(n46131), .O(\o_Rx_DV_N_3261[6] )) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2544_12 (.CI(n46336), .I0(n1968), .I1(n2013), .CO(n46337));
    SB_LUT4 add_2544_11_lut (.I0(GND_net), .I1(n1969), .I2(n1879), .I3(n46335), 
            .O(n7546[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2544_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i48175_4_lut (.I0(n61300), .I1(n62763), .I2(n43_adj_4852), 
            .I3(n60714), .O(n62888));   // verilog/uart_rx.v(119[33:55])
    defparam i48175_4_lut.LUT_INIT = 16'hccca;
    SB_CARRY add_2544_11 (.CI(n46335), .I0(n1969), .I1(n1879), .CO(n46336));
    SB_LUT4 add_2544_10_lut (.I0(GND_net), .I1(n1970), .I2(n1742), .I3(n46334), 
            .O(n7546[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2544_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_38_add_2_8 (.CI(n46131), .I0(n294[6]), .I1(VCC_net), 
            .CO(n46132));
    SB_CARRY add_2544_10 (.CI(n46334), .I0(n1970), .I1(n1742), .CO(n46335));
    SB_LUT4 sub_38_add_2_7_lut (.I0(GND_net), .I1(n294[5]), .I2(VCC_net), 
            .I3(n46130), .O(\o_Rx_DV_N_3261[5] )) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2544_9_lut (.I0(GND_net), .I1(n1971), .I2(n1602), .I3(n46333), 
            .O(n7546[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2544_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i48130_3_lut (.I0(n62842), .I1(baudrate[10]), .I2(n37_adj_4897), 
            .I3(GND_net), .O(n62843));   // verilog/uart_rx.v(119[33:55])
    defparam i48130_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i48061_3_lut (.I0(n62843), .I1(baudrate[11]), .I2(n39_adj_4898), 
            .I3(GND_net), .O(n62774));   // verilog/uart_rx.v(119[33:55])
    defparam i48061_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_2544_9 (.CI(n46333), .I0(n1971), .I1(n1602), .CO(n46334));
    SB_LUT4 i47481_4_lut (.I0(n39_adj_4898), .I1(n37_adj_4897), .I2(n35_adj_4894), 
            .I3(n60091), .O(n62194));
    defparam i47481_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i46585_3_lut (.I0(n62532), .I1(baudrate[12]), .I2(n33_adj_4859), 
            .I3(GND_net), .O(n61298));   // verilog/uart_rx.v(119[33:55])
    defparam i46585_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i48286_4_lut (.I0(n61298), .I1(n62888), .I2(n43_adj_4852), 
            .I3(n62477), .O(n62999));   // verilog/uart_rx.v(119[33:55])
    defparam i48286_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i48287_3_lut (.I0(n62999), .I1(baudrate[18]), .I2(n2828), 
            .I3(GND_net), .O(n63000));   // verilog/uart_rx.v(119[33:55])
    defparam i48287_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i48131_4_lut (.I0(n28), .I1(n20_adj_4885), .I2(n31_adj_4873), 
            .I3(n60109), .O(n62844));   // verilog/uart_rx.v(119[33:55])
    defparam i48131_4_lut.LUT_INIT = 16'haaac;
    SB_CARRY sub_38_add_2_7 (.CI(n46130), .I0(n294[5]), .I1(VCC_net), 
            .CO(n46131));
    SB_LUT4 div_37_i745_4_lut (.I0(n961), .I1(n40_adj_4882), .I2(n294[18]), 
            .I3(baudrate[2]), .O(n1114));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i745_4_lut.LUT_INIT = 16'h6a9a;
    SB_LUT4 div_37_i846_3_lut (.I0(n1114), .I1(n7390[20]), .I2(n294[17]), 
            .I3(GND_net), .O(n1264));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i846_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i642_4_lut (.I0(n805), .I1(baudrate[1]), .I2(n294[19]), 
            .I3(baudrate[0]), .O(n961));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i642_4_lut.LUT_INIT = 16'h9a6a;
    SB_LUT4 i4_2_lut (.I0(baudrate[6]), .I1(baudrate[7]), .I2(GND_net), 
            .I3(GND_net), .O(n22_adj_4899));
    defparam i4_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i5_2_lut (.I0(baudrate[8]), .I1(baudrate[9]), .I2(GND_net), 
            .I3(GND_net), .O(n23_adj_4900));
    defparam i5_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i1_2_lut_adj_955 (.I0(baudrate[4]), .I1(baudrate[5]), .I2(GND_net), 
            .I3(GND_net), .O(n56292));
    defparam i1_2_lut_adj_955.LUT_INIT = 16'heeee;
    SB_LUT4 i1_2_lut_adj_956 (.I0(baudrate[28]), .I1(baudrate[31]), .I2(GND_net), 
            .I3(GND_net), .O(n56264));
    defparam i1_2_lut_adj_956.LUT_INIT = 16'heeee;
    SB_LUT4 i1_4_lut_adj_957 (.I0(n56264), .I1(n56274), .I2(n56376), .I3(n56456), 
            .O(n22501));
    defparam i1_4_lut_adj_957.LUT_INIT = 16'hfffe;
    SB_LUT4 i15_4_lut (.I0(n56292), .I1(n23_adj_4900), .I2(n22_adj_4899), 
            .I3(n24_adj_4901), .O(n33));
    defparam i15_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 div_37_LessThan_450_i46_4_lut (.I0(n59864), .I1(baudrate[2]), 
            .I2(n644), .I3(n48_adj_4774), .O(n46_adj_4903));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_450_i46_4_lut.LUT_INIT = 16'h0c8e;
    SB_LUT4 div_37_LessThan_450_i48_3_lut (.I0(n46_adj_4903), .I1(baudrate[3]), 
            .I2(n53644), .I3(GND_net), .O(n48_adj_4904));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_450_i48_3_lut.LUT_INIT = 16'he8e8;
    SB_LUT4 i1_4_lut_adj_958 (.I0(n33), .I1(n22501), .I2(n31_adj_4905), 
            .I3(n56416), .O(n22484));
    defparam i1_4_lut_adj_958.LUT_INIT = 16'hfffe;
    SB_LUT4 i21959_2_lut (.I0(baudrate[1]), .I1(baudrate[0]), .I2(GND_net), 
            .I3(GND_net), .O(n35471));
    defparam i21959_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1_3_lut_adj_959 (.I0(n22484), .I1(n48_adj_4904), .I2(baudrate[0]), 
            .I3(GND_net), .O(n805));
    defparam i1_3_lut_adj_959.LUT_INIT = 16'hefef;
    SB_LUT4 i21957_2_lut (.I0(baudrate[1]), .I1(baudrate[0]), .I2(GND_net), 
            .I3(GND_net), .O(n35469));
    defparam i21957_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i47511_3_lut (.I0(n16_adj_4889), .I1(baudrate[13]), .I2(n39_adj_4849), 
            .I3(GND_net), .O(n62224));   // verilog/uart_rx.v(119[33:55])
    defparam i47511_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i47512_3_lut (.I0(n62224), .I1(baudrate[14]), .I2(n41_adj_4848), 
            .I3(GND_net), .O(n62225));   // verilog/uart_rx.v(119[33:55])
    defparam i47512_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i47072_4_lut (.I0(n41_adj_4848), .I1(n39_adj_4849), .I2(n27_adj_4861), 
            .I3(n59963), .O(n61785));
    defparam i47072_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i47621_3_lut (.I0(n22_adj_4906), .I1(baudrate[7]), .I2(n27_adj_4861), 
            .I3(GND_net), .O(n62334));   // verilog/uart_rx.v(119[33:55])
    defparam i47621_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i46569_3_lut (.I0(n62225), .I1(baudrate[15]), .I2(n43_adj_4847), 
            .I3(GND_net), .O(n61282));   // verilog/uart_rx.v(119[33:55])
    defparam i46569_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1766_i28_3_lut (.I0(n20_adj_4907), .I1(baudrate[9]), 
            .I2(n31_adj_4853), .I3(GND_net), .O(n28_adj_4908));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1766_i28_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i48135_4_lut (.I0(n28_adj_4908), .I1(n18_adj_4909), .I2(n31_adj_4853), 
            .I3(n59955), .O(n62848));   // verilog/uart_rx.v(119[33:55])
    defparam i48135_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i48136_3_lut (.I0(n62848), .I1(baudrate[10]), .I2(n33_adj_4855), 
            .I3(GND_net), .O(n62849));   // verilog/uart_rx.v(119[33:55])
    defparam i48136_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i48053_3_lut (.I0(n62849), .I1(baudrate[11]), .I2(n35_adj_4857), 
            .I3(GND_net), .O(n62766));   // verilog/uart_rx.v(119[33:55])
    defparam i48053_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i46219_4_lut (.I0(n41_adj_4848), .I1(n39_adj_4849), .I2(n37_adj_4846), 
            .I3(n62164), .O(n60931));
    defparam i46219_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i47828_4_lut (.I0(n61282), .I1(n62334), .I2(n43_adj_4847), 
            .I3(n61785), .O(n62541));   // verilog/uart_rx.v(119[33:55])
    defparam i47828_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i47911_3_lut (.I0(n62766), .I1(baudrate[12]), .I2(n37_adj_4846), 
            .I3(GND_net), .O(n36_adj_4910));   // verilog/uart_rx.v(119[33:55])
    defparam i47911_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i48030_4_lut (.I0(n36_adj_4910), .I1(n62541), .I2(n43_adj_4847), 
            .I3(n60931), .O(n62743));   // verilog/uart_rx.v(119[33:55])
    defparam i48030_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i48031_3_lut (.I0(n62743), .I1(baudrate[16]), .I2(n2597), 
            .I3(GND_net), .O(n62744));   // verilog/uart_rx.v(119[33:55])
    defparam i48031_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_i2173_1_lut (.I0(baudrate[2]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n698));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2173_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_37_i1916_3_lut (.I0(n2730), .I1(n7702[6]), .I2(n294[5]), 
            .I3(GND_net), .O(n2844));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1916_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1685_i39_2_lut (.I0(n2480), .I1(baudrate[12]), 
            .I2(GND_net), .I3(GND_net), .O(n39_adj_4911));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1685_i39_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1685_i45_2_lut (.I0(n2477), .I1(baudrate[15]), 
            .I2(GND_net), .I3(GND_net), .O(n45_adj_4912));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1685_i45_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1685_i43_2_lut (.I0(n2478), .I1(baudrate[14]), 
            .I2(GND_net), .I3(GND_net), .O(n43_adj_4913));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1685_i43_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1685_i41_2_lut (.I0(n2479), .I1(baudrate[13]), 
            .I2(GND_net), .I3(GND_net), .O(n41_adj_4914));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1685_i41_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1685_i33_2_lut (.I0(n2483), .I1(baudrate[9]), 
            .I2(GND_net), .I3(GND_net), .O(n33_adj_4915));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1685_i33_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1685_i35_2_lut (.I0(n2482), .I1(baudrate[10]), 
            .I2(GND_net), .I3(GND_net), .O(n35_adj_4916));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1685_i35_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1685_i37_2_lut (.I0(n2481), .I1(baudrate[11]), 
            .I2(GND_net), .I3(GND_net), .O(n37_adj_4917));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1685_i37_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1685_i27_2_lut (.I0(n2486), .I1(baudrate[6]), 
            .I2(GND_net), .I3(GND_net), .O(n27_adj_4918));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1685_i27_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1685_i29_2_lut (.I0(n2485), .I1(baudrate[7]), 
            .I2(GND_net), .I3(GND_net), .O(n29_adj_4919));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1685_i29_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1685_i31_2_lut (.I0(n2484), .I1(baudrate[8]), 
            .I2(GND_net), .I3(GND_net), .O(n31_adj_4920));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1685_i31_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1685_i21_2_lut (.I0(n2489), .I1(baudrate[3]), 
            .I2(GND_net), .I3(GND_net), .O(n21_adj_4921));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1685_i21_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_2544_8_lut (.I0(GND_net), .I1(n1972), .I2(n1459), .I3(n46332), 
            .O(n7546[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2544_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2544_8 (.CI(n46332), .I0(n1972), .I1(n1459), .CO(n46333));
    SB_LUT4 add_2544_7_lut (.I0(GND_net), .I1(n1973), .I2(n1460), .I3(n46331), 
            .O(n7546[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2544_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2544_7 (.CI(n46331), .I0(n1973), .I1(n1460), .CO(n46332));
    SB_LUT4 sub_38_add_2_6_lut (.I0(GND_net), .I1(n294[4]), .I2(VCC_net), 
            .I3(n46129), .O(\o_Rx_DV_N_3261[4] )) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2544_6_lut (.I0(GND_net), .I1(n1974), .I2(n1011), .I3(n46330), 
            .O(n7546[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2544_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2544_6 (.CI(n46330), .I0(n1974), .I1(n1011), .CO(n46331));
    SB_LUT4 add_2544_5_lut (.I0(GND_net), .I1(n1975), .I2(n856), .I3(n46329), 
            .O(n7546[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2544_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_38_add_2_6 (.CI(n46129), .I0(n294[4]), .I1(VCC_net), 
            .CO(n46130));
    SB_CARRY add_2544_5 (.CI(n46329), .I0(n1975), .I1(n856), .CO(n46330));
    SB_LUT4 sub_38_add_2_5_lut (.I0(GND_net), .I1(n294[3]), .I2(VCC_net), 
            .I3(n46128), .O(\o_Rx_DV_N_3261[3] )) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2544_4_lut (.I0(GND_net), .I1(n1976), .I2(n698), .I3(n46328), 
            .O(n7546[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2544_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2544_4 (.CI(n46328), .I0(n1976), .I1(n698), .CO(n46329));
    SB_LUT4 add_2544_3_lut (.I0(GND_net), .I1(n1977), .I2(n858), .I3(n46327), 
            .O(n7546[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2544_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2544_3 (.CI(n46327), .I0(n1977), .I1(n858), .CO(n46328));
    SB_LUT4 add_2544_2_lut (.I0(GND_net), .I1(GND_net), .I2(n538), .I3(VCC_net), 
            .O(n7546[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2544_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_38_add_2_5 (.CI(n46128), .I0(n294[3]), .I1(VCC_net), 
            .CO(n46129));
    SB_CARRY add_2544_2 (.CI(VCC_net), .I0(GND_net), .I1(n538), .CO(n46327));
    SB_LUT4 sub_38_add_2_4_lut (.I0(GND_net), .I1(n294[2]), .I2(VCC_net), 
            .I3(n46127), .O(\o_Rx_DV_N_3261[2] )) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2543_13_lut (.I0(GND_net), .I1(n1831), .I2(n2144), .I3(n46326), 
            .O(n7520[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2543_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2543_12_lut (.I0(GND_net), .I1(n1832), .I2(n2013), .I3(n46325), 
            .O(n7520[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2543_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2543_12 (.CI(n46325), .I0(n1832), .I1(n2013), .CO(n46326));
    SB_LUT4 add_2543_11_lut (.I0(GND_net), .I1(n1833), .I2(n1879), .I3(n46324), 
            .O(n7520[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2543_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2543_11 (.CI(n46324), .I0(n1833), .I1(n1879), .CO(n46325));
    SB_LUT4 i5705_4_lut (.I0(n961), .I1(baudrate[2]), .I2(n962), .I3(baudrate[1]), 
            .O(n19008));   // verilog/uart_rx.v(119[33:55])
    defparam i5705_4_lut.LUT_INIT = 16'ha2aa;
    SB_LUT4 div_37_LessThan_1685_i23_2_lut (.I0(n2488), .I1(baudrate[4]), 
            .I2(GND_net), .I3(GND_net), .O(n23_adj_4922));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1685_i23_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY sub_38_add_2_4 (.CI(n46127), .I0(n294[2]), .I1(VCC_net), 
            .CO(n46128));
    SB_LUT4 sub_38_add_2_3_lut (.I0(GND_net), .I1(n294[1]), .I2(VCC_net), 
            .I3(n46126), .O(\o_Rx_DV_N_3261[1] )) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_38_add_2_3 (.CI(n46126), .I0(n294[1]), .I1(VCC_net), 
            .CO(n46127));
    SB_LUT4 add_2543_10_lut (.I0(GND_net), .I1(n1834), .I2(n1742), .I3(n46323), 
            .O(n7520[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2543_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2543_10 (.CI(n46323), .I0(n1834), .I1(n1742), .CO(n46324));
    SB_LUT4 add_2543_9_lut (.I0(GND_net), .I1(n1835), .I2(n1602), .I3(n46322), 
            .O(n7520[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2543_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_38_add_2_2_lut (.I0(GND_net), .I1(n54733), .I2(GND_net), 
            .I3(VCC_net), .O(\o_Rx_DV_N_3261[0] )) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2543_9 (.CI(n46322), .I0(n1835), .I1(n1602), .CO(n46323));
    SB_LUT4 add_2543_8_lut (.I0(GND_net), .I1(n1836), .I2(n1459), .I3(n46321), 
            .O(n7520[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2543_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2543_8 (.CI(n46321), .I0(n1836), .I1(n1459), .CO(n46322));
    SB_CARRY sub_38_add_2_2 (.CI(VCC_net), .I0(n54733), .I1(GND_net), 
            .CO(n46126));
    SB_LUT4 add_2543_7_lut (.I0(GND_net), .I1(n1837), .I2(n1460), .I3(n46320), 
            .O(n7520[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2543_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2543_7 (.CI(n46320), .I0(n1837), .I1(n1460), .CO(n46321));
    SB_LUT4 add_2543_6_lut (.I0(GND_net), .I1(n1838), .I2(n1011), .I3(n46319), 
            .O(n7520[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2543_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2543_6 (.CI(n46319), .I0(n1838), .I1(n1011), .CO(n46320));
    SB_LUT4 add_2543_5_lut (.I0(GND_net), .I1(n1839), .I2(n856), .I3(n46318), 
            .O(n7520[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2543_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_i1414_3_lut (.I0(n1973), .I1(n7546[16]), .I2(n294[11]), 
            .I3(GND_net), .O(n2105));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1414_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_2543_5 (.CI(n46318), .I0(n1839), .I1(n856), .CO(n46319));
    SB_LUT4 add_2543_4_lut (.I0(GND_net), .I1(n1840), .I2(n698), .I3(n46317), 
            .O(n7520[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2543_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2543_4 (.CI(n46317), .I0(n1840), .I1(n698), .CO(n46318));
    SB_LUT4 div_37_i1501_3_lut (.I0(n2105), .I1(n7572[16]), .I2(n294[10]), 
            .I3(GND_net), .O(n2234));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1501_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1685_i25_2_lut (.I0(n2487), .I1(baudrate[5]), 
            .I2(GND_net), .I3(GND_net), .O(n25_adj_4923));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1685_i25_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_2543_3_lut (.I0(GND_net), .I1(n1841), .I2(n858), .I3(n46316), 
            .O(n7520[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2543_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_i1586_3_lut (.I0(n2234), .I1(n7598[16]), .I2(n294[9]), 
            .I3(GND_net), .O(n2360));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1586_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_2543_3 (.CI(n46316), .I0(n1841), .I1(n858), .CO(n46317));
    SB_LUT4 add_2543_2_lut (.I0(n53900), .I1(GND_net), .I2(n538), .I3(VCC_net), 
            .O(n55678)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2543_2_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_2543_2 (.CI(VCC_net), .I0(GND_net), .I1(n538), .CO(n46316));
    SB_LUT4 add_2542_11_lut (.I0(GND_net), .I1(n1693), .I2(n2013), .I3(n46315), 
            .O(n7494[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2542_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2542_10_lut (.I0(GND_net), .I1(n1694), .I2(n1879), .I3(n46314), 
            .O(n7494[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2542_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2542_10 (.CI(n46314), .I0(n1694), .I1(n1879), .CO(n46315));
    SB_LUT4 add_2542_9_lut (.I0(GND_net), .I1(n1695), .I2(n1742), .I3(n46313), 
            .O(n7494[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2542_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2542_9 (.CI(n46313), .I0(n1695), .I1(n1742), .CO(n46314));
    SB_LUT4 add_2542_8_lut (.I0(GND_net), .I1(n1696), .I2(n1602), .I3(n46312), 
            .O(n7494[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2542_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_i1669_3_lut (.I0(n2360), .I1(n7624[16]), .I2(n294[8]), 
            .I3(GND_net), .O(n2483));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1669_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i47899_3_lut (.I0(n62774), .I1(baudrate[12]), .I2(n41_adj_4924), 
            .I3(GND_net), .O(n62612));   // verilog/uart_rx.v(119[33:55])
    defparam i47899_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_2542_8 (.CI(n46312), .I0(n1696), .I1(n1602), .CO(n46313));
    SB_LUT4 add_2542_7_lut (.I0(GND_net), .I1(n1697), .I2(n1459), .I3(n46311), 
            .O(n7494[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2542_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2542_7 (.CI(n46311), .I0(n1697), .I1(n1459), .CO(n46312));
    SB_LUT4 add_2542_6_lut (.I0(GND_net), .I1(n1698), .I2(n1460), .I3(n46310), 
            .O(n7494[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2542_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2542_6 (.CI(n46310), .I0(n1698), .I1(n1460), .CO(n46311));
    SB_LUT4 add_2542_5_lut (.I0(GND_net), .I1(n1699), .I2(n1011), .I3(n46309), 
            .O(n7494[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2542_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2542_5 (.CI(n46309), .I0(n1699), .I1(n1011), .CO(n46310));
    SB_LUT4 add_2542_4_lut (.I0(GND_net), .I1(n1700), .I2(n856), .I3(n46308), 
            .O(n7494[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2542_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2542_4 (.CI(n46308), .I0(n1700), .I1(n856), .CO(n46309));
    SB_LUT4 div_37_i1750_3_lut (.I0(n2483), .I1(n7650[16]), .I2(n294[7]), 
            .I3(GND_net), .O(n2603));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1750_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1685_i19_2_lut (.I0(n2490), .I1(baudrate[2]), 
            .I2(GND_net), .I3(GND_net), .O(n19_adj_4925));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1685_i19_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i48191_4_lut (.I0(n62612), .I1(n62844), .I2(n41_adj_4924), 
            .I3(n62194), .O(n62904));   // verilog/uart_rx.v(119[33:55])
    defparam i48191_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 div_37_i1829_3_lut (.I0(n2603), .I1(n7676[16]), .I2(n294[6]), 
            .I3(GND_net), .O(n2720));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1829_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i45316_4_lut (.I0(n25_adj_4923), .I1(n23_adj_4922), .I2(n21_adj_4921), 
            .I3(n19_adj_4925), .O(n60028));
    defparam i45316_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i45300_4_lut (.I0(n31_adj_4920), .I1(n29_adj_4919), .I2(n27_adj_4918), 
            .I3(n60028), .O(n60012));
    defparam i45300_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i47461_4_lut (.I0(n37_adj_4917), .I1(n35_adj_4916), .I2(n33_adj_4915), 
            .I3(n60012), .O(n62174));
    defparam i47461_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 add_2542_3_lut (.I0(GND_net), .I1(n1701), .I2(n698), .I3(n46307), 
            .O(n7494[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2542_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_LessThan_1685_i18_3_lut (.I0(baudrate[0]), .I1(baudrate[1]), 
            .I2(n2491), .I3(GND_net), .O(n18_adj_4926));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1685_i18_3_lut.LUT_INIT = 16'h8e8e;
    SB_CARRY add_2542_3 (.CI(n46307), .I0(n1701), .I1(n698), .CO(n46308));
    SB_LUT4 add_2542_2_lut (.I0(GND_net), .I1(n1702), .I2(n858), .I3(VCC_net), 
            .O(n7494[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2542_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2542_2 (.CI(VCC_net), .I0(n1702), .I1(n858), .CO(n46307));
    SB_LUT4 i47693_3_lut (.I0(n18_adj_4926), .I1(baudrate[13]), .I2(n41_adj_4914), 
            .I3(GND_net), .O(n62406));   // verilog/uart_rx.v(119[33:55])
    defparam i47693_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i47694_3_lut (.I0(n62406), .I1(baudrate[14]), .I2(n43_adj_4913), 
            .I3(GND_net), .O(n62407));   // verilog/uart_rx.v(119[33:55])
    defparam i47694_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i46267_4_lut (.I0(n43_adj_4913), .I1(n41_adj_4914), .I2(n29_adj_4919), 
            .I3(n60021), .O(n60979));
    defparam i46267_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 add_2541_11_lut (.I0(GND_net), .I1(n1552), .I2(n1879), .I3(n46306), 
            .O(n7468[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2541_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_LessThan_1845_i33_2_lut (.I0(n2720), .I1(baudrate[11]), 
            .I2(GND_net), .I3(GND_net), .O(n33_adj_4927));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1845_i33_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1685_i26_3_lut (.I0(n24_adj_4928), .I1(baudrate[7]), 
            .I2(n29_adj_4919), .I3(GND_net), .O(n26_adj_4929));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1685_i26_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF r_Rx_Byte_i6 (.Q(rx_data[6]), .C(clk16MHz), .D(n27051));   // verilog/uart_rx.v(50[10] 145[8])
    SB_LUT4 div_37_LessThan_341_i48_4_lut (.I0(n56818), .I1(baudrate[2]), 
            .I2(n54397), .I3(n35471), .O(n48_adj_4774));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_341_i48_4_lut.LUT_INIT = 16'hd4c0;
    SB_LUT4 i47616_3_lut (.I0(n62407), .I1(baudrate[15]), .I2(n45_adj_4912), 
            .I3(GND_net), .O(n42_adj_4930));   // verilog/uart_rx.v(119[33:55])
    defparam i47616_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_2541_10_lut (.I0(GND_net), .I1(n1553), .I2(n1742), .I3(n46305), 
            .O(n7468[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2541_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2541_10 (.CI(n46305), .I0(n1553), .I1(n1742), .CO(n46306));
    SB_LUT4 add_2541_9_lut (.I0(GND_net), .I1(n1554), .I2(n1602), .I3(n46304), 
            .O(n7468[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2541_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2541_9 (.CI(n46304), .I0(n1554), .I1(n1602), .CO(n46305));
    SB_LUT4 add_2541_8_lut (.I0(GND_net), .I1(n1555), .I2(n1459), .I3(n46303), 
            .O(n7468[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2541_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i5_3_lut (.I0(r_SM_Main[0]), .I1(\o_Rx_DV_N_3261[24] ), .I2(n27), 
            .I3(GND_net), .O(n14_adj_4931));
    defparam i5_3_lut.LUT_INIT = 16'h0202;
    SB_DFF r_Rx_Byte_i5 (.Q(rx_data[5]), .C(clk16MHz), .D(n26970));   // verilog/uart_rx.v(50[10] 145[8])
    SB_LUT4 i6_4_lut (.I0(n29), .I1(\o_Rx_DV_N_3261[12] ), .I2(n23), .I3(n4834), 
            .O(n15_adj_4932));
    defparam i6_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 i8_4_lut (.I0(n15_adj_4932), .I1(\o_Rx_DV_N_3261[8] ), .I2(n14_adj_4931), 
            .I3(n52823), .O(n63689));
    defparam i8_4_lut.LUT_INIT = 16'h2000;
    SB_LUT4 i1_4_lut_adj_960 (.I0(baudrate[11]), .I1(n56176), .I2(n56710), 
            .I3(baudrate[12]), .O(n56184));
    defparam i1_4_lut_adj_960.LUT_INIT = 16'hfffe;
    SB_CARRY add_2541_8 (.CI(n46303), .I0(n1555), .I1(n1459), .CO(n46304));
    SB_LUT4 add_2541_7_lut (.I0(GND_net), .I1(n1556), .I2(n1460), .I3(n46302), 
            .O(n7468[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2541_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_LessThan_1685_i30_3_lut (.I0(n22_adj_4933), .I1(baudrate[9]), 
            .I2(n33_adj_4915), .I3(GND_net), .O(n30_adj_4934));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1685_i30_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_2541_7 (.CI(n46302), .I0(n1556), .I1(n1460), .CO(n46303));
    SB_LUT4 add_2541_6_lut (.I0(GND_net), .I1(n1557), .I2(n1011), .I3(n46301), 
            .O(n7468[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2541_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i48133_4_lut (.I0(n30_adj_4934), .I1(n20_adj_4935), .I2(n33_adj_4915), 
            .I3(n60008), .O(n62846));   // verilog/uart_rx.v(119[33:55])
    defparam i48133_4_lut.LUT_INIT = 16'haaac;
    SB_CARRY add_2541_6 (.CI(n46301), .I0(n1557), .I1(n1011), .CO(n46302));
    SB_LUT4 add_2541_5_lut (.I0(GND_net), .I1(n1558), .I2(n856), .I3(n46300), 
            .O(n7468[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2541_5_lut.LUT_INIT = 16'hC33C;
    SB_DFF r_Rx_Byte_i0 (.Q(rx_data[0]), .C(clk16MHz), .D(n26836));   // verilog/uart_rx.v(50[10] 145[8])
    SB_DFFE r_Rx_DV_58 (.Q(rx_data_ready), .C(clk16MHz), .E(VCC_net), 
            .D(n48959));   // verilog/uart_rx.v(50[10] 145[8])
    SB_DFFE r_Bit_Index_i0 (.Q(\r_Bit_Index[0] ), .C(clk16MHz), .E(VCC_net), 
            .D(n26832));   // verilog/uart_rx.v(50[10] 145[8])
    SB_LUT4 i42090_1_lut (.I0(n56792), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n53900));
    defparam i42090_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_2541_5 (.CI(n46300), .I0(n1558), .I1(n856), .CO(n46301));
    SB_LUT4 add_2541_4_lut (.I0(GND_net), .I1(n1559), .I2(n698), .I3(n46299), 
            .O(n7468[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2541_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2541_4 (.CI(n46299), .I0(n1559), .I1(n698), .CO(n46300));
    SB_LUT4 add_2541_3_lut (.I0(GND_net), .I1(n1560), .I2(n858), .I3(n46298), 
            .O(n7468[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2541_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i48134_3_lut (.I0(n62846), .I1(baudrate[10]), .I2(n35_adj_4916), 
            .I3(GND_net), .O(n62847));   // verilog/uart_rx.v(119[33:55])
    defparam i48134_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_2541_3 (.CI(n46298), .I0(n1560), .I1(n858), .CO(n46299));
    SB_LUT4 add_2541_2_lut (.I0(GND_net), .I1(GND_net), .I2(n538), .I3(VCC_net), 
            .O(n7468[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2541_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2541_2 (.CI(VCC_net), .I0(GND_net), .I1(n538), .CO(n46298));
    SB_LUT4 add_2540_10_lut (.I0(GND_net), .I1(n1408), .I2(n1742), .I3(n46297), 
            .O(n7442[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2540_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i48055_3_lut (.I0(n62847), .I1(baudrate[11]), .I2(n37_adj_4917), 
            .I3(GND_net), .O(n62768));   // verilog/uart_rx.v(119[33:55])
    defparam i48055_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i46271_4_lut (.I0(n43_adj_4913), .I1(n41_adj_4914), .I2(n39_adj_4911), 
            .I3(n62174), .O(n60983));
    defparam i46271_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 add_2540_9_lut (.I0(GND_net), .I1(n1409), .I2(n1602), .I3(n46296), 
            .O(n7442[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2540_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i47222_4_lut (.I0(n42_adj_4930), .I1(n26_adj_4929), .I2(n45_adj_4912), 
            .I3(n60979), .O(n61935));   // verilog/uart_rx.v(119[33:55])
    defparam i47222_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i47907_3_lut (.I0(n62768), .I1(baudrate[12]), .I2(n39_adj_4911), 
            .I3(GND_net), .O(n62620));   // verilog/uart_rx.v(119[33:55])
    defparam i47907_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i47224_4_lut (.I0(n62620), .I1(n61935), .I2(n45_adj_4912), 
            .I3(n60983), .O(n61937));   // verilog/uart_rx.v(119[33:55])
    defparam i47224_4_lut.LUT_INIT = 16'hccca;
    SB_CARRY add_2540_9 (.CI(n46296), .I0(n1409), .I1(n1602), .CO(n46297));
    SB_LUT4 add_2540_8_lut (.I0(GND_net), .I1(n1410), .I2(n1459), .I3(n46295), 
            .O(n7442[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2540_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2540_8 (.CI(n46295), .I0(n1410), .I1(n1459), .CO(n46296));
    SB_LUT4 add_2540_7_lut (.I0(GND_net), .I1(n1411), .I2(n1460), .I3(n46294), 
            .O(n7442[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2540_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i48192_3_lut (.I0(n62904), .I1(baudrate[13]), .I2(n2355), 
            .I3(GND_net), .O(n62905));   // verilog/uart_rx.v(119[33:55])
    defparam i48192_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i48155_3_lut (.I0(n62905), .I1(baudrate[14]), .I2(n2354), 
            .I3(GND_net), .O(n62868));   // verilog/uart_rx.v(119[33:55])
    defparam i48155_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i1_4_lut_adj_961 (.I0(n56182), .I1(n22498), .I2(n56184), .I3(n56180), 
            .O(n22504));
    defparam i1_4_lut_adj_961.LUT_INIT = 16'hfffe;
    SB_LUT4 div_37_i1758_3_lut (.I0(n2491), .I1(n7650[8]), .I2(n294[7]), 
            .I3(GND_net), .O(n2611));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1758_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_adj_962 (.I0(baudrate[25]), .I1(baudrate[31]), .I2(GND_net), 
            .I3(GND_net), .O(n56430));
    defparam i1_2_lut_adj_962.LUT_INIT = 16'heeee;
    SB_LUT4 div_37_i1837_3_lut (.I0(n2611), .I1(n7676[8]), .I2(n294[6]), 
            .I3(GND_net), .O(n2728));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1837_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1845_i17_2_lut (.I0(n2728), .I1(baudrate[3]), 
            .I2(GND_net), .I3(GND_net), .O(n17_adj_4936));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1845_i17_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1845_i19_2_lut (.I0(n2727), .I1(baudrate[4]), 
            .I2(GND_net), .I3(GND_net), .O(n19_adj_4937));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1845_i19_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1845_i27_2_lut (.I0(n2723), .I1(baudrate[8]), 
            .I2(GND_net), .I3(GND_net), .O(n27_adj_4938));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1845_i27_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_4_lut_adj_963 (.I0(n56470), .I1(n56156), .I2(n56308), .I3(baudrate[19]), 
            .O(n22498));
    defparam i1_4_lut_adj_963.LUT_INIT = 16'hfffe;
    SB_LUT4 i46105_4_lut (.I0(n37_adj_4939), .I1(n25_adj_4940), .I2(n23_adj_4941), 
            .I3(n21_adj_4942), .O(n60817));
    defparam i46105_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i47054_4_lut (.I0(n19_adj_4937), .I1(n17_adj_4936), .I2(n2729), 
            .I3(baudrate[2]), .O(n61767));
    defparam i47054_4_lut.LUT_INIT = 16'heffe;
    SB_LUT4 i47435_4_lut (.I0(n25_adj_4940), .I1(n23_adj_4941), .I2(n21_adj_4942), 
            .I3(n61767), .O(n62148));
    defparam i47435_4_lut.LUT_INIT = 16'hfeff;
    SB_CARRY add_2540_7 (.CI(n46294), .I0(n1411), .I1(n1460), .CO(n46295));
    SB_LUT4 add_2540_6_lut (.I0(GND_net), .I1(n1412), .I2(n1011), .I3(n46293), 
            .O(n7442[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2540_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_LessThan_2210_i41_4_lut (.I0(n3154), .I1(baudrate[20]), 
            .I2(n7806[20]), .I3(n294[1]), .O(n41));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i41_4_lut.LUT_INIT = 16'h3c66;
    SB_LUT4 i47431_4_lut (.I0(n31_adj_4943), .I1(n29_adj_4944), .I2(n27_adj_4938), 
            .I3(n62148), .O(n62144));
    defparam i47431_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 div_37_LessThan_2210_i39_4_lut (.I0(n3155), .I1(baudrate[19]), 
            .I2(n7806[19]), .I3(n294[1]), .O(n39));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i39_4_lut.LUT_INIT = 16'h3c66;
    SB_LUT4 i46107_4_lut (.I0(n37_adj_4939), .I1(n35_adj_4945), .I2(n33_adj_4927), 
            .I3(n62144), .O(n60819));
    defparam i46107_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 div_37_LessThan_2210_i37_4_lut (.I0(n3156), .I1(baudrate[18]), 
            .I2(n7806[18]), .I3(n294[1]), .O(n37));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i37_4_lut.LUT_INIT = 16'h3c66;
    SB_LUT4 i46063_4_lut (.I0(n22504), .I1(n60180), .I2(n48_adj_4774), 
            .I3(baudrate[0]), .O(n804));
    defparam i46063_4_lut.LUT_INIT = 16'h3633;
    SB_LUT4 div_37_LessThan_2210_i29_4_lut (.I0(n3160), .I1(baudrate[14]), 
            .I2(n7806[14]), .I3(n294[1]), .O(n29_c));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i29_4_lut.LUT_INIT = 16'h3c66;
    SB_LUT4 div_37_LessThan_2210_i31_4_lut (.I0(n3159), .I1(baudrate[15]), 
            .I2(n7806[15]), .I3(n294[1]), .O(n31));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i31_4_lut.LUT_INIT = 16'h3c66;
    SB_LUT4 div_37_LessThan_2210_i23_4_lut (.I0(n3163), .I1(baudrate[11]), 
            .I2(n7806[11]), .I3(n294[1]), .O(n23_c));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i23_4_lut.LUT_INIT = 16'h3c66;
    SB_LUT4 div_37_LessThan_2210_i25_4_lut (.I0(n3162), .I1(baudrate[12]), 
            .I2(n7806[12]), .I3(n294[1]), .O(n25));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i25_4_lut.LUT_INIT = 16'h3c66;
    SB_LUT4 div_37_LessThan_2210_i7_4_lut (.I0(n3171), .I1(baudrate[3]), 
            .I2(n7806[3]), .I3(n294[1]), .O(n7));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i7_4_lut.LUT_INIT = 16'h3c66;
    SB_LUT4 div_37_LessThan_1845_i14_3_lut (.I0(baudrate[0]), .I1(baudrate[1]), 
            .I2(n2730), .I3(GND_net), .O(n14_adj_4946));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1845_i14_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i47491_3_lut (.I0(n14_adj_4946), .I1(baudrate[13]), .I2(n37_adj_4939), 
            .I3(GND_net), .O(n62204));   // verilog/uart_rx.v(119[33:55])
    defparam i47491_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i47492_3_lut (.I0(n62204), .I1(baudrate[14]), .I2(n39_adj_4801), 
            .I3(GND_net), .O(n62205));   // verilog/uart_rx.v(119[33:55])
    defparam i47492_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_2210_i45_4_lut (.I0(n3152), .I1(baudrate[22]), 
            .I2(n7806[22]), .I3(n294[1]), .O(n45_adj_4766));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i45_4_lut.LUT_INIT = 16'h3c66;
    SB_LUT4 div_37_LessThan_557_i42_3_lut (.I0(baudrate[0]), .I1(baudrate[1]), 
            .I2(n805), .I3(GND_net), .O(n42_adj_4947));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_557_i42_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i47541_3_lut (.I0(n42_adj_4947), .I1(baudrate[2]), .I2(n804), 
            .I3(GND_net), .O(n62254));   // verilog/uart_rx.v(119[33:55])
    defparam i47541_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i47542_3_lut (.I0(n62254), .I1(baudrate[3]), .I2(n803), .I3(GND_net), 
            .O(n62255));   // verilog/uart_rx.v(119[33:55])
    defparam i47542_3_lut.LUT_INIT = 16'h8e8e;
    SB_CARRY add_2540_6 (.CI(n46293), .I0(n1412), .I1(n1011), .CO(n46294));
    SB_LUT4 i42084_1_lut (.I0(n56786), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n53891));
    defparam i42084_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_37_LessThan_2210_i43_4_lut (.I0(n3153), .I1(baudrate[21]), 
            .I2(n7806[21]), .I3(n294[1]), .O(n43));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i43_4_lut.LUT_INIT = 16'h3c66;
    SB_LUT4 add_2540_5_lut (.I0(GND_net), .I1(n1413), .I2(n856), .I3(n46292), 
            .O(n7442[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2540_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2540_5 (.CI(n46292), .I0(n1413), .I1(n856), .CO(n46293));
    SB_LUT4 div_37_LessThan_2210_i9_4_lut (.I0(n3170), .I1(baudrate[4]), 
            .I2(n7806[4]), .I3(n294[1]), .O(n9));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i9_4_lut.LUT_INIT = 16'h3c66;
    SB_LUT4 add_2540_4_lut (.I0(GND_net), .I1(n1414), .I2(n698), .I3(n46291), 
            .O(n7442[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2540_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_LessThan_2210_i17_4_lut (.I0(n3166), .I1(baudrate[8]), 
            .I2(n7806[8]), .I3(n294[1]), .O(n17));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i17_4_lut.LUT_INIT = 16'h3c66;
    SB_LUT4 div_37_LessThan_2210_i19_4_lut (.I0(n3165), .I1(baudrate[9]), 
            .I2(n7806[9]), .I3(n294[1]), .O(n19));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i19_4_lut.LUT_INIT = 16'h3c66;
    SB_CARRY add_2540_4 (.CI(n46291), .I0(n1414), .I1(n698), .CO(n46292));
    SB_LUT4 add_2540_3_lut (.I0(GND_net), .I1(n1415), .I2(n858), .I3(n46290), 
            .O(n7442[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2540_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_LessThan_2210_i21_4_lut (.I0(n3164), .I1(baudrate[10]), 
            .I2(n7806[10]), .I3(n294[1]), .O(n21));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i21_4_lut.LUT_INIT = 16'h3c66;
    SB_CARRY add_2540_3 (.CI(n46290), .I0(n1415), .I1(n858), .CO(n46291));
    SB_LUT4 div_37_LessThan_2210_i35_4_lut (.I0(n3157), .I1(baudrate[17]), 
            .I2(n7806[17]), .I3(n294[1]), .O(n35));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i35_4_lut.LUT_INIT = 16'h3c66;
    SB_LUT4 div_37_LessThan_2210_i33_4_lut (.I0(n3158), .I1(baudrate[16]), 
            .I2(n7806[16]), .I3(n294[1]), .O(n33_c));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i33_4_lut.LUT_INIT = 16'h3c66;
    SB_LUT4 add_2540_2_lut (.I0(n53909), .I1(GND_net), .I2(n538), .I3(VCC_net), 
            .O(n55676)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2540_2_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_2540_2 (.CI(VCC_net), .I0(GND_net), .I1(n538), .CO(n46290));
    SB_LUT4 div_37_LessThan_557_i48_3_lut (.I0(n62255), .I1(baudrate[4]), 
            .I2(n53646), .I3(GND_net), .O(n48_adj_4948));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_557_i48_3_lut.LUT_INIT = 16'he8e8;
    SB_LUT4 div_37_i1838_3_lut (.I0(n2612), .I1(n7676[7]), .I2(n294[6]), 
            .I3(GND_net), .O(n2729));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1838_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_3_lut_4_lut_adj_964 (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[2]), 
            .I2(\r_Bit_Index[0] ), .I3(n4_adj_4821), .O(n55964));   // verilog/uart_rx.v(98[17:39])
    defparam i1_3_lut_4_lut_adj_964.LUT_INIT = 16'hffbf;
    SB_LUT4 i1_3_lut_4_lut_adj_965 (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[2]), 
            .I2(\r_Bit_Index[0] ), .I3(n4_adj_4821), .O(n55996));   // verilog/uart_rx.v(98[17:39])
    defparam i1_3_lut_4_lut_adj_965.LUT_INIT = 16'hfffb;
    SB_LUT4 i1_3_lut_adj_966 (.I0(n56814), .I1(n48_adj_4948), .I2(baudrate[0]), 
            .I3(GND_net), .O(n962));
    defparam i1_3_lut_adj_966.LUT_INIT = 16'h1010;
    SB_LUT4 i46057_3_lut (.I0(n962), .I1(baudrate[1]), .I2(n294[18]), 
            .I3(GND_net), .O(n1115));
    defparam i46057_3_lut.LUT_INIT = 16'h6a6a;
    SB_LUT4 div_37_i2172_1_lut (.I0(baudrate[3]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n856));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2172_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_37_i847_3_lut (.I0(n1115), .I1(n7390[19]), .I2(n294[17]), 
            .I3(GND_net), .O(n1265));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i847_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1915_3_lut (.I0(n2729), .I1(n7702[7]), .I2(n294[5]), 
            .I3(GND_net), .O(n2843));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1915_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i946_3_lut (.I0(n1265), .I1(n7416[19]), .I2(n294[16]), 
            .I3(GND_net), .O(n1412));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i946_3_lut.LUT_INIT = 16'hcaca;
    SB_DFFSR r_SM_Main_i1 (.Q(\r_SM_Main[1] ), .C(clk16MHz), .D(n3_adj_4949), 
            .R(\r_SM_Main[2] ));   // verilog/uart_rx.v(50[10] 145[8])
    SB_LUT4 div_37_i2171_1_lut (.I0(baudrate[4]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n1011));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2171_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_37_i1914_3_lut (.I0(n2728), .I1(n7702[8]), .I2(n294[5]), 
            .I3(GND_net), .O(n2842));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1914_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1517_i43_2_lut (.I0(n2229), .I1(baudrate[12]), 
            .I2(GND_net), .I3(GND_net), .O(n43_adj_4950));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1517_i43_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1517_i41_2_lut (.I0(n2230), .I1(baudrate[11]), 
            .I2(GND_net), .I3(GND_net), .O(n41_adj_4951));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1517_i41_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_2539_9_lut (.I0(GND_net), .I1(n1261), .I2(n1602), .I3(n46289), 
            .O(n7416[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2539_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2539_8_lut (.I0(GND_net), .I1(n1262), .I2(n1459), .I3(n46288), 
            .O(n7416[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2539_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2539_8 (.CI(n46288), .I0(n1262), .I1(n1459), .CO(n46289));
    SB_LUT4 add_2539_7_lut (.I0(GND_net), .I1(n1263), .I2(n1460), .I3(n46287), 
            .O(n7416[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2539_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2539_7 (.CI(n46287), .I0(n1263), .I1(n1460), .CO(n46288));
    SB_LUT4 add_2539_6_lut (.I0(GND_net), .I1(n1264), .I2(n1011), .I3(n46286), 
            .O(n7416[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2539_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2539_6 (.CI(n46286), .I0(n1264), .I1(n1011), .CO(n46287));
    SB_LUT4 div_37_LessThan_1517_i39_2_lut (.I0(n2231), .I1(baudrate[10]), 
            .I2(GND_net), .I3(GND_net), .O(n39_adj_4952));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1517_i39_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1517_i37_2_lut (.I0(n2232), .I1(baudrate[9]), 
            .I2(GND_net), .I3(GND_net), .O(n37_adj_4953));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1517_i37_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1517_i33_2_lut (.I0(n2234), .I1(baudrate[7]), 
            .I2(GND_net), .I3(GND_net), .O(n33_adj_4954));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1517_i33_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_2539_5_lut (.I0(GND_net), .I1(n1265), .I2(n856), .I3(n46285), 
            .O(n7416[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2539_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2539_5 (.CI(n46285), .I0(n1265), .I1(n856), .CO(n46286));
    SB_LUT4 div_37_LessThan_1517_i35_2_lut (.I0(n2233), .I1(baudrate[8]), 
            .I2(GND_net), .I3(GND_net), .O(n35_adj_4955));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1517_i35_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_4_lut_adj_967 (.I0(n56274), .I1(n56208), .I2(n56206), .I3(n56464), 
            .O(n22385));
    defparam i1_4_lut_adj_967.LUT_INIT = 16'hfffe;
    SB_LUT4 div_37_LessThan_1517_i25_2_lut (.I0(n2238), .I1(baudrate[3]), 
            .I2(GND_net), .I3(GND_net), .O(n25_adj_4956));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1517_i25_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1517_i27_2_lut (.I0(n2237), .I1(baudrate[4]), 
            .I2(GND_net), .I3(GND_net), .O(n27_adj_4957));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1517_i27_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1517_i29_2_lut (.I0(n2236), .I1(baudrate[5]), 
            .I2(GND_net), .I3(GND_net), .O(n29_adj_4958));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1517_i29_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_2539_4_lut (.I0(GND_net), .I1(n1266), .I2(n698), .I3(n46284), 
            .O(n7416[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2539_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2539_4 (.CI(n46284), .I0(n1266), .I1(n698), .CO(n46285));
    SB_LUT4 div_37_LessThan_1517_i31_2_lut (.I0(n2235), .I1(baudrate[6]), 
            .I2(GND_net), .I3(GND_net), .O(n31_adj_4959));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1517_i31_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1517_i23_2_lut (.I0(n2239), .I1(baudrate[2]), 
            .I2(GND_net), .I3(GND_net), .O(n23_adj_4960));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1517_i23_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i45483_4_lut (.I0(n29_adj_4958), .I1(n27_adj_4957), .I2(n25_adj_4956), 
            .I3(n23_adj_4960), .O(n60195));
    defparam i45483_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i45460_4_lut (.I0(n35_adj_4955), .I1(n33_adj_4954), .I2(n31_adj_4959), 
            .I3(n60195), .O(n60172));
    defparam i45460_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 add_2539_3_lut (.I0(GND_net), .I1(n1267), .I2(n858), .I3(n46283), 
            .O(n7416[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2539_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2539_3 (.CI(n46283), .I0(n1267), .I1(n858), .CO(n46284));
    SB_LUT4 div_37_LessThan_1517_i22_3_lut (.I0(baudrate[0]), .I1(baudrate[1]), 
            .I2(n2240), .I3(GND_net), .O(n22_adj_4961));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1517_i22_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_LessThan_1517_i30_3_lut (.I0(n28_adj_4962), .I1(baudrate[7]), 
            .I2(n33_adj_4954), .I3(GND_net), .O(n30_adj_4963));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1517_i30_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_2539_2_lut (.I0(n53913), .I1(GND_net), .I2(n538), .I3(VCC_net), 
            .O(n55674)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2539_2_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_2539_2 (.CI(VCC_net), .I0(GND_net), .I1(n538), .CO(n46283));
    SB_LUT4 add_2538_8_lut (.I0(GND_net), .I1(n1111), .I2(n1459), .I3(n46282), 
            .O(n7390[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2538_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2538_7_lut (.I0(GND_net), .I1(n1112), .I2(n1460), .I3(n46281), 
            .O(n7390[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2538_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_LessThan_1517_i34_3_lut (.I0(n26_adj_4964), .I1(baudrate[9]), 
            .I2(n37_adj_4953), .I3(GND_net), .O(n34_adj_4965));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1517_i34_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i48095_4_lut (.I0(n34_adj_4965), .I1(n24_adj_4966), .I2(n37_adj_4953), 
            .I3(n60166), .O(n62808));   // verilog/uart_rx.v(119[33:55])
    defparam i48095_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i48096_3_lut (.I0(n62808), .I1(baudrate[10]), .I2(n39_adj_4952), 
            .I3(GND_net), .O(n62809));   // verilog/uart_rx.v(119[33:55])
    defparam i48096_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i48065_3_lut (.I0(n62809), .I1(baudrate[11]), .I2(n41_adj_4951), 
            .I3(GND_net), .O(n62778));   // verilog/uart_rx.v(119[33:55])
    defparam i48065_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i47531_4_lut (.I0(n41_adj_4951), .I1(n39_adj_4952), .I2(n37_adj_4953), 
            .I3(n60172), .O(n62244));
    defparam i47531_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i47701_4_lut (.I0(n30_adj_4963), .I1(n22_adj_4961), .I2(n33_adj_4954), 
            .I3(n60187), .O(n62414));   // verilog/uart_rx.v(119[33:55])
    defparam i47701_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i1_2_lut_adj_968 (.I0(baudrate[26]), .I1(baudrate[27]), .I2(GND_net), 
            .I3(GND_net), .O(n56456));
    defparam i1_2_lut_adj_968.LUT_INIT = 16'heeee;
    SB_LUT4 i47895_3_lut (.I0(n62778), .I1(baudrate[12]), .I2(n43_adj_4950), 
            .I3(GND_net), .O(n42_adj_4967));   // verilog/uart_rx.v(119[33:55])
    defparam i47895_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_adj_969 (.I0(baudrate[30]), .I1(baudrate[31]), .I2(GND_net), 
            .I3(GND_net), .O(n56458));
    defparam i1_2_lut_adj_969.LUT_INIT = 16'heeee;
    SB_LUT4 i47962_4_lut (.I0(n42_adj_4967), .I1(n62414), .I2(n43_adj_4950), 
            .I3(n62244), .O(n62675));   // verilog/uart_rx.v(119[33:55])
    defparam i47962_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i1_4_lut_adj_970 (.I0(n56458), .I1(n56456), .I2(baudrate[17]), 
            .I3(n56484), .O(n56474));
    defparam i1_4_lut_adj_970.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_3_lut_adj_971 (.I0(n56472), .I1(n56474), .I2(n56470), .I3(GND_net), 
            .O(n22473));
    defparam i1_3_lut_adj_971.LUT_INIT = 16'hfefe;
    SB_LUT4 i39218_1_lut (.I0(n22473), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n53883));
    defparam i39218_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i47963_3_lut (.I0(n62675), .I1(baudrate[13]), .I2(n2228), 
            .I3(GND_net), .O(n62676));   // verilog/uart_rx.v(119[33:55])
    defparam i47963_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_i1232_3_lut (.I0(n1698), .I1(n7494[18]), .I2(n294[13]), 
            .I3(GND_net), .O(n1836));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1232_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_2538_7 (.CI(n46281), .I0(n1112), .I1(n1460), .CO(n46282));
    SB_LUT4 div_37_i1323_3_lut (.I0(n1836), .I1(n7520[18]), .I2(n294[12]), 
            .I3(GND_net), .O(n1971));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1323_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_2538_6_lut (.I0(GND_net), .I1(n1113), .I2(n1011), .I3(n46280), 
            .O(n7390[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2538_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2538_6 (.CI(n46280), .I0(n1113), .I1(n1011), .CO(n46281));
    SB_LUT4 div_37_i1412_3_lut (.I0(n1971), .I1(n7546[18]), .I2(n294[11]), 
            .I3(GND_net), .O(n2103));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1412_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1499_3_lut (.I0(n2103), .I1(n7572[18]), .I2(n294[10]), 
            .I3(GND_net), .O(n2232));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1499_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1676_3_lut (.I0(n2367), .I1(n7624[9]), .I2(n294[8]), 
            .I3(GND_net), .O(n2490));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1676_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1757_3_lut (.I0(n2490), .I1(n7650[9]), .I2(n294[7]), 
            .I3(GND_net), .O(n2610));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1757_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1836_3_lut (.I0(n2610), .I1(n7676[9]), .I2(n294[6]), 
            .I3(GND_net), .O(n2727));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1836_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1584_3_lut (.I0(n2232), .I1(n7598[18]), .I2(n294[9]), 
            .I3(GND_net), .O(n2358));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1584_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1667_3_lut (.I0(n2358), .I1(n7624[18]), .I2(n294[8]), 
            .I3(GND_net), .O(n2481));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1667_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2170_1_lut (.I0(baudrate[5]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n1460));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2170_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_37_i1913_3_lut (.I0(n2727), .I1(n7702[9]), .I2(n294[5]), 
            .I3(GND_net), .O(n2841));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1913_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_2538_5_lut (.I0(GND_net), .I1(n1114), .I2(n856), .I3(n46279), 
            .O(n7390[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2538_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2538_5 (.CI(n46279), .I0(n1114), .I1(n856), .CO(n46280));
    SB_LUT4 add_2538_4_lut (.I0(GND_net), .I1(n1115), .I2(n698), .I3(n46278), 
            .O(n7390[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2538_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_i1748_3_lut (.I0(n2481), .I1(n7650[18]), .I2(n294[7]), 
            .I3(GND_net), .O(n2601));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1748_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1662_3_lut (.I0(n2353), .I1(n7624[23]), .I2(n294[8]), 
            .I3(GND_net), .O(n2476));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1662_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1430_i37_2_lut (.I0(n2103), .I1(baudrate[8]), 
            .I2(GND_net), .I3(GND_net), .O(n37_adj_4968));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1430_i37_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1430_i35_2_lut (.I0(n2104), .I1(baudrate[7]), 
            .I2(GND_net), .I3(GND_net), .O(n35_adj_4969));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1430_i35_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_2538_4 (.CI(n46278), .I0(n1115), .I1(n698), .CO(n46279));
    SB_LUT4 add_2538_3_lut (.I0(GND_net), .I1(n1116), .I2(n858), .I3(n46277), 
            .O(n7390[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2538_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_i1743_3_lut (.I0(n2476), .I1(n7650[23]), .I2(n294[7]), 
            .I3(GND_net), .O(n2596));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1743_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1822_3_lut (.I0(n2596), .I1(n7676[23]), .I2(n294[6]), 
            .I3(GND_net), .O(n2713));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1822_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1430_i41_2_lut (.I0(n2101), .I1(baudrate[10]), 
            .I2(GND_net), .I3(GND_net), .O(n41_adj_4970));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1430_i41_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1430_i39_2_lut (.I0(n2102), .I1(baudrate[9]), 
            .I2(GND_net), .I3(GND_net), .O(n39_adj_4971));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1430_i39_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1430_i29_2_lut (.I0(n2107), .I1(baudrate[4]), 
            .I2(GND_net), .I3(GND_net), .O(n29_adj_4972));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1430_i29_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_2538_3 (.CI(n46277), .I0(n1116), .I1(n858), .CO(n46278));
    SB_LUT4 add_2538_2_lut (.I0(n53917), .I1(GND_net), .I2(n538), .I3(VCC_net), 
            .O(n55672)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2538_2_lut.LUT_INIT = 16'h8228;
    SB_LUT4 div_37_LessThan_1430_i31_2_lut (.I0(n2106), .I1(baudrate[5]), 
            .I2(GND_net), .I3(GND_net), .O(n31_adj_4973));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1430_i31_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_765_i43_2_lut (.I0(n1113), .I1(baudrate[4]), 
            .I2(GND_net), .I3(GND_net), .O(n43_adj_4974));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_765_i43_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1430_i33_2_lut (.I0(n2105), .I1(baudrate[6]), 
            .I2(GND_net), .I3(GND_net), .O(n33_adj_4975));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1430_i33_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1430_i27_2_lut (.I0(n2108), .I1(baudrate[3]), 
            .I2(GND_net), .I3(GND_net), .O(n27_adj_4976));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1430_i27_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i45550_4_lut (.I0(n33_adj_4975), .I1(n31_adj_4973), .I2(n29_adj_4972), 
            .I3(n27_adj_4976), .O(n60262));
    defparam i45550_4_lut.LUT_INIT = 16'haaab;
    SB_CARRY add_2538_2 (.CI(VCC_net), .I0(GND_net), .I1(n538), .CO(n46277));
    SB_LUT4 i42059_4_lut (.I0(baudrate[1]), .I1(n56346), .I2(n56292), 
            .I3(baudrate[3]), .O(n56762));
    defparam i42059_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 div_37_LessThan_765_i38_3_lut (.I0(baudrate[0]), .I1(baudrate[1]), 
            .I2(n1116), .I3(GND_net), .O(n38_adj_4977));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_765_i38_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_LessThan_765_i42_3_lut (.I0(n40_adj_4978), .I1(baudrate[4]), 
            .I2(n43_adj_4974), .I3(GND_net), .O(n42_adj_4979));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_765_i42_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1430_i38_3_lut (.I0(n30_adj_4980), .I1(baudrate[10]), 
            .I2(n41_adj_4970), .I3(GND_net), .O(n38_adj_4981));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1430_i38_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i21982_rep_6_2_lut (.I0(n7546[11]), .I1(n294[11]), .I2(GND_net), 
            .I3(GND_net), .O(n53894));   // verilog/uart_rx.v(119[33:55])
    defparam i21982_rep_6_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i48072_4_lut (.I0(n42_adj_4979), .I1(n38_adj_4977), .I2(n43_adj_4974), 
            .I3(n60469), .O(n62785));   // verilog/uart_rx.v(119[33:55])
    defparam i48072_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i48073_3_lut (.I0(n62785), .I1(baudrate[5]), .I2(n1112), .I3(GND_net), 
            .O(n62786));   // verilog/uart_rx.v(119[33:55])
    defparam i48073_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_LessThan_1430_i26_4_lut (.I0(n53894), .I1(baudrate[2]), 
            .I2(n2109), .I3(baudrate[1]), .O(n26_adj_4982));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1430_i26_4_lut.LUT_INIT = 16'h4d0c;
    SB_LUT4 i47707_3_lut (.I0(n26_adj_4982), .I1(baudrate[6]), .I2(n33_adj_4975), 
            .I3(GND_net), .O(n62420));   // verilog/uart_rx.v(119[33:55])
    defparam i47707_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i47708_3_lut (.I0(n62420), .I1(baudrate[7]), .I2(n35_adj_4969), 
            .I3(GND_net), .O(n62421));   // verilog/uart_rx.v(119[33:55])
    defparam i47708_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i45521_4_lut (.I0(n39_adj_4971), .I1(n37_adj_4968), .I2(n35_adj_4969), 
            .I3(n60262), .O(n60233));
    defparam i45521_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i48093_4_lut (.I0(n38_adj_4981), .I1(n28_adj_4983), .I2(n41_adj_4970), 
            .I3(n60227), .O(n62806));   // verilog/uart_rx.v(119[33:55])
    defparam i48093_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i47600_3_lut (.I0(n62421), .I1(baudrate[8]), .I2(n37_adj_4968), 
            .I3(GND_net), .O(n62313));   // verilog/uart_rx.v(119[33:55])
    defparam i47600_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i948_3_lut (.I0(n1267), .I1(n7416[17]), .I2(n294[16]), 
            .I3(GND_net), .O(n1414));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i948_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i48258_4_lut (.I0(n62313), .I1(n62806), .I2(n41_adj_4970), 
            .I3(n60233), .O(n62971));   // verilog/uart_rx.v(119[33:55])
    defparam i48258_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i48259_3_lut (.I0(n62971), .I1(baudrate[11]), .I2(n2100), 
            .I3(GND_net), .O(n62972));   // verilog/uart_rx.v(119[33:55])
    defparam i48259_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_i1045_3_lut (.I0(n1414), .I1(n7442[17]), .I2(n294[15]), 
            .I3(GND_net), .O(n1558));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1045_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i48178_3_lut (.I0(n62972), .I1(baudrate[12]), .I2(n2099), 
            .I3(GND_net), .O(n62891));   // verilog/uart_rx.v(119[33:55])
    defparam i48178_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i48171_3_lut (.I0(n62891), .I1(baudrate[13]), .I2(n2098), 
            .I3(GND_net), .O(n48_adj_4984));   // verilog/uart_rx.v(119[33:55])
    defparam i48171_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_i1140_3_lut (.I0(n1558), .I1(n7468[17]), .I2(n294[14]), 
            .I3(GND_net), .O(n1699));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1140_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1233_3_lut (.I0(n1699), .I1(n7494[17]), .I2(n294[13]), 
            .I3(GND_net), .O(n1837));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1233_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_972 (.I0(baudrate[27]), .I1(baudrate[24]), .I2(baudrate[29]), 
            .I3(baudrate[30]), .O(n56410));
    defparam i1_4_lut_adj_972.LUT_INIT = 16'hfffe;
    SB_LUT4 div_37_i1324_3_lut (.I0(n1837), .I1(n7520[17]), .I2(n294[12]), 
            .I3(GND_net), .O(n1972));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1324_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_973 (.I0(n56418), .I1(n56274), .I2(n56416), .I3(n56410), 
            .O(n22464));
    defparam i1_4_lut_adj_973.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_3_lut_adj_974 (.I0(n22464), .I1(n48_adj_4984), .I2(baudrate[0]), 
            .I3(GND_net), .O(n2240));
    defparam i1_3_lut_adj_974.LUT_INIT = 16'hefef;
    SB_LUT4 i48503_4_lut_4_lut (.I0(\r_SM_Main_2__N_3219[1] ), .I1(\r_SM_Main[1] ), 
            .I2(n6_adj_4985), .I3(n55461), .O(n53789));
    defparam i48503_4_lut_4_lut.LUT_INIT = 16'h0703;
    SB_LUT4 div_37_i1413_3_lut (.I0(n1972), .I1(n7546[17]), .I2(n294[11]), 
            .I3(GND_net), .O(n2104));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1413_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1592_3_lut (.I0(n2240), .I1(n7598[10]), .I2(n294[9]), 
            .I3(GND_net), .O(n2366));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1592_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_3_lut_4_lut_adj_975 (.I0(baudrate[2]), .I1(baudrate[3]), 
            .I2(n56292), .I3(n56346), .O(n56242));
    defparam i1_3_lut_4_lut_adj_975.LUT_INIT = 16'hfffe;
    SB_LUT4 div_37_i1500_3_lut (.I0(n2104), .I1(n7572[17]), .I2(n294[10]), 
            .I3(GND_net), .O(n2233));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1500_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_976 (.I0(n56762), .I1(n56786), .I2(n56344), .I3(n56118), 
            .O(n48_adj_4986));
    defparam i1_4_lut_adj_976.LUT_INIT = 16'h0100;
    SB_LUT4 i1_2_lut_3_lut_4_lut (.I0(baudrate[16]), .I1(baudrate[17]), 
            .I2(baudrate[15]), .I3(baudrate[14]), .O(n56382));
    defparam i1_2_lut_3_lut_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 div_37_i1675_3_lut (.I0(n2366), .I1(n7624[10]), .I2(n294[8]), 
            .I3(GND_net), .O(n2489));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1675_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1585_3_lut (.I0(n2233), .I1(n7598[17]), .I2(n294[9]), 
            .I3(GND_net), .O(n2359));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1585_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF r_Rx_Byte_i4 (.Q(rx_data[4]), .C(clk16MHz), .D(n26587));   // verilog/uart_rx.v(50[10] 145[8])
    SB_LUT4 div_37_i1756_3_lut (.I0(n2489), .I1(n7650[10]), .I2(n294[7]), 
            .I3(GND_net), .O(n2609));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1756_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1668_3_lut (.I0(n2359), .I1(n7624[17]), .I2(n294[8]), 
            .I3(GND_net), .O(n2482));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1668_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1749_3_lut (.I0(n2482), .I1(n7650[17]), .I2(n294[7]), 
            .I3(GND_net), .O(n2602));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1749_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1835_3_lut (.I0(n2609), .I1(n7676[10]), .I2(n294[6]), 
            .I3(GND_net), .O(n2726));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1835_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF r_Rx_Byte_i7 (.Q(rx_data[7]), .C(clk16MHz), .D(n26062));   // verilog/uart_rx.v(50[10] 145[8])
    SB_LUT4 div_37_i1828_3_lut (.I0(n2602), .I1(n7676[17]), .I2(n294[6]), 
            .I3(GND_net), .O(n2719));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1828_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2169_1_lut (.I0(baudrate[6]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n1459));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2169_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_37_i1912_3_lut (.I0(n2726), .I1(n7702[10]), .I2(n294[5]), 
            .I3(GND_net), .O(n2840));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1912_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1845_i35_2_lut (.I0(n2719), .I1(baudrate[12]), 
            .I2(GND_net), .I3(GND_net), .O(n35_adj_4945));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1845_i35_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_977 (.I0(baudrate[24]), .I1(baudrate[29]), .I2(GND_net), 
            .I3(GND_net), .O(n56484));
    defparam i1_2_lut_adj_977.LUT_INIT = 16'heeee;
    SB_LUT4 i1_2_lut_adj_978 (.I0(baudrate[30]), .I1(baudrate[25]), .I2(GND_net), 
            .I3(GND_net), .O(n56354));
    defparam i1_2_lut_adj_978.LUT_INIT = 16'heeee;
    SB_LUT4 add_2554_25_lut (.I0(GND_net), .I1(n3151), .I2(n3186), .I3(n46513), 
            .O(n7806[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2554_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2554_24_lut (.I0(GND_net), .I1(n3152), .I2(n3082), .I3(n46512), 
            .O(n7806[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2554_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2554_24 (.CI(n46512), .I0(n3152), .I1(n3082), .CO(n46513));
    SB_LUT4 add_2554_23_lut (.I0(GND_net), .I1(n3153), .I2(n3188), .I3(n46511), 
            .O(n7806[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2554_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2554_23 (.CI(n46511), .I0(n3153), .I1(n3188), .CO(n46512));
    SB_LUT4 add_2554_22_lut (.I0(GND_net), .I1(n3154), .I2(n3084), .I3(n46510), 
            .O(n7806[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2554_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2554_22 (.CI(n46510), .I0(n3154), .I1(n3084), .CO(n46511));
    SB_LUT4 add_2554_21_lut (.I0(GND_net), .I1(n3155), .I2(n2977), .I3(n46509), 
            .O(n7806[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2554_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2554_21 (.CI(n46509), .I0(n3155), .I1(n2977), .CO(n46510));
    SB_LUT4 add_2554_20_lut (.I0(GND_net), .I1(n3156), .I2(n2867), .I3(n46508), 
            .O(n7806[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2554_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2554_20 (.CI(n46508), .I0(n3156), .I1(n2867), .CO(n46509));
    SB_LUT4 add_2554_19_lut (.I0(GND_net), .I1(n3157), .I2(n2754), .I3(n46507), 
            .O(n7806[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2554_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2554_19 (.CI(n46507), .I0(n3157), .I1(n2754), .CO(n46508));
    SB_LUT4 add_2554_18_lut (.I0(GND_net), .I1(n3158), .I2(n2638), .I3(n46506), 
            .O(n7806[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2554_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2554_18 (.CI(n46506), .I0(n3158), .I1(n2638), .CO(n46507));
    SB_LUT4 i7_2_lut (.I0(baudrate[12]), .I1(baudrate[13]), .I2(GND_net), 
            .I3(GND_net), .O(n25_adj_4987));
    defparam i7_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 add_2554_17_lut (.I0(GND_net), .I1(n3159), .I2(n2519), .I3(n46505), 
            .O(n7806[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2554_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2554_17 (.CI(n46505), .I0(n3159), .I1(n2519), .CO(n46506));
    SB_LUT4 add_2554_16_lut (.I0(GND_net), .I1(n3160), .I2(n2397), .I3(n46504), 
            .O(n7806[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2554_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2554_16 (.CI(n46504), .I0(n3160), .I1(n2397), .CO(n46505));
    SB_LUT4 add_2554_15_lut (.I0(GND_net), .I1(n3161), .I2(n2272), .I3(n46503), 
            .O(n7806[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2554_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2554_15 (.CI(n46503), .I0(n3161), .I1(n2272), .CO(n46504));
    SB_LUT4 add_2554_14_lut (.I0(GND_net), .I1(n3162), .I2(n2144), .I3(n46502), 
            .O(n7806[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2554_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2554_14 (.CI(n46502), .I0(n3162), .I1(n2144), .CO(n46503));
    SB_LUT4 add_2554_13_lut (.I0(GND_net), .I1(n3163), .I2(n2013), .I3(n46501), 
            .O(n7806[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2554_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2554_13 (.CI(n46501), .I0(n3163), .I1(n2013), .CO(n46502));
    SB_LUT4 add_2554_12_lut (.I0(GND_net), .I1(n3164), .I2(n1879), .I3(n46500), 
            .O(n7806[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2554_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2554_12 (.CI(n46500), .I0(n3164), .I1(n1879), .CO(n46501));
    SB_LUT4 add_2554_11_lut (.I0(GND_net), .I1(n3165), .I2(n1742), .I3(n46499), 
            .O(n7806[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2554_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2554_11 (.CI(n46499), .I0(n3165), .I1(n1742), .CO(n46500));
    SB_LUT4 add_2554_10_lut (.I0(GND_net), .I1(n3166), .I2(n1602), .I3(n46498), 
            .O(n7806[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2554_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2554_10 (.CI(n46498), .I0(n3166), .I1(n1602), .CO(n46499));
    SB_LUT4 add_2554_9_lut (.I0(GND_net), .I1(n3167), .I2(n1459), .I3(n46497), 
            .O(n7806[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2554_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2554_9 (.CI(n46497), .I0(n3167), .I1(n1459), .CO(n46498));
    SB_LUT4 add_2554_8_lut (.I0(GND_net), .I1(n3168), .I2(n1460), .I3(n46496), 
            .O(n7806[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2554_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2554_8 (.CI(n46496), .I0(n3168), .I1(n1460), .CO(n46497));
    SB_LUT4 add_2554_7_lut (.I0(GND_net), .I1(n3169), .I2(n1011), .I3(n46495), 
            .O(n7806[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2554_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2554_7 (.CI(n46495), .I0(n3169), .I1(n1011), .CO(n46496));
    SB_LUT4 add_2554_6_lut (.I0(GND_net), .I1(n3170), .I2(n856), .I3(n46494), 
            .O(n7806[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2554_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2554_6 (.CI(n46494), .I0(n3170), .I1(n856), .CO(n46495));
    SB_LUT4 add_2554_5_lut (.I0(GND_net), .I1(n3171), .I2(n698), .I3(n46493), 
            .O(n7806[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2554_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2554_5 (.CI(n46493), .I0(n3171), .I1(n698), .CO(n46494));
    SB_LUT4 add_2554_4_lut (.I0(GND_net), .I1(n3172), .I2(n858), .I3(n46492), 
            .O(n7806[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2554_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2554_4 (.CI(n46492), .I0(n3172), .I1(n858), .CO(n46493));
    SB_LUT4 add_2554_3_lut (.I0(n53859), .I1(GND_net), .I2(n538), .I3(n46491), 
            .O(n55696)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2554_3_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_2554_3 (.CI(n46491), .I0(GND_net), .I1(n538), .CO(n46492));
    SB_CARRY add_2554_2 (.CI(VCC_net), .I0(GND_net), .I1(VCC_net), .CO(n46491));
    SB_LUT4 add_2553_23_lut (.I0(GND_net), .I1(n3046), .I2(n3082), .I3(n46490), 
            .O(n7780[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2553_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2553_22_lut (.I0(GND_net), .I1(n3047), .I2(n3188), .I3(n46489), 
            .O(n7780[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2553_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2553_22 (.CI(n46489), .I0(n3047), .I1(n3188), .CO(n46490));
    SB_LUT4 add_2553_21_lut (.I0(GND_net), .I1(n3048), .I2(n3084), .I3(n46488), 
            .O(n7780[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2553_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2553_21 (.CI(n46488), .I0(n3048), .I1(n3084), .CO(n46489));
    SB_LUT4 add_2553_20_lut (.I0(GND_net), .I1(n3049), .I2(n2977), .I3(n46487), 
            .O(n7780[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2553_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2553_20 (.CI(n46487), .I0(n3049), .I1(n2977), .CO(n46488));
    SB_LUT4 add_2553_19_lut (.I0(GND_net), .I1(n3050), .I2(n2867), .I3(n46486), 
            .O(n7780[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2553_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2553_19 (.CI(n46486), .I0(n3050), .I1(n2867), .CO(n46487));
    SB_LUT4 add_2553_18_lut (.I0(GND_net), .I1(n3051), .I2(n2754), .I3(n46485), 
            .O(n7780[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2553_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2553_18 (.CI(n46485), .I0(n3051), .I1(n2754), .CO(n46486));
    SB_LUT4 add_2553_17_lut (.I0(GND_net), .I1(n3052), .I2(n2638), .I3(n46484), 
            .O(n7780[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2553_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2553_17 (.CI(n46484), .I0(n3052), .I1(n2638), .CO(n46485));
    SB_LUT4 add_2553_16_lut (.I0(GND_net), .I1(n3053), .I2(n2519), .I3(n46483), 
            .O(n7780[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2553_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2553_16 (.CI(n46483), .I0(n3053), .I1(n2519), .CO(n46484));
    SB_LUT4 add_2553_15_lut (.I0(GND_net), .I1(n3054), .I2(n2397), .I3(n46482), 
            .O(n7780[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2553_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2553_15 (.CI(n46482), .I0(n3054), .I1(n2397), .CO(n46483));
    SB_LUT4 add_2553_14_lut (.I0(GND_net), .I1(n3055), .I2(n2272), .I3(n46481), 
            .O(n7780[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2553_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2553_14 (.CI(n46481), .I0(n3055), .I1(n2272), .CO(n46482));
    SB_LUT4 add_2553_13_lut (.I0(GND_net), .I1(n3056), .I2(n2144), .I3(n46480), 
            .O(n7780[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2553_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2553_13 (.CI(n46480), .I0(n3056), .I1(n2144), .CO(n46481));
    SB_LUT4 add_2553_12_lut (.I0(GND_net), .I1(n3057), .I2(n2013), .I3(n46479), 
            .O(n7780[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2553_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2553_12 (.CI(n46479), .I0(n3057), .I1(n2013), .CO(n46480));
    SB_LUT4 add_2553_11_lut (.I0(GND_net), .I1(n3058), .I2(n1879), .I3(n46478), 
            .O(n7780[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2553_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2553_11 (.CI(n46478), .I0(n3058), .I1(n1879), .CO(n46479));
    SB_LUT4 add_2553_10_lut (.I0(GND_net), .I1(n3059), .I2(n1742), .I3(n46477), 
            .O(n7780[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2553_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2553_10 (.CI(n46477), .I0(n3059), .I1(n1742), .CO(n46478));
    SB_LUT4 add_2553_9_lut (.I0(GND_net), .I1(n3060), .I2(n1602), .I3(n46476), 
            .O(n7780[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2553_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2553_9 (.CI(n46476), .I0(n3060), .I1(n1602), .CO(n46477));
    SB_LUT4 add_2553_8_lut (.I0(GND_net), .I1(n3061), .I2(n1459), .I3(n46475), 
            .O(n7780[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2553_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2553_8 (.CI(n46475), .I0(n3061), .I1(n1459), .CO(n46476));
    SB_LUT4 add_2553_7_lut (.I0(GND_net), .I1(n3062), .I2(n1460), .I3(n46474), 
            .O(n7780[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2553_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2553_7 (.CI(n46474), .I0(n3062), .I1(n1460), .CO(n46475));
    SB_LUT4 add_2553_6_lut (.I0(GND_net), .I1(n3063), .I2(n1011), .I3(n46473), 
            .O(n7780[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2553_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2553_6 (.CI(n46473), .I0(n3063), .I1(n1011), .CO(n46474));
    SB_LUT4 add_2553_5_lut (.I0(GND_net), .I1(n3064), .I2(n856), .I3(n46472), 
            .O(n7780[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2553_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2553_5 (.CI(n46472), .I0(n3064), .I1(n856), .CO(n46473));
    SB_LUT4 add_2553_4_lut (.I0(GND_net), .I1(n3065), .I2(n698), .I3(n46471), 
            .O(n7780[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2553_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2553_4 (.CI(n46471), .I0(n3065), .I1(n698), .CO(n46472));
    SB_LUT4 add_2553_3_lut (.I0(GND_net), .I1(n3066), .I2(n858), .I3(n46470), 
            .O(n7780[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2553_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2553_3 (.CI(n46470), .I0(n3066), .I1(n858), .CO(n46471));
    SB_LUT4 add_2553_2_lut (.I0(n53863), .I1(GND_net), .I2(n538), .I3(VCC_net), 
            .O(n55694)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2553_2_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_2553_2 (.CI(VCC_net), .I0(GND_net), .I1(n538), .CO(n46470));
    SB_LUT4 add_2552_22_lut (.I0(GND_net), .I1(n2938), .I2(n3188), .I3(n46469), 
            .O(n7754[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2552_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_2_lut_adj_979 (.I0(baudrate[31]), .I1(baudrate[26]), .I2(GND_net), 
            .I3(GND_net), .O(n56358));
    defparam i1_2_lut_adj_979.LUT_INIT = 16'heeee;
    SB_LUT4 i1_2_lut_adj_980 (.I0(baudrate[27]), .I1(baudrate[30]), .I2(GND_net), 
            .I3(GND_net), .O(n56308));
    defparam i1_2_lut_adj_980.LUT_INIT = 16'heeee;
    SB_LUT4 add_2552_21_lut (.I0(GND_net), .I1(n2939), .I2(n3084), .I3(n46468), 
            .O(n7754[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2552_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2552_21 (.CI(n46468), .I0(n2939), .I1(n3084), .CO(n46469));
    SB_LUT4 add_2552_20_lut (.I0(GND_net), .I1(n2940), .I2(n2977), .I3(n46467), 
            .O(n7754[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2552_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2552_20 (.CI(n46467), .I0(n2940), .I1(n2977), .CO(n46468));
    SB_LUT4 add_2552_19_lut (.I0(GND_net), .I1(n2941), .I2(n2867), .I3(n46466), 
            .O(n7754[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2552_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2552_19 (.CI(n46466), .I0(n2941), .I1(n2867), .CO(n46467));
    SB_LUT4 add_2552_18_lut (.I0(GND_net), .I1(n2942), .I2(n2754), .I3(n46465), 
            .O(n7754[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2552_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2552_18 (.CI(n46465), .I0(n2942), .I1(n2754), .CO(n46466));
    SB_LUT4 add_2552_17_lut (.I0(GND_net), .I1(n2943), .I2(n2638), .I3(n46464), 
            .O(n7754[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2552_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_2_lut_adj_981 (.I0(baudrate[25]), .I1(baudrate[28]), .I2(GND_net), 
            .I3(GND_net), .O(n56452));
    defparam i1_2_lut_adj_981.LUT_INIT = 16'heeee;
    SB_CARRY add_2552_17 (.CI(n46464), .I0(n2943), .I1(n2638), .CO(n46465));
    SB_LUT4 i42069_4_lut (.I0(n56486), .I1(baudrate[16]), .I2(baudrate[15]), 
            .I3(n56452), .O(n56772));
    defparam i42069_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 add_2552_16_lut (.I0(GND_net), .I1(n2944), .I2(n2519), .I3(n46463), 
            .O(n7754[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2552_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2552_16 (.CI(n46463), .I0(n2944), .I1(n2519), .CO(n46464));
    SB_LUT4 add_2552_15_lut (.I0(GND_net), .I1(n2945), .I2(n2397), .I3(n46462), 
            .O(n7754[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2552_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2552_15 (.CI(n46462), .I0(n2945), .I1(n2397), .CO(n46463));
    SB_LUT4 add_2552_14_lut (.I0(GND_net), .I1(n2946), .I2(n2272), .I3(n46461), 
            .O(n7754[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2552_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2552_14 (.CI(n46461), .I0(n2946), .I1(n2272), .CO(n46462));
    SB_LUT4 add_2552_13_lut (.I0(GND_net), .I1(n2947), .I2(n2144), .I3(n46460), 
            .O(n7754[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2552_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2552_13 (.CI(n46460), .I0(n2947), .I1(n2144), .CO(n46461));
    SB_LUT4 add_2552_12_lut (.I0(GND_net), .I1(n2948), .I2(n2013), .I3(n46459), 
            .O(n7754[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2552_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2552_12 (.CI(n46459), .I0(n2948), .I1(n2013), .CO(n46460));
    SB_LUT4 add_2552_11_lut (.I0(GND_net), .I1(n2949), .I2(n1879), .I3(n46458), 
            .O(n7754[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2552_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2552_11 (.CI(n46458), .I0(n2949), .I1(n1879), .CO(n46459));
    SB_LUT4 add_2552_10_lut (.I0(GND_net), .I1(n2950), .I2(n1742), .I3(n46457), 
            .O(n7754[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2552_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2552_10 (.CI(n46457), .I0(n2950), .I1(n1742), .CO(n46458));
    SB_LUT4 i42071_4_lut (.I0(n56358), .I1(n56484), .I2(n56308), .I3(baudrate[17]), 
            .O(n56774));
    defparam i42071_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 add_2552_9_lut (.I0(GND_net), .I1(n2951), .I2(n1602), .I3(n46456), 
            .O(n7754[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2552_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i42083_3_lut (.I0(n56774), .I1(n56772), .I2(n56472), .I3(GND_net), 
            .O(n56786));
    defparam i42083_3_lut.LUT_INIT = 16'hfefe;
    SB_CARRY add_2552_9 (.CI(n46456), .I0(n2951), .I1(n1602), .CO(n46457));
    SB_LUT4 add_2552_8_lut (.I0(GND_net), .I1(n2952), .I2(n1459), .I3(n46455), 
            .O(n7754[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2552_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2552_8 (.CI(n46455), .I0(n2952), .I1(n1459), .CO(n46456));
    SB_LUT4 add_2552_7_lut (.I0(GND_net), .I1(n2953), .I2(n1460), .I3(n46454), 
            .O(n7754[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2552_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2552_7 (.CI(n46454), .I0(n2953), .I1(n1460), .CO(n46455));
    SB_LUT4 add_2552_6_lut (.I0(GND_net), .I1(n2954), .I2(n1011), .I3(n46453), 
            .O(n7754[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2552_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_3_lut_4_lut_adj_982 (.I0(n24_adj_4901), .I1(n56792), .I2(n7468[14]), 
            .I3(n48_adj_4988), .O(n1702));
    defparam i1_3_lut_4_lut_adj_982.LUT_INIT = 16'h0010;
    SB_CARRY add_2552_6 (.CI(n46453), .I0(n2954), .I1(n1011), .CO(n46454));
    SB_LUT4 i1_3_lut_4_lut_adj_983 (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[2]), 
            .I2(\r_Bit_Index[0] ), .I3(n4_adj_4821), .O(n55884));   // verilog/uart_rx.v(98[17:39])
    defparam i1_3_lut_4_lut_adj_983.LUT_INIT = 16'hffdf;
    SB_LUT4 add_2552_5_lut (.I0(GND_net), .I1(n2955), .I2(n856), .I3(n46452), 
            .O(n7754[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2552_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2552_5 (.CI(n46452), .I0(n2955), .I1(n856), .CO(n46453));
    SB_LUT4 add_2552_4_lut (.I0(GND_net), .I1(n2956), .I2(n698), .I3(n46451), 
            .O(n7754[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2552_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i42007_2_lut (.I0(baudrate[13]), .I1(baudrate[14]), .I2(GND_net), 
            .I3(GND_net), .O(n56710));
    defparam i42007_2_lut.LUT_INIT = 16'heeee;
    SB_CARRY add_2552_4 (.CI(n46451), .I0(n2956), .I1(n698), .CO(n46452));
    SB_LUT4 add_2552_3_lut (.I0(GND_net), .I1(n2957), .I2(n858), .I3(n46450), 
            .O(n7754[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2552_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_3_lut_4_lut_adj_984 (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[2]), 
            .I2(\r_Bit_Index[0] ), .I3(n4_adj_4821), .O(n55900));   // verilog/uart_rx.v(98[17:39])
    defparam i1_3_lut_4_lut_adj_984.LUT_INIT = 16'hfffd;
    SB_CARRY add_2552_3 (.CI(n46450), .I0(n2957), .I1(n858), .CO(n46451));
    SB_LUT4 add_2552_2_lut (.I0(n53867), .I1(GND_net), .I2(n538), .I3(VCC_net), 
            .O(n55692)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2552_2_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_2552_2 (.CI(VCC_net), .I0(GND_net), .I1(n538), .CO(n46450));
    SB_LUT4 add_2551_21_lut (.I0(GND_net), .I1(n2827), .I2(n3084), .I3(n46449), 
            .O(n7728[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2551_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2551_20_lut (.I0(GND_net), .I1(n2828), .I2(n2977), .I3(n46448), 
            .O(n7728[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2551_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2551_20 (.CI(n46448), .I0(n2828), .I1(n2977), .CO(n46449));
    SB_LUT4 add_2551_19_lut (.I0(GND_net), .I1(n2829), .I2(n2867), .I3(n46447), 
            .O(n7728[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2551_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_2_lut_adj_985 (.I0(baudrate[27]), .I1(baudrate[28]), .I2(GND_net), 
            .I3(GND_net), .O(n56356));
    defparam i1_2_lut_adj_985.LUT_INIT = 16'heeee;
    SB_CARRY add_2551_19 (.CI(n46447), .I0(n2829), .I1(n2867), .CO(n46448));
    SB_LUT4 add_2551_18_lut (.I0(GND_net), .I1(n2830), .I2(n2754), .I3(n46446), 
            .O(n7728[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2551_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2551_18 (.CI(n46446), .I0(n2830), .I1(n2754), .CO(n46447));
    SB_LUT4 div_37_LessThan_1341_i37_2_lut (.I0(n1971), .I1(baudrate[7]), 
            .I2(GND_net), .I3(GND_net), .O(n37_adj_4989));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1341_i37_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_2551_17_lut (.I0(GND_net), .I1(n2831), .I2(n2638), .I3(n46445), 
            .O(n7728[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2551_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2551_17 (.CI(n46445), .I0(n2831), .I1(n2638), .CO(n46446));
    SB_LUT4 add_2551_16_lut (.I0(GND_net), .I1(n2832), .I2(n2519), .I3(n46444), 
            .O(n7728[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2551_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_LessThan_1341_i35_2_lut (.I0(n1972), .I1(baudrate[6]), 
            .I2(GND_net), .I3(GND_net), .O(n35_adj_4990));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1341_i35_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_986 (.I0(baudrate[22]), .I1(baudrate[23]), .I2(GND_net), 
            .I3(GND_net), .O(n56486));
    defparam i1_2_lut_adj_986.LUT_INIT = 16'heeee;
    SB_LUT4 div_37_LessThan_1341_i41_2_lut (.I0(n1969), .I1(baudrate[9]), 
            .I2(GND_net), .I3(GND_net), .O(n41_adj_4991));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1341_i41_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1157_i43_2_lut (.I0(n1695), .I1(baudrate[8]), 
            .I2(GND_net), .I3(GND_net), .O(n43_adj_4992));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1157_i43_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1341_i29_2_lut (.I0(n1975), .I1(baudrate[3]), 
            .I2(GND_net), .I3(GND_net), .O(n29_adj_4993));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1341_i29_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1157_i39_2_lut (.I0(n1697), .I1(baudrate[6]), 
            .I2(GND_net), .I3(GND_net), .O(n39_adj_4994));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1157_i39_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1341_i31_2_lut (.I0(n1974), .I1(baudrate[4]), 
            .I2(GND_net), .I3(GND_net), .O(n31_adj_4995));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1341_i31_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1341_i33_2_lut (.I0(n1973), .I1(baudrate[5]), 
            .I2(GND_net), .I3(GND_net), .O(n33_adj_4996));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1341_i33_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1341_i39_2_lut (.I0(n1970), .I1(baudrate[8]), 
            .I2(GND_net), .I3(GND_net), .O(n39_adj_4997));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1341_i39_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_987 (.I0(n56382), .I1(n56472), .I2(GND_net), 
            .I3(GND_net), .O(n56388));
    defparam i1_2_lut_adj_987.LUT_INIT = 16'heeee;
    SB_LUT4 div_37_LessThan_1341_i27_2_lut (.I0(n1976), .I1(baudrate[2]), 
            .I2(GND_net), .I3(GND_net), .O(n27_adj_4998));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1341_i27_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i45616_4_lut (.I0(n33_adj_4996), .I1(n31_adj_4995), .I2(n29_adj_4993), 
            .I3(n27_adj_4998), .O(n60328));
    defparam i45616_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i1_2_lut_4_lut (.I0(n62676), .I1(baudrate[14]), .I2(n2227), 
            .I3(n55680), .O(n2367));   // verilog/uart_rx.v(119[33:55])
    defparam i1_2_lut_4_lut.LUT_INIT = 16'h7100;
    SB_LUT4 div_37_LessThan_1341_i38_3_lut (.I0(n30_adj_4999), .I1(baudrate[9]), 
            .I2(n41_adj_4991), .I3(GND_net), .O(n38_adj_5000));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1341_i38_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1341_i26_3_lut (.I0(baudrate[0]), .I1(baudrate[1]), 
            .I2(n1977), .I3(GND_net), .O(n26_adj_5001));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1341_i26_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i48523_2_lut_4_lut (.I0(n62676), .I1(baudrate[14]), .I2(n2227), 
            .I3(n56786), .O(n294[9]));   // verilog/uart_rx.v(119[33:55])
    defparam i48523_2_lut_4_lut.LUT_INIT = 16'h0071;
    SB_LUT4 i47711_3_lut (.I0(n26_adj_5001), .I1(baudrate[5]), .I2(n33_adj_4996), 
            .I3(GND_net), .O(n62424));   // verilog/uart_rx.v(119[33:55])
    defparam i47711_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i47712_3_lut (.I0(n62424), .I1(baudrate[6]), .I2(n35_adj_4990), 
            .I3(GND_net), .O(n62425));   // verilog/uart_rx.v(119[33:55])
    defparam i47712_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_988 (.I0(n56556), .I1(n56318), .I2(n56486), .I3(n56308), 
            .O(n22481));
    defparam i1_4_lut_adj_988.LUT_INIT = 16'hfffe;
    SB_LUT4 i21967_rep_8_2_lut (.I0(baudrate[0]), .I1(n294[19]), .I2(GND_net), 
            .I3(GND_net), .O(n53920));   // verilog/uart_rx.v(119[33:55])
    defparam i21967_rep_8_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i45605_4_lut (.I0(n39_adj_4997), .I1(n37_adj_4989), .I2(n35_adj_4990), 
            .I3(n60328), .O(n60317));
    defparam i45605_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 div_37_LessThan_662_i42_4_lut (.I0(n53920), .I1(baudrate[2]), 
            .I2(n961), .I3(baudrate[1]), .O(n42_adj_5002));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_662_i42_4_lut.LUT_INIT = 16'h4d0c;
    SB_LUT4 i48156_4_lut (.I0(n38_adj_5000), .I1(n28_adj_5003), .I2(n41_adj_4991), 
            .I3(n60315), .O(n62869));   // verilog/uart_rx.v(119[33:55])
    defparam i48156_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i47596_3_lut (.I0(n62425), .I1(baudrate[7]), .I2(n37_adj_4989), 
            .I3(GND_net), .O(n62309));   // verilog/uart_rx.v(119[33:55])
    defparam i47596_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_989 (.I0(n56242), .I1(n22385), .I2(n56344), .I3(n56382), 
            .O(n22444));
    defparam i1_4_lut_adj_989.LUT_INIT = 16'hfffe;
    SB_LUT4 i47579_3_lut (.I0(n42_adj_5002), .I1(baudrate[3]), .I2(n960), 
            .I3(GND_net), .O(n62292));   // verilog/uart_rx.v(119[33:55])
    defparam i47579_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_LessThan_1845_i40_3_lut (.I0(n22_adj_5004), .I1(baudrate[17]), 
            .I2(n45_adj_4858), .I3(GND_net), .O(n40_adj_5005));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1845_i40_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i47580_3_lut (.I0(n62292), .I1(baudrate[4]), .I2(n959), .I3(GND_net), 
            .O(n62293));   // verilog/uart_rx.v(119[33:55])
    defparam i47580_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_LessThan_662_i48_3_lut (.I0(n62293), .I1(baudrate[5]), 
            .I2(n53648), .I3(GND_net), .O(n48_adj_5006));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_662_i48_3_lut.LUT_INIT = 16'he8e8;
    SB_LUT4 i46093_4_lut (.I0(n43_adj_4809), .I1(n41_adj_4808), .I2(n39_adj_4801), 
            .I3(n60817), .O(n60805));
    defparam i46093_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i48254_4_lut (.I0(n62309), .I1(n62869), .I2(n41_adj_4991), 
            .I3(n60317), .O(n62967));   // verilog/uart_rx.v(119[33:55])
    defparam i48254_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i1_4_lut_adj_990 (.I0(n56346), .I1(n22481), .I2(n56388), .I3(n56344), 
            .O(n22507));
    defparam i1_4_lut_adj_990.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_3_lut_adj_991 (.I0(n22507), .I1(n48_adj_5006), .I2(baudrate[0]), 
            .I3(GND_net), .O(n1116));
    defparam i1_3_lut_adj_991.LUT_INIT = 16'hefef;
    SB_LUT4 i48255_3_lut (.I0(n62967), .I1(baudrate[10]), .I2(n1968), 
            .I3(GND_net), .O(n62968));   // verilog/uart_rx.v(119[33:55])
    defparam i48255_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i1_2_lut_4_lut_adj_992 (.I0(n61937), .I1(baudrate[16]), .I2(n2476), 
            .I3(n55684), .O(n2612));   // verilog/uart_rx.v(119[33:55])
    defparam i1_2_lut_4_lut_adj_992.LUT_INIT = 16'h7100;
    SB_LUT4 i48529_2_lut_4_lut (.I0(n61937), .I1(baudrate[16]), .I2(n2476), 
            .I3(n22473), .O(n294[7]));   // verilog/uart_rx.v(119[33:55])
    defparam i48529_2_lut_4_lut.LUT_INIT = 16'h0071;
    SB_LUT4 div_37_i848_3_lut (.I0(n1116), .I1(n7390[18]), .I2(n294[17]), 
            .I3(GND_net), .O(n1266));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i848_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i947_3_lut (.I0(n1266), .I1(n7416[18]), .I2(n294[16]), 
            .I3(GND_net), .O(n1413));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i947_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1044_3_lut (.I0(n1413), .I1(n7442[18]), .I2(n294[15]), 
            .I3(GND_net), .O(n1557));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1044_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1139_3_lut (.I0(n1557), .I1(n7468[18]), .I2(n294[14]), 
            .I3(GND_net), .O(n1698));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1139_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i48182_3_lut (.I0(n62968), .I1(baudrate[11]), .I2(n1967), 
            .I3(GND_net), .O(n62895));   // verilog/uart_rx.v(119[33:55])
    defparam i48182_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_LessThan_1157_i37_2_lut (.I0(n1698), .I1(baudrate[5]), 
            .I2(GND_net), .I3(GND_net), .O(n37_adj_5007));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1157_i37_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i48169_3_lut (.I0(n62895), .I1(baudrate[12]), .I2(n1966), 
            .I3(GND_net), .O(n48_adj_5008));   // verilog/uart_rx.v(119[33:55])
    defparam i48169_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i48526_2_lut_4_lut (.I0(n62868), .I1(baudrate[15]), .I2(n2353), 
            .I3(n22470), .O(n294[8]));   // verilog/uart_rx.v(119[33:55])
    defparam i48526_2_lut_4_lut.LUT_INIT = 16'h0071;
    SB_LUT4 i47625_4_lut (.I0(n40_adj_5005), .I1(n20_adj_5009), .I2(n45_adj_4858), 
            .I3(n60792), .O(n62338));   // verilog/uart_rx.v(119[33:55])
    defparam i47625_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i1_2_lut_4_lut_adj_993 (.I0(n62868), .I1(baudrate[15]), .I2(n2353), 
            .I3(n55682), .O(n2491));   // verilog/uart_rx.v(119[33:55])
    defparam i1_2_lut_4_lut_adj_993.LUT_INIT = 16'h7100;
    SB_LUT4 div_37_LessThan_1157_i41_2_lut (.I0(n1696), .I1(baudrate[7]), 
            .I2(GND_net), .I3(GND_net), .O(n41_adj_5010));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1157_i41_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1506_3_lut (.I0(n2110), .I1(n7572[11]), .I2(n294[10]), 
            .I3(GND_net), .O(n2239));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1506_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1591_3_lut (.I0(n2239), .I1(n7598[11]), .I2(n294[9]), 
            .I3(GND_net), .O(n2365));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1591_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1674_3_lut (.I0(n2365), .I1(n7624[11]), .I2(n294[8]), 
            .I3(GND_net), .O(n2488));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1674_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1755_3_lut (.I0(n2488), .I1(n7650[11]), .I2(n294[7]), 
            .I3(GND_net), .O(n2608));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1755_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i46066_4_lut (.I0(n22444), .I1(n60170), .I2(n48_adj_4986), 
            .I3(baudrate[0]), .O(n644));
    defparam i46066_4_lut.LUT_INIT = 16'h3633;
    SB_LUT4 i21975_rep_7_2_lut (.I0(n7468[14]), .I1(n294[14]), .I2(GND_net), 
            .I3(GND_net), .O(n53903));   // verilog/uart_rx.v(119[33:55])
    defparam i21975_rep_7_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 div_37_i1834_3_lut (.I0(n2608), .I1(n7676[11]), .I2(n294[6]), 
            .I3(GND_net), .O(n2725));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1834_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_3_lut_4_lut_adj_994 (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[2]), 
            .I2(\r_Bit_Index[0] ), .I3(n4_adj_4821), .O(n55916));   // verilog/uart_rx.v(98[17:39])
    defparam i1_3_lut_4_lut_adj_994.LUT_INIT = 16'hfffe;
    SB_LUT4 div_37_i2168_1_lut (.I0(baudrate[7]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n1602));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2168_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_37_LessThan_1157_i32_4_lut (.I0(n53903), .I1(baudrate[2]), 
            .I2(n1701), .I3(baudrate[1]), .O(n32_adj_5011));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1157_i32_4_lut.LUT_INIT = 16'h4d0c;
    SB_LUT4 i47515_3_lut (.I0(n32_adj_5011), .I1(baudrate[6]), .I2(n39_adj_4994), 
            .I3(GND_net), .O(n62228));   // verilog/uart_rx.v(119[33:55])
    defparam i47515_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1911_3_lut (.I0(n2725), .I1(n7702[11]), .I2(n294[5]), 
            .I3(GND_net), .O(n2839));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1911_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_3_lut_4_lut_adj_995 (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[2]), 
            .I2(\r_Bit_Index[0] ), .I3(n4_adj_4821), .O(n55932));   // verilog/uart_rx.v(98[17:39])
    defparam i1_3_lut_4_lut_adj_995.LUT_INIT = 16'hffef;
    SB_LUT4 i47516_3_lut (.I0(n62228), .I1(baudrate[7]), .I2(n41_adj_5010), 
            .I3(GND_net), .O(n62229));   // verilog/uart_rx.v(119[33:55])
    defparam i47516_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i46579_3_lut (.I0(n62205), .I1(baudrate[15]), .I2(n41_adj_4808), 
            .I3(GND_net), .O(n61292));   // verilog/uart_rx.v(119[33:55])
    defparam i46579_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i46660_4_lut (.I0(n41_adj_5010), .I1(n39_adj_4994), .I2(n37_adj_5007), 
            .I3(n60410), .O(n61373));
    defparam i46660_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i47591_3_lut (.I0(n34_adj_5012), .I1(baudrate[5]), .I2(n37_adj_5007), 
            .I3(GND_net), .O(n62304));   // verilog/uart_rx.v(119[33:55])
    defparam i47591_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1250_i39_2_lut (.I0(n1835), .I1(baudrate[7]), 
            .I2(GND_net), .I3(GND_net), .O(n39_adj_5013));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1250_i39_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i46558_3_lut (.I0(n62229), .I1(baudrate[8]), .I2(n43_adj_4992), 
            .I3(GND_net), .O(n61271));   // verilog/uart_rx.v(119[33:55])
    defparam i46558_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1250_i43_2_lut (.I0(n1833), .I1(baudrate[9]), 
            .I2(GND_net), .I3(GND_net), .O(n43_adj_5014));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1250_i43_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1250_i37_2_lut (.I0(n1836), .I1(baudrate[6]), 
            .I2(GND_net), .I3(GND_net), .O(n37_adj_5015));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1250_i37_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i47832_4_lut (.I0(n61271), .I1(n62304), .I2(n43_adj_4992), 
            .I3(n61373), .O(n62545));   // verilog/uart_rx.v(119[33:55])
    defparam i47832_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 div_37_LessThan_1250_i31_2_lut (.I0(n1839), .I1(baudrate[3]), 
            .I2(GND_net), .I3(GND_net), .O(n31_adj_5016));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1250_i31_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1250_i35_2_lut (.I0(n1837), .I1(baudrate[5]), 
            .I2(GND_net), .I3(GND_net), .O(n35_adj_5017));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1250_i35_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i47833_3_lut (.I0(n62545), .I1(baudrate[9]), .I2(n1694), .I3(GND_net), 
            .O(n62546));   // verilog/uart_rx.v(119[33:55])
    defparam i47833_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i41997_2_lut (.I0(\o_Rx_DV_N_3261[12] ), .I1(n52650), .I2(GND_net), 
            .I3(GND_net), .O(n56700));
    defparam i41997_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 div_37_LessThan_1250_i33_2_lut (.I0(n1838), .I1(baudrate[4]), 
            .I2(GND_net), .I3(GND_net), .O(n33_adj_5018));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1250_i33_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1250_i41_2_lut (.I0(n1834), .I1(baudrate[8]), 
            .I2(GND_net), .I3(GND_net), .O(n41_adj_5019));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1250_i41_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i42077_4_lut (.I0(\o_Rx_DV_N_3261[24] ), .I1(n29), .I2(n23), 
            .I3(n56700), .O(n56780));
    defparam i42077_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 r_SM_Main_2__I_0_62_Mux_0_i2_4_lut (.I0(n55814), .I1(\r_SM_Main_2__N_3219[1] ), 
            .I2(r_SM_Main[0]), .I3(n27), .O(n2));   // verilog/uart_rx.v(53[7] 144[14])
    defparam r_SM_Main_2__I_0_62_Mux_0_i2_4_lut.LUT_INIT = 16'hc0c5;
    SB_LUT4 r_SM_Main_2__I_0_62_Mux_0_i1_4_lut (.I0(r_Rx_Data), .I1(n56780), 
            .I2(r_SM_Main[0]), .I3(n27), .O(n9473));   // verilog/uart_rx.v(53[7] 144[14])
    defparam r_SM_Main_2__I_0_62_Mux_0_i1_4_lut.LUT_INIT = 16'h0a3a;
    SB_LUT4 div_37_LessThan_1250_i29_2_lut (.I0(n1840), .I1(baudrate[2]), 
            .I2(GND_net), .I3(GND_net), .O(n29_adj_5020));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1250_i29_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 r_SM_Main_2__I_0_62_Mux_0_i3_3_lut (.I0(n9473), .I1(n2), .I2(\r_SM_Main[1] ), 
            .I3(GND_net), .O(n3));   // verilog/uart_rx.v(53[7] 144[14])
    defparam r_SM_Main_2__I_0_62_Mux_0_i3_3_lut.LUT_INIT = 16'hc5c5;
    SB_LUT4 i45652_4_lut (.I0(n35_adj_5017), .I1(n33_adj_5018), .I2(n31_adj_5016), 
            .I3(n29_adj_5020), .O(n60364));
    defparam i45652_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 div_37_LessThan_965_i41_2_lut (.I0(n1411), .I1(baudrate[5]), 
            .I2(GND_net), .I3(GND_net), .O(n41_adj_5021));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_965_i41_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_965_i43_2_lut (.I0(n1410), .I1(baudrate[6]), 
            .I2(GND_net), .I3(GND_net), .O(n43_adj_5022));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_965_i43_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1062_i39_2_lut (.I0(n1556), .I1(baudrate[5]), 
            .I2(GND_net), .I3(GND_net), .O(n39_adj_5023));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1062_i39_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1062_i41_2_lut (.I0(n1555), .I1(baudrate[6]), 
            .I2(GND_net), .I3(GND_net), .O(n41_adj_5024));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1062_i41_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1062_i37_2_lut (.I0(n1557), .I1(baudrate[4]), 
            .I2(GND_net), .I3(GND_net), .O(n37_adj_5025));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1062_i37_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1062_i43_2_lut (.I0(n1554), .I1(baudrate[7]), 
            .I2(GND_net), .I3(GND_net), .O(n43_adj_5026));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1062_i43_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_996 (.I0(baudrate[17]), .I1(baudrate[18]), .I2(GND_net), 
            .I3(GND_net), .O(n56160));
    defparam i1_2_lut_adj_996.LUT_INIT = 16'heeee;
    SB_LUT4 div_37_i535_4_lut (.I0(n644), .I1(n44), .I2(n294[20]), .I3(baudrate[2]), 
            .O(n803));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i535_4_lut.LUT_INIT = 16'h6a9a;
    SB_LUT4 i5659_4_lut (.I0(n804), .I1(n35469), .I2(n18896), .I3(baudrate[2]), 
            .O(n18960));   // verilog/uart_rx.v(119[33:55])
    defparam i5659_4_lut.LUT_INIT = 16'ha2aa;
    SB_LUT4 div_37_LessThan_1602_i27_2_lut (.I0(n2363), .I1(baudrate[5]), 
            .I2(GND_net), .I3(GND_net), .O(n27_adj_4868));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1602_i27_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1602_i29_2_lut (.I0(n2362), .I1(baudrate[6]), 
            .I2(GND_net), .I3(GND_net), .O(n29_adj_4874));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1602_i29_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1602_i25_2_lut (.I0(n2364), .I1(baudrate[4]), 
            .I2(GND_net), .I3(GND_net), .O(n25_adj_4869));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1602_i25_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1602_i33_2_lut (.I0(n2360), .I1(baudrate[8]), 
            .I2(GND_net), .I3(GND_net), .O(n33_adj_4872));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1602_i33_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1157_i48_3_lut (.I0(n62546), .I1(baudrate[10]), 
            .I2(n1693), .I3(GND_net), .O(n48_adj_5027));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1157_i48_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_LessThan_1602_i23_2_lut (.I0(n2365), .I1(baudrate[3]), 
            .I2(GND_net), .I3(GND_net), .O(n23_adj_4870));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1602_i23_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1250_i40_3_lut (.I0(n32_adj_5028), .I1(baudrate[9]), 
            .I2(n43_adj_5014), .I3(GND_net), .O(n40_adj_5029));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1250_i40_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1602_i35_2_lut (.I0(n2359), .I1(baudrate[9]), 
            .I2(GND_net), .I3(GND_net), .O(n35_adj_4894));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1602_i35_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1602_i37_2_lut (.I0(n2358), .I1(baudrate[10]), 
            .I2(GND_net), .I3(GND_net), .O(n37_adj_4897));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1602_i37_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_4_lut_adj_997 (.I0(n56486), .I1(n56356), .I2(n56358), .I3(baudrate[11]), 
            .O(n56386));
    defparam i1_4_lut_adj_997.LUT_INIT = 16'hfffe;
    SB_LUT4 div_37_LessThan_1602_i39_2_lut (.I0(n2357), .I1(baudrate[11]), 
            .I2(GND_net), .I3(GND_net), .O(n39_adj_4898));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1602_i39_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1602_i31_2_lut (.I0(n2361), .I1(baudrate[7]), 
            .I2(GND_net), .I3(GND_net), .O(n31_adj_4873));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1602_i31_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1602_i41_2_lut (.I0(n2356), .I1(baudrate[12]), 
            .I2(GND_net), .I3(GND_net), .O(n41_adj_4924));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1602_i41_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1845_i21_2_lut (.I0(n2726), .I1(baudrate[5]), 
            .I2(GND_net), .I3(GND_net), .O(n21_adj_4942));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1845_i21_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1845_i37_2_lut (.I0(n2718), .I1(baudrate[13]), 
            .I2(GND_net), .I3(GND_net), .O(n37_adj_4939));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1845_i37_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1845_i25_2_lut (.I0(n2724), .I1(baudrate[7]), 
            .I2(GND_net), .I3(GND_net), .O(n25_adj_4940));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1845_i25_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1845_i23_2_lut (.I0(n2725), .I1(baudrate[6]), 
            .I2(GND_net), .I3(GND_net), .O(n23_adj_4941));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1845_i23_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1250_i28_3_lut (.I0(baudrate[0]), .I1(baudrate[1]), 
            .I2(n1841), .I3(GND_net), .O(n28_adj_5030));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1250_i28_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i47513_3_lut (.I0(n28_adj_5030), .I1(baudrate[5]), .I2(n35_adj_5017), 
            .I3(GND_net), .O(n62226));   // verilog/uart_rx.v(119[33:55])
    defparam i47513_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i47514_3_lut (.I0(n62226), .I1(baudrate[6]), .I2(n37_adj_5015), 
            .I3(GND_net), .O(n62227));   // verilog/uart_rx.v(119[33:55])
    defparam i47514_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i45637_4_lut (.I0(n41_adj_5019), .I1(n39_adj_5013), .I2(n37_adj_5015), 
            .I3(n60364), .O(n60349));
    defparam i45637_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i47713_4_lut (.I0(n40_adj_5029), .I1(n30_adj_5031), .I2(n43_adj_5014), 
            .I3(n60347), .O(n62426));   // verilog/uart_rx.v(119[33:55])
    defparam i47713_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i46561_3_lut (.I0(n62227), .I1(baudrate[7]), .I2(n39_adj_5013), 
            .I3(GND_net), .O(n61274));   // verilog/uart_rx.v(119[33:55])
    defparam i46561_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i48091_4_lut (.I0(n61274), .I1(n62426), .I2(n43_adj_5014), 
            .I3(n60349), .O(n62804));   // verilog/uart_rx.v(119[33:55])
    defparam i48091_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i3834_2_lut (.I0(n18960), .I1(n9112), .I2(GND_net), .I3(GND_net), 
            .O(n44_adj_5032));   // verilog/uart_rx.v(119[33:55])
    defparam i3834_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i48092_3_lut (.I0(n62804), .I1(baudrate[10]), .I2(n1832), 
            .I3(GND_net), .O(n62805));   // verilog/uart_rx.v(119[33:55])
    defparam i48092_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i1_4_lut_adj_998 (.I0(n56386), .I1(n56388), .I2(n56376), .I3(n25_adj_4987), 
            .O(n22492));
    defparam i1_4_lut_adj_998.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_3_lut_adj_999 (.I0(n22492), .I1(n48_adj_5027), .I2(baudrate[0]), 
            .I3(GND_net), .O(n1841));
    defparam i1_3_lut_adj_999.LUT_INIT = 16'hefef;
    SB_LUT4 div_37_i1328_3_lut (.I0(n1841), .I1(n7520[13]), .I2(n294[12]), 
            .I3(GND_net), .O(n1976));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1328_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1418_3_lut (.I0(n1977), .I1(n7546[12]), .I2(n294[11]), 
            .I3(GND_net), .O(n2109));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1418_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1505_3_lut (.I0(n2109), .I1(n7572[12]), .I2(n294[10]), 
            .I3(GND_net), .O(n2238));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1505_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i640_4_lut (.I0(n803), .I1(baudrate[3]), .I2(n294[19]), 
            .I3(n44_adj_5032), .O(n959));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i640_4_lut.LUT_INIT = 16'h6a9a;
    SB_LUT4 div_37_i1417_3_lut (.I0(n1976), .I1(n7546[13]), .I2(n294[11]), 
            .I3(GND_net), .O(n2108));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1417_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1590_3_lut (.I0(n2238), .I1(n7598[12]), .I2(n294[9]), 
            .I3(GND_net), .O(n2364));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1590_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1673_3_lut (.I0(n2364), .I1(n7624[12]), .I2(n294[8]), 
            .I3(GND_net), .O(n2487));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1673_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1504_3_lut (.I0(n2108), .I1(n7572[13]), .I2(n294[10]), 
            .I3(GND_net), .O(n2237));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1504_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1589_3_lut (.I0(n2237), .I1(n7598[13]), .I2(n294[9]), 
            .I3(GND_net), .O(n2363));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1589_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1672_3_lut (.I0(n2363), .I1(n7624[13]), .I2(n294[8]), 
            .I3(GND_net), .O(n2486));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1672_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1753_3_lut (.I0(n2486), .I1(n7650[13]), .I2(n294[7]), 
            .I3(GND_net), .O(n2606));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1753_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i39198_1_lut (.I0(n22481), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n53863));
    defparam i39198_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_37_i1832_3_lut (.I0(n2606), .I1(n7676[13]), .I2(n294[6]), 
            .I3(GND_net), .O(n2723));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1832_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1754_3_lut (.I0(n2487), .I1(n7650[12]), .I2(n294[7]), 
            .I3(GND_net), .O(n2607));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1754_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i944_3_lut (.I0(n1263), .I1(n7416[21]), .I2(n294[16]), 
            .I3(GND_net), .O(n1410));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i944_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1041_3_lut (.I0(n1410), .I1(n7442[21]), .I2(n294[15]), 
            .I3(GND_net), .O(n1554));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1041_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1136_3_lut (.I0(n1554), .I1(n7468[21]), .I2(n294[14]), 
            .I3(GND_net), .O(n1695));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1136_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1833_3_lut (.I0(n2607), .I1(n7676[12]), .I2(n294[6]), 
            .I3(GND_net), .O(n2724));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1833_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2167_1_lut (.I0(baudrate[8]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n1742));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2167_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_37_i1910_3_lut (.I0(n2724), .I1(n7702[12]), .I2(n294[5]), 
            .I3(GND_net), .O(n2838));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1910_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2166_1_lut (.I0(baudrate[9]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n1879));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2166_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_37_i1909_3_lut (.I0(n2723), .I1(n7702[13]), .I2(n294[5]), 
            .I3(GND_net), .O(n2837));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1909_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1229_3_lut (.I0(n1695), .I1(n7494[21]), .I2(n294[13]), 
            .I3(GND_net), .O(n1833));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1229_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2165_1_lut (.I0(baudrate[10]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n2013));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2165_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_37_i2156_1_lut (.I0(baudrate[19]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n3084));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2156_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_37_i1908_3_lut (.I0(n2722), .I1(n7702[14]), .I2(n294[5]), 
            .I3(GND_net), .O(n2836));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1908_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2155_1_lut (.I0(baudrate[20]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n3188));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2155_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_37_i2083_1_lut (.I0(baudrate[21]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n3082));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2083_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_37_i2153_1_lut (.I0(baudrate[22]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n3186));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2153_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_37_i2164_1_lut (.I0(baudrate[11]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n2144));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2164_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_37_i1907_3_lut (.I0(n2721), .I1(n7702[15]), .I2(n294[5]), 
            .I3(GND_net), .O(n2835));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1907_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1320_3_lut (.I0(n1833), .I1(n7520[21]), .I2(n294[12]), 
            .I3(GND_net), .O(n1968));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1320_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1409_3_lut (.I0(n1968), .I1(n7546[21]), .I2(n294[11]), 
            .I3(GND_net), .O(n2100));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1409_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i743_4_lut (.I0(n959), .I1(baudrate[4]), .I2(n294[18]), 
            .I3(n44_adj_5033), .O(n1112));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i743_4_lut.LUT_INIT = 16'h6a9a;
    SB_LUT4 div_37_i1496_3_lut (.I0(n2100), .I1(n7572[21]), .I2(n294[10]), 
            .I3(GND_net), .O(n2229));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1496_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1581_3_lut (.I0(n2229), .I1(n7598[21]), .I2(n294[9]), 
            .I3(GND_net), .O(n2355));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1581_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1664_3_lut (.I0(n2355), .I1(n7624[21]), .I2(n294[8]), 
            .I3(GND_net), .O(n2478));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1664_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1745_3_lut (.I0(n2478), .I1(n7650[21]), .I2(n294[7]), 
            .I3(GND_net), .O(n2598));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1745_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2163_1_lut (.I0(baudrate[12]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n2272));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2163_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_37_i1906_3_lut (.I0(n2720), .I1(n7702[16]), .I2(n294[5]), 
            .I3(GND_net), .O(n2834));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1906_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i945_3_lut (.I0(n1264), .I1(n7416[20]), .I2(n294[16]), 
            .I3(GND_net), .O(n1411));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i945_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1042_3_lut (.I0(n1411), .I1(n7442[20]), .I2(n294[15]), 
            .I3(GND_net), .O(n1555));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1042_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2162_1_lut (.I0(baudrate[13]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n2397));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2162_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_37_i1137_3_lut (.I0(n1555), .I1(n7468[20]), .I2(n294[14]), 
            .I3(GND_net), .O(n1696));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1137_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1230_3_lut (.I0(n1696), .I1(n7494[20]), .I2(n294[13]), 
            .I3(GND_net), .O(n1834));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1230_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1905_3_lut (.I0(n2719), .I1(n7702[17]), .I2(n294[5]), 
            .I3(GND_net), .O(n2833));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1905_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i844_3_lut (.I0(n1112), .I1(n7390[22]), .I2(n294[17]), 
            .I3(GND_net), .O(n1262));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i844_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1321_3_lut (.I0(n1834), .I1(n7520[20]), .I2(n294[12]), 
            .I3(GND_net), .O(n1969));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1321_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4005_2_lut_4_lut (.I0(n960), .I1(n9276), .I2(n19008), .I3(baudrate[3]), 
            .O(n44_adj_5033));   // verilog/uart_rx.v(119[33:55])
    defparam i4005_2_lut_4_lut.LUT_INIT = 16'ha8fe;
    SB_LUT4 div_37_i1410_3_lut (.I0(n1969), .I1(n7546[20]), .I2(n294[11]), 
            .I3(GND_net), .O(n2101));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1410_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1497_3_lut (.I0(n2101), .I1(n7572[20]), .I2(n294[10]), 
            .I3(GND_net), .O(n2230));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1497_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1582_3_lut (.I0(n2230), .I1(n7598[20]), .I2(n294[9]), 
            .I3(GND_net), .O(n2356));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1582_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1665_3_lut (.I0(n2356), .I1(n7624[20]), .I2(n294[8]), 
            .I3(GND_net), .O(n2479));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1665_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1746_3_lut (.I0(n2479), .I1(n7650[20]), .I2(n294[7]), 
            .I3(GND_net), .O(n2599));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1746_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13_2_lut_3_lut_4_lut (.I0(baudrate[14]), .I1(baudrate[15]), 
            .I2(baudrate[12]), .I3(baudrate[13]), .O(n31_adj_4905));
    defparam i13_2_lut_3_lut_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_3_lut (.I0(baudrate[0]), .I1(baudrate[1]), .I2(n56818), 
            .I3(GND_net), .O(n35725));
    defparam i1_2_lut_3_lut.LUT_INIT = 16'h0202;
    SB_LUT4 i42115_3_lut_4_lut (.I0(baudrate[3]), .I1(baudrate[4]), .I2(n56814), 
            .I3(baudrate[2]), .O(n56818));
    defparam i42115_3_lut_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 div_37_i943_3_lut (.I0(n1262), .I1(n7416[22]), .I2(n294[16]), 
            .I3(GND_net), .O(n1409));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i943_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1000 (.I0(baudrate[20]), .I1(baudrate[21]), 
            .I2(baudrate[18]), .I3(baudrate[19]), .O(n56472));
    defparam i1_2_lut_3_lut_4_lut_adj_1000.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1001 (.I0(baudrate[20]), .I1(baudrate[21]), 
            .I2(baudrate[22]), .I3(baudrate[23]), .O(n56274));
    defparam i1_2_lut_3_lut_4_lut_adj_1001.LUT_INIT = 16'hfffe;
    SB_LUT4 i48454_3_lut_4_lut_3_lut (.I0(n56818), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n56822));
    defparam i48454_3_lut_4_lut_3_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i48520_2_lut_3_lut_4_lut (.I0(baudrate[13]), .I1(baudrate[14]), 
            .I2(n56786), .I3(n48_adj_5008), .O(n294[11]));
    defparam i48520_2_lut_3_lut_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 i42089_2_lut_3_lut_4_lut (.I0(baudrate[13]), .I1(baudrate[14]), 
            .I2(n56786), .I3(baudrate[12]), .O(n56792));
    defparam i42089_2_lut_3_lut_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1002 (.I0(baudrate[5]), .I1(baudrate[6]), 
            .I2(baudrate[3]), .I3(baudrate[4]), .O(n56182));
    defparam i1_2_lut_3_lut_4_lut_adj_1002.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_3_lut_adj_1003 (.I0(\r_SM_Main[1] ), .I1(r_SM_Main[0]), 
            .I2(\r_SM_Main[2] ), .I3(GND_net), .O(n4_adj_4821));
    defparam i1_2_lut_3_lut_adj_1003.LUT_INIT = 16'hfdfd;
    SB_LUT4 i42102_1_lut (.I0(n56804), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n53917));
    defparam i42102_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_37_LessThan_965_i45_2_lut (.I0(n1409), .I1(baudrate[7]), 
            .I2(GND_net), .I3(GND_net), .O(n45_adj_5034));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_965_i45_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_965_i39_2_lut (.I0(n1412), .I1(baudrate[4]), 
            .I2(GND_net), .I3(GND_net), .O(n39_adj_5035));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_965_i39_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i42099_2_lut (.I0(baudrate[8]), .I1(n56800), .I2(GND_net), 
            .I3(GND_net), .O(n56802));
    defparam i42099_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i1_2_lut_4_lut_adj_1004 (.I0(n62744), .I1(baudrate[17]), .I2(n2596), 
            .I3(n55686), .O(n2730));   // verilog/uart_rx.v(119[33:55])
    defparam i1_2_lut_4_lut_adj_1004.LUT_INIT = 16'h7100;
    SB_LUT4 i48532_2_lut_4_lut (.I0(n62744), .I1(baudrate[17]), .I2(n2596), 
            .I3(n22385), .O(n294[6]));   // verilog/uart_rx.v(119[33:55])
    defparam i48532_2_lut_4_lut.LUT_INIT = 16'h0071;
    SB_LUT4 div_37_LessThan_965_i34_3_lut (.I0(baudrate[0]), .I1(baudrate[1]), 
            .I2(n1415), .I3(GND_net), .O(n34_adj_5036));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_965_i34_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_LessThan_1845_i16_3_lut_3_lut (.I0(baudrate[2]), .I1(baudrate[3]), 
            .I2(n2728), .I3(GND_net), .O(n16_adj_5037));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1845_i16_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_LessThan_1845_i26_3_lut (.I0(n18_adj_5038), .I1(baudrate[9]), 
            .I2(n29_adj_4944), .I3(GND_net), .O(n26_adj_5039));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1845_i26_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i47537_3_lut (.I0(n34_adj_5036), .I1(baudrate[5]), .I2(n41_adj_5021), 
            .I3(GND_net), .O(n62250));   // verilog/uart_rx.v(119[33:55])
    defparam i47537_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i47936_4_lut (.I0(n26_adj_5039), .I1(n16_adj_5037), .I2(n29_adj_4944), 
            .I3(n60840), .O(n62649));   // verilog/uart_rx.v(119[33:55])
    defparam i47936_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i47538_3_lut (.I0(n62250), .I1(baudrate[6]), .I2(n43_adj_5022), 
            .I3(GND_net), .O(n62251));   // verilog/uart_rx.v(119[33:55])
    defparam i47538_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i47937_3_lut (.I0(n62649), .I1(baudrate[10]), .I2(n31_adj_4943), 
            .I3(GND_net), .O(n62650));   // verilog/uart_rx.v(119[33:55])
    defparam i47937_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i46692_4_lut (.I0(n43_adj_5022), .I1(n41_adj_5021), .I2(n39_adj_5035), 
            .I3(n60449), .O(n61405));
    defparam i46692_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 div_37_LessThan_965_i38_3_lut (.I0(n36_adj_5040), .I1(baudrate[4]), 
            .I2(n39_adj_5035), .I3(GND_net), .O(n38_adj_5041));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_965_i38_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i47821_3_lut (.I0(n62650), .I1(baudrate[11]), .I2(n33_adj_4927), 
            .I3(GND_net), .O(n62534));   // verilog/uart_rx.v(119[33:55])
    defparam i47821_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i46551_3_lut (.I0(n62251), .I1(baudrate[7]), .I2(n45_adj_5034), 
            .I3(GND_net), .O(n61264));   // verilog/uart_rx.v(119[33:55])
    defparam i46551_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i47778_4_lut (.I0(n43_adj_4809), .I1(n41_adj_4808), .I2(n39_adj_4801), 
            .I3(n60819), .O(n62491));
    defparam i47778_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i47585_4_lut (.I0(n61264), .I1(n38_adj_5041), .I2(n45_adj_5034), 
            .I3(n61405), .O(n62298));   // verilog/uart_rx.v(119[33:55])
    defparam i47585_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i46087_4_lut (.I0(r_SM_Main[0]), .I1(\o_Rx_DV_N_3261[12] ), 
            .I2(n4834), .I3(\o_Rx_DV_N_3261[8] ), .O(n59759));   // verilog/uart_rx.v(53[7] 144[14])
    defparam i46087_4_lut.LUT_INIT = 16'hfffd;
    SB_LUT4 i46140_4_lut (.I0(r_Rx_Data), .I1(\o_Rx_DV_N_3261[12] ), .I2(n52650), 
            .I3(r_SM_Main[0]), .O(n59765));   // verilog/uart_rx.v(53[7] 144[14])
    defparam i46140_4_lut.LUT_INIT = 16'h0100;
    SB_LUT4 i46084_4_lut (.I0(n59759), .I1(\o_Rx_DV_N_3261[24] ), .I2(n29), 
            .I3(n23), .O(n59756));   // verilog/uart_rx.v(53[7] 144[14])
    defparam i46084_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i46090_4_lut (.I0(n59765), .I1(\o_Rx_DV_N_3261[24] ), .I2(n29), 
            .I3(n23), .O(n59762));   // verilog/uart_rx.v(53[7] 144[14])
    defparam i46090_4_lut.LUT_INIT = 16'h0002;
    SB_LUT4 r_SM_Main_2__I_0_62_Mux_1_i3_4_lut (.I0(n59762), .I1(n59756), 
            .I2(\r_SM_Main[1] ), .I3(n27), .O(n3_adj_4949));   // verilog/uart_rx.v(53[7] 144[14])
    defparam r_SM_Main_2__I_0_62_Mux_1_i3_4_lut.LUT_INIT = 16'hf0ca;
    SB_LUT4 i42100_1_lut_2_lut (.I0(baudrate[8]), .I1(n56800), .I2(GND_net), 
            .I3(GND_net), .O(n53913));
    defparam i42100_1_lut_2_lut.LUT_INIT = 16'h1111;
    SB_LUT4 i42101_2_lut_3_lut (.I0(baudrate[7]), .I1(baudrate[8]), .I2(n56800), 
            .I3(GND_net), .O(n56804));
    defparam i42101_2_lut_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i48535_2_lut_4_lut (.I0(n62799), .I1(baudrate[18]), .I2(n2713), 
            .I3(n22498), .O(n294[5]));   // verilog/uart_rx.v(119[33:55])
    defparam i48535_2_lut_4_lut.LUT_INIT = 16'h0071;
    SB_LUT4 i1_2_lut_4_lut_adj_1005 (.I0(n62799), .I1(baudrate[18]), .I2(n2713), 
            .I3(n55688), .O(n2845));   // verilog/uart_rx.v(119[33:55])
    defparam i1_2_lut_4_lut_adj_1005.LUT_INIT = 16'h7100;
    SB_LUT4 i48506_2_lut_4_lut (.I0(n62298), .I1(baudrate[8]), .I2(n1408), 
            .I3(n56800), .O(n294[15]));   // verilog/uart_rx.v(119[33:55])
    defparam i48506_2_lut_4_lut.LUT_INIT = 16'h0071;
    SB_LUT4 i48084_4_lut (.I0(n61292), .I1(n62338), .I2(n45_adj_4858), 
            .I3(n60805), .O(n62797));   // verilog/uart_rx.v(119[33:55])
    defparam i48084_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i1_2_lut_4_lut_adj_1006 (.I0(n62298), .I1(baudrate[8]), .I2(n1408), 
            .I3(n55676), .O(n1560));   // verilog/uart_rx.v(119[33:55])
    defparam i1_2_lut_4_lut_adj_1006.LUT_INIT = 16'h7100;
    SB_LUT4 i46577_3_lut (.I0(n62534), .I1(baudrate[12]), .I2(n35_adj_4945), 
            .I3(GND_net), .O(n61290));   // verilog/uart_rx.v(119[33:55])
    defparam i46577_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1142_3_lut (.I0(n1560), .I1(n7468[15]), .I2(n294[14]), 
            .I3(GND_net), .O(n1701));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1142_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i48086_4_lut (.I0(n61290), .I1(n62797), .I2(n45_adj_4858), 
            .I3(n62491), .O(n62799));   // verilog/uart_rx.v(119[33:55])
    defparam i48086_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 div_37_i1235_3_lut (.I0(n1701), .I1(n7494[15]), .I2(n294[13]), 
            .I3(GND_net), .O(n1839));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1235_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1326_3_lut (.I0(n1839), .I1(n7520[15]), .I2(n294[12]), 
            .I3(GND_net), .O(n1974));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1326_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1415_3_lut (.I0(n1974), .I1(n7546[15]), .I2(n294[11]), 
            .I3(GND_net), .O(n2106));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1415_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1827_3_lut (.I0(n2601), .I1(n7676[18]), .I2(n294[6]), 
            .I3(GND_net), .O(n2718));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1827_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1502_3_lut (.I0(n2106), .I1(n7572[15]), .I2(n294[10]), 
            .I3(GND_net), .O(n2235));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1502_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2161_1_lut (.I0(baudrate[14]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n2519));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2161_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_37_i1587_3_lut (.I0(n2235), .I1(n7598[15]), .I2(n294[9]), 
            .I3(GND_net), .O(n2361));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1587_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1904_3_lut (.I0(n2718), .I1(n7702[18]), .I2(n294[5]), 
            .I3(GND_net), .O(n2832));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1904_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1670_3_lut (.I0(n2361), .I1(n7624[15]), .I2(n294[8]), 
            .I3(GND_net), .O(n2484));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1670_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1751_3_lut (.I0(n2484), .I1(n7650[15]), .I2(n294[7]), 
            .I3(GND_net), .O(n2604));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1751_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1830_3_lut (.I0(n2604), .I1(n7676[15]), .I2(n294[6]), 
            .I3(GND_net), .O(n2721));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1830_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1845_i31_2_lut (.I0(n2721), .I1(baudrate[10]), 
            .I2(GND_net), .I3(GND_net), .O(n31_adj_4943));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1845_i31_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i6_2_lut (.I0(baudrate[10]), .I1(baudrate[11]), .I2(GND_net), 
            .I3(GND_net), .O(n24_adj_4901));
    defparam i6_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i2108_3_lut (.I0(r_Bit_Index[2]), .I1(r_Bit_Index[1]), .I2(\r_Bit_Index[0] ), 
            .I3(GND_net), .O(n479[2]));   // verilog/uart_rx.v(103[36:51])
    defparam i2108_3_lut.LUT_INIT = 16'h6a6a;
    SB_LUT4 i39194_1_lut_4_lut (.I0(n56558), .I1(n56560), .I2(n56356), 
            .I3(n56556), .O(n53859));
    defparam i39194_1_lut_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 div_37_LessThan_1062_i32_3_lut (.I0(baudrate[0]), .I1(baudrate[1]), 
            .I2(n1560), .I3(GND_net), .O(n32_adj_5042));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1062_i32_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i47535_3_lut (.I0(n32_adj_5042), .I1(baudrate[5]), .I2(n39_adj_5023), 
            .I3(GND_net), .O(n62248));   // verilog/uart_rx.v(119[33:55])
    defparam i47535_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i46128_2_lut_4_lut (.I0(n2723), .I1(baudrate[8]), .I2(n2727), 
            .I3(baudrate[4]), .O(n60840));
    defparam i46128_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 i1_4_lut_adj_1007 (.I0(r_Clock_Count[1]), .I1(r_Clock_Count[0]), 
            .I2(\o_Rx_DV_N_3261[2] ), .I3(\o_Rx_DV_N_3261[1] ), .O(n56246));   // verilog/uart_rx.v(69[17:62])
    defparam i1_4_lut_adj_1007.LUT_INIT = 16'h7bde;
    SB_LUT4 i42098_1_lut (.I0(n56800), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n53909));
    defparam i42098_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 equal_257_i3_2_lut (.I0(r_Clock_Count[2]), .I1(\o_Rx_DV_N_3261[3] ), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_5043));   // verilog/uart_rx.v(69[17:62])
    defparam equal_257_i3_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_4_lut_adj_1008 (.I0(r_Clock_Count[3]), .I1(n3_adj_5043), 
            .I2(\o_Rx_DV_N_3261[4] ), .I3(n56246), .O(n56250));   // verilog/uart_rx.v(69[17:62])
    defparam i1_4_lut_adj_1008.LUT_INIT = 16'hffde;
    SB_LUT4 equal_257_i5_2_lut (.I0(r_Clock_Count[4]), .I1(\o_Rx_DV_N_3261[5] ), 
            .I2(GND_net), .I3(GND_net), .O(n5));   // verilog/uart_rx.v(69[17:62])
    defparam equal_257_i5_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i47536_3_lut (.I0(n62248), .I1(baudrate[6]), .I2(n41_adj_5024), 
            .I3(GND_net), .O(n62249));   // verilog/uart_rx.v(119[33:55])
    defparam i47536_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_1009 (.I0(r_Clock_Count[5]), .I1(n5), .I2(\o_Rx_DV_N_3261[6] ), 
            .I3(n56250), .O(n56254));   // verilog/uart_rx.v(69[17:62])
    defparam i1_4_lut_adj_1009.LUT_INIT = 16'hffde;
    SB_LUT4 i39214_1_lut (.I0(n22385), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n53879));
    defparam i39214_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 equal_257_i8_2_lut (.I0(r_Clock_Count[7]), .I1(\o_Rx_DV_N_3261[8] ), 
            .I2(GND_net), .I3(GND_net), .O(n8_adj_5044));   // verilog/uart_rx.v(69[17:62])
    defparam equal_257_i8_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_4_lut_adj_1010 (.I0(r_Clock_Count[6]), .I1(n8_adj_5044), 
            .I2(n56254), .I3(\o_Rx_DV_N_3261[7] ), .O(n52650));   // verilog/uart_rx.v(69[17:62])
    defparam i1_4_lut_adj_1010.LUT_INIT = 16'hfdfe;
    SB_LUT4 i48538_2_lut_4_lut (.I0(n63000), .I1(baudrate[19]), .I2(n2827), 
            .I3(n22501), .O(n294[4]));   // verilog/uart_rx.v(119[33:55])
    defparam i48538_2_lut_4_lut.LUT_INIT = 16'h0071;
    SB_LUT4 i1_2_lut_4_lut_adj_1011 (.I0(n63000), .I1(baudrate[19]), .I2(n2827), 
            .I3(n55690), .O(n2957));   // verilog/uart_rx.v(119[33:55])
    defparam i1_2_lut_4_lut_adj_1011.LUT_INIT = 16'h7100;
    SB_LUT4 i46176_2_lut (.I0(n52650), .I1(r_Rx_Data), .I2(GND_net), .I3(GND_net), 
            .O(n59788));
    defparam i46176_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i46173_4_lut (.I0(n59788), .I1(n29), .I2(n23), .I3(\o_Rx_DV_N_3261[12] ), 
            .O(n59785));
    defparam i46173_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i48499_2_lut_4_lut (.I0(n62568), .I1(baudrate[7]), .I2(n1261), 
            .I3(n56802), .O(n294[16]));   // verilog/uart_rx.v(119[33:55])
    defparam i48499_2_lut_4_lut.LUT_INIT = 16'h0071;
    SB_LUT4 i46678_4_lut (.I0(n41_adj_5024), .I1(n39_adj_5023), .I2(n37_adj_5025), 
            .I3(n60433), .O(n61391));
    defparam i46678_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i45467_4_lut (.I0(n59785), .I1(r_SM_Main[0]), .I2(n27), .I3(\o_Rx_DV_N_3261[24] ), 
            .O(n59782));
    defparam i45467_4_lut.LUT_INIT = 16'hccc8;
    SB_LUT4 i1_2_lut_4_lut_adj_1012 (.I0(n62568), .I1(baudrate[7]), .I2(n1261), 
            .I3(n55674), .O(n1415));   // verilog/uart_rx.v(119[33:55])
    defparam i1_2_lut_4_lut_adj_1012.LUT_INIT = 16'h7100;
    SB_LUT4 i1_2_lut_4_lut_adj_1013 (.I0(n63004), .I1(baudrate[20]), .I2(n2938), 
            .I3(n55692), .O(n3066));   // verilog/uart_rx.v(119[33:55])
    defparam i1_2_lut_4_lut_adj_1013.LUT_INIT = 16'h7100;
    SB_LUT4 i1_2_lut_4_lut_adj_1014 (.I0(n62805), .I1(baudrate[11]), .I2(n1831), 
            .I3(n55678), .O(n1977));   // verilog/uart_rx.v(119[33:55])
    defparam i1_2_lut_4_lut_adj_1014.LUT_INIT = 16'h7100;
    SB_LUT4 i48517_2_lut_4_lut (.I0(n62805), .I1(baudrate[11]), .I2(n1831), 
            .I3(n56792), .O(n294[12]));   // verilog/uart_rx.v(119[33:55])
    defparam i48517_2_lut_4_lut.LUT_INIT = 16'h0071;
    SB_LUT4 i48543_2_lut_4_lut (.I0(n63004), .I1(baudrate[20]), .I2(n2938), 
            .I3(n22476), .O(n294[3]));   // verilog/uart_rx.v(119[33:55])
    defparam i48543_2_lut_4_lut.LUT_INIT = 16'h0071;
    SB_LUT4 i47589_3_lut (.I0(n34_adj_5045), .I1(baudrate[4]), .I2(n37_adj_5025), 
            .I3(GND_net), .O(n62302));   // verilog/uart_rx.v(119[33:55])
    defparam i47589_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i39202_1_lut_4_lut (.I0(n56488), .I1(n56486), .I2(n56490), 
            .I3(n56354), .O(n53867));
    defparam i39202_1_lut_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 i48422_4_lut (.I0(\r_SM_Main[2] ), .I1(n59782), .I2(\r_SM_Main_2__N_3219[1] ), 
            .I3(\r_SM_Main[1] ), .O(n25950));
    defparam i48422_4_lut.LUT_INIT = 16'h0511;
    SB_LUT4 i1_4_lut_adj_1015 (.I0(n52650), .I1(\r_SM_Main[1] ), .I2(r_Rx_Data), 
            .I3(r_SM_Main[0]), .O(n55766));
    defparam i1_4_lut_adj_1015.LUT_INIT = 16'h1000;
    SB_LUT4 i4003_2_lut_3_lut (.I0(baudrate[3]), .I1(n19008), .I2(n9276), 
            .I3(GND_net), .O(n9283));   // verilog/uart_rx.v(119[33:55])
    defparam i4003_2_lut_3_lut.LUT_INIT = 16'h5454;
    SB_LUT4 i3832_2_lut_4_lut (.I0(baudrate[2]), .I1(n805), .I2(baudrate[1]), 
            .I3(baudrate[0]), .O(n9112));   // verilog/uart_rx.v(119[33:55])
    defparam i3832_2_lut_4_lut.LUT_INIT = 16'h0445;
    SB_LUT4 div_37_LessThan_1250_i30_3_lut_3_lut (.I0(baudrate[2]), .I1(baudrate[3]), 
            .I2(n1839), .I3(GND_net), .O(n30_adj_5031));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1250_i30_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i45635_2_lut_4_lut (.I0(n1834), .I1(baudrate[8]), .I2(n1838), 
            .I3(baudrate[4]), .O(n60347));
    defparam i45635_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 div_37_LessThan_1250_i32_3_lut_3_lut (.I0(baudrate[4]), .I1(baudrate[8]), 
            .I2(n1834), .I3(GND_net), .O(n32_adj_5028));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1250_i32_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_LessThan_1845_i18_3_lut_3_lut (.I0(baudrate[4]), .I1(baudrate[8]), 
            .I2(n2723), .I3(GND_net), .O(n18_adj_5038));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1845_i18_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i46555_3_lut (.I0(n62249), .I1(baudrate[7]), .I2(n43_adj_5026), 
            .I3(GND_net), .O(n61268));   // verilog/uart_rx.v(119[33:55])
    defparam i46555_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i47836_4_lut (.I0(n61268), .I1(n62302), .I2(n43_adj_5026), 
            .I3(n61391), .O(n62549));   // verilog/uart_rx.v(119[33:55])
    defparam i47836_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i45458_2_lut_3_lut (.I0(baudrate[1]), .I1(n48_adj_4774), .I2(n22504), 
            .I3(GND_net), .O(n60170));   // verilog/uart_rx.v(119[33:55])
    defparam i45458_2_lut_3_lut.LUT_INIT = 16'h0202;
    SB_LUT4 i1_4_lut_adj_1016 (.I0(n29), .I1(n23), .I2(\o_Rx_DV_N_3261[12] ), 
            .I3(n55766), .O(n55772));
    defparam i1_4_lut_adj_1016.LUT_INIT = 16'h0100;
    SB_LUT4 i48322_4_lut (.I0(\r_SM_Main[2] ), .I1(\o_Rx_DV_N_3261[24] ), 
            .I2(n27), .I3(n55772), .O(n24619));   // verilog/uart_rx.v(53[7] 144[14])
    defparam i48322_4_lut.LUT_INIT = 16'h5455;
    SB_LUT4 i1_3_lut_4_lut_adj_1017 (.I0(n22504), .I1(n48_adj_4774), .I2(baudrate[1]), 
            .I3(baudrate[0]), .O(n44));
    defparam i1_3_lut_4_lut_adj_1017.LUT_INIT = 16'hefff;
    SB_LUT4 i47837_3_lut (.I0(n62549), .I1(baudrate[8]), .I2(n1553), .I3(GND_net), 
            .O(n62550));   // verilog/uart_rx.v(119[33:55])
    defparam i47837_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_LessThan_1062_i48_3_lut (.I0(n62550), .I1(baudrate[9]), 
            .I2(n1552), .I3(GND_net), .O(n48_adj_4988));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1062_i48_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i1_2_lut_4_lut_adj_1018 (.I0(baudrate[6]), .I1(baudrate[7]), 
            .I2(baudrate[8]), .I3(baudrate[9]), .O(n56346));
    defparam i1_2_lut_4_lut_adj_1018.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_4_lut_adj_1019 (.I0(baudrate[28]), .I1(baudrate[26]), 
            .I2(baudrate[24]), .I3(baudrate[31]), .O(n56318));
    defparam i1_2_lut_4_lut_adj_1019.LUT_INIT = 16'hfffe;
    SB_LUT4 div_37_LessThan_1341_i28_3_lut_3_lut (.I0(baudrate[2]), .I1(baudrate[3]), 
            .I2(n1975), .I3(GND_net), .O(n28_adj_5003));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1341_i28_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_i1236_3_lut (.I0(n1702), .I1(n7494[14]), .I2(n294[13]), 
            .I3(GND_net), .O(n1840));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1236_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_4_lut_adj_1020 (.I0(n62401), .I1(baudrate[21]), .I2(n3046), 
            .I3(n55694), .O(n3172));   // verilog/uart_rx.v(119[33:55])
    defparam i1_2_lut_4_lut_adj_1020.LUT_INIT = 16'h7100;
    SB_LUT4 i45603_2_lut_4_lut (.I0(n1970), .I1(baudrate[8]), .I2(n1974), 
            .I3(baudrate[4]), .O(n60315));
    defparam i45603_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 div_37_LessThan_1341_i30_3_lut_3_lut (.I0(baudrate[4]), .I1(baudrate[8]), 
            .I2(n1970), .I3(GND_net), .O(n30_adj_4999));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1341_i30_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_i1327_3_lut (.I0(n1840), .I1(n7520[14]), .I2(n294[12]), 
            .I3(GND_net), .O(n1975));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1327_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i48550_2_lut_4_lut (.I0(n62401), .I1(baudrate[21]), .I2(n3046), 
            .I3(n22481), .O(n294[2]));   // verilog/uart_rx.v(119[33:55])
    defparam i48550_2_lut_4_lut.LUT_INIT = 16'h0071;
    SB_LUT4 div_37_i1416_3_lut (.I0(n1975), .I1(n7546[14]), .I2(n294[11]), 
            .I3(GND_net), .O(n2107));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1416_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i42035_2_lut_3_lut_4_lut (.I0(baudrate[5]), .I1(baudrate[6]), 
            .I2(baudrate[8]), .I3(baudrate[7]), .O(n56738));
    defparam i42035_2_lut_3_lut_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i48509_2_lut_3_lut_4_lut (.I0(baudrate[10]), .I1(baudrate[11]), 
            .I2(n56792), .I3(n48_adj_4988), .O(n294[14]));
    defparam i48509_2_lut_3_lut_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 i42097_2_lut_3_lut_4_lut (.I0(baudrate[10]), .I1(baudrate[11]), 
            .I2(n56792), .I3(baudrate[9]), .O(n56800));
    defparam i42097_2_lut_3_lut_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i42111_2_lut_3_lut (.I0(baudrate[5]), .I1(baudrate[6]), .I2(n56804), 
            .I3(GND_net), .O(n56814));
    defparam i42111_2_lut_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i1_2_lut_4_lut_adj_1021 (.I0(baudrate[30]), .I1(baudrate[25]), 
            .I2(baudrate[24]), .I3(baudrate[29]), .O(n56376));
    defparam i1_2_lut_4_lut_adj_1021.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_3_lut_4_lut_adj_1022 (.I0(baudrate[7]), .I1(baudrate[8]), 
            .I2(baudrate[10]), .I3(baudrate[9]), .O(n56180));
    defparam i1_3_lut_4_lut_adj_1022.LUT_INIT = 16'hfffe;
    SB_LUT4 i45721_3_lut_4_lut (.I0(n1558), .I1(baudrate[3]), .I2(baudrate[2]), 
            .I3(n1559), .O(n60433));   // verilog/uart_rx.v(119[33:55])
    defparam i45721_3_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 div_37_LessThan_1062_i34_3_lut_3_lut (.I0(n1558), .I1(baudrate[3]), 
            .I2(baudrate[2]), .I3(GND_net), .O(n34_adj_5045));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1062_i34_3_lut_3_lut.LUT_INIT = 16'hd4d4;
    SB_LUT4 i45737_3_lut_4_lut (.I0(n1413), .I1(baudrate[3]), .I2(baudrate[2]), 
            .I3(n1414), .O(n60449));   // verilog/uart_rx.v(119[33:55])
    defparam i45737_3_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 div_37_LessThan_965_i36_3_lut_3_lut (.I0(n1413), .I1(baudrate[3]), 
            .I2(baudrate[2]), .I3(GND_net), .O(n36_adj_5040));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_965_i36_3_lut_3_lut.LUT_INIT = 16'hd4d4;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1023 (.I0(baudrate[16]), .I1(baudrate[17]), 
            .I2(baudrate[18]), .I3(baudrate[19]), .O(n56416));
    defparam i1_2_lut_3_lut_4_lut_adj_1023.LUT_INIT = 16'hfffe;
    SB_LUT4 i10_2_lut_3_lut_4_lut (.I0(baudrate[2]), .I1(baudrate[3]), .I2(baudrate[1]), 
            .I3(baudrate[0]), .O(n28_adj_5046));
    defparam i10_2_lut_3_lut_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 div_37_LessThan_866_i38_3_lut_3_lut (.I0(n1265), .I1(baudrate[3]), 
            .I2(baudrate[2]), .I3(GND_net), .O(n38_adj_4822));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_866_i38_3_lut_3_lut.LUT_INIT = 16'hd4d4;
    SB_LUT4 i45747_3_lut_4_lut (.I0(n1265), .I1(baudrate[3]), .I2(baudrate[2]), 
            .I3(n1266), .O(n60459));   // verilog/uart_rx.v(119[33:55])
    defparam i45747_3_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 i48319_2_lut_3_lut_4_lut (.I0(\r_SM_Main_2__N_3219[1] ), .I1(\r_SM_Main[1] ), 
            .I2(r_SM_Main[0]), .I3(\r_SM_Main[2] ), .O(n24621));
    defparam i48319_2_lut_3_lut_4_lut.LUT_INIT = 16'h0007;
    SB_LUT4 i45698_3_lut_4_lut (.I0(n1699), .I1(baudrate[4]), .I2(baudrate[3]), 
            .I3(n1700), .O(n60410));   // verilog/uart_rx.v(119[33:55])
    defparam i45698_3_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 i1_2_lut_adj_1024 (.I0(baudrate[18]), .I1(baudrate[19]), .I2(GND_net), 
            .I3(GND_net), .O(n56464));
    defparam i1_2_lut_adj_1024.LUT_INIT = 16'heeee;
    SB_LUT4 i46154_4_lut (.I0(\o_Rx_DV_N_3261[8] ), .I1(\o_Rx_DV_N_3261[12] ), 
            .I2(n4834), .I3(n52823), .O(n59876));
    defparam i46154_4_lut.LUT_INIT = 16'h0100;
    SB_LUT4 i46145_4_lut (.I0(n59876), .I1(\o_Rx_DV_N_3261[24] ), .I2(n29), 
            .I3(n23), .O(n59873));
    defparam i46145_4_lut.LUT_INIT = 16'h0002;
    SB_LUT4 i14_4_lut (.I0(\r_SM_Main[1] ), .I1(n59873), .I2(r_SM_Main[0]), 
            .I3(n27), .O(n24535));
    defparam i14_4_lut.LUT_INIT = 16'h05c5;
    SB_LUT4 div_37_LessThan_1157_i34_3_lut_3_lut (.I0(n1699), .I1(baudrate[4]), 
            .I2(baudrate[3]), .I3(GND_net), .O(n34_adj_5012));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1157_i34_3_lut_3_lut.LUT_INIT = 16'hd4d4;
    SB_LUT4 div_37_LessThan_1430_i28_3_lut_3_lut (.I0(baudrate[3]), .I1(baudrate[4]), 
            .I2(n2107), .I3(GND_net), .O(n28_adj_4983));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1430_i28_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i45515_2_lut_4_lut (.I0(n2102), .I1(baudrate[9]), .I2(n2106), 
            .I3(baudrate[5]), .O(n60227));
    defparam i45515_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 div_37_LessThan_1430_i30_3_lut_3_lut (.I0(baudrate[5]), .I1(baudrate[9]), 
            .I2(n2102), .I3(GND_net), .O(n30_adj_4980));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1430_i30_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i16_4_lut (.I0(n31_adj_4905), .I1(baudrate[16]), .I2(n28_adj_5046), 
            .I3(n22473), .O(n34));
    defparam i16_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 div_37_LessThan_1845_i20_3_lut_3_lut (.I0(baudrate[5]), .I1(baudrate[6]), 
            .I2(n2725), .I3(GND_net), .O(n20_adj_5009));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1845_i20_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i1_3_lut_4_lut_adj_1025 (.I0(baudrate[14]), .I1(baudrate[2]), 
            .I2(baudrate[1]), .I3(baudrate[0]), .O(n56118));
    defparam i1_3_lut_4_lut_adj_1025.LUT_INIT = 16'h1000;
    SB_LUT4 i2_3_lut (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[2]), .I2(\r_Bit_Index[0] ), 
            .I3(GND_net), .O(n55461));
    defparam i2_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 i1_4_lut_adj_1026 (.I0(n56428), .I1(n56430), .I2(n56308), 
            .I3(n56484), .O(n56448));
    defparam i1_4_lut_adj_1026.LUT_INIT = 16'hfffe;
    SB_LUT4 i2_2_lut (.I0(r_SM_Main[0]), .I1(\r_SM_Main[2] ), .I2(GND_net), 
            .I3(GND_net), .O(n6_adj_4985));
    defparam i2_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i1_3_lut_4_lut_adj_1027 (.I0(n56710), .I1(n56786), .I2(n7546[11]), 
            .I3(n48_adj_5008), .O(n2110));
    defparam i1_3_lut_4_lut_adj_1027.LUT_INIT = 16'h0010;
    SB_LUT4 i1_3_lut_adj_1028 (.I0(n56416), .I1(n56448), .I2(n56274), 
            .I3(GND_net), .O(n22470));
    defparam i1_3_lut_adj_1028.LUT_INIT = 16'hfefe;
    SB_LUT4 i1_2_lut_4_lut_adj_1029 (.I0(baudrate[22]), .I1(baudrate[23]), 
            .I2(baudrate[25]), .I3(baudrate[28]), .O(n56470));
    defparam i1_2_lut_4_lut_adj_1029.LUT_INIT = 16'hfffe;
    SB_LUT4 div_37_i1503_3_lut (.I0(n2107), .I1(n7572[14]), .I2(n294[10]), 
            .I3(GND_net), .O(n2236));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1503_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1517_i24_3_lut_3_lut (.I0(baudrate[2]), .I1(baudrate[3]), 
            .I2(n2238), .I3(GND_net), .O(n24_adj_4966));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1517_i24_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i45454_2_lut_4_lut (.I0(n2233), .I1(baudrate[8]), .I2(n2237), 
            .I3(baudrate[4]), .O(n60166));
    defparam i45454_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 i5706_4_lut_4_lut (.I0(n960), .I1(n9276), .I2(n19008), .I3(baudrate[3]), 
            .O(n19010));   // verilog/uart_rx.v(119[33:55])
    defparam i5706_4_lut_4_lut.LUT_INIT = 16'ha8aa;
    SB_LUT4 div_37_LessThan_1517_i26_3_lut_3_lut (.I0(baudrate[4]), .I1(baudrate[8]), 
            .I2(n2233), .I3(GND_net), .O(n26_adj_4964));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1517_i26_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i1_3_lut_4_lut_adj_1030 (.I0(baudrate[20]), .I1(baudrate[21]), 
            .I2(n56484), .I3(n56358), .O(n56156));
    defparam i1_3_lut_4_lut_adj_1030.LUT_INIT = 16'hfffe;
    SB_LUT4 div_37_i1588_3_lut (.I0(n2236), .I1(n7598[14]), .I2(n294[9]), 
            .I3(GND_net), .O(n2362));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1588_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1671_3_lut (.I0(n2362), .I1(n7624[14]), .I2(n294[8]), 
            .I3(GND_net), .O(n2485));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1671_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i45475_2_lut_4_lut (.I0(n2235), .I1(baudrate[6]), .I2(n2236), 
            .I3(baudrate[5]), .O(n60187));
    defparam i45475_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 div_37_LessThan_1517_i28_3_lut_3_lut (.I0(baudrate[5]), .I1(baudrate[6]), 
            .I2(n2235), .I3(GND_net), .O(n28_adj_4962));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1517_i28_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_i1752_3_lut (.I0(n2485), .I1(n7650[14]), .I2(n294[7]), 
            .I3(GND_net), .O(n2605));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1752_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_3_lut_4_lut_adj_1031 (.I0(baudrate[25]), .I1(baudrate[28]), 
            .I2(baudrate[26]), .I3(baudrate[29]), .O(n56208));
    defparam i1_3_lut_4_lut_adj_1031.LUT_INIT = 16'hfffe;
    SB_LUT4 i39222_1_lut_3_lut (.I0(n56416), .I1(n56448), .I2(n56274), 
            .I3(GND_net), .O(n53887));
    defparam i39222_1_lut_3_lut.LUT_INIT = 16'h0101;
    SB_LUT4 i1_3_lut_4_lut_adj_1032 (.I0(baudrate[30]), .I1(baudrate[31]), 
            .I2(baudrate[24]), .I3(baudrate[27]), .O(n56206));
    defparam i1_3_lut_4_lut_adj_1032.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_4_lut_adj_1033 (.I0(baudrate[10]), .I1(baudrate[11]), 
            .I2(baudrate[12]), .I3(baudrate[13]), .O(n56344));
    defparam i1_2_lut_4_lut_adj_1033.LUT_INIT = 16'hfffe;
    SB_LUT4 i46080_2_lut_4_lut (.I0(n2715), .I1(baudrate[16]), .I2(n2724), 
            .I3(baudrate[7]), .O(n60792));
    defparam i46080_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 div_37_LessThan_1845_i22_3_lut_3_lut (.I0(baudrate[7]), .I1(baudrate[16]), 
            .I2(n2715), .I3(GND_net), .O(n22_adj_5004));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1845_i22_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i45468_2_lut_3_lut (.I0(baudrate[1]), .I1(n48_adj_4904), .I2(n22484), 
            .I3(GND_net), .O(n60180));   // verilog/uart_rx.v(119[33:55])
    defparam i45468_2_lut_3_lut.LUT_INIT = 16'h0202;
    SB_LUT4 div_37_LessThan_1685_i20_3_lut_3_lut (.I0(baudrate[2]), .I1(baudrate[3]), 
            .I2(n2489), .I3(GND_net), .O(n20_adj_4935));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1685_i20_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i45296_2_lut_4_lut (.I0(n2484), .I1(baudrate[8]), .I2(n2488), 
            .I3(baudrate[4]), .O(n60008));
    defparam i45296_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 i1_3_lut_4_lut_adj_1034 (.I0(baudrate[15]), .I1(baudrate[17]), 
            .I2(baudrate[18]), .I3(baudrate[16]), .O(n56176));
    defparam i1_3_lut_4_lut_adj_1034.LUT_INIT = 16'hfffe;
    SB_LUT4 div_37_LessThan_1685_i22_3_lut_3_lut (.I0(baudrate[4]), .I1(baudrate[8]), 
            .I2(n2484), .I3(GND_net), .O(n22_adj_4933));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1685_i22_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_i1831_3_lut (.I0(n2605), .I1(n7676[14]), .I2(n294[6]), 
            .I3(GND_net), .O(n2722));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1831_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1845_i29_2_lut (.I0(n2722), .I1(baudrate[9]), 
            .I2(GND_net), .I3(GND_net), .O(n29_adj_4944));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1845_i29_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1685_i24_3_lut_3_lut (.I0(baudrate[5]), .I1(baudrate[6]), 
            .I2(n2486), .I3(GND_net), .O(n24_adj_4928));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1685_i24_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i45309_2_lut_4_lut (.I0(n2486), .I1(baudrate[6]), .I2(n2487), 
            .I3(baudrate[5]), .O(n60021));
    defparam i45309_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 i3996_2_lut_3_lut (.I0(baudrate[2]), .I1(n962), .I2(baudrate[1]), 
            .I3(GND_net), .O(n9276));   // verilog/uart_rx.v(119[33:55])
    defparam i3996_2_lut_3_lut.LUT_INIT = 16'h4545;
    SB_LUT4 i3827_2_lut_3_lut (.I0(n805), .I1(baudrate[1]), .I2(baudrate[0]), 
            .I3(GND_net), .O(n42));   // verilog/uart_rx.v(119[33:55])
    defparam i3827_2_lut_3_lut.LUT_INIT = 16'h2b2b;
    SB_LUT4 i1_2_lut_adj_1035 (.I0(baudrate[3]), .I1(baudrate[4]), .I2(GND_net), 
            .I3(GND_net), .O(n56174));
    defparam i1_2_lut_adj_1035.LUT_INIT = 16'heeee;
    SB_LUT4 i2101_2_lut (.I0(r_Bit_Index[1]), .I1(\r_Bit_Index[0] ), .I2(GND_net), 
            .I3(GND_net), .O(n479[1]));   // verilog/uart_rx.v(103[36:51])
    defparam i2101_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i48437_2_lut (.I0(baudrate[1]), .I1(n56818), .I2(GND_net), 
            .I3(GND_net), .O(n294[23]));
    defparam i48437_2_lut.LUT_INIT = 16'h1111;
    SB_LUT4 i48496_2_lut_4_lut (.I0(n62786), .I1(baudrate[6]), .I2(n1111), 
            .I3(n56804), .O(n294[17]));   // verilog/uart_rx.v(119[33:55])
    defparam i48496_2_lut_4_lut.LUT_INIT = 16'h0071;
    SB_LUT4 i1_2_lut_4_lut_adj_1036 (.I0(n62786), .I1(baudrate[6]), .I2(n1111), 
            .I3(n55672), .O(n1267));   // verilog/uart_rx.v(119[33:55])
    defparam i1_2_lut_4_lut_adj_1036.LUT_INIT = 16'h7100;
    SB_LUT4 i48428_2_lut (.I0(n48_adj_4774), .I1(n22504), .I2(GND_net), 
            .I3(GND_net), .O(n294[21]));
    defparam i48428_2_lut.LUT_INIT = 16'h1111;
    SB_LUT4 i42045_4_lut (.I0(baudrate[29]), .I1(baudrate[25]), .I2(baudrate[31]), 
            .I3(baudrate[24]), .O(n56748));
    defparam i42045_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 div_37_LessThan_1766_i18_3_lut_3_lut (.I0(baudrate[2]), .I1(baudrate[3]), 
            .I2(n2610), .I3(GND_net), .O(n18_adj_4909));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1766_i18_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_LessThan_765_i40_3_lut_3_lut (.I0(n1114), .I1(baudrate[3]), 
            .I2(baudrate[2]), .I3(GND_net), .O(n40_adj_4978));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_765_i40_3_lut_3_lut.LUT_INIT = 16'hd4d4;
    SB_LUT4 i45243_2_lut_4_lut (.I0(n2605), .I1(baudrate[8]), .I2(n2609), 
            .I3(baudrate[4]), .O(n59955));
    defparam i45243_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 div_37_LessThan_1766_i20_3_lut_3_lut (.I0(baudrate[4]), .I1(baudrate[8]), 
            .I2(n2605), .I3(GND_net), .O(n20_adj_4907));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1766_i20_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i45757_3_lut_4_lut (.I0(n1114), .I1(baudrate[3]), .I2(baudrate[2]), 
            .I3(n1115), .O(n60469));   // verilog/uart_rx.v(119[33:55])
    defparam i45757_3_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 div_37_LessThan_1766_i22_3_lut_3_lut (.I0(baudrate[5]), .I1(baudrate[6]), 
            .I2(n2607), .I3(GND_net), .O(n22_adj_4906));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1766_i22_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i1_4_lut_adj_1037 (.I0(baudrate[28]), .I1(n56160), .I2(n56554), 
            .I3(baudrate[1]), .O(n56080));
    defparam i1_4_lut_adj_1037.LUT_INIT = 16'h0100;
    SB_LUT4 i5600_2_lut_3_lut (.I0(n805), .I1(baudrate[1]), .I2(baudrate[0]), 
            .I3(GND_net), .O(n18896));   // verilog/uart_rx.v(119[33:55])
    defparam i5600_2_lut_3_lut.LUT_INIT = 16'h2a2a;
    SB_LUT4 i46170_2_lut_3_lut (.I0(n22504), .I1(baudrate[1]), .I2(baudrate[0]), 
            .I3(GND_net), .O(n59864));   // verilog/uart_rx.v(119[33:55])
    defparam i46170_2_lut_3_lut.LUT_INIT = 16'h4040;
    SB_LUT4 div_37_LessThan_1602_i22_3_lut_3_lut (.I0(baudrate[2]), .I1(baudrate[3]), 
            .I2(n2365), .I3(GND_net), .O(n22_adj_4896));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1602_i22_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i42065_4_lut (.I0(baudrate[16]), .I1(n56748), .I2(baudrate[23]), 
            .I3(baudrate[27]), .O(n56768));
    defparam i42065_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_3_lut_4_lut_adj_1038 (.I0(baudrate[14]), .I1(baudrate[15]), 
            .I2(n56452), .I3(n56358), .O(n56418));
    defparam i1_3_lut_4_lut_adj_1038.LUT_INIT = 16'hfffe;
    SB_LUT4 i42063_4_lut (.I0(baudrate[9]), .I1(n24_adj_4901), .I2(baudrate[21]), 
            .I3(baudrate[22]), .O(n56766));
    defparam i42063_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i45373_2_lut_4_lut (.I0(n2360), .I1(baudrate[8]), .I2(n2364), 
            .I3(baudrate[4]), .O(n60085));
    defparam i45373_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 i42061_4_lut (.I0(baudrate[2]), .I1(n56174), .I2(baudrate[19]), 
            .I3(baudrate[20]), .O(n56764));
    defparam i42061_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1039 (.I0(n56766), .I1(n56768), .I2(n31_adj_4905), 
            .I3(n56080), .O(n56098));
    defparam i1_4_lut_adj_1039.LUT_INIT = 16'h0100;
    SB_LUT4 div_37_LessThan_1602_i24_3_lut_3_lut (.I0(baudrate[4]), .I1(baudrate[8]), 
            .I2(n2360), .I3(GND_net), .O(n24_adj_4893));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1602_i24_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i1_rep_33_4_lut (.I0(n35725), .I1(n56098), .I2(n56764), .I3(n56738), 
            .O(n54397));   // verilog/uart_rx.v(119[33:55])
    defparam i1_rep_33_4_lut.LUT_INIT = 16'haaae;
    SB_LUT4 div_37_LessThan_1922_i14_3_lut_3_lut (.I0(baudrate[2]), .I1(baudrate[3]), 
            .I2(n2843), .I3(GND_net), .O(n14_adj_4892));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1922_i14_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i46043_2_lut_4_lut (.I0(n2838), .I1(baudrate[8]), .I2(n2842), 
            .I3(baudrate[4]), .O(n60755));
    defparam i46043_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 div_37_LessThan_1922_i16_3_lut_3_lut (.I0(baudrate[4]), .I1(baudrate[8]), 
            .I2(n2838), .I3(GND_net), .O(n16_adj_4890));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1922_i16_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_LessThan_1922_i18_3_lut_3_lut (.I0(baudrate[5]), .I1(baudrate[6]), 
            .I2(n2840), .I3(GND_net), .O(n18_adj_4888));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1922_i18_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i46000_2_lut_4_lut (.I0(n2830), .I1(baudrate[16]), .I2(n2839), 
            .I3(baudrate[7]), .O(n60712));
    defparam i46000_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 div_37_LessThan_1922_i20_3_lut_3_lut (.I0(baudrate[7]), .I1(baudrate[16]), 
            .I2(n2830), .I3(GND_net), .O(n20_adj_4886));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1922_i20_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i45251_2_lut_4_lut (.I0(n2607), .I1(baudrate[6]), .I2(n2608), 
            .I3(baudrate[5]), .O(n59963));
    defparam i45251_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 i45397_2_lut_4_lut (.I0(n2362), .I1(baudrate[6]), .I2(n2363), 
            .I3(baudrate[5]), .O(n60109));
    defparam i45397_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 div_37_LessThan_1602_i26_3_lut_3_lut (.I0(baudrate[5]), .I1(baudrate[6]), 
            .I2(n2362), .I3(GND_net), .O(n26));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1602_i26_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i48431_2_lut_4_lut (.I0(n62891), .I1(baudrate[13]), .I2(n2098), 
            .I3(n22464), .O(n294[10]));   // verilog/uart_rx.v(119[33:55])
    defparam i48431_2_lut_4_lut.LUT_INIT = 16'h0071;
    SB_LUT4 div_37_LessThan_1997_i12_3_lut_3_lut (.I0(baudrate[2]), .I1(baudrate[3]), 
            .I2(n2955), .I3(GND_net), .O(n12_adj_4845));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1997_i12_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i48413_2_lut (.I0(n48_adj_4904), .I1(n22484), .I2(GND_net), 
            .I3(GND_net), .O(n294[20]));   // verilog/uart_rx.v(119[33:55])
    defparam i48413_2_lut.LUT_INIT = 16'h1111;
    SB_LUT4 i45963_2_lut_4_lut (.I0(n2950), .I1(baudrate[8]), .I2(n2954), 
            .I3(baudrate[4]), .O(n60675));
    defparam i45963_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 div_37_LessThan_1997_i14_3_lut_3_lut (.I0(baudrate[4]), .I1(baudrate[8]), 
            .I2(n2950), .I3(GND_net), .O(n14_adj_4844));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1997_i14_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_LessThan_1997_i16_3_lut_3_lut (.I0(baudrate[5]), .I1(baudrate[6]), 
            .I2(n2952), .I3(GND_net), .O(n16_adj_4843));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1997_i16_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i45906_2_lut_4_lut (.I0(n2942), .I1(baudrate[16]), .I2(n2951), 
            .I3(baudrate[7]), .O(n60618));
    defparam i45906_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 div_37_LessThan_1997_i18_3_lut_3_lut (.I0(baudrate[7]), .I1(baudrate[16]), 
            .I2(n2942), .I3(GND_net), .O(n18));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1997_i18_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i1_2_lut_4_lut_adj_1040 (.I0(baudrate[28]), .I1(baudrate[26]), 
            .I2(baudrate[24]), .I3(baudrate[29]), .O(n56490));
    defparam i1_2_lut_4_lut_adj_1040.LUT_INIT = 16'hfffe;
    SB_LUT4 i48425_2_lut_4_lut (.I0(n62546), .I1(baudrate[10]), .I2(n1693), 
            .I3(n22492), .O(n294[13]));   // verilog/uart_rx.v(119[33:55])
    defparam i48425_2_lut_4_lut.LUT_INIT = 16'h0071;
    SB_LUT4 div_37_LessThan_2070_i10_3_lut_3_lut (.I0(baudrate[2]), .I1(baudrate[3]), 
            .I2(n3064), .I3(GND_net), .O(n10_adj_4818));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2070_i10_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_LessThan_2070_i14_3_lut_3_lut (.I0(baudrate[5]), .I1(baudrate[6]), 
            .I2(n3061), .I3(GND_net), .O(n14_adj_4817));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2070_i14_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i45827_2_lut_4_lut (.I0(n3051), .I1(baudrate[16]), .I2(n3060), 
            .I3(baudrate[7]), .O(n60539));
    defparam i45827_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 div_37_LessThan_2070_i16_3_lut_3_lut (.I0(baudrate[7]), .I1(baudrate[16]), 
            .I2(n3051), .I3(GND_net), .O(n16_adj_4815));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2070_i16_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i3998_2_lut (.I0(n19008), .I1(n9276), .I2(GND_net), .I3(GND_net), 
            .O(n42_adj_4787));   // verilog/uart_rx.v(119[33:55])
    defparam i3998_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 div_37_LessThan_2070_i12_3_lut_3_lut (.I0(baudrate[4]), .I1(baudrate[8]), 
            .I2(n3059), .I3(GND_net), .O(n12_adj_4819));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2070_i12_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i45867_2_lut_4_lut (.I0(n3059), .I1(baudrate[8]), .I2(n3063), 
            .I3(baudrate[4]), .O(n60579));
    defparam i45867_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 i1_3_lut_adj_1041 (.I0(n22444), .I1(n48_adj_4986), .I2(n35471), 
            .I3(GND_net), .O(n54439));
    defparam i1_3_lut_adj_1041.LUT_INIT = 16'hefef;
    SB_LUT4 i39210_1_lut (.I0(n22498), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n53875));
    defparam i39210_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i48553_2_lut_4_lut (.I0(n62762), .I1(baudrate[22]), .I2(n3151), 
            .I3(n22434), .O(n294[1]));
    defparam i48553_2_lut_4_lut.LUT_INIT = 16'h0071;
    SB_LUT4 div_37_LessThan_2141_i8_3_lut_3_lut (.I0(baudrate[2]), .I1(baudrate[3]), 
            .I2(n3170), .I3(GND_net), .O(n8_adj_4793));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2141_i8_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_LessThan_2141_i12_3_lut_3_lut (.I0(baudrate[5]), .I1(baudrate[6]), 
            .I2(n3167), .I3(GND_net), .O(n12_adj_4792));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2141_i12_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i45751_2_lut_4_lut (.I0(n3157), .I1(baudrate[16]), .I2(n3166), 
            .I3(baudrate[7]), .O(n60463));
    defparam i45751_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 div_37_LessThan_2141_i14_3_lut_3_lut (.I0(baudrate[7]), .I1(baudrate[16]), 
            .I2(n3157), .I3(GND_net), .O(n14));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2141_i14_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_i427_4_lut (.I0(n54397), .I1(n54439), .I2(n294[21]), 
            .I3(baudrate[2]), .O(n53644));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i427_4_lut.LUT_INIT = 16'h6a9a;
    SB_LUT4 i48416_2_lut_4_lut (.I0(n62293), .I1(baudrate[5]), .I2(n53648), 
            .I3(n22507), .O(n294[18]));   // verilog/uart_rx.v(119[33:55])
    defparam i48416_2_lut_4_lut.LUT_INIT = 16'h0017;
    SB_LUT4 div_37_LessThan_2141_i10_3_lut_3_lut (.I0(baudrate[4]), .I1(baudrate[8]), 
            .I2(n3165), .I3(GND_net), .O(n10_adj_4794));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2141_i10_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i45791_2_lut_4_lut (.I0(n3165), .I1(baudrate[8]), .I2(n3169), 
            .I3(baudrate[4]), .O(n60503));
    defparam i45791_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 i1_2_lut_3_lut_adj_1042 (.I0(baudrate[26]), .I1(baudrate[30]), 
            .I2(baudrate[23]), .I3(GND_net), .O(n56560));
    defparam i1_2_lut_3_lut_adj_1042.LUT_INIT = 16'hfefe;
    SB_LUT4 i48493_2_lut_4_lut (.I0(n62255), .I1(baudrate[4]), .I2(n53646), 
            .I3(n56814), .O(n294[19]));
    defparam i48493_2_lut_4_lut.LUT_INIT = 16'h0017;
    
endmodule
//
// Verilog Description of module \quadrature_decoder(0) 
//

module \quadrature_decoder(0)  (ENCODER1_B_N_keep, n1543, ENCODER1_A_N_keep, 
            n26242, n1548, n26211, b_prev, n26186, a_prev, position_31__N_3609, 
            encoder1_position, \a_new[1] , \b_new[1] , GND_net, VCC_net, 
            debounce_cnt_N_3606) /* synthesis lattice_noprune=1 */ ;
    input ENCODER1_B_N_keep;
    input n1543;
    input ENCODER1_A_N_keep;
    input n26242;
    output n1548;
    input n26211;
    output b_prev;
    input n26186;
    output a_prev;
    output position_31__N_3609;
    output [31:0]encoder1_position;
    output \a_new[1] ;
    output \b_new[1] ;
    input GND_net;
    input VCC_net;
    output debounce_cnt_N_3606;
    
    wire [1:0]b_new;   // vhdl/quadrature_decoder.vhd(40[9:14])
    wire [1:0]a_new;   // vhdl/quadrature_decoder.vhd(39[9:14])
    wire [31:0]n133;
    
    wire direction_N_3613, n46574, n46573, n46572, n46571, n46570, 
        n46569, n46568, n46567, n46566, n46565, n46564, n46563, 
        n46562, n46561, n46560, n46559, n46558, n46557, n46556, 
        n46555, n46554, n46553, n46552, n46551, n46550, n46549, 
        n46548, n46547, n46546, n46545, n46544;
    
    SB_DFF b_new_i0 (.Q(b_new[0]), .C(n1543), .D(ENCODER1_B_N_keep));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    SB_DFF a_new_i0 (.Q(a_new[0]), .C(n1543), .D(ENCODER1_A_N_keep));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    SB_DFF direction_42 (.Q(n1548), .C(n1543), .D(n26242));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    SB_DFF b_prev_41 (.Q(b_prev), .C(n1543), .D(n26211));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    SB_DFF a_prev_40 (.Q(a_prev), .C(n1543), .D(n26186));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    SB_DFFE position_1936__i0 (.Q(encoder1_position[0]), .C(n1543), .E(position_31__N_3609), 
            .D(n133[0]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFF a_new_i1 (.Q(\a_new[1] ), .C(n1543), .D(a_new[0]));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    SB_DFF b_new_i1 (.Q(\b_new[1] ), .C(n1543), .D(b_new[0]));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    SB_LUT4 position_1936_add_4_33_lut (.I0(GND_net), .I1(direction_N_3613), 
            .I2(encoder1_position[31]), .I3(n46574), .O(n133[31])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1936_add_4_33_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 position_1936_add_4_32_lut (.I0(GND_net), .I1(direction_N_3613), 
            .I2(encoder1_position[30]), .I3(n46573), .O(n133[30])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1936_add_4_32_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1936_add_4_32 (.CI(n46573), .I0(direction_N_3613), 
            .I1(encoder1_position[30]), .CO(n46574));
    SB_LUT4 position_1936_add_4_31_lut (.I0(GND_net), .I1(direction_N_3613), 
            .I2(encoder1_position[29]), .I3(n46572), .O(n133[29])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1936_add_4_31_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1936_add_4_31 (.CI(n46572), .I0(direction_N_3613), 
            .I1(encoder1_position[29]), .CO(n46573));
    SB_LUT4 position_1936_add_4_30_lut (.I0(GND_net), .I1(direction_N_3613), 
            .I2(encoder1_position[28]), .I3(n46571), .O(n133[28])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1936_add_4_30_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1936_add_4_30 (.CI(n46571), .I0(direction_N_3613), 
            .I1(encoder1_position[28]), .CO(n46572));
    SB_LUT4 position_1936_add_4_29_lut (.I0(GND_net), .I1(direction_N_3613), 
            .I2(encoder1_position[27]), .I3(n46570), .O(n133[27])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1936_add_4_29_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1936_add_4_29 (.CI(n46570), .I0(direction_N_3613), 
            .I1(encoder1_position[27]), .CO(n46571));
    SB_LUT4 position_1936_add_4_28_lut (.I0(GND_net), .I1(direction_N_3613), 
            .I2(encoder1_position[26]), .I3(n46569), .O(n133[26])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1936_add_4_28_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1936_add_4_28 (.CI(n46569), .I0(direction_N_3613), 
            .I1(encoder1_position[26]), .CO(n46570));
    SB_LUT4 position_1936_add_4_27_lut (.I0(GND_net), .I1(direction_N_3613), 
            .I2(encoder1_position[25]), .I3(n46568), .O(n133[25])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1936_add_4_27_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1936_add_4_27 (.CI(n46568), .I0(direction_N_3613), 
            .I1(encoder1_position[25]), .CO(n46569));
    SB_LUT4 position_1936_add_4_26_lut (.I0(GND_net), .I1(direction_N_3613), 
            .I2(encoder1_position[24]), .I3(n46567), .O(n133[24])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1936_add_4_26_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1936_add_4_26 (.CI(n46567), .I0(direction_N_3613), 
            .I1(encoder1_position[24]), .CO(n46568));
    SB_LUT4 position_1936_add_4_25_lut (.I0(GND_net), .I1(direction_N_3613), 
            .I2(encoder1_position[23]), .I3(n46566), .O(n133[23])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1936_add_4_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1936_add_4_25 (.CI(n46566), .I0(direction_N_3613), 
            .I1(encoder1_position[23]), .CO(n46567));
    SB_LUT4 position_1936_add_4_24_lut (.I0(GND_net), .I1(direction_N_3613), 
            .I2(encoder1_position[22]), .I3(n46565), .O(n133[22])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1936_add_4_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1936_add_4_24 (.CI(n46565), .I0(direction_N_3613), 
            .I1(encoder1_position[22]), .CO(n46566));
    SB_LUT4 position_1936_add_4_23_lut (.I0(GND_net), .I1(direction_N_3613), 
            .I2(encoder1_position[21]), .I3(n46564), .O(n133[21])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1936_add_4_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1936_add_4_23 (.CI(n46564), .I0(direction_N_3613), 
            .I1(encoder1_position[21]), .CO(n46565));
    SB_LUT4 position_1936_add_4_22_lut (.I0(GND_net), .I1(direction_N_3613), 
            .I2(encoder1_position[20]), .I3(n46563), .O(n133[20])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1936_add_4_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1936_add_4_22 (.CI(n46563), .I0(direction_N_3613), 
            .I1(encoder1_position[20]), .CO(n46564));
    SB_DFFE position_1936__i1 (.Q(encoder1_position[1]), .C(n1543), .E(position_31__N_3609), 
            .D(n133[1]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1936__i2 (.Q(encoder1_position[2]), .C(n1543), .E(position_31__N_3609), 
            .D(n133[2]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_LUT4 position_1936_add_4_21_lut (.I0(GND_net), .I1(direction_N_3613), 
            .I2(encoder1_position[19]), .I3(n46562), .O(n133[19])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1936_add_4_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1936_add_4_21 (.CI(n46562), .I0(direction_N_3613), 
            .I1(encoder1_position[19]), .CO(n46563));
    SB_LUT4 position_1936_add_4_20_lut (.I0(GND_net), .I1(direction_N_3613), 
            .I2(encoder1_position[18]), .I3(n46561), .O(n133[18])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1936_add_4_20_lut.LUT_INIT = 16'hC33C;
    SB_DFFE position_1936__i3 (.Q(encoder1_position[3]), .C(n1543), .E(position_31__N_3609), 
            .D(n133[3]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1936__i4 (.Q(encoder1_position[4]), .C(n1543), .E(position_31__N_3609), 
            .D(n133[4]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1936__i5 (.Q(encoder1_position[5]), .C(n1543), .E(position_31__N_3609), 
            .D(n133[5]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1936__i6 (.Q(encoder1_position[6]), .C(n1543), .E(position_31__N_3609), 
            .D(n133[6]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1936__i7 (.Q(encoder1_position[7]), .C(n1543), .E(position_31__N_3609), 
            .D(n133[7]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1936__i8 (.Q(encoder1_position[8]), .C(n1543), .E(position_31__N_3609), 
            .D(n133[8]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1936__i9 (.Q(encoder1_position[9]), .C(n1543), .E(position_31__N_3609), 
            .D(n133[9]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1936__i10 (.Q(encoder1_position[10]), .C(n1543), .E(position_31__N_3609), 
            .D(n133[10]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1936__i11 (.Q(encoder1_position[11]), .C(n1543), .E(position_31__N_3609), 
            .D(n133[11]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1936__i12 (.Q(encoder1_position[12]), .C(n1543), .E(position_31__N_3609), 
            .D(n133[12]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1936__i13 (.Q(encoder1_position[13]), .C(n1543), .E(position_31__N_3609), 
            .D(n133[13]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1936__i14 (.Q(encoder1_position[14]), .C(n1543), .E(position_31__N_3609), 
            .D(n133[14]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1936__i15 (.Q(encoder1_position[15]), .C(n1543), .E(position_31__N_3609), 
            .D(n133[15]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1936__i16 (.Q(encoder1_position[16]), .C(n1543), .E(position_31__N_3609), 
            .D(n133[16]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1936__i17 (.Q(encoder1_position[17]), .C(n1543), .E(position_31__N_3609), 
            .D(n133[17]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1936__i18 (.Q(encoder1_position[18]), .C(n1543), .E(position_31__N_3609), 
            .D(n133[18]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1936__i19 (.Q(encoder1_position[19]), .C(n1543), .E(position_31__N_3609), 
            .D(n133[19]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1936__i20 (.Q(encoder1_position[20]), .C(n1543), .E(position_31__N_3609), 
            .D(n133[20]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1936__i21 (.Q(encoder1_position[21]), .C(n1543), .E(position_31__N_3609), 
            .D(n133[21]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1936__i22 (.Q(encoder1_position[22]), .C(n1543), .E(position_31__N_3609), 
            .D(n133[22]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1936__i23 (.Q(encoder1_position[23]), .C(n1543), .E(position_31__N_3609), 
            .D(n133[23]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1936__i24 (.Q(encoder1_position[24]), .C(n1543), .E(position_31__N_3609), 
            .D(n133[24]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1936__i25 (.Q(encoder1_position[25]), .C(n1543), .E(position_31__N_3609), 
            .D(n133[25]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1936__i26 (.Q(encoder1_position[26]), .C(n1543), .E(position_31__N_3609), 
            .D(n133[26]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1936__i27 (.Q(encoder1_position[27]), .C(n1543), .E(position_31__N_3609), 
            .D(n133[27]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1936__i28 (.Q(encoder1_position[28]), .C(n1543), .E(position_31__N_3609), 
            .D(n133[28]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1936__i29 (.Q(encoder1_position[29]), .C(n1543), .E(position_31__N_3609), 
            .D(n133[29]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1936__i30 (.Q(encoder1_position[30]), .C(n1543), .E(position_31__N_3609), 
            .D(n133[30]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1936__i31 (.Q(encoder1_position[31]), .C(n1543), .E(position_31__N_3609), 
            .D(n133[31]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_CARRY position_1936_add_4_20 (.CI(n46561), .I0(direction_N_3613), 
            .I1(encoder1_position[18]), .CO(n46562));
    SB_LUT4 position_1936_add_4_19_lut (.I0(GND_net), .I1(direction_N_3613), 
            .I2(encoder1_position[17]), .I3(n46560), .O(n133[17])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1936_add_4_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1936_add_4_19 (.CI(n46560), .I0(direction_N_3613), 
            .I1(encoder1_position[17]), .CO(n46561));
    SB_LUT4 position_1936_add_4_18_lut (.I0(GND_net), .I1(direction_N_3613), 
            .I2(encoder1_position[16]), .I3(n46559), .O(n133[16])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1936_add_4_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1936_add_4_18 (.CI(n46559), .I0(direction_N_3613), 
            .I1(encoder1_position[16]), .CO(n46560));
    SB_LUT4 position_1936_add_4_17_lut (.I0(GND_net), .I1(direction_N_3613), 
            .I2(encoder1_position[15]), .I3(n46558), .O(n133[15])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1936_add_4_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1936_add_4_17 (.CI(n46558), .I0(direction_N_3613), 
            .I1(encoder1_position[15]), .CO(n46559));
    SB_LUT4 position_1936_add_4_16_lut (.I0(GND_net), .I1(direction_N_3613), 
            .I2(encoder1_position[14]), .I3(n46557), .O(n133[14])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1936_add_4_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1936_add_4_16 (.CI(n46557), .I0(direction_N_3613), 
            .I1(encoder1_position[14]), .CO(n46558));
    SB_LUT4 position_1936_add_4_15_lut (.I0(GND_net), .I1(direction_N_3613), 
            .I2(encoder1_position[13]), .I3(n46556), .O(n133[13])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1936_add_4_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1936_add_4_15 (.CI(n46556), .I0(direction_N_3613), 
            .I1(encoder1_position[13]), .CO(n46557));
    SB_LUT4 position_1936_add_4_14_lut (.I0(GND_net), .I1(direction_N_3613), 
            .I2(encoder1_position[12]), .I3(n46555), .O(n133[12])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1936_add_4_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1936_add_4_14 (.CI(n46555), .I0(direction_N_3613), 
            .I1(encoder1_position[12]), .CO(n46556));
    SB_LUT4 position_1936_add_4_13_lut (.I0(GND_net), .I1(direction_N_3613), 
            .I2(encoder1_position[11]), .I3(n46554), .O(n133[11])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1936_add_4_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1936_add_4_13 (.CI(n46554), .I0(direction_N_3613), 
            .I1(encoder1_position[11]), .CO(n46555));
    SB_LUT4 position_1936_add_4_12_lut (.I0(GND_net), .I1(direction_N_3613), 
            .I2(encoder1_position[10]), .I3(n46553), .O(n133[10])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1936_add_4_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1936_add_4_12 (.CI(n46553), .I0(direction_N_3613), 
            .I1(encoder1_position[10]), .CO(n46554));
    SB_LUT4 position_1936_add_4_11_lut (.I0(GND_net), .I1(direction_N_3613), 
            .I2(encoder1_position[9]), .I3(n46552), .O(n133[9])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1936_add_4_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1936_add_4_11 (.CI(n46552), .I0(direction_N_3613), 
            .I1(encoder1_position[9]), .CO(n46553));
    SB_LUT4 position_1936_add_4_10_lut (.I0(GND_net), .I1(direction_N_3613), 
            .I2(encoder1_position[8]), .I3(n46551), .O(n133[8])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1936_add_4_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1936_add_4_10 (.CI(n46551), .I0(direction_N_3613), 
            .I1(encoder1_position[8]), .CO(n46552));
    SB_LUT4 position_1936_add_4_9_lut (.I0(GND_net), .I1(direction_N_3613), 
            .I2(encoder1_position[7]), .I3(n46550), .O(n133[7])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1936_add_4_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1936_add_4_9 (.CI(n46550), .I0(direction_N_3613), 
            .I1(encoder1_position[7]), .CO(n46551));
    SB_LUT4 position_1936_add_4_8_lut (.I0(GND_net), .I1(direction_N_3613), 
            .I2(encoder1_position[6]), .I3(n46549), .O(n133[6])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1936_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1936_add_4_8 (.CI(n46549), .I0(direction_N_3613), 
            .I1(encoder1_position[6]), .CO(n46550));
    SB_LUT4 position_1936_add_4_7_lut (.I0(GND_net), .I1(direction_N_3613), 
            .I2(encoder1_position[5]), .I3(n46548), .O(n133[5])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1936_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1936_add_4_7 (.CI(n46548), .I0(direction_N_3613), 
            .I1(encoder1_position[5]), .CO(n46549));
    SB_LUT4 position_1936_add_4_6_lut (.I0(GND_net), .I1(direction_N_3613), 
            .I2(encoder1_position[4]), .I3(n46547), .O(n133[4])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1936_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1936_add_4_6 (.CI(n46547), .I0(direction_N_3613), 
            .I1(encoder1_position[4]), .CO(n46548));
    SB_LUT4 position_1936_add_4_5_lut (.I0(GND_net), .I1(direction_N_3613), 
            .I2(encoder1_position[3]), .I3(n46546), .O(n133[3])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1936_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1936_add_4_5 (.CI(n46546), .I0(direction_N_3613), 
            .I1(encoder1_position[3]), .CO(n46547));
    SB_LUT4 position_1936_add_4_4_lut (.I0(GND_net), .I1(direction_N_3613), 
            .I2(encoder1_position[2]), .I3(n46545), .O(n133[2])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1936_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1936_add_4_4 (.CI(n46545), .I0(direction_N_3613), 
            .I1(encoder1_position[2]), .CO(n46546));
    SB_LUT4 position_1936_add_4_3_lut (.I0(GND_net), .I1(direction_N_3613), 
            .I2(encoder1_position[1]), .I3(n46544), .O(n133[1])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1936_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1936_add_4_3 (.CI(n46544), .I0(direction_N_3613), 
            .I1(encoder1_position[1]), .CO(n46545));
    SB_LUT4 position_1936_add_4_2_lut (.I0(GND_net), .I1(GND_net), .I2(encoder1_position[0]), 
            .I3(VCC_net), .O(n133[0])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1936_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1936_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(encoder1_position[0]), 
            .CO(n46544));
    SB_LUT4 debounce_cnt_I_920_4_lut (.I0(a_new[0]), .I1(b_new[0]), .I2(\a_new[1] ), 
            .I3(\b_new[1] ), .O(debounce_cnt_N_3606));   // vhdl/quadrature_decoder.vhd(53[8:58])
    defparam debounce_cnt_I_920_4_lut.LUT_INIT = 16'h7bde;
    SB_LUT4 position_31__I_921_4_lut (.I0(a_prev), .I1(b_prev), .I2(\a_new[1] ), 
            .I3(\b_new[1] ), .O(position_31__N_3609));   // vhdl/quadrature_decoder.vhd(63[11:57])
    defparam position_31__I_921_4_lut.LUT_INIT = 16'h7bde;
    SB_LUT4 b_prev_I_0_48_2_lut (.I0(b_prev), .I1(\a_new[1] ), .I2(GND_net), 
            .I3(GND_net), .O(direction_N_3613));   // vhdl/quadrature_decoder.vhd(64[18:37])
    defparam b_prev_I_0_48_2_lut.LUT_INIT = 16'h9999;
    
endmodule
//
// Verilog Description of module pwm
//

module pwm (n2568, pwm_out, clk32MHz, reset, pwm_setpoint, GND_net, 
            VCC_net, \PWMLimit[7] , \setpoint[7] , n15) /* synthesis syn_module_defined=1 */ ;
    input n2568;
    output pwm_out;
    input clk32MHz;
    input reset;
    input [23:0]pwm_setpoint;
    input GND_net;
    input VCC_net;
    input \PWMLimit[7] ;
    input \setpoint[7] ;
    output n15;
    
    wire clk32MHz /* synthesis SET_AS_NETWORK=clk32MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(31[16:24])
    
    wire pwm_out_N_412, n52381;
    wire [23:0]pwm_counter;   // verilog/pwm.v(11[19:30])
    
    wire n39, n41, n45, n43, n37, n29, n31, n23, n25, n35, 
        n33, n11, n13, n15_c, n27, n9, n17, n19, n21, n60376, 
        n59985, n12, n30, n60789, n61583, n61357, n62519, n61811, 
        n62735, n6, n62451, n62452, n16, n24, n60873, n8, n60845, 
        n62212, n62223, n4, n62457, n62458, n59957, n10, n59947, 
        n62645, n28, n62933, n62934, n62823, n60896, n62741, n62215, 
        n62861, n52391, n52393, n52395, n52279, n52119, n52059, 
        n52013, n51971, n51927, n51889, n51857, n51819, n51783, 
        n51751, n51709, n51669, n51629, n51591, n51551, n51511, 
        n51471, n51439, n51399, n46543, n45_adj_4762, n46542, n46541, 
        n46540, n46539, n46538, n46537, n46536, n46535, n46534, 
        n46533, n46532, n46531, n46530, n46529, n46528, n46527, 
        n46526, n46525, n46524, n46523, n46522, n46521, n55155, 
        n16_adj_4764, n55170, n14, n18, n13_adj_4765;
    
    SB_DFFE pwm_out_12 (.Q(pwm_out), .C(clk32MHz), .E(n2568), .D(pwm_out_N_412));   // verilog/pwm.v(16[12] 26[6])
    SB_DFFR pwm_counter_1935__i0 (.Q(pwm_counter[0]), .C(clk32MHz), .D(n52381), 
            .R(reset));   // verilog/pwm.v(17[20:33])
    SB_LUT4 duty_23__I_0_i39_2_lut (.I0(pwm_counter[19]), .I1(pwm_setpoint[19]), 
            .I2(GND_net), .I3(GND_net), .O(n39));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i39_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i41_2_lut (.I0(pwm_counter[20]), .I1(pwm_setpoint[20]), 
            .I2(GND_net), .I3(GND_net), .O(n41));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i41_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i45_2_lut (.I0(pwm_counter[22]), .I1(pwm_setpoint[22]), 
            .I2(GND_net), .I3(GND_net), .O(n45));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i45_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i43_2_lut (.I0(pwm_counter[21]), .I1(pwm_setpoint[21]), 
            .I2(GND_net), .I3(GND_net), .O(n43));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i43_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i37_2_lut (.I0(pwm_counter[18]), .I1(pwm_setpoint[18]), 
            .I2(GND_net), .I3(GND_net), .O(n37));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i37_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i29_2_lut (.I0(pwm_counter[14]), .I1(pwm_setpoint[14]), 
            .I2(GND_net), .I3(GND_net), .O(n29));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i29_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i31_2_lut (.I0(pwm_counter[15]), .I1(pwm_setpoint[15]), 
            .I2(GND_net), .I3(GND_net), .O(n31));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i31_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i23_2_lut (.I0(pwm_counter[11]), .I1(pwm_setpoint[11]), 
            .I2(GND_net), .I3(GND_net), .O(n23));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i23_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i25_2_lut (.I0(pwm_counter[12]), .I1(pwm_setpoint[12]), 
            .I2(GND_net), .I3(GND_net), .O(n25));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i25_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i35_2_lut (.I0(pwm_counter[17]), .I1(pwm_setpoint[17]), 
            .I2(GND_net), .I3(GND_net), .O(n35));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i35_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i33_2_lut (.I0(pwm_counter[16]), .I1(pwm_setpoint[16]), 
            .I2(GND_net), .I3(GND_net), .O(n33));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i33_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i11_2_lut (.I0(pwm_counter[5]), .I1(pwm_setpoint[5]), 
            .I2(GND_net), .I3(GND_net), .O(n11));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i11_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i13_2_lut (.I0(pwm_counter[6]), .I1(pwm_setpoint[6]), 
            .I2(GND_net), .I3(GND_net), .O(n13));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i13_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i15_2_lut (.I0(pwm_counter[7]), .I1(pwm_setpoint[7]), 
            .I2(GND_net), .I3(GND_net), .O(n15_c));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i15_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i27_2_lut (.I0(pwm_counter[13]), .I1(pwm_setpoint[13]), 
            .I2(GND_net), .I3(GND_net), .O(n27));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i27_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i9_2_lut (.I0(pwm_counter[4]), .I1(pwm_setpoint[4]), 
            .I2(GND_net), .I3(GND_net), .O(n9));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i9_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i17_2_lut (.I0(pwm_counter[8]), .I1(pwm_setpoint[8]), 
            .I2(GND_net), .I3(GND_net), .O(n17));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i17_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i19_2_lut (.I0(pwm_counter[9]), .I1(pwm_setpoint[9]), 
            .I2(GND_net), .I3(GND_net), .O(n19));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i19_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i21_2_lut (.I0(pwm_counter[10]), .I1(pwm_setpoint[10]), 
            .I2(GND_net), .I3(GND_net), .O(n21));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i21_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i45664_4_lut (.I0(n21), .I1(n19), .I2(n17), .I3(n9), .O(n60376));
    defparam i45664_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i45273_4_lut (.I0(n27), .I1(n15_c), .I2(n13), .I3(n11), 
            .O(n59985));
    defparam i45273_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 duty_23__I_0_i30_3_lut (.I0(n12), .I1(pwm_setpoint[17]), .I2(n35), 
            .I3(GND_net), .O(n30));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i30_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i46870_4_lut (.I0(n13), .I1(n11), .I2(n9), .I3(n60789), 
            .O(n61583));
    defparam i46870_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i46644_4_lut (.I0(n19), .I1(n17), .I2(n15_c), .I3(n61583), 
            .O(n61357));
    defparam i46644_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i47806_4_lut (.I0(n25), .I1(n23), .I2(n21), .I3(n61357), 
            .O(n62519));
    defparam i47806_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i47098_4_lut (.I0(n31), .I1(n29), .I2(n27), .I3(n62519), 
            .O(n61811));
    defparam i47098_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i48022_4_lut (.I0(n37), .I1(n35), .I2(n33), .I3(n61811), 
            .O(n62735));
    defparam i48022_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i47738_3_lut (.I0(n6), .I1(pwm_setpoint[10]), .I2(n21), .I3(GND_net), 
            .O(n62451));   // verilog/pwm.v(21[8:24])
    defparam i47738_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i47739_3_lut (.I0(n62451), .I1(pwm_setpoint[11]), .I2(n23), 
            .I3(GND_net), .O(n62452));   // verilog/pwm.v(21[8:24])
    defparam i47739_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_i24_3_lut (.I0(n16), .I1(pwm_setpoint[22]), .I2(n45), 
            .I3(GND_net), .O(n24));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i24_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i46161_4_lut (.I0(n43), .I1(n25), .I2(n23), .I3(n60376), 
            .O(n60873));
    defparam i46161_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i47499_4_lut (.I0(n24), .I1(n8), .I2(n45), .I3(n60845), 
            .O(n62212));   // verilog/pwm.v(21[8:24])
    defparam i47499_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i47510_3_lut (.I0(n62452), .I1(pwm_setpoint[12]), .I2(n25), 
            .I3(GND_net), .O(n62223));   // verilog/pwm.v(21[8:24])
    defparam i47510_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_i4_4_lut (.I0(pwm_counter[0]), .I1(pwm_setpoint[1]), 
            .I2(pwm_counter[1]), .I3(pwm_setpoint[0]), .O(n4));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i4_4_lut.LUT_INIT = 16'h4d0c;
    SB_LUT4 i47744_3_lut (.I0(n4), .I1(pwm_setpoint[13]), .I2(n27), .I3(GND_net), 
            .O(n62457));   // verilog/pwm.v(21[8:24])
    defparam i47744_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i47745_3_lut (.I0(n62457), .I1(pwm_setpoint[14]), .I2(n29), 
            .I3(GND_net), .O(n62458));   // verilog/pwm.v(21[8:24])
    defparam i47745_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i45245_4_lut (.I0(n33), .I1(n31), .I2(n29), .I3(n59985), 
            .O(n59957));
    defparam i45245_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i47932_4_lut (.I0(n30), .I1(n10), .I2(n35), .I3(n59947), 
            .O(n62645));   // verilog/pwm.v(21[8:24])
    defparam i47932_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i47504_3_lut (.I0(n62458), .I1(pwm_setpoint[15]), .I2(n31), 
            .I3(GND_net), .O(n28));   // verilog/pwm.v(21[8:24])
    defparam i47504_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i48220_4_lut (.I0(n28), .I1(n62645), .I2(n35), .I3(n59957), 
            .O(n62933));   // verilog/pwm.v(21[8:24])
    defparam i48220_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i48221_3_lut (.I0(n62933), .I1(pwm_setpoint[18]), .I2(n37), 
            .I3(GND_net), .O(n62934));   // verilog/pwm.v(21[8:24])
    defparam i48221_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i48110_3_lut (.I0(n62934), .I1(pwm_setpoint[19]), .I2(n39), 
            .I3(GND_net), .O(n62823));   // verilog/pwm.v(21[8:24])
    defparam i48110_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i46184_4_lut (.I0(n43), .I1(n41), .I2(n39), .I3(n62735), 
            .O(n60896));
    defparam i46184_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i48028_4_lut (.I0(n62223), .I1(n62212), .I2(n45), .I3(n60873), 
            .O(n62741));   // verilog/pwm.v(21[8:24])
    defparam i48028_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i47502_3_lut (.I0(n62823), .I1(pwm_setpoint[20]), .I2(n41), 
            .I3(GND_net), .O(n62215));   // verilog/pwm.v(21[8:24])
    defparam i47502_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i48148_4_lut (.I0(n62215), .I1(n62741), .I2(n45), .I3(n60896), 
            .O(n62861));   // verilog/pwm.v(21[8:24])
    defparam i48148_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i48149_3_lut (.I0(n62861), .I1(pwm_counter[23]), .I2(pwm_setpoint[23]), 
            .I3(GND_net), .O(pwm_out_N_412));   // verilog/pwm.v(21[8:24])
    defparam i48149_3_lut.LUT_INIT = 16'h8e8e;
    SB_DFFR pwm_counter_1935__i1 (.Q(pwm_counter[1]), .C(clk32MHz), .D(n52391), 
            .R(reset));   // verilog/pwm.v(17[20:33])
    SB_DFFR pwm_counter_1935__i2 (.Q(pwm_counter[2]), .C(clk32MHz), .D(n52393), 
            .R(reset));   // verilog/pwm.v(17[20:33])
    SB_DFFR pwm_counter_1935__i3 (.Q(pwm_counter[3]), .C(clk32MHz), .D(n52395), 
            .R(reset));   // verilog/pwm.v(17[20:33])
    SB_DFFR pwm_counter_1935__i4 (.Q(pwm_counter[4]), .C(clk32MHz), .D(n52279), 
            .R(reset));   // verilog/pwm.v(17[20:33])
    SB_DFFR pwm_counter_1935__i5 (.Q(pwm_counter[5]), .C(clk32MHz), .D(n52119), 
            .R(reset));   // verilog/pwm.v(17[20:33])
    SB_DFFR pwm_counter_1935__i6 (.Q(pwm_counter[6]), .C(clk32MHz), .D(n52059), 
            .R(reset));   // verilog/pwm.v(17[20:33])
    SB_DFFR pwm_counter_1935__i7 (.Q(pwm_counter[7]), .C(clk32MHz), .D(n52013), 
            .R(reset));   // verilog/pwm.v(17[20:33])
    SB_DFFR pwm_counter_1935__i8 (.Q(pwm_counter[8]), .C(clk32MHz), .D(n51971), 
            .R(reset));   // verilog/pwm.v(17[20:33])
    SB_DFFR pwm_counter_1935__i9 (.Q(pwm_counter[9]), .C(clk32MHz), .D(n51927), 
            .R(reset));   // verilog/pwm.v(17[20:33])
    SB_DFFR pwm_counter_1935__i10 (.Q(pwm_counter[10]), .C(clk32MHz), .D(n51889), 
            .R(reset));   // verilog/pwm.v(17[20:33])
    SB_DFFR pwm_counter_1935__i11 (.Q(pwm_counter[11]), .C(clk32MHz), .D(n51857), 
            .R(reset));   // verilog/pwm.v(17[20:33])
    SB_DFFR pwm_counter_1935__i12 (.Q(pwm_counter[12]), .C(clk32MHz), .D(n51819), 
            .R(reset));   // verilog/pwm.v(17[20:33])
    SB_DFFR pwm_counter_1935__i13 (.Q(pwm_counter[13]), .C(clk32MHz), .D(n51783), 
            .R(reset));   // verilog/pwm.v(17[20:33])
    SB_DFFR pwm_counter_1935__i14 (.Q(pwm_counter[14]), .C(clk32MHz), .D(n51751), 
            .R(reset));   // verilog/pwm.v(17[20:33])
    SB_DFFR pwm_counter_1935__i15 (.Q(pwm_counter[15]), .C(clk32MHz), .D(n51709), 
            .R(reset));   // verilog/pwm.v(17[20:33])
    SB_DFFR pwm_counter_1935__i16 (.Q(pwm_counter[16]), .C(clk32MHz), .D(n51669), 
            .R(reset));   // verilog/pwm.v(17[20:33])
    SB_DFFR pwm_counter_1935__i17 (.Q(pwm_counter[17]), .C(clk32MHz), .D(n51629), 
            .R(reset));   // verilog/pwm.v(17[20:33])
    SB_DFFR pwm_counter_1935__i18 (.Q(pwm_counter[18]), .C(clk32MHz), .D(n51591), 
            .R(reset));   // verilog/pwm.v(17[20:33])
    SB_DFFR pwm_counter_1935__i19 (.Q(pwm_counter[19]), .C(clk32MHz), .D(n51551), 
            .R(reset));   // verilog/pwm.v(17[20:33])
    SB_DFFR pwm_counter_1935__i20 (.Q(pwm_counter[20]), .C(clk32MHz), .D(n51511), 
            .R(reset));   // verilog/pwm.v(17[20:33])
    SB_DFFR pwm_counter_1935__i21 (.Q(pwm_counter[21]), .C(clk32MHz), .D(n51471), 
            .R(reset));   // verilog/pwm.v(17[20:33])
    SB_DFFR pwm_counter_1935__i22 (.Q(pwm_counter[22]), .C(clk32MHz), .D(n51439), 
            .R(reset));   // verilog/pwm.v(17[20:33])
    SB_DFFR pwm_counter_1935__i23 (.Q(pwm_counter[23]), .C(clk32MHz), .D(n51399), 
            .R(reset));   // verilog/pwm.v(17[20:33])
    SB_LUT4 pwm_counter_1935_add_4_25_lut (.I0(n45_adj_4762), .I1(GND_net), 
            .I2(pwm_counter[23]), .I3(n46543), .O(n51399)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1935_add_4_25_lut.LUT_INIT = 16'h8228;
    SB_LUT4 pwm_counter_1935_add_4_24_lut (.I0(n45_adj_4762), .I1(GND_net), 
            .I2(pwm_counter[22]), .I3(n46542), .O(n51439)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1935_add_4_24_lut.LUT_INIT = 16'h8228;
    SB_CARRY pwm_counter_1935_add_4_24 (.CI(n46542), .I0(GND_net), .I1(pwm_counter[22]), 
            .CO(n46543));
    SB_LUT4 pwm_counter_1935_add_4_23_lut (.I0(n45_adj_4762), .I1(GND_net), 
            .I2(pwm_counter[21]), .I3(n46541), .O(n51471)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1935_add_4_23_lut.LUT_INIT = 16'h8228;
    SB_CARRY pwm_counter_1935_add_4_23 (.CI(n46541), .I0(GND_net), .I1(pwm_counter[21]), 
            .CO(n46542));
    SB_LUT4 pwm_counter_1935_add_4_22_lut (.I0(n45_adj_4762), .I1(GND_net), 
            .I2(pwm_counter[20]), .I3(n46540), .O(n51511)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1935_add_4_22_lut.LUT_INIT = 16'h8228;
    SB_CARRY pwm_counter_1935_add_4_22 (.CI(n46540), .I0(GND_net), .I1(pwm_counter[20]), 
            .CO(n46541));
    SB_LUT4 pwm_counter_1935_add_4_21_lut (.I0(n45_adj_4762), .I1(GND_net), 
            .I2(pwm_counter[19]), .I3(n46539), .O(n51551)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1935_add_4_21_lut.LUT_INIT = 16'h8228;
    SB_CARRY pwm_counter_1935_add_4_21 (.CI(n46539), .I0(GND_net), .I1(pwm_counter[19]), 
            .CO(n46540));
    SB_LUT4 pwm_counter_1935_add_4_20_lut (.I0(n45_adj_4762), .I1(GND_net), 
            .I2(pwm_counter[18]), .I3(n46538), .O(n51591)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1935_add_4_20_lut.LUT_INIT = 16'h8228;
    SB_CARRY pwm_counter_1935_add_4_20 (.CI(n46538), .I0(GND_net), .I1(pwm_counter[18]), 
            .CO(n46539));
    SB_LUT4 pwm_counter_1935_add_4_19_lut (.I0(n45_adj_4762), .I1(GND_net), 
            .I2(pwm_counter[17]), .I3(n46537), .O(n51629)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1935_add_4_19_lut.LUT_INIT = 16'h8228;
    SB_CARRY pwm_counter_1935_add_4_19 (.CI(n46537), .I0(GND_net), .I1(pwm_counter[17]), 
            .CO(n46538));
    SB_LUT4 pwm_counter_1935_add_4_18_lut (.I0(n45_adj_4762), .I1(GND_net), 
            .I2(pwm_counter[16]), .I3(n46536), .O(n51669)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1935_add_4_18_lut.LUT_INIT = 16'h8228;
    SB_CARRY pwm_counter_1935_add_4_18 (.CI(n46536), .I0(GND_net), .I1(pwm_counter[16]), 
            .CO(n46537));
    SB_LUT4 pwm_counter_1935_add_4_17_lut (.I0(n45_adj_4762), .I1(GND_net), 
            .I2(pwm_counter[15]), .I3(n46535), .O(n51709)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1935_add_4_17_lut.LUT_INIT = 16'h8228;
    SB_CARRY pwm_counter_1935_add_4_17 (.CI(n46535), .I0(GND_net), .I1(pwm_counter[15]), 
            .CO(n46536));
    SB_LUT4 pwm_counter_1935_add_4_16_lut (.I0(n45_adj_4762), .I1(GND_net), 
            .I2(pwm_counter[14]), .I3(n46534), .O(n51751)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1935_add_4_16_lut.LUT_INIT = 16'h8228;
    SB_CARRY pwm_counter_1935_add_4_16 (.CI(n46534), .I0(GND_net), .I1(pwm_counter[14]), 
            .CO(n46535));
    SB_LUT4 pwm_counter_1935_add_4_15_lut (.I0(n45_adj_4762), .I1(GND_net), 
            .I2(pwm_counter[13]), .I3(n46533), .O(n51783)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1935_add_4_15_lut.LUT_INIT = 16'h8228;
    SB_CARRY pwm_counter_1935_add_4_15 (.CI(n46533), .I0(GND_net), .I1(pwm_counter[13]), 
            .CO(n46534));
    SB_LUT4 pwm_counter_1935_add_4_14_lut (.I0(n45_adj_4762), .I1(GND_net), 
            .I2(pwm_counter[12]), .I3(n46532), .O(n51819)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1935_add_4_14_lut.LUT_INIT = 16'h8228;
    SB_CARRY pwm_counter_1935_add_4_14 (.CI(n46532), .I0(GND_net), .I1(pwm_counter[12]), 
            .CO(n46533));
    SB_LUT4 pwm_counter_1935_add_4_13_lut (.I0(n45_adj_4762), .I1(GND_net), 
            .I2(pwm_counter[11]), .I3(n46531), .O(n51857)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1935_add_4_13_lut.LUT_INIT = 16'h8228;
    SB_CARRY pwm_counter_1935_add_4_13 (.CI(n46531), .I0(GND_net), .I1(pwm_counter[11]), 
            .CO(n46532));
    SB_LUT4 pwm_counter_1935_add_4_12_lut (.I0(n45_adj_4762), .I1(GND_net), 
            .I2(pwm_counter[10]), .I3(n46530), .O(n51889)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1935_add_4_12_lut.LUT_INIT = 16'h8228;
    SB_CARRY pwm_counter_1935_add_4_12 (.CI(n46530), .I0(GND_net), .I1(pwm_counter[10]), 
            .CO(n46531));
    SB_LUT4 pwm_counter_1935_add_4_11_lut (.I0(n45_adj_4762), .I1(GND_net), 
            .I2(pwm_counter[9]), .I3(n46529), .O(n51927)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1935_add_4_11_lut.LUT_INIT = 16'h8228;
    SB_CARRY pwm_counter_1935_add_4_11 (.CI(n46529), .I0(GND_net), .I1(pwm_counter[9]), 
            .CO(n46530));
    SB_LUT4 pwm_counter_1935_add_4_10_lut (.I0(n45_adj_4762), .I1(GND_net), 
            .I2(pwm_counter[8]), .I3(n46528), .O(n51971)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1935_add_4_10_lut.LUT_INIT = 16'h8228;
    SB_CARRY pwm_counter_1935_add_4_10 (.CI(n46528), .I0(GND_net), .I1(pwm_counter[8]), 
            .CO(n46529));
    SB_LUT4 pwm_counter_1935_add_4_9_lut (.I0(n45_adj_4762), .I1(GND_net), 
            .I2(pwm_counter[7]), .I3(n46527), .O(n52013)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1935_add_4_9_lut.LUT_INIT = 16'h8228;
    SB_CARRY pwm_counter_1935_add_4_9 (.CI(n46527), .I0(GND_net), .I1(pwm_counter[7]), 
            .CO(n46528));
    SB_LUT4 pwm_counter_1935_add_4_8_lut (.I0(n45_adj_4762), .I1(GND_net), 
            .I2(pwm_counter[6]), .I3(n46526), .O(n52059)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1935_add_4_8_lut.LUT_INIT = 16'h8228;
    SB_CARRY pwm_counter_1935_add_4_8 (.CI(n46526), .I0(GND_net), .I1(pwm_counter[6]), 
            .CO(n46527));
    SB_LUT4 pwm_counter_1935_add_4_7_lut (.I0(n45_adj_4762), .I1(GND_net), 
            .I2(pwm_counter[5]), .I3(n46525), .O(n52119)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1935_add_4_7_lut.LUT_INIT = 16'h8228;
    SB_CARRY pwm_counter_1935_add_4_7 (.CI(n46525), .I0(GND_net), .I1(pwm_counter[5]), 
            .CO(n46526));
    SB_LUT4 pwm_counter_1935_add_4_6_lut (.I0(n45_adj_4762), .I1(GND_net), 
            .I2(pwm_counter[4]), .I3(n46524), .O(n52279)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1935_add_4_6_lut.LUT_INIT = 16'h8228;
    SB_CARRY pwm_counter_1935_add_4_6 (.CI(n46524), .I0(GND_net), .I1(pwm_counter[4]), 
            .CO(n46525));
    SB_LUT4 pwm_counter_1935_add_4_5_lut (.I0(n45_adj_4762), .I1(GND_net), 
            .I2(pwm_counter[3]), .I3(n46523), .O(n52395)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1935_add_4_5_lut.LUT_INIT = 16'h8228;
    SB_CARRY pwm_counter_1935_add_4_5 (.CI(n46523), .I0(GND_net), .I1(pwm_counter[3]), 
            .CO(n46524));
    SB_LUT4 pwm_counter_1935_add_4_4_lut (.I0(n45_adj_4762), .I1(GND_net), 
            .I2(pwm_counter[2]), .I3(n46522), .O(n52393)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1935_add_4_4_lut.LUT_INIT = 16'h8228;
    SB_CARRY pwm_counter_1935_add_4_4 (.CI(n46522), .I0(GND_net), .I1(pwm_counter[2]), 
            .CO(n46523));
    SB_LUT4 pwm_counter_1935_add_4_3_lut (.I0(n45_adj_4762), .I1(GND_net), 
            .I2(pwm_counter[1]), .I3(n46521), .O(n52391)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1935_add_4_3_lut.LUT_INIT = 16'h8228;
    SB_CARRY pwm_counter_1935_add_4_3 (.CI(n46521), .I0(GND_net), .I1(pwm_counter[1]), 
            .CO(n46522));
    SB_LUT4 pwm_counter_1935_add_4_2_lut (.I0(n45_adj_4762), .I1(GND_net), 
            .I2(pwm_counter[0]), .I3(VCC_net), .O(n52381)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1935_add_4_2_lut.LUT_INIT = 16'h8228;
    SB_CARRY pwm_counter_1935_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(pwm_counter[0]), 
            .CO(n46521));
    SB_LUT4 i46077_3_lut_4_lut (.I0(pwm_counter[3]), .I1(pwm_setpoint[3]), 
            .I2(pwm_setpoint[2]), .I3(pwm_counter[2]), .O(n60789));   // verilog/pwm.v(21[8:24])
    defparam i46077_3_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 duty_23__I_0_i6_3_lut_3_lut (.I0(pwm_counter[3]), .I1(pwm_setpoint[3]), 
            .I2(pwm_setpoint[2]), .I3(GND_net), .O(n6));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i6_3_lut_3_lut.LUT_INIT = 16'hd4d4;
    SB_LUT4 i8_2_lut (.I0(\PWMLimit[7] ), .I1(\setpoint[7] ), .I2(GND_net), 
            .I3(GND_net), .O(n15));   // verilog/TinyFPGA_B.v(230[22:30])
    defparam i8_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut (.I0(pwm_counter[16]), .I1(pwm_counter[13]), .I2(pwm_counter[19]), 
            .I3(pwm_counter[18]), .O(n55155));
    defparam i3_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i6_4_lut (.I0(pwm_counter[22]), .I1(pwm_counter[11]), .I2(n55155), 
            .I3(pwm_counter[17]), .O(n16_adj_4764));
    defparam i6_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i2_3_lut (.I0(pwm_counter[6]), .I1(pwm_counter[8]), .I2(pwm_counter[7]), 
            .I3(GND_net), .O(n55170));
    defparam i2_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i4_2_lut (.I0(pwm_counter[15]), .I1(pwm_counter[14]), .I2(GND_net), 
            .I3(GND_net), .O(n14));
    defparam i4_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i8_3_lut (.I0(pwm_counter[20]), .I1(n16_adj_4764), .I2(pwm_counter[12]), 
            .I3(GND_net), .O(n18));
    defparam i8_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i3_4_lut_adj_947 (.I0(n55170), .I1(pwm_counter[21]), .I2(pwm_counter[10]), 
            .I3(pwm_counter[9]), .O(n13_adj_4765));
    defparam i3_4_lut_adj_947.LUT_INIT = 16'heccc;
    SB_LUT4 i1_4_lut (.I0(pwm_counter[23]), .I1(n13_adj_4765), .I2(n18), 
            .I3(n14), .O(n45_adj_4762));   // verilog/pwm.v(17[20:33])
    defparam i1_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 duty_23__I_0_i8_3_lut_3_lut (.I0(pwm_setpoint[4]), .I1(pwm_setpoint[8]), 
            .I2(pwm_counter[8]), .I3(GND_net), .O(n8));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i8_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i46133_2_lut_4_lut (.I0(pwm_counter[21]), .I1(pwm_setpoint[21]), 
            .I2(pwm_counter[9]), .I3(pwm_setpoint[9]), .O(n60845));
    defparam i46133_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 duty_23__I_0_i16_3_lut_3_lut (.I0(pwm_setpoint[9]), .I1(pwm_setpoint[21]), 
            .I2(pwm_counter[21]), .I3(GND_net), .O(n16));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i16_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 duty_23__I_0_i10_3_lut_3_lut (.I0(pwm_setpoint[5]), .I1(pwm_setpoint[6]), 
            .I2(pwm_counter[6]), .I3(GND_net), .O(n10));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i10_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i45235_2_lut_4_lut (.I0(pwm_counter[16]), .I1(pwm_setpoint[16]), 
            .I2(pwm_counter[7]), .I3(pwm_setpoint[7]), .O(n59947));
    defparam i45235_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 duty_23__I_0_i12_3_lut_3_lut (.I0(pwm_setpoint[7]), .I1(pwm_setpoint[16]), 
            .I2(pwm_counter[16]), .I3(GND_net), .O(n12));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i12_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    
endmodule
//
// Verilog Description of module motorControl
//

module motorControl (GND_net, \Kp[12] , \Ki[3] , n348, n32007, \Kp[13] , 
            VCC_net, \PID_CONTROLLER.integral , n292, \Ki[4] , \Kp[6] , 
            IntegralLimit, \Ki[7] , n344, \Ki[0] , n341, \Kp[1] , 
            \Kp[0] , \Ki[5] , \Ki[6] , \Kp[7] , \Ki[8] , \Kp[8] , 
            \Ki[9] , \Kp[9] , \Ki[10] , \Kp[10] , control_update, 
            duty, clk16MHz, reset, n240, \Kp[2] , setpoint, \Kp[3] , 
            \Ki[11] , \Ki[12] , n284, n258, \Kp[4] , \Ki[1] , n349, 
            n53, \Ki[2] , \Kp[11] , \deadband[0] , n339, n338, n336, 
            n337, n340, \Kp[14] , \Kp[5] , n490, n417, n344_adj_1, 
            n271, n198, n125, n35, n26870, n26869, n26868, n26867, 
            n26866, n26865, n26864, n26863, n26862, n26861, n26860, 
            n26859, n26858, n26857, n26856, n26855, n26854, n26853, 
            n26852, n26851, n26850, n26849, n26780, \Kp[15] , n343, 
            \deadband[1] , n26085, \motor_state[23] , \motor_state[22] , 
            \motor_state[21] , \motor_state[20] , \motor_state[19] , \motor_state[18] , 
            \motor_state[17] , \motor_state[16] , \motor_state[15] , \motor_state[14] , 
            \motor_state[13] , \motor_state[12] , n35211, \motor_state[10] , 
            \motor_state[9] , \motor_state[8] , \motor_state[7] , n33792, 
            \motor_state[5] , \motor_state[4] , \motor_state[3] , \motor_state[2] , 
            n1, \motor_state[0] , n350, \Ki[13] , \Ki[14] , n351, 
            \deadband[5] , n345, \Ki[15] , \deadband[6] , \deadband[7] , 
            \deadband[8] , \deadband[9] , \deadband[10] , \deadband[11] , 
            \deadband[12] , \deadband[13] , \deadband[14] , \deadband[15] , 
            \deadband[16] , n352, \deadband[17] , \deadband[18] , PWMLimit, 
            \deadband[19] , \deadband[20] , \deadband[21] , \deadband[22] , 
            \deadband[23] , n359, n353, n346, n35713, n354, \control_mode[0] , 
            \control_mode[5] , \control_mode[4] , n1_adj_2, n355, \control_mode[6] , 
            \control_mode[7] , \control_mode[1] , n19, n15, n356, 
            \deadband[3] , \deadband[4] , n357, n358, n347) /* synthesis syn_module_defined=1 */ ;
    input GND_net;
    input \Kp[12] ;
    input \Ki[3] ;
    output n348;
    input n32007;
    input \Kp[13] ;
    input VCC_net;
    output [23:0]\PID_CONTROLLER.integral ;
    output n292;
    input \Ki[4] ;
    input \Kp[6] ;
    input [23:0]IntegralLimit;
    input \Ki[7] ;
    output n344;
    input \Ki[0] ;
    output n341;
    input \Kp[1] ;
    input \Kp[0] ;
    input \Ki[5] ;
    input \Ki[6] ;
    input \Kp[7] ;
    input \Ki[8] ;
    input \Kp[8] ;
    input \Ki[9] ;
    input \Kp[9] ;
    input \Ki[10] ;
    input \Kp[10] ;
    output control_update;
    output [23:0]duty;
    input clk16MHz;
    input reset;
    output n240;
    input \Kp[2] ;
    input [23:0]setpoint;
    input \Kp[3] ;
    input \Ki[11] ;
    input \Ki[12] ;
    output n284;
    output n258;
    input \Kp[4] ;
    input \Ki[1] ;
    output n349;
    input n53;
    input \Ki[2] ;
    input \Kp[11] ;
    input \deadband[0] ;
    output n339;
    output n338;
    output n336;
    output n337;
    output n340;
    input \Kp[14] ;
    input \Kp[5] ;
    input n490;
    input n417;
    input n344_adj_1;
    input n271;
    input n198;
    input n125;
    input n35;
    input n26870;
    input n26869;
    input n26868;
    input n26867;
    input n26866;
    input n26865;
    input n26864;
    input n26863;
    input n26862;
    input n26861;
    input n26860;
    input n26859;
    input n26858;
    input n26857;
    input n26856;
    input n26855;
    input n26854;
    input n26853;
    input n26852;
    input n26851;
    input n26850;
    input n26849;
    input n26780;
    input \Kp[15] ;
    output n343;
    input \deadband[1] ;
    input n26085;
    input \motor_state[23] ;
    input \motor_state[22] ;
    input \motor_state[21] ;
    input \motor_state[20] ;
    input \motor_state[19] ;
    input \motor_state[18] ;
    input \motor_state[17] ;
    input \motor_state[16] ;
    input \motor_state[15] ;
    input \motor_state[14] ;
    input \motor_state[13] ;
    input \motor_state[12] ;
    input n35211;
    input \motor_state[10] ;
    input \motor_state[9] ;
    input \motor_state[8] ;
    input \motor_state[7] ;
    input n33792;
    input \motor_state[5] ;
    input \motor_state[4] ;
    input \motor_state[3] ;
    input \motor_state[2] ;
    input n1;
    input \motor_state[0] ;
    output n350;
    input \Ki[13] ;
    input \Ki[14] ;
    output n351;
    input \deadband[5] ;
    output n345;
    input \Ki[15] ;
    input \deadband[6] ;
    input \deadband[7] ;
    input \deadband[8] ;
    input \deadband[9] ;
    input \deadband[10] ;
    input \deadband[11] ;
    input \deadband[12] ;
    input \deadband[13] ;
    input \deadband[14] ;
    input \deadband[15] ;
    input \deadband[16] ;
    output n352;
    input \deadband[17] ;
    input \deadband[18] ;
    input [23:0]PWMLimit;
    input \deadband[19] ;
    input \deadband[20] ;
    input \deadband[21] ;
    input \deadband[22] ;
    input \deadband[23] ;
    output n359;
    output n353;
    output n346;
    output n35713;
    output n354;
    input \control_mode[0] ;
    input \control_mode[5] ;
    input \control_mode[4] ;
    input n1_adj_2;
    output n355;
    input \control_mode[6] ;
    input \control_mode[7] ;
    input \control_mode[1] ;
    input n19;
    input n15;
    output n356;
    input \deadband[3] ;
    input \deadband[4] ;
    output n357;
    output n358;
    output n347;
    
    wire clk16MHz /* synthesis SET_AS_NETWORK=clk16MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(31[6:14])
    
    wire n46176;
    wire [23:0]n28;
    
    wire n46177;
    wire [23:0]n207;
    
    wire n907;
    wire [7:0]n17669;
    wire [6:0]n17795;
    
    wire n411, n46732;
    wire [7:0]n17609;
    wire [6:0]n17750;
    
    wire n630, n47053, n557, n47052, n46733, n484, n47051, n338_c, 
        n46731;
    wire [23:0]n34;
    
    wire n46175, n253, n46174, n411_adj_4203, n47050, n338_adj_4204, 
        n47049, n265, n46730, n265_adj_4205, n47048, n192, n46729, 
        n50, n119, n980, n192_adj_4206, n47047;
    wire [12:0]n16284;
    wire [11:0]n16645;
    
    wire n980_adj_4207, n46728, n50_adj_4208, n119_adj_4209;
    wire [17:0]n13879;
    wire [16:0]n14525;
    
    wire n47046, n907_adj_4210, n46727, n47045, n834, n46726, n47044, 
        n761, n46725, n688, n46724, n1111, n47043, n46173, n615, 
        n46723, n1038, n47042, n542, n46722, n45, n31995;
    wire [23:0]n285;
    wire [23:0]n36;
    
    wire n46172, n965, n47041, n469, n46721, n892, n47040, n46171, 
        n396, n46720, n323, n46719, n819, n47039, n250, n46718, 
        n46170, n177, n46717;
    wire [23:0]n233;
    
    wire n46059, n46169, n35_c, n104, n46060;
    wire [10:0]n16954;
    
    wire n910, n46716, n837, n46715, n746, n47038, n764, n46714, 
        n46168, n673, n47037, n691, n46713, n46167, n600, n47036, 
        n46058, n618, n46712, n527, n47035, n545, n46711, n46166, 
        n472, n46710, n399, n46709, n46165, n454, n47034, n326, 
        n46708, n46707, n180, n46706, n46057, n381, n47033, n38, 
        n107, n46164;
    wire [5:0]n17891;
    
    wire n560, n46705, n308, n47032, n487, n46704, n414, n46703, 
        n341_c, n46702, n268, n46701, n235, n47031, n195, n46700, 
        n46163, n53_c, n122, n162, n47030;
    wire [9:0]n17215;
    
    wire n840, n46699, n20, n89, n767, n46698, n694, n46697;
    wire [15:0]n15101;
    
    wire n47029, n47028, n621, n46696, n1114, n47027, n46056, 
        n1041, n47026, n548, n46695, n968, n47025, n475, n46694, 
        n46162, n46055, n895, n47024, n402, n46693, n822, n47023, 
        n329, n46692, n46161, n749, n47022, n256, n46691, n676, 
        n47021, n183, n46690, n41, n110, n46160, n46054, n603, 
        n47020, n530, n47019, n46159, n457, n47018, n46158, n384, 
        n47017, n311, n47016, n46157, n46053, n238, n47015, n46052, 
        n46156, n56, n101, n32, n46155, n165, n47014, n23, n92;
    wire [5:0]n17859;
    
    wire n560_adj_4214, n47013, n45_adj_4216, n39, n46154, n41_adj_4219, 
        n43, n37, n487_adj_4220, n47012, n63680, n46153, n35_adj_4222, 
        n174, n46051, counter_31__N_3487, n414_adj_4223, n47011, n9440, 
        n59906, n4357, n63485, n247_adj_4224, n46152, n341_adj_4226, 
        n47010, n46151;
    wire [23:0]n310;
    wire [23:0]n535;
    wire [23:0]n455;
    
    wire n63488, n27, n268_adj_4229, n47009, n46150, n320, n59905, 
        n63479, n31, n195_adj_4233, n47008, n63482, n33, n46050, 
        n29, n21_adj_4235, n19_adj_4236, n17_adj_4237, n9_adj_4238, 
        n60366, n122_adj_4240;
    wire [14:0]n15611;
    
    wire n47007, n1117, n47006, n1044, n47005, n15_adj_4241, n13_adj_4242, 
        n11_adj_4243, n60326, n971, n47004, n898, n47003, n825, 
        n47002, n59904, n63467, n63470, n752, n47001, n12_adj_4244, 
        n10_adj_4245, n30, n679, n47000, n60399, n61363, n61351, 
        n25_adj_4246, n23_adj_4247, n62631, n606, n46999, n61917, 
        n62769, n16_adj_4248, n533, n46998, n460_adj_4249, n46997, 
        n387, n46996, n6_adj_4250, n61956, n61957, n8_adj_4251, 
        n24_adj_4252, n314, n46995, n60182, n241_adj_4253, n46994, 
        n168, n46993, n26, n95;
    wire [13:0]n16059;
    
    wire n1120, n46992, n60177, n61877, n1047, n46991, n974, n46990, 
        n901, n46989, n828, n46988, n755, n46987, n61119, n4_adj_4254, 
        n61954, n682, n46986, n61955, n609, n46985, n536, n46984, 
        n60235, n463, n46983, n390, n46982, n317, n46981, n244_adj_4255, 
        n46980, n60223, n62402, n171, n46979, n29_adj_4256, n98, 
        n61121, n62802, n62803;
    wire [3:0]n17997;
    
    wire n6_adj_4257;
    wire [4:0]n17940;
    
    wire n62801, n60193, n62553, n61127, n62753, n45_adj_4258, n41_adj_4259;
    wire [1:0]n18055;
    
    wire n45772;
    wire [2:0]n18034;
    
    wire n43_adj_4260, n39_adj_4261, n37_adj_4264, n31_adj_4266, n33_adj_4267, 
        n29_adj_4268, n56496, n56500, n56498, n59903, n63461, n27_adj_4269, 
        n45721, n56506, n4_adj_4270, n21_adj_4271, n19_adj_4272, n17_adj_4273, 
        n9_adj_4274, n60087, n8_adj_4275, n6_adj_4276, n55441, n15_adj_4277, 
        n13_adj_4278, n11_adj_4279, n60051, n12_adj_4280, n393, n46978, 
        n10_adj_4281, n46977, n46976, n46975, n466, n46974, n59930, 
        n63677;
    wire [12:0]n16449;
    
    wire n1050, n46973, n977, n46972, n904, n46971, n831, n46970, 
        n758, n46969, n63464, n59902, n63455, n63458, n685, n46968, 
        n612, n46967;
    wire [13:0]n61;
    wire [31:0]counter;   // verilog/motorControl.v(22[11:18])
    
    wire n46625, n59901, n63449, n46624, n46623, n539_adj_4285, 
        n46966, n30_adj_4287, n46622, n46965, n46964, n46621, n63452, 
        n46963, n46620, n46962, n46619, n46618, n46961, n46617, 
        n46616, n60168, n61076, n59900, n63443, n61056, n63446, 
        n25_adj_4289, n23_adj_4290, n62529, n59899, n63437;
    wire [11:0]n16785;
    
    wire n46960, n46615, n63440, n61833, n62737, n46959, n834_adj_4292, 
        n46958, n761_adj_4293, n46957, n46614, n688_adj_4294, n46956, 
        n46613, n59898, n63431, n615_adj_4295, n46955, n63434, n542_adj_4296, 
        n46954, n16_adj_4297, n59897, n63425, n469_adj_4298, n46953, 
        n63428, n396_adj_4300, n46952, n6_adj_4301, n62449, n62450, 
        n323_adj_4302, n46951, n59896, n63419, n63422, n8_adj_4304, 
        n250_adj_4305, n46950, n24_adj_4306, n59983, n177_adj_4307, 
        n46949, n59981, n61879, n35_adj_4308, n104_adj_4309, n62233, 
        n59886, n63407, n63410, n59885, n63401;
    wire [10:0]n17071;
    
    wire n910_adj_4310, n46948, n837_adj_4311, n46947, n764_adj_4312, 
        n46946, n4_adj_4313, n691_adj_4314, n46945, n62447, n63404, 
        n62448, n618_adj_4315, n46944, n59884, n63395, n545_adj_4316, 
        n46943, n472_adj_4317, n46942, n63398, n399_adj_4319, n46941, 
        n326_adj_4320, n46940, n253_adj_4321, n46939, n180_adj_4322, 
        n46938, n38_adj_4323, n107_adj_4324;
    wire [0:0]n9524;
    wire [21:0]n10031;
    
    wire n46937;
    wire [47:0]n42;
    
    wire n46936, n60019, n46935, n46934, n46933, n60010, n62775, 
        n46932, n46931, n46930, n1096, n46929, n1023, n46928, 
        n62235, n950, n46927, n877, n46926, n804, n46925, n731, 
        n46924, n658, n46923, n585, n46922, n512, n46921, n59883, 
        n63389, n439_adj_4325, n46920, n366, n46919, n293_adj_4326, 
        n46918, n220_adj_4327, n46917, n147, n46916, n5_adj_4328, 
        n74_adj_4329;
    wire [20:0]n11044;
    
    wire n46915, n46914, n46913, n46912, n46911, n46910, n46909, 
        n1099, n46908, n1026, n46907, n953, n46906, n880, n46905, 
        n807, n46904, n734, n46903, n661, n46902, n588, n46901, 
        n515, n46900, n442_adj_4330, n46899, n369, n46898, n62963, 
        n296_adj_4331, n46897, n62964, n223_adj_4332, n46896, n150, 
        n46895, n8_adj_4333, n77, n62909;
    wire [19:0]n11965;
    
    wire n46894, n46893, n46892, n46891, n59987, n46890, n62238, 
        n46889, n40, n1102, n46888, n1029, n46887, n62557, n956, 
        n46886, n883, n46885, n810, n46884, n737, n46883, n664, 
        n46882, n591, n46881, n518, n46880, n445_adj_4334, n46879, 
        n372, n46878, n63392, n299_adj_4335, n46877, n226_adj_4336, 
        n46876, n153, n46875, n11_adj_4337, n80;
    wire [18:0]n12802;
    
    wire n46874, n46873, n46872, n46871, n46870, n1105, n46869, 
        n1032, n46868, n959, n46867, n886, n46866, n813, n46865, 
        n63554, n63512, n63506, n63380, n63368, n63356, n63344, 
        n63278, n740, n46864, n667, n46863, n594, n46862, n521, 
        n46861, n448_adj_4338, n46860, n375, n46859, n302_adj_4339, 
        n46858, n229, n46857, n156, n46856, n14_adj_4340, n83;
    wire [9:0]n17311;
    
    wire n840_adj_4341, n46855, n767_adj_4342, n46854, n694_adj_4343, 
        n46853, n621_adj_4344, n46852, n548_adj_4345, n46851, n475_adj_4346, 
        n46850, n402_adj_4347, n46849, n329_adj_4348, n46848;
    wire [0:0]n10055;
    
    wire n46095, n256_adj_4349, n46847;
    wire [43:0]n360;
    
    wire n46094, n46093, n183_adj_4351, n46846, n41_adj_4352, n110_adj_4353;
    wire [17:0]n13559;
    
    wire n46845, n46844, n46092, n46091, n46843, n46842, n1108, 
        n46841, n1035, n46840, n962, n46839, n889, n46838, n816, 
        n46837, n743, n46836, n670, n46835, n597, n46834, n524, 
        n46833, n451_adj_4355, n46832, n378, n46831, n305_adj_4356, 
        n46830, n232, n46829, n159, n46828, n17_adj_4357, n86;
    wire [16:0]n14240;
    
    wire n46827, n46826, n46825, n1111_adj_4358, n46824, n1038_adj_4359, 
        n46823, n965_adj_4360, n46822, n892_adj_4361, n46821, n819_adj_4362, 
        n46820, n746_adj_4363, n46819, n673_adj_4364, n46818, n600_adj_4365, 
        n46817, n527_adj_4366, n46816, n454_adj_4367, n46815, n381_adj_4368, 
        n46814, n308_adj_4369, n46813, n235_adj_4370, n46812, n162_adj_4371, 
        n46811, n20_adj_4372, n89_adj_4373;
    wire [8:0]n17509;
    
    wire n770, n46810, n697, n46809, n46090, n46089, n46241, n46240, 
        n46088, n624, n46808, n551_adj_4375, n46807, n46239;
    wire [8:0]n17432;
    
    wire n770_adj_4376, n47175, n697_adj_4377, n47174, n478, n46806, 
        n624_adj_4378, n47173, n46238, n46237, n46087, n46236, n551_adj_4379, 
        n47172, n478_adj_4380, n47171, n405, n46805, n405_adj_4381, 
        n47170, n332, n46804, n332_adj_4382, n47169, n259, n46803, 
        n259_adj_4383, n47168, n186, n47167, n46235, n46234, n46233, 
        n46232, n186_adj_4384, n46802, n44, n113, n44_adj_4385, 
        n113_adj_4386;
    wire [21:0]n10514;
    
    wire n47166, n47165;
    wire [15:0]n14849;
    
    wire n46801, n46086, n47164, n46800, n46231, n46230, n46085, 
        n1114_adj_4388, n46799, n47163, n1041_adj_4389, n46798, n47162, 
        n968_adj_4390, n46797, n47161, n46229, n47160, n46228, n46227, 
        n46226, n47159, n1096_adj_4391, n47158, n895_adj_4392, n46796, 
        n1023_adj_4393, n47157, n822_adj_4394, n46795, n950_adj_4395, 
        n47156, n877_adj_4396, n47155, n749_adj_4397, n46794, n46225, 
        n804_adj_4399, n47154, n46224, n731_adj_4400, n47153, n46223, 
        n46222, n46221, n46220, n658_adj_4401, n47152, n585_adj_4403, 
        n47151, n676_adj_4404, n46793, n512_adj_4405, n47150, n46084, 
        n603_adj_4406, n46792, n46219;
    wire [23:0]n46;
    
    wire n46218, n439_adj_4409, n47149, n46217, n366_adj_4412, n47148, 
        n293_adj_4413, n47147, n530_adj_4414, n46791, n220_adj_4415, 
        n47146, n46216, n147_adj_4418, n47145, n457_adj_4419, n46790, 
        n5_adj_4420, n74_adj_4421, n384_adj_4422, n46789, n46215, 
        n46214, n46213, n46212, n46083, n46211, n46082;
    wire [20:0]n11481;
    
    wire n47144, n46081, n46210, n47143, n311_adj_4429, n46788, 
        n47142, n238_adj_4430, n46787, n47141, n165_adj_4431, n46786, 
        n47140, n47139, n23_adj_4432, n92_adj_4433, n47138;
    wire [14:0]n15390;
    
    wire n46785, n1099_adj_4434, n47137, n46209, n46208, n46207, 
        n46206, n46080, n46079, n1026_adj_4439, n47136, n1117_adj_4440, 
        n46784, n953_adj_4441, n47135, n1044_adj_4442, n46783, n880_adj_4443, 
        n47134, n46205, n971_adj_4445, n46782, n807_adj_4446, n47133, 
        n898_adj_4447, n46781, n734_adj_4448, n47132, n46204, n661_adj_4450, 
        n47131, n46203, n46202, n46078, n588_adj_4453, n47130, n515_adj_4454, 
        n47129, n442_adj_4455, n47128, n825_adj_4456, n46780, n369_adj_4457, 
        n47127, n752_adj_4458, n46779, n296_adj_4459, n47126, n679_adj_4460, 
        n46778, n223_adj_4461, n47125, n46077, n46201, n46200, n46199, 
        n46076, n46198, n150_adj_4467, n47124, n46075, n46074, n46073, 
        n606_adj_4469, n46777, n533_adj_4470, n46776, n8_adj_4471, 
        n77_adj_4472, n460_adj_4473, n46775, n54612, n490_adj_4474, 
        n47123, n46197;
    wire [4:0]n17961;
    
    wire n417_adj_4477, n47122, n344_adj_4478, n47121, n271_adj_4479, 
        n47120, n46196, n198_adj_4481, n47119, n46072, n46071, n47, 
        n46195, n56_adj_4484, n125_adj_4485, n46194;
    wire [19:0]n12361;
    
    wire n47118, n47117, n46070, n46193, n47116, n46192, n47115, 
        n46069, n46191, n387_adj_4491, n46774, n47114, n47113, n46068, 
        n1102_adj_4492, n47112, n314_adj_4493, n46773, n46190, n1029_adj_4496, 
        n47111, n46067, n241_adj_4497, n46772, n46189, n956_adj_4499, 
        n47110, n168_adj_4500, n46771, n883_adj_4501, n47109, n26_adj_4502, 
        n95_adj_4503, n810_adj_4504, n47108, n700, n46770, n46188, 
        n46066, n737_adj_4506, n47107, n46187, n46065, n46186, n664_adj_4510, 
        n47106, n591_adj_4511, n47105, n627, n46769, n518_adj_4512, 
        n47104, n46185, n46064, n445_adj_4514, n47103, n554_adj_4515, 
        n46768, n372_adj_4516, n47102, n481, n46767, n46184, n46063, 
        n46183, n299_adj_4519, n47101, n226_adj_4520, n47100, n153_adj_4521, 
        n47099, n408, n46766, n11_adj_4522, n80_adj_4523, n335, 
        n46765, n46182, n46181, n46062, n262, n46764, n700_adj_4526, 
        n47098, n627_adj_4527, n47097, n189, n46763, n46180, n46061, 
        n554_adj_4529, n47096, n46179, n46178, n481_adj_4532, n47095, 
        n47_adj_4533, n116, n408_adj_4534, n47094, n335_adj_4535, 
        n47093;
    wire [13:0]n15867;
    
    wire n1120_adj_4536, n46762, n262_adj_4537, n47092, n1047_adj_4538, 
        n46761, n189_adj_4539, n47091, n974_adj_4540, n46760, n47_adj_4541, 
        n116_adj_4542, n901_adj_4543, n46759;
    wire [18:0]n13159;
    
    wire n47090, n47089, n828_adj_4544, n46758, n47088, n755_adj_4545, 
        n46757, n682_adj_4546, n46756, n47087, n609_adj_4548, n46755, 
        n47086, n536_adj_4549, n46754, n1105_adj_4550, n47085, n463_adj_4551, 
        n46753, n390_adj_4552, n46752, n1032_adj_4553, n47084, n959_adj_4554, 
        n47083, n886_adj_4555, n47082, n317_adj_4556, n46751, n813_adj_4557, 
        n47081, n244_adj_4558, n46750, n740_adj_4559, n47080, n171_adj_4560, 
        n46749, n667_adj_4561, n47079, n594_adj_4562, n47078, n29_adj_4563, 
        n98_adj_4564, n1050_adj_4565, n46748, n977_adj_4566, n46747, 
        n521_adj_4567, n47077, n904_adj_4568, n46746, n448_adj_4569, 
        n47076, n375_adj_4570, n47075, n302_adj_4571, n47074, n831_adj_4572, 
        n46745, n229_adj_4573, n47073, n758_adj_4574, n46744, n685_adj_4575, 
        n46743, n156_adj_4576, n47072, n612_adj_4577, n46742, n14_adj_4578, 
        n83_adj_4579, n47071, n539_adj_4580, n46741, n47070, n466_adj_4581, 
        n46740, n47069, n47068, n1108_adj_4582, n47067, n1035_adj_4583, 
        n47066, n962_adj_4584, n47065, n393_adj_4585, n46739, n889_adj_4586, 
        n47064, n320_adj_4587, n46738, n247_adj_4588, n46737, n816_adj_4589, 
        n47063, n174_adj_4590, n46736, n32_adj_4591, n101_adj_4592, 
        n743_adj_4593, n47062, n630_adj_4594, n46735, n670_adj_4595, 
        n47061, n557_adj_4596, n46734, n597_adj_4597, n47060, n524_adj_4598, 
        n47059, n451_adj_4599, n47058, n378_adj_4600, n47057, n305_adj_4601, 
        n47056, n232_adj_4602, n47055, n59882, n63377, n159_adj_4603, 
        n47054, n17_adj_4604, n86_adj_4605, n484_adj_4606, n41_adj_4607, 
        n39_adj_4608, n45_adj_4609, n43_adj_4610, n21_adj_4611, n23_adj_4612, 
        n25_adj_4613, n17_adj_4614, n19_adj_4615, n37_adj_4616, n35_adj_4617, 
        n27_adj_4618, n29_adj_4619, n31_adj_4620, n9_adj_4621, n11_adj_4622, 
        n13_adj_4623, n15_adj_4624, n41_adj_4625, n39_adj_4626, n45_adj_4627, 
        n43_adj_4628, n29_adj_4629, n31_adj_4630, n23_adj_4631, n25_adj_4632, 
        n37_adj_4633, n35_adj_4634, n33_adj_4635, n11_adj_4636, n13_adj_4637, 
        n15_adj_4638, n27_adj_4639, n9_adj_4640, n17_adj_4641, n19_adj_4642, 
        n21_adj_4643, n60501, n60479, n12_adj_4644, n10_adj_4645, 
        n30_adj_4646, n60553, n61495, n61487, n62667, n61994, n62810, 
        n16_adj_4647, n6_adj_4648, n62364, n62365, n8_adj_4649, n24_adj_4650, 
        n60405, n60401, n61875, n61109, n4_adj_4651, n62360, n62361, 
        n60445, n60441, n62747, n61111, n62965, n62966, n62907, 
        n60412, n62551, n61117, n62751, n131, n41_adj_4652, n39_adj_4653, 
        n45_adj_4654, n43_adj_4655, n37_adj_4656, n45802, n56550, 
        n23_adj_4657;
    wire [3:0]n18009;
    
    wire n4_adj_4658, n25_adj_4659, n347_c, n6_adj_4660, n53040, n29_adj_4661, 
        n56546, n68_adj_4662, n31_adj_4663, n45797, n47176, n56536, 
        n64292, n56540, n8_adj_4664, n6_adj_4665, n35_adj_4666, n33_adj_4667, 
        n11_adj_4668, n13_adj_4669, n15_adj_4670, n27_adj_4671, n9_adj_4672, 
        n17_adj_4673, n19_adj_4674, n21_adj_4675, n60710, n60700, 
        n12_adj_4676, n10_adj_4677, n30_adj_4678, n60732, n61663, 
        n61657, n62709, n62090, n62826, n16_adj_4679, n6_adj_4680, 
        n62284, n62285, n8_adj_4681, n24_adj_4682, n60654, n60650, 
        n61885, n61147, n4_adj_4683, n62282, n62283, n60687, n60683, 
        n62790, n61149, n62900, n62901, n62876, n60656, n62563, 
        n61155, n62755, n41_adj_4684, n39_adj_4685, n45_adj_4686, 
        n43_adj_4687, n37_adj_4688, n29_adj_4689, n31_adj_4690, n23_adj_4691, 
        n25_adj_4692, n35_adj_4693, n33_adj_4694, n11_adj_4695, n13_adj_4696, 
        n27_adj_4697, n9_adj_4698, n17_adj_4699, n21_adj_4700, n12_adj_4702, 
        n52622, n60652, n60630, n12_adj_4705, n30_adj_4706, n60673, 
        n61613, n61605, n62695, n62060, n62820, n6_adj_4707, n62370, 
        n62371, n16_adj_4708, n24_adj_4709, n60569, n8_adj_4710, n60561, 
        n61873, n61099, n4_adj_4711, n62368, n62369, n60611, n59911, 
        n63551, n10_adj_4712, n60601, n62745, n61101, n62961, n62962, 
        n62913, n60577, n62547, n61107, n62749, n105, n33_adj_4713, 
        n43_adj_4714, n37_adj_4715, n33_adj_4716, n31_adj_4717, n4_adj_4718, 
        n35_adj_4719, n21_adj_4720, n23_adj_4721, n25_adj_4722, n27_adj_4723, 
        n29_adj_4724, n13_adj_4725, n15_adj_4726, n17_adj_4727, n9_adj_4728, 
        n11_adj_4729, n19_adj_4730, n60813, n61729, n63839, n60821, 
        n61739, n63853, n61713, n63818, n14_adj_4731, n60763, n12_adj_4732, 
        n32_adj_4733, n60830, n61745, n63860, n61743, n63849, n60815, 
        n63829, n62136, n63838, n62727, n61719, n10_adj_4734, n60967, 
        n61805, n61801, n59938, n14_adj_4735, n6_adj_4736, n62336, 
        n62337, n59932, n12_adj_4737, n32_adj_4738, n60898, n60894, 
        n62781, n61129, n8_adj_4739, n62296, n62297, n10_adj_4740, 
        n61727, n63834, n61883, n61137, n6_adj_4741, n62290, n62291, 
        n60771, n63827, n62788, n61139, n62487, n62898, n62435, 
        n62995, n62996, n62787, n62595, n62596, n8_adj_4742, n62443, 
        n62444, n59961, n60941, n61881, n62241, n62160, n62896, 
        n62439, n63007, n63008, n63002, n62599, n62562, n62600, 
        n35399, n6646, n6648, n22268, n35687, n60603, n12_adj_4743, 
        n10_adj_4744, n30_adj_4745, n60648, n61581, n61571, n62691, 
        n62046, n62818, n6_adj_4746, n62276, n62277, n16_adj_4747, 
        n8_adj_4748, n24_adj_4749, n60613, n60559, n60555, n61887, 
        n61157, n4_adj_4750, n62272, n62273, n59851, n63365, n60589, 
        n60585, n62583, n61159, n62902, n62903, n62874, n60565, 
        n62565, n61165, n62757, n4_adj_4751, n54971, n22302, n56609, 
        n23_adj_4752, n22_adj_4753, n26_adj_4754, n4_adj_4755, n45825, 
        n59843, n63353, n22266, n4_adj_4756, n45885, n59737, n63341, 
        n59908, n63509, n59723, n59907, n63503, n63275;
    
    SB_CARRY unary_minus_27_add_3_6 (.CI(n46176), .I0(GND_net), .I1(n28[4]), 
            .CO(n46177));
    SB_LUT4 mult_23_i610_2_lut (.I0(\Kp[12] ), .I1(n207[14]), .I2(GND_net), 
            .I3(GND_net), .O(n907));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i610_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_4732_6_lut (.I0(GND_net), .I1(n17795[3]), .I2(n411), .I3(n46732), 
            .O(n17669[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4732_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4726_9_lut (.I0(GND_net), .I1(n17750[6]), .I2(n630), .I3(n47053), 
            .O(n17609[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4726_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4726_8_lut (.I0(GND_net), .I1(n17750[5]), .I2(n557), .I3(n47052), 
            .O(n17609[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4726_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4726_8 (.CI(n47052), .I0(n17750[5]), .I1(n557), .CO(n47053));
    SB_CARRY add_4732_6 (.CI(n46732), .I0(n17795[3]), .I1(n411), .CO(n46733));
    SB_LUT4 add_4726_7_lut (.I0(GND_net), .I1(n17750[4]), .I2(n484), .I3(n47051), 
            .O(n17609[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4726_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4732_5_lut (.I0(GND_net), .I1(n17795[2]), .I2(n338_c), 
            .I3(n46731), .O(n17669[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4732_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_27_add_3_5_lut (.I0(GND_net), .I1(GND_net), .I2(n28[3]), 
            .I3(n46175), .O(n34[3])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_27_add_3_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_27_add_3_5 (.CI(n46175), .I0(GND_net), .I1(n28[3]), 
            .CO(n46176));
    SB_LUT4 mult_24_i171_2_lut (.I0(\Ki[3] ), .I1(n348), .I2(GND_net), 
            .I3(GND_net), .O(n253));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i171_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_27_add_3_4_lut (.I0(GND_net), .I1(GND_net), .I2(n32007), 
            .I3(n46174), .O(n34[2])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_27_add_3_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4726_7 (.CI(n47051), .I0(n17750[4]), .I1(n484), .CO(n47052));
    SB_CARRY unary_minus_27_add_3_4 (.CI(n46174), .I0(GND_net), .I1(n32007), 
            .CO(n46175));
    SB_CARRY add_4732_5 (.CI(n46731), .I0(n17795[2]), .I1(n338_c), .CO(n46732));
    SB_LUT4 add_4726_6_lut (.I0(GND_net), .I1(n17750[3]), .I2(n411_adj_4203), 
            .I3(n47050), .O(n17609[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4726_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4726_6 (.CI(n47050), .I0(n17750[3]), .I1(n411_adj_4203), 
            .CO(n47051));
    SB_LUT4 add_4726_5_lut (.I0(GND_net), .I1(n17750[2]), .I2(n338_adj_4204), 
            .I3(n47049), .O(n17609[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4726_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4732_4_lut (.I0(GND_net), .I1(n17795[1]), .I2(n265), .I3(n46730), 
            .O(n17669[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4732_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4726_5 (.CI(n47049), .I0(n17750[2]), .I1(n338_adj_4204), 
            .CO(n47050));
    SB_CARRY add_4732_4 (.CI(n46730), .I0(n17795[1]), .I1(n265), .CO(n46731));
    SB_LUT4 add_4726_4_lut (.I0(GND_net), .I1(n17750[1]), .I2(n265_adj_4205), 
            .I3(n47048), .O(n17609[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4726_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4732_3_lut (.I0(GND_net), .I1(n17795[0]), .I2(n192), .I3(n46729), 
            .O(n17669[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4732_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4726_4 (.CI(n47048), .I0(n17750[1]), .I1(n265_adj_4205), 
            .CO(n47049));
    SB_CARRY add_4732_3 (.CI(n46729), .I0(n17795[0]), .I1(n192), .CO(n46730));
    SB_LUT4 add_4732_2_lut (.I0(GND_net), .I1(n50), .I2(n119), .I3(GND_net), 
            .O(n17669[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4732_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_23_i659_2_lut (.I0(\Kp[13] ), .I1(n207[14]), .I2(GND_net), 
            .I3(GND_net), .O(n980));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i659_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_4726_3_lut (.I0(GND_net), .I1(n17750[0]), .I2(n192_adj_4206), 
            .I3(n47047), .O(n17609[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4726_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4732_2 (.CI(GND_net), .I0(n50), .I1(n119), .CO(n46729));
    SB_CARRY add_4726_3 (.CI(n47047), .I0(n17750[0]), .I1(n192_adj_4206), 
            .CO(n47048));
    SB_LUT4 add_4621_14_lut (.I0(GND_net), .I1(n16645[11]), .I2(n980_adj_4207), 
            .I3(n46728), .O(n16284[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4621_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4726_2_lut (.I0(GND_net), .I1(n50_adj_4208), .I2(n119_adj_4209), 
            .I3(GND_net), .O(n17609[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4726_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4726_2 (.CI(GND_net), .I0(n50_adj_4208), .I1(n119_adj_4209), 
            .CO(n47047));
    SB_LUT4 add_4482_19_lut (.I0(GND_net), .I1(n14525[16]), .I2(GND_net), 
            .I3(n47046), .O(n13879[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4482_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4621_13_lut (.I0(GND_net), .I1(n16645[10]), .I2(n907_adj_4210), 
            .I3(n46727), .O(n16284[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4621_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4621_13 (.CI(n46727), .I0(n16645[10]), .I1(n907_adj_4210), 
            .CO(n46728));
    SB_LUT4 add_4482_18_lut (.I0(GND_net), .I1(n14525[15]), .I2(GND_net), 
            .I3(n47045), .O(n13879[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4482_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4482_18 (.CI(n47045), .I0(n14525[15]), .I1(GND_net), 
            .CO(n47046));
    SB_LUT4 add_4621_12_lut (.I0(GND_net), .I1(n16645[9]), .I2(n834), 
            .I3(n46726), .O(n16284[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4621_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4621_12 (.CI(n46726), .I0(n16645[9]), .I1(n834), .CO(n46727));
    SB_LUT4 add_4482_17_lut (.I0(GND_net), .I1(n14525[14]), .I2(GND_net), 
            .I3(n47044), .O(n13879[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4482_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4621_11_lut (.I0(GND_net), .I1(n16645[8]), .I2(n761), 
            .I3(n46725), .O(n16284[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4621_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4482_17 (.CI(n47044), .I0(n14525[14]), .I1(GND_net), 
            .CO(n47045));
    SB_CARRY add_4621_11 (.CI(n46725), .I0(n16645[8]), .I1(n761), .CO(n46726));
    SB_LUT4 add_4621_10_lut (.I0(GND_net), .I1(n16645[7]), .I2(n688), 
            .I3(n46724), .O(n16284[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4621_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4482_16_lut (.I0(GND_net), .I1(n14525[13]), .I2(n1111), 
            .I3(n47043), .O(n13879[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4482_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_27_add_3_3_lut (.I0(GND_net), .I1(GND_net), .I2(n28[1]), 
            .I3(n46173), .O(n34[1])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_27_add_3_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_27_add_3_3 (.CI(n46173), .I0(GND_net), .I1(n28[1]), 
            .CO(n46174));
    SB_CARRY add_4621_10 (.CI(n46724), .I0(n16645[7]), .I1(n688), .CO(n46725));
    SB_LUT4 add_4621_9_lut (.I0(GND_net), .I1(n16645[6]), .I2(n615), .I3(n46723), 
            .O(n16284[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4621_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4482_16 (.CI(n47043), .I0(n14525[13]), .I1(n1111), .CO(n47044));
    SB_LUT4 add_4482_15_lut (.I0(GND_net), .I1(n14525[12]), .I2(n1038), 
            .I3(n47042), .O(n13879[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4482_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4621_9 (.CI(n46723), .I0(n16645[6]), .I1(n615), .CO(n46724));
    SB_LUT4 add_4621_8_lut (.I0(GND_net), .I1(n16645[5]), .I2(n542), .I3(n46722), 
            .O(n16284[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4621_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4621_8 (.CI(n46722), .I0(n16645[5]), .I1(n542), .CO(n46723));
    SB_LUT4 unary_minus_27_add_3_2_lut (.I0(n31995), .I1(GND_net), .I2(n28[0]), 
            .I3(VCC_net), .O(n45)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_27_add_3_2_lut.LUT_INIT = 16'h8228;
    SB_CARRY unary_minus_27_add_3_2 (.CI(VCC_net), .I0(GND_net), .I1(n28[0]), 
            .CO(n46173));
    SB_CARRY add_4482_15 (.CI(n47042), .I0(n14525[12]), .I1(n1038), .CO(n47043));
    SB_LUT4 unary_minus_20_add_3_25_lut (.I0(GND_net), .I1(GND_net), .I2(n36[23]), 
            .I3(n46172), .O(n285[23])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4482_14_lut (.I0(GND_net), .I1(n14525[11]), .I2(n965), 
            .I3(n47041), .O(n13879[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4482_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4482_14 (.CI(n47041), .I0(n14525[11]), .I1(n965), .CO(n47042));
    SB_LUT4 add_4621_7_lut (.I0(GND_net), .I1(n16645[4]), .I2(n469), .I3(n46721), 
            .O(n16284[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4621_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4482_13_lut (.I0(GND_net), .I1(n14525[10]), .I2(n892), 
            .I3(n47040), .O(n13879[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4482_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_20_add_3_24_lut (.I0(GND_net), .I1(GND_net), .I2(n36[22]), 
            .I3(n46171), .O(n285[22])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4621_7 (.CI(n46721), .I0(n16645[4]), .I1(n469), .CO(n46722));
    SB_LUT4 add_4621_6_lut (.I0(GND_net), .I1(n16645[3]), .I2(n396), .I3(n46720), 
            .O(n16284[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4621_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4621_6 (.CI(n46720), .I0(n16645[3]), .I1(n396), .CO(n46721));
    SB_CARRY add_4482_13 (.CI(n47040), .I0(n14525[10]), .I1(n892), .CO(n47041));
    SB_LUT4 add_4621_5_lut (.I0(GND_net), .I1(n16645[2]), .I2(n323), .I3(n46719), 
            .O(n16284[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4621_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4621_5 (.CI(n46719), .I0(n16645[2]), .I1(n323), .CO(n46720));
    SB_LUT4 add_4482_12_lut (.I0(GND_net), .I1(n14525[9]), .I2(n819), 
            .I3(n47039), .O(n13879[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4482_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4621_4_lut (.I0(GND_net), .I1(n16645[1]), .I2(n250), .I3(n46718), 
            .O(n16284[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4621_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4621_4 (.CI(n46718), .I0(n16645[1]), .I1(n250), .CO(n46719));
    SB_CARRY unary_minus_20_add_3_24 (.CI(n46171), .I0(GND_net), .I1(n36[22]), 
            .CO(n46172));
    SB_LUT4 unary_minus_20_add_3_23_lut (.I0(GND_net), .I1(GND_net), .I2(n36[21]), 
            .I3(n46170), .O(n285[21])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4621_3_lut (.I0(GND_net), .I1(n16645[0]), .I2(n177), .I3(n46717), 
            .O(n16284[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4621_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4621_3 (.CI(n46717), .I0(n16645[0]), .I1(n177), .CO(n46718));
    SB_LUT4 add_16_12_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [10]), 
            .I2(n207[14]), .I3(n46059), .O(n233[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_16_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_20_add_3_23 (.CI(n46170), .I0(GND_net), .I1(n36[21]), 
            .CO(n46171));
    SB_LUT4 unary_minus_20_add_3_22_lut (.I0(GND_net), .I1(GND_net), .I2(n36[20]), 
            .I3(n46169), .O(n285[20])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4621_2_lut (.I0(GND_net), .I1(n35_c), .I2(n104), .I3(GND_net), 
            .O(n16284[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4621_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4621_2 (.CI(GND_net), .I0(n35_c), .I1(n104), .CO(n46717));
    SB_CARRY add_16_12 (.CI(n46059), .I0(\PID_CONTROLLER.integral [10]), 
            .I1(n207[14]), .CO(n46060));
    SB_CARRY add_4482_12 (.CI(n47039), .I0(n14525[9]), .I1(n819), .CO(n47040));
    SB_LUT4 add_4646_13_lut (.I0(GND_net), .I1(n16954[10]), .I2(n910), 
            .I3(n46716), .O(n16645[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4646_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4646_12_lut (.I0(GND_net), .I1(n16954[9]), .I2(n837), 
            .I3(n46715), .O(n16645[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4646_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4482_11_lut (.I0(GND_net), .I1(n14525[8]), .I2(n746), 
            .I3(n47038), .O(n13879[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4482_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4646_12 (.CI(n46715), .I0(n16954[9]), .I1(n837), .CO(n46716));
    SB_CARRY add_4482_11 (.CI(n47038), .I0(n14525[8]), .I1(n746), .CO(n47039));
    SB_CARRY unary_minus_20_add_3_22 (.CI(n46169), .I0(GND_net), .I1(n36[20]), 
            .CO(n46170));
    SB_LUT4 add_4646_11_lut (.I0(GND_net), .I1(n16954[8]), .I2(n764), 
            .I3(n46714), .O(n16645[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4646_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4646_11 (.CI(n46714), .I0(n16954[8]), .I1(n764), .CO(n46715));
    SB_LUT4 unary_minus_20_add_3_21_lut (.I0(GND_net), .I1(GND_net), .I2(n36[19]), 
            .I3(n46168), .O(n285[19])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4482_10_lut (.I0(GND_net), .I1(n14525[7]), .I2(n673), 
            .I3(n47037), .O(n13879[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4482_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_20_add_3_21 (.CI(n46168), .I0(GND_net), .I1(n36[19]), 
            .CO(n46169));
    SB_LUT4 add_4646_10_lut (.I0(GND_net), .I1(n16954[7]), .I2(n691), 
            .I3(n46713), .O(n16645[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4646_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_20_add_3_20_lut (.I0(GND_net), .I1(GND_net), .I2(n36[18]), 
            .I3(n46167), .O(n285[18])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4482_10 (.CI(n47037), .I0(n14525[7]), .I1(n673), .CO(n47038));
    SB_LUT4 add_4482_9_lut (.I0(GND_net), .I1(n14525[6]), .I2(n600), .I3(n47036), 
            .O(n13879[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4482_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4482_9 (.CI(n47036), .I0(n14525[6]), .I1(n600), .CO(n47037));
    SB_LUT4 add_16_11_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [9]), 
            .I2(n207[13]), .I3(n46058), .O(n233[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_16_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4646_10 (.CI(n46713), .I0(n16954[7]), .I1(n691), .CO(n46714));
    SB_LUT4 add_4646_9_lut (.I0(GND_net), .I1(n16954[6]), .I2(n618), .I3(n46712), 
            .O(n16645[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4646_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4646_9 (.CI(n46712), .I0(n16954[6]), .I1(n618), .CO(n46713));
    SB_CARRY unary_minus_20_add_3_20 (.CI(n46167), .I0(GND_net), .I1(n36[18]), 
            .CO(n46168));
    SB_LUT4 add_4482_8_lut (.I0(GND_net), .I1(n14525[5]), .I2(n527), .I3(n47035), 
            .O(n13879[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4482_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4646_8_lut (.I0(GND_net), .I1(n16954[5]), .I2(n545), .I3(n46711), 
            .O(n16645[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4646_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4646_8 (.CI(n46711), .I0(n16954[5]), .I1(n545), .CO(n46712));
    SB_LUT4 unary_minus_20_add_3_19_lut (.I0(GND_net), .I1(GND_net), .I2(n36[17]), 
            .I3(n46166), .O(n292)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4482_8 (.CI(n47035), .I0(n14525[5]), .I1(n527), .CO(n47036));
    SB_LUT4 add_4646_7_lut (.I0(GND_net), .I1(n16954[4]), .I2(n472), .I3(n46710), 
            .O(n16645[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4646_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4646_7 (.CI(n46710), .I0(n16954[4]), .I1(n472), .CO(n46711));
    SB_CARRY unary_minus_20_add_3_19 (.CI(n46166), .I0(GND_net), .I1(n36[17]), 
            .CO(n46167));
    SB_LUT4 add_4646_6_lut (.I0(GND_net), .I1(n16954[3]), .I2(n399), .I3(n46709), 
            .O(n16645[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4646_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_20_add_3_18_lut (.I0(GND_net), .I1(GND_net), .I2(n36[16]), 
            .I3(n46165), .O(n285[16])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4646_6 (.CI(n46709), .I0(n16954[3]), .I1(n399), .CO(n46710));
    SB_CARRY add_16_11 (.CI(n46058), .I0(\PID_CONTROLLER.integral [9]), 
            .I1(n207[13]), .CO(n46059));
    SB_LUT4 add_4482_7_lut (.I0(GND_net), .I1(n14525[4]), .I2(n454), .I3(n47034), 
            .O(n13879[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4482_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4646_5_lut (.I0(GND_net), .I1(n16954[2]), .I2(n326), .I3(n46708), 
            .O(n16645[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4646_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4646_5 (.CI(n46708), .I0(n16954[2]), .I1(n326), .CO(n46709));
    SB_CARRY add_4482_7 (.CI(n47034), .I0(n14525[4]), .I1(n454), .CO(n47035));
    SB_LUT4 add_4646_4_lut (.I0(GND_net), .I1(n16954[1]), .I2(n253), .I3(n46707), 
            .O(n16645[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4646_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4646_4 (.CI(n46707), .I0(n16954[1]), .I1(n253), .CO(n46708));
    SB_CARRY unary_minus_20_add_3_18 (.CI(n46165), .I0(GND_net), .I1(n36[16]), 
            .CO(n46166));
    SB_LUT4 add_4646_3_lut (.I0(GND_net), .I1(n16954[0]), .I2(n180), .I3(n46706), 
            .O(n16645[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4646_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_16_10_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [8]), 
            .I2(n207[12]), .I3(n46057), .O(n233[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_16_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4646_3 (.CI(n46706), .I0(n16954[0]), .I1(n180), .CO(n46707));
    SB_LUT4 add_4482_6_lut (.I0(GND_net), .I1(n14525[3]), .I2(n381), .I3(n47033), 
            .O(n13879[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4482_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4646_2_lut (.I0(GND_net), .I1(n38), .I2(n107), .I3(GND_net), 
            .O(n16645[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4646_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4646_2 (.CI(GND_net), .I0(n38), .I1(n107), .CO(n46706));
    SB_LUT4 unary_minus_20_add_3_17_lut (.I0(GND_net), .I1(GND_net), .I2(n36[15]), 
            .I3(n46164), .O(n285[15])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4746_8_lut (.I0(GND_net), .I1(n17891[5]), .I2(n560), .I3(n46705), 
            .O(n17795[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4746_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4482_6 (.CI(n47033), .I0(n14525[3]), .I1(n381), .CO(n47034));
    SB_LUT4 add_4482_5_lut (.I0(GND_net), .I1(n14525[2]), .I2(n308), .I3(n47032), 
            .O(n13879[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4482_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4746_7_lut (.I0(GND_net), .I1(n17891[4]), .I2(n487), .I3(n46704), 
            .O(n17795[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4746_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4482_5 (.CI(n47032), .I0(n14525[2]), .I1(n308), .CO(n47033));
    SB_CARRY add_4746_7 (.CI(n46704), .I0(n17891[4]), .I1(n487), .CO(n46705));
    SB_LUT4 add_4746_6_lut (.I0(GND_net), .I1(n17891[3]), .I2(n414), .I3(n46703), 
            .O(n17795[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4746_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4746_6 (.CI(n46703), .I0(n17891[3]), .I1(n414), .CO(n46704));
    SB_LUT4 add_4746_5_lut (.I0(GND_net), .I1(n17891[2]), .I2(n341_c), 
            .I3(n46702), .O(n17795[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4746_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4746_5 (.CI(n46702), .I0(n17891[2]), .I1(n341_c), .CO(n46703));
    SB_LUT4 add_4746_4_lut (.I0(GND_net), .I1(n17891[1]), .I2(n268), .I3(n46701), 
            .O(n17795[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4746_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4482_4_lut (.I0(GND_net), .I1(n14525[1]), .I2(n235), .I3(n47031), 
            .O(n13879[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4482_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4746_4 (.CI(n46701), .I0(n17891[1]), .I1(n268), .CO(n46702));
    SB_LUT4 add_4746_3_lut (.I0(GND_net), .I1(n17891[0]), .I2(n195), .I3(n46700), 
            .O(n17795[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4746_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4482_4 (.CI(n47031), .I0(n14525[1]), .I1(n235), .CO(n47032));
    SB_CARRY unary_minus_20_add_3_17 (.CI(n46164), .I0(GND_net), .I1(n36[15]), 
            .CO(n46165));
    SB_CARRY add_4746_3 (.CI(n46700), .I0(n17891[0]), .I1(n195), .CO(n46701));
    SB_LUT4 unary_minus_20_add_3_16_lut (.I0(GND_net), .I1(GND_net), .I2(n36[14]), 
            .I3(n46163), .O(n285[14])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4746_2_lut (.I0(GND_net), .I1(n53_c), .I2(n122), .I3(GND_net), 
            .O(n17795[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4746_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4746_2 (.CI(GND_net), .I0(n53_c), .I1(n122), .CO(n46700));
    SB_LUT4 add_4482_3_lut (.I0(GND_net), .I1(n14525[0]), .I2(n162), .I3(n47030), 
            .O(n13879[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4482_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4669_12_lut (.I0(GND_net), .I1(n17215[9]), .I2(n840), 
            .I3(n46699), .O(n16954[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4669_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4482_3 (.CI(n47030), .I0(n14525[0]), .I1(n162), .CO(n47031));
    SB_LUT4 add_4482_2_lut (.I0(GND_net), .I1(n20), .I2(n89), .I3(GND_net), 
            .O(n13879[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4482_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4669_11_lut (.I0(GND_net), .I1(n17215[8]), .I2(n767), 
            .I3(n46698), .O(n16954[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4669_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4669_11 (.CI(n46698), .I0(n17215[8]), .I1(n767), .CO(n46699));
    SB_CARRY add_4482_2 (.CI(GND_net), .I0(n20), .I1(n89), .CO(n47030));
    SB_LUT4 add_4669_10_lut (.I0(GND_net), .I1(n17215[7]), .I2(n694), 
            .I3(n46697), .O(n16954[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4669_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_24_i220_2_lut (.I0(\Ki[4] ), .I1(n348), .I2(GND_net), 
            .I3(GND_net), .O(n326));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i220_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i306_2_lut (.I0(\Kp[6] ), .I1(n207[9]), .I2(GND_net), 
            .I3(GND_net), .O(n454));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i306_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_4516_18_lut (.I0(GND_net), .I1(n15101[15]), .I2(GND_net), 
            .I3(n47029), .O(n14525[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4516_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4516_17_lut (.I0(GND_net), .I1(n15101[14]), .I2(GND_net), 
            .I3(n47028), .O(n14525[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4516_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4669_10 (.CI(n46697), .I0(n17215[7]), .I1(n694), .CO(n46698));
    SB_CARRY add_4516_17 (.CI(n47028), .I0(n15101[14]), .I1(GND_net), 
            .CO(n47029));
    SB_LUT4 add_4669_9_lut (.I0(GND_net), .I1(n17215[6]), .I2(n621), .I3(n46696), 
            .O(n16954[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4669_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4516_16_lut (.I0(GND_net), .I1(n15101[13]), .I2(n1114), 
            .I3(n47027), .O(n14525[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4516_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4516_16 (.CI(n47027), .I0(n15101[13]), .I1(n1114), .CO(n47028));
    SB_CARRY add_4669_9 (.CI(n46696), .I0(n17215[6]), .I1(n621), .CO(n46697));
    SB_CARRY unary_minus_20_add_3_16 (.CI(n46163), .I0(GND_net), .I1(n36[14]), 
            .CO(n46164));
    SB_LUT4 add_16_9_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [7]), 
            .I2(n207[11]), .I3(n46056), .O(n233[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_16_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_20_inv_0_i17_1_lut (.I0(IntegralLimit[16]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n36[16]));   // verilog/motorControl.v(59[24:38])
    defparam unary_minus_20_inv_0_i17_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_4516_15_lut (.I0(GND_net), .I1(n15101[12]), .I2(n1041), 
            .I3(n47026), .O(n14525[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4516_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4669_8_lut (.I0(GND_net), .I1(n17215[5]), .I2(n548), .I3(n46695), 
            .O(n16954[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4669_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4516_15 (.CI(n47026), .I0(n15101[12]), .I1(n1041), .CO(n47027));
    SB_CARRY add_4669_8 (.CI(n46695), .I0(n17215[5]), .I1(n548), .CO(n46696));
    SB_LUT4 add_4516_14_lut (.I0(GND_net), .I1(n15101[11]), .I2(n968), 
            .I3(n47025), .O(n14525[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4516_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4669_7_lut (.I0(GND_net), .I1(n17215[4]), .I2(n475), .I3(n46694), 
            .O(n16954[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4669_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_20_add_3_15_lut (.I0(GND_net), .I1(GND_net), .I2(n36[13]), 
            .I3(n46162), .O(n285[13])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_16_9 (.CI(n46056), .I0(\PID_CONTROLLER.integral [7]), .I1(n207[11]), 
            .CO(n46057));
    SB_CARRY add_4516_14 (.CI(n47025), .I0(n15101[11]), .I1(n968), .CO(n47026));
    SB_CARRY add_4669_7 (.CI(n46694), .I0(n17215[4]), .I1(n475), .CO(n46695));
    SB_CARRY unary_minus_20_add_3_15 (.CI(n46162), .I0(GND_net), .I1(n36[13]), 
            .CO(n46163));
    SB_LUT4 add_16_8_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [6]), 
            .I2(n207[10]), .I3(n46055), .O(n233[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_16_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4516_13_lut (.I0(GND_net), .I1(n15101[10]), .I2(n895), 
            .I3(n47024), .O(n14525[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4516_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4516_13 (.CI(n47024), .I0(n15101[10]), .I1(n895), .CO(n47025));
    SB_LUT4 add_4669_6_lut (.I0(GND_net), .I1(n17215[3]), .I2(n402), .I3(n46693), 
            .O(n16954[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4669_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4516_12_lut (.I0(GND_net), .I1(n15101[9]), .I2(n822), 
            .I3(n47023), .O(n14525[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4516_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4669_6 (.CI(n46693), .I0(n17215[3]), .I1(n402), .CO(n46694));
    SB_CARRY add_4516_12 (.CI(n47023), .I0(n15101[9]), .I1(n822), .CO(n47024));
    SB_LUT4 add_4669_5_lut (.I0(GND_net), .I1(n17215[2]), .I2(n329), .I3(n46692), 
            .O(n16954[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4669_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_20_add_3_14_lut (.I0(GND_net), .I1(GND_net), .I2(n36[12]), 
            .I3(n46161), .O(n285[12])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4669_5 (.CI(n46692), .I0(n17215[2]), .I1(n329), .CO(n46693));
    SB_LUT4 add_4516_11_lut (.I0(GND_net), .I1(n15101[8]), .I2(n749), 
            .I3(n47022), .O(n14525[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4516_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4669_4_lut (.I0(GND_net), .I1(n17215[1]), .I2(n256), .I3(n46691), 
            .O(n16954[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4669_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4516_11 (.CI(n47022), .I0(n15101[8]), .I1(n749), .CO(n47023));
    SB_CARRY add_4669_4 (.CI(n46691), .I0(n17215[1]), .I1(n256), .CO(n46692));
    SB_LUT4 add_4516_10_lut (.I0(GND_net), .I1(n15101[7]), .I2(n676), 
            .I3(n47021), .O(n14525[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4516_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4669_3_lut (.I0(GND_net), .I1(n17215[0]), .I2(n183), .I3(n46690), 
            .O(n16954[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4669_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_20_add_3_14 (.CI(n46161), .I0(GND_net), .I1(n36[12]), 
            .CO(n46162));
    SB_CARRY add_4669_3 (.CI(n46690), .I0(n17215[0]), .I1(n183), .CO(n46691));
    SB_CARRY add_4516_10 (.CI(n47021), .I0(n15101[7]), .I1(n676), .CO(n47022));
    SB_LUT4 add_4669_2_lut (.I0(GND_net), .I1(n41), .I2(n110), .I3(GND_net), 
            .O(n16954[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4669_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_20_add_3_13_lut (.I0(GND_net), .I1(GND_net), .I2(n36[11]), 
            .I3(n46160), .O(n285[11])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_16_8 (.CI(n46055), .I0(\PID_CONTROLLER.integral [6]), .I1(n207[10]), 
            .CO(n46056));
    SB_LUT4 add_16_7_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [5]), 
            .I2(n207[9]), .I3(n46054), .O(n233[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_16_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4669_2 (.CI(GND_net), .I0(n41), .I1(n110), .CO(n46690));
    SB_LUT4 add_4516_9_lut (.I0(GND_net), .I1(n15101[6]), .I2(n603), .I3(n47020), 
            .O(n14525[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4516_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4516_9 (.CI(n47020), .I0(n15101[6]), .I1(n603), .CO(n47021));
    SB_LUT4 add_4516_8_lut (.I0(GND_net), .I1(n15101[5]), .I2(n530), .I3(n47019), 
            .O(n14525[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4516_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_20_add_3_13 (.CI(n46160), .I0(GND_net), .I1(n36[11]), 
            .CO(n46161));
    SB_CARRY add_4516_8 (.CI(n47019), .I0(n15101[5]), .I1(n530), .CO(n47020));
    SB_LUT4 unary_minus_20_add_3_12_lut (.I0(GND_net), .I1(GND_net), .I2(n36[10]), 
            .I3(n46159), .O(n285[10])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_24_i375_2_lut (.I0(\Ki[7] ), .I1(n344), .I2(GND_net), 
            .I3(GND_net), .O(n557));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i375_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_4516_7_lut (.I0(GND_net), .I1(n15101[4]), .I2(n457), .I3(n47018), 
            .O(n14525[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4516_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4516_7 (.CI(n47018), .I0(n15101[4]), .I1(n457), .CO(n47019));
    SB_CARRY unary_minus_20_add_3_12 (.CI(n46159), .I0(GND_net), .I1(n36[10]), 
            .CO(n46160));
    SB_LUT4 unary_minus_20_add_3_11_lut (.I0(GND_net), .I1(GND_net), .I2(n36[9]), 
            .I3(n46158), .O(n285[9])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4516_6_lut (.I0(GND_net), .I1(n15101[3]), .I2(n384), .I3(n47017), 
            .O(n14525[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4516_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4516_6 (.CI(n47017), .I0(n15101[3]), .I1(n384), .CO(n47018));
    SB_LUT4 add_4516_5_lut (.I0(GND_net), .I1(n15101[2]), .I2(n311), .I3(n47016), 
            .O(n14525[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4516_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_20_add_3_11 (.CI(n46158), .I0(GND_net), .I1(n36[9]), 
            .CO(n46159));
    SB_CARRY add_16_7 (.CI(n46054), .I0(\PID_CONTROLLER.integral [5]), .I1(n207[9]), 
            .CO(n46055));
    SB_CARRY add_4516_5 (.CI(n47016), .I0(n15101[2]), .I1(n311), .CO(n47017));
    SB_LUT4 unary_minus_20_add_3_10_lut (.I0(GND_net), .I1(GND_net), .I2(n36[8]), 
            .I3(n46157), .O(n285[8])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_16_6_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [4]), 
            .I2(n207[8]), .I3(n46053), .O(n233[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_16_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_16_6 (.CI(n46053), .I0(\PID_CONTROLLER.integral [4]), .I1(n207[8]), 
            .CO(n46054));
    SB_LUT4 add_4516_4_lut (.I0(GND_net), .I1(n15101[1]), .I2(n238), .I3(n47015), 
            .O(n14525[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4516_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_20_add_3_10 (.CI(n46157), .I0(GND_net), .I1(n36[8]), 
            .CO(n46158));
    SB_LUT4 add_16_5_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [3]), 
            .I2(n207[7]), .I3(n46052), .O(n233[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_16_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4516_4 (.CI(n47015), .I0(n15101[1]), .I1(n238), .CO(n47016));
    SB_LUT4 unary_minus_20_add_3_9_lut (.I0(GND_net), .I1(GND_net), .I2(n36[7]), 
            .I3(n46156), .O(n285[7])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_24_i38_2_lut (.I0(\Ki[0] ), .I1(n341), .I2(GND_net), 
            .I3(GND_net), .O(n56));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i38_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i69_2_lut (.I0(\Kp[1] ), .I1(n207[13]), .I2(GND_net), 
            .I3(GND_net), .O(n101));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i69_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i22_2_lut (.I0(\Kp[0] ), .I1(n207[14]), .I2(GND_net), 
            .I3(GND_net), .O(n32));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i22_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i269_2_lut (.I0(\Ki[5] ), .I1(n348), .I2(GND_net), 
            .I3(GND_net), .O(n399));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i269_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_16_5 (.CI(n46052), .I0(\PID_CONTROLLER.integral [3]), .I1(n207[7]), 
            .CO(n46053));
    SB_CARRY unary_minus_20_add_3_9 (.CI(n46156), .I0(GND_net), .I1(n36[7]), 
            .CO(n46157));
    SB_LUT4 unary_minus_20_add_3_8_lut (.I0(GND_net), .I1(GND_net), .I2(n36[6]), 
            .I3(n46155), .O(n285[6])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_24_i318_2_lut (.I0(\Ki[6] ), .I1(n348), .I2(GND_net), 
            .I3(GND_net), .O(n472));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i318_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_20_inv_0_i18_1_lut (.I0(IntegralLimit[17]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n36[17]));   // verilog/motorControl.v(59[24:38])
    defparam unary_minus_20_inv_0_i18_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_24_i367_2_lut (.I0(\Ki[7] ), .I1(n348), .I2(GND_net), 
            .I3(GND_net), .O(n545));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i367_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i355_2_lut (.I0(\Kp[7] ), .I1(n207[9]), .I2(GND_net), 
            .I3(GND_net), .O(n527));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i355_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_4516_3_lut (.I0(GND_net), .I1(n15101[0]), .I2(n165), .I3(n47014), 
            .O(n14525[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4516_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4516_3 (.CI(n47014), .I0(n15101[0]), .I1(n165), .CO(n47015));
    SB_LUT4 mult_24_i416_2_lut (.I0(\Ki[8] ), .I1(n348), .I2(GND_net), 
            .I3(GND_net), .O(n618));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i416_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_4516_2_lut (.I0(GND_net), .I1(n23), .I2(n92), .I3(GND_net), 
            .O(n14525[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4516_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_23_i404_2_lut (.I0(\Kp[8] ), .I1(n207[9]), .I2(GND_net), 
            .I3(GND_net), .O(n600));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i404_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_4516_2 (.CI(GND_net), .I0(n23), .I1(n92), .CO(n47014));
    SB_LUT4 add_4741_8_lut (.I0(GND_net), .I1(n17859[5]), .I2(n560_adj_4214), 
            .I3(n47013), .O(n17750[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4741_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_20_add_3_8 (.CI(n46155), .I0(GND_net), .I1(n36[6]), 
            .CO(n46156));
    SB_LUT4 LessThan_17_i45_2_lut (.I0(IntegralLimit[22]), .I1(n233[22]), 
            .I2(GND_net), .I3(GND_net), .O(n45_adj_4216));   // verilog/motorControl.v(56[14:36])
    defparam LessThan_17_i45_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_17_i39_2_lut (.I0(IntegralLimit[19]), .I1(n233[19]), 
            .I2(GND_net), .I3(GND_net), .O(n39));   // verilog/motorControl.v(56[14:36])
    defparam LessThan_17_i39_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 unary_minus_20_add_3_7_lut (.I0(GND_net), .I1(GND_net), .I2(n36[5]), 
            .I3(n46154), .O(n285[5])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_20_inv_0_i19_1_lut (.I0(IntegralLimit[18]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n36[18]));   // verilog/motorControl.v(59[24:38])
    defparam unary_minus_20_inv_0_i19_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_24_i465_2_lut (.I0(\Ki[9] ), .I1(n348), .I2(GND_net), 
            .I3(GND_net), .O(n691));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i465_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i453_2_lut (.I0(\Kp[9] ), .I1(n207[9]), .I2(GND_net), 
            .I3(GND_net), .O(n673));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i453_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_17_i41_2_lut (.I0(IntegralLimit[20]), .I1(n233[20]), 
            .I2(GND_net), .I3(GND_net), .O(n41_adj_4219));   // verilog/motorControl.v(56[14:36])
    defparam LessThan_17_i41_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_17_i43_2_lut (.I0(IntegralLimit[21]), .I1(n233[21]), 
            .I2(GND_net), .I3(GND_net), .O(n43));   // verilog/motorControl.v(56[14:36])
    defparam LessThan_17_i43_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_17_i37_2_lut (.I0(IntegralLimit[18]), .I1(n233[18]), 
            .I2(GND_net), .I3(GND_net), .O(n37));   // verilog/motorControl.v(56[14:36])
    defparam LessThan_17_i37_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 unary_minus_20_inv_0_i20_1_lut (.I0(IntegralLimit[19]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n36[19]));   // verilog/motorControl.v(59[24:38])
    defparam unary_minus_20_inv_0_i20_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_24_i514_2_lut (.I0(\Ki[10] ), .I1(n348), .I2(GND_net), 
            .I3(GND_net), .O(n764));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i514_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_4741_7_lut (.I0(GND_net), .I1(n17859[4]), .I2(n487_adj_4220), 
            .I3(n47012), .O(n17750[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4741_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_23_i502_2_lut (.I0(\Kp[10] ), .I1(n207[9]), .I2(GND_net), 
            .I3(GND_net), .O(n746));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i502_2_lut.LUT_INIT = 16'h8888;
    SB_DFFER result_i0_i0 (.Q(duty[0]), .C(clk16MHz), .E(control_update), 
            .D(n63680), .R(reset));   // verilog/motorControl.v(42[14] 73[8])
    SB_CARRY unary_minus_20_add_3_7 (.CI(n46154), .I0(GND_net), .I1(n36[5]), 
            .CO(n46155));
    SB_LUT4 unary_minus_20_add_3_6_lut (.I0(GND_net), .I1(GND_net), .I2(n36[4]), 
            .I3(n46153), .O(n285[4])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_17_i35_2_lut (.I0(IntegralLimit[17]), .I1(n240), .I2(GND_net), 
            .I3(GND_net), .O(n35_adj_4222));   // verilog/motorControl.v(56[14:36])
    defparam LessThan_17_i35_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY unary_minus_20_add_3_6 (.CI(n46153), .I0(GND_net), .I1(n36[4]), 
            .CO(n46154));
    SB_LUT4 mult_23_i118_2_lut (.I0(\Kp[2] ), .I1(n207[13]), .I2(GND_net), 
            .I3(GND_net), .O(n174));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i118_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_16_4_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [2]), 
            .I2(n207[6]), .I3(n46051), .O(n233[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_16_4_lut.LUT_INIT = 16'hC33C;
    SB_DFF control_update_46 (.Q(control_update), .C(clk16MHz), .D(counter_31__N_3487));   // verilog/motorControl.v(24[10] 31[6])
    SB_CARRY add_4741_7 (.CI(n47012), .I0(n17859[4]), .I1(n487_adj_4220), 
            .CO(n47013));
    SB_LUT4 add_4741_6_lut (.I0(GND_net), .I1(n17859[3]), .I2(n414_adj_4223), 
            .I3(n47011), .O(n17750[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4741_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 n9440_bdd_4_lut_48748 (.I0(n9440), .I1(n59906), .I2(setpoint[20]), 
            .I3(n4357), .O(n63485));
    defparam n9440_bdd_4_lut_48748.LUT_INIT = 16'he4aa;
    SB_LUT4 mult_23_i167_2_lut (.I0(\Kp[3] ), .I1(n207[13]), .I2(GND_net), 
            .I3(GND_net), .O(n247_adj_4224));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i167_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i563_2_lut (.I0(\Ki[11] ), .I1(n348), .I2(GND_net), 
            .I3(GND_net), .O(n837));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i563_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_4741_6 (.CI(n47011), .I0(n17859[3]), .I1(n414_adj_4223), 
            .CO(n47012));
    SB_LUT4 unary_minus_20_add_3_5_lut (.I0(GND_net), .I1(GND_net), .I2(n36[3]), 
            .I3(n46152), .O(n285[3])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_24_i612_2_lut (.I0(\Ki[12] ), .I1(n348), .I2(GND_net), 
            .I3(GND_net), .O(n910));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i612_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY unary_minus_20_add_3_5 (.CI(n46152), .I0(GND_net), .I1(n36[3]), 
            .CO(n46153));
    SB_LUT4 add_4741_5_lut (.I0(GND_net), .I1(n17859[2]), .I2(n341_adj_4226), 
            .I3(n47010), .O(n17750[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4741_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_20_add_3_4_lut (.I0(GND_net), .I1(GND_net), .I2(n36[2]), 
            .I3(n46151), .O(n285[2])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4741_5 (.CI(n47010), .I0(n17859[2]), .I1(n341_adj_4226), 
            .CO(n47011));
    SB_LUT4 mux_21_i12_3_lut (.I0(n233[11]), .I1(n285[11]), .I2(n284), 
            .I3(GND_net), .O(n310[11]));   // verilog/motorControl.v(58[20] 60[14])
    defparam mux_21_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 n63485_bdd_4_lut (.I0(n63485), .I1(n535[20]), .I2(n455[20]), 
            .I3(n4357), .O(n63488));
    defparam n63485_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 LessThan_17_i27_2_lut (.I0(IntegralLimit[13]), .I1(n233[13]), 
            .I2(GND_net), .I3(GND_net), .O(n27));   // verilog/motorControl.v(56[14:36])
    defparam LessThan_17_i27_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mux_22_i12_3_lut (.I0(n310[11]), .I1(IntegralLimit[11]), .I2(n258), 
            .I3(GND_net), .O(n348));   // verilog/motorControl.v(58[20] 60[14])
    defparam mux_22_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_4741_4_lut (.I0(GND_net), .I1(n17859[1]), .I2(n268_adj_4229), 
            .I3(n47009), .O(n17750[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4741_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_20_add_3_4 (.CI(n46151), .I0(GND_net), .I1(n36[2]), 
            .CO(n46152));
    SB_CARRY add_4741_4 (.CI(n47009), .I0(n17859[1]), .I1(n268_adj_4229), 
            .CO(n47010));
    SB_LUT4 unary_minus_20_add_3_3_lut (.I0(GND_net), .I1(GND_net), .I2(n36[1]), 
            .I3(n46150), .O(n285[1])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_16_4 (.CI(n46051), .I0(\PID_CONTROLLER.integral [2]), .I1(n207[6]), 
            .CO(n46052));
    SB_LUT4 mult_23_i216_2_lut (.I0(\Kp[4] ), .I1(n207[13]), .I2(GND_net), 
            .I3(GND_net), .O(n320));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i216_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY unary_minus_20_add_3_3 (.CI(n46150), .I0(GND_net), .I1(n36[1]), 
            .CO(n46151));
    SB_LUT4 n9440_bdd_4_lut_48733 (.I0(n9440), .I1(n59905), .I2(setpoint[19]), 
            .I3(n4357), .O(n63479));
    defparam n9440_bdd_4_lut_48733.LUT_INIT = 16'he4aa;
    SB_LUT4 unary_minus_20_add_3_2_lut (.I0(GND_net), .I1(GND_net), .I2(n36[0]), 
            .I3(VCC_net), .O(n285[0])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_20_add_3_2 (.CI(VCC_net), .I0(GND_net), .I1(n36[0]), 
            .CO(n46150));
    SB_LUT4 LessThan_17_i31_2_lut (.I0(IntegralLimit[15]), .I1(n233[15]), 
            .I2(GND_net), .I3(GND_net), .O(n31));   // verilog/motorControl.v(56[14:36])
    defparam LessThan_17_i31_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_4741_3_lut (.I0(GND_net), .I1(n17859[0]), .I2(n195_adj_4233), 
            .I3(n47008), .O(n17750[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4741_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4741_3 (.CI(n47008), .I0(n17859[0]), .I1(n195_adj_4233), 
            .CO(n47009));
    SB_LUT4 n63479_bdd_4_lut (.I0(n63479), .I1(n535[19]), .I2(n455[19]), 
            .I3(n4357), .O(n63482));
    defparam n63479_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 LessThan_17_i33_2_lut (.I0(IntegralLimit[16]), .I1(n233[16]), 
            .I2(GND_net), .I3(GND_net), .O(n33));   // verilog/motorControl.v(56[14:36])
    defparam LessThan_17_i33_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_24_i71_2_lut (.I0(\Ki[1] ), .I1(n349), .I2(GND_net), 
            .I3(GND_net), .O(n104));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i71_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_16_3_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [1]), 
            .I2(n207[5]), .I3(n46050), .O(n233[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_16_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_17_i29_2_lut (.I0(IntegralLimit[14]), .I1(n233[14]), 
            .I2(GND_net), .I3(GND_net), .O(n29));   // verilog/motorControl.v(56[14:36])
    defparam LessThan_17_i29_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i45654_4_lut (.I0(n21_adj_4235), .I1(n19_adj_4236), .I2(n17_adj_4237), 
            .I3(n9_adj_4238), .O(n60366));
    defparam i45654_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 mult_24_i24_2_lut (.I0(\Ki[0] ), .I1(n348), .I2(GND_net), 
            .I3(GND_net), .O(n35_c));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i24_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_4741_2_lut (.I0(GND_net), .I1(n53), .I2(n122_adj_4240), 
            .I3(GND_net), .O(n17750[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4741_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_20_inv_0_i21_1_lut (.I0(IntegralLimit[20]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n36[20]));   // verilog/motorControl.v(59[24:38])
    defparam unary_minus_20_inv_0_i21_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_4741_2 (.CI(GND_net), .I0(n53), .I1(n122_adj_4240), .CO(n47008));
    SB_LUT4 add_4548_17_lut (.I0(GND_net), .I1(n15611[14]), .I2(GND_net), 
            .I3(n47007), .O(n15101[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4548_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_16_3 (.CI(n46050), .I0(\PID_CONTROLLER.integral [1]), .I1(n207[5]), 
            .CO(n46051));
    SB_LUT4 add_4548_16_lut (.I0(GND_net), .I1(n15611[13]), .I2(n1117), 
            .I3(n47006), .O(n15101[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4548_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4548_16 (.CI(n47006), .I0(n15611[13]), .I1(n1117), .CO(n47007));
    SB_LUT4 add_4548_15_lut (.I0(GND_net), .I1(n15611[12]), .I2(n1044), 
            .I3(n47005), .O(n15101[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4548_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i45614_4_lut (.I0(n27), .I1(n15_adj_4241), .I2(n13_adj_4242), 
            .I3(n11_adj_4243), .O(n60326));
    defparam i45614_4_lut.LUT_INIT = 16'haaab;
    SB_CARRY add_4548_15 (.CI(n47005), .I0(n15611[12]), .I1(n1044), .CO(n47006));
    SB_LUT4 add_4548_14_lut (.I0(GND_net), .I1(n15611[11]), .I2(n971), 
            .I3(n47004), .O(n15101[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4548_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_24_i120_2_lut (.I0(\Ki[2] ), .I1(n349), .I2(GND_net), 
            .I3(GND_net), .O(n177));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i120_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_20_inv_0_i22_1_lut (.I0(IntegralLimit[21]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n36[21]));   // verilog/motorControl.v(59[24:38])
    defparam unary_minus_20_inv_0_i22_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_4548_14 (.CI(n47004), .I0(n15611[11]), .I1(n971), .CO(n47005));
    SB_LUT4 add_4548_13_lut (.I0(GND_net), .I1(n15611[10]), .I2(n898), 
            .I3(n47003), .O(n15101[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4548_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_16_10 (.CI(n46057), .I0(\PID_CONTROLLER.integral [8]), 
            .I1(n207[12]), .CO(n46058));
    SB_LUT4 mult_24_i169_2_lut (.I0(\Ki[3] ), .I1(n349), .I2(GND_net), 
            .I3(GND_net), .O(n250));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i169_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_4548_13 (.CI(n47003), .I0(n15611[10]), .I1(n898), .CO(n47004));
    SB_LUT4 add_4548_12_lut (.I0(GND_net), .I1(n15611[9]), .I2(n825), 
            .I3(n47002), .O(n15101[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4548_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 n9440_bdd_4_lut_48728 (.I0(n9440), .I1(n59904), .I2(setpoint[18]), 
            .I3(n4357), .O(n63467));
    defparam n9440_bdd_4_lut_48728.LUT_INIT = 16'he4aa;
    SB_LUT4 mult_23_i551_2_lut (.I0(\Kp[11] ), .I1(n207[9]), .I2(GND_net), 
            .I3(GND_net), .O(n819));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i551_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 n63467_bdd_4_lut (.I0(n63467), .I1(n535[18]), .I2(n455[18]), 
            .I3(n4357), .O(n63470));
    defparam n63467_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 add_16_2_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [0]), 
            .I2(n207[4]), .I3(GND_net), .O(n233[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_16_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4548_12 (.CI(n47002), .I0(n15611[9]), .I1(n825), .CO(n47003));
    SB_LUT4 add_4548_11_lut (.I0(GND_net), .I1(n15611[8]), .I2(n752), 
            .I3(n47001), .O(n15101[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4548_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_16_2 (.CI(GND_net), .I0(\PID_CONTROLLER.integral [0]), 
            .I1(n207[4]), .CO(n46050));
    SB_LUT4 LessThan_17_i12_3_lut (.I0(n233[7]), .I1(n233[16]), .I2(n33), 
            .I3(GND_net), .O(n12_adj_4244));   // verilog/motorControl.v(56[14:36])
    defparam LessThan_17_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_24_i218_2_lut (.I0(\Ki[4] ), .I1(n349), .I2(GND_net), 
            .I3(GND_net), .O(n323));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i218_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_4548_11 (.CI(n47001), .I0(n15611[8]), .I1(n752), .CO(n47002));
    SB_LUT4 LessThan_17_i10_3_lut (.I0(n233[5]), .I1(n233[6]), .I2(n13_adj_4242), 
            .I3(GND_net), .O(n10_adj_4245));   // verilog/motorControl.v(56[14:36])
    defparam LessThan_17_i10_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_17_i30_3_lut (.I0(n12_adj_4244), .I1(n240), .I2(n35_adj_4222), 
            .I3(GND_net), .O(n30));   // verilog/motorControl.v(56[14:36])
    defparam LessThan_17_i30_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_4548_10_lut (.I0(GND_net), .I1(n15611[7]), .I2(n679), 
            .I3(n47000), .O(n15101[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4548_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4548_10 (.CI(n47000), .I0(n15611[7]), .I1(n679), .CO(n47001));
    SB_LUT4 i46650_4_lut (.I0(n13_adj_4242), .I1(n11_adj_4243), .I2(n9_adj_4238), 
            .I3(n60399), .O(n61363));
    defparam i46650_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 mult_24_i267_2_lut (.I0(\Ki[5] ), .I1(n349), .I2(GND_net), 
            .I3(GND_net), .O(n396));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i267_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_20_inv_0_i23_1_lut (.I0(IntegralLimit[22]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n36[22]));   // verilog/motorControl.v(59[24:38])
    defparam unary_minus_20_inv_0_i23_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i46638_4_lut (.I0(n19_adj_4236), .I1(n17_adj_4237), .I2(n15_adj_4241), 
            .I3(n61363), .O(n61351));
    defparam i46638_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i47918_4_lut (.I0(n25_adj_4246), .I1(n23_adj_4247), .I2(n21_adj_4235), 
            .I3(n61351), .O(n62631));
    defparam i47918_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 add_4548_9_lut (.I0(GND_net), .I1(n15611[6]), .I2(n606), .I3(n46999), 
            .O(n15101[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4548_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_23_i600_2_lut (.I0(\Kp[12] ), .I1(n207[9]), .I2(GND_net), 
            .I3(GND_net), .O(n892));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i600_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i47204_4_lut (.I0(n31), .I1(n29), .I2(n27), .I3(n62631), 
            .O(n61917));
    defparam i47204_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 mult_24_i316_2_lut (.I0(\Ki[6] ), .I1(n349), .I2(GND_net), 
            .I3(GND_net), .O(n469));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i316_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i649_2_lut (.I0(\Kp[13] ), .I1(n207[9]), .I2(GND_net), 
            .I3(GND_net), .O(n965));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i649_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i48056_4_lut (.I0(n37), .I1(n35_adj_4222), .I2(n33), .I3(n61917), 
            .O(n62769));
    defparam i48056_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 unary_minus_20_inv_0_i24_1_lut (.I0(IntegralLimit[23]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n36[23]));   // verilog/motorControl.v(59[24:38])
    defparam unary_minus_20_inv_0_i24_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_4548_9 (.CI(n46999), .I0(n15611[6]), .I1(n606), .CO(n47000));
    SB_LUT4 LessThan_17_i16_3_lut (.I0(n233[9]), .I1(n233[21]), .I2(n43), 
            .I3(GND_net), .O(n16_adj_4248));   // verilog/motorControl.v(56[14:36])
    defparam LessThan_17_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_4548_8_lut (.I0(GND_net), .I1(n15611[5]), .I2(n533), .I3(n46998), 
            .O(n15101[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4548_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i18440_1_lut (.I0(n455[0]), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n31995));   // verilog/motorControl.v(61[20:40])
    defparam i18440_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_27_inv_0_i1_1_lut (.I0(\deadband[0] ), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n28[0]));   // verilog/motorControl.v(62[45:54])
    defparam unary_minus_27_inv_0_i1_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_4548_8 (.CI(n46998), .I0(n15611[5]), .I1(n533), .CO(n46999));
    SB_LUT4 add_4548_7_lut (.I0(GND_net), .I1(n15611[4]), .I2(n460_adj_4249), 
            .I3(n46997), .O(n15101[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4548_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4548_7 (.CI(n46997), .I0(n15611[4]), .I1(n460_adj_4249), 
            .CO(n46998));
    SB_LUT4 add_4548_6_lut (.I0(GND_net), .I1(n15611[3]), .I2(n387), .I3(n46996), 
            .O(n15101[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4548_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4548_6 (.CI(n46996), .I0(n15611[3]), .I1(n387), .CO(n46997));
    SB_LUT4 i47243_3_lut (.I0(n6_adj_4250), .I1(n233[10]), .I2(n21_adj_4235), 
            .I3(GND_net), .O(n61956));   // verilog/motorControl.v(56[14:36])
    defparam i47243_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i47244_3_lut (.I0(n61956), .I1(n233[11]), .I2(n23_adj_4247), 
            .I3(GND_net), .O(n61957));   // verilog/motorControl.v(56[14:36])
    defparam i47244_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_17_i8_3_lut (.I0(n233[4]), .I1(n233[8]), .I2(n17_adj_4237), 
            .I3(GND_net), .O(n8_adj_4251));   // verilog/motorControl.v(56[14:36])
    defparam LessThan_17_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_17_i24_3_lut (.I0(n16_adj_4248), .I1(n233[22]), .I2(n45_adj_4216), 
            .I3(GND_net), .O(n24_adj_4252));   // verilog/motorControl.v(56[14:36])
    defparam LessThan_17_i24_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_4548_5_lut (.I0(GND_net), .I1(n15611[2]), .I2(n314), .I3(n46995), 
            .O(n15101[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4548_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i45470_4_lut (.I0(n43), .I1(n25_adj_4246), .I2(n23_adj_4247), 
            .I3(n60366), .O(n60182));
    defparam i45470_4_lut.LUT_INIT = 16'haaab;
    SB_CARRY add_4548_5 (.CI(n46995), .I0(n15611[2]), .I1(n314), .CO(n46996));
    SB_LUT4 add_4548_4_lut (.I0(GND_net), .I1(n15611[1]), .I2(n241_adj_4253), 
            .I3(n46994), .O(n15101[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4548_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4548_4 (.CI(n46994), .I0(n15611[1]), .I1(n241_adj_4253), 
            .CO(n46995));
    SB_LUT4 add_4548_3_lut (.I0(GND_net), .I1(n15611[0]), .I2(n168), .I3(n46993), 
            .O(n15101[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4548_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4548_3 (.CI(n46993), .I0(n15611[0]), .I1(n168), .CO(n46994));
    SB_LUT4 add_4548_2_lut (.I0(GND_net), .I1(n26), .I2(n95), .I3(GND_net), 
            .O(n15101[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4548_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4548_2 (.CI(GND_net), .I0(n26), .I1(n95), .CO(n46993));
    SB_LUT4 add_4578_16_lut (.I0(GND_net), .I1(n16059[13]), .I2(n1120), 
            .I3(n46992), .O(n15611[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4578_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i47164_4_lut (.I0(n24_adj_4252), .I1(n8_adj_4251), .I2(n45_adj_4216), 
            .I3(n60177), .O(n61877));   // verilog/motorControl.v(56[14:36])
    defparam i47164_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 add_4578_15_lut (.I0(GND_net), .I1(n16059[12]), .I2(n1047), 
            .I3(n46991), .O(n15611[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4578_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4578_15 (.CI(n46991), .I0(n16059[12]), .I1(n1047), .CO(n46992));
    SB_LUT4 add_4578_14_lut (.I0(GND_net), .I1(n16059[11]), .I2(n974), 
            .I3(n46990), .O(n15611[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4578_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4578_14 (.CI(n46990), .I0(n16059[11]), .I1(n974), .CO(n46991));
    SB_LUT4 add_4578_13_lut (.I0(GND_net), .I1(n16059[10]), .I2(n901), 
            .I3(n46989), .O(n15611[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4578_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4578_13 (.CI(n46989), .I0(n16059[10]), .I1(n901), .CO(n46990));
    SB_LUT4 add_4578_12_lut (.I0(GND_net), .I1(n16059[9]), .I2(n828), 
            .I3(n46988), .O(n15611[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4578_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4578_12 (.CI(n46988), .I0(n16059[9]), .I1(n828), .CO(n46989));
    SB_LUT4 add_4578_11_lut (.I0(GND_net), .I1(n16059[8]), .I2(n755), 
            .I3(n46987), .O(n15611[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4578_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4578_11 (.CI(n46987), .I0(n16059[8]), .I1(n755), .CO(n46988));
    SB_LUT4 i46406_3_lut (.I0(n61957), .I1(n233[12]), .I2(n25_adj_4246), 
            .I3(GND_net), .O(n61119));   // verilog/motorControl.v(56[14:36])
    defparam i46406_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_17_i4_4_lut (.I0(n233[0]), .I1(n233[1]), .I2(IntegralLimit[1]), 
            .I3(IntegralLimit[0]), .O(n4_adj_4254));   // verilog/motorControl.v(56[14:36])
    defparam LessThan_17_i4_4_lut.LUT_INIT = 16'h0c8e;
    SB_LUT4 i47241_3_lut (.I0(n4_adj_4254), .I1(n233[13]), .I2(n27), .I3(GND_net), 
            .O(n61954));   // verilog/motorControl.v(56[14:36])
    defparam i47241_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_4578_10_lut (.I0(GND_net), .I1(n16059[7]), .I2(n682), 
            .I3(n46986), .O(n15611[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4578_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4578_10 (.CI(n46986), .I0(n16059[7]), .I1(n682), .CO(n46987));
    SB_LUT4 i47242_3_lut (.I0(n61954), .I1(n233[14]), .I2(n29), .I3(GND_net), 
            .O(n61955));   // verilog/motorControl.v(56[14:36])
    defparam i47242_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_4578_9_lut (.I0(GND_net), .I1(n16059[6]), .I2(n609), .I3(n46985), 
            .O(n15611[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4578_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4578_9 (.CI(n46985), .I0(n16059[6]), .I1(n609), .CO(n46986));
    SB_LUT4 add_4578_8_lut (.I0(GND_net), .I1(n16059[5]), .I2(n536), .I3(n46984), 
            .O(n15611[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4578_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4578_8 (.CI(n46984), .I0(n16059[5]), .I1(n536), .CO(n46985));
    SB_LUT4 i45523_4_lut (.I0(n33), .I1(n31), .I2(n29), .I3(n60326), 
            .O(n60235));
    defparam i45523_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 add_4578_7_lut (.I0(GND_net), .I1(n16059[4]), .I2(n463), .I3(n46983), 
            .O(n15611[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4578_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4578_7 (.CI(n46983), .I0(n16059[4]), .I1(n463), .CO(n46984));
    SB_LUT4 add_4578_6_lut (.I0(GND_net), .I1(n16059[3]), .I2(n390), .I3(n46982), 
            .O(n15611[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4578_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4578_6 (.CI(n46982), .I0(n16059[3]), .I1(n390), .CO(n46983));
    SB_LUT4 add_4578_5_lut (.I0(GND_net), .I1(n16059[2]), .I2(n317), .I3(n46981), 
            .O(n15611[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4578_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4578_5 (.CI(n46981), .I0(n16059[2]), .I1(n317), .CO(n46982));
    SB_LUT4 add_4578_4_lut (.I0(GND_net), .I1(n16059[1]), .I2(n244_adj_4255), 
            .I3(n46980), .O(n15611[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4578_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4578_4 (.CI(n46980), .I0(n16059[1]), .I1(n244_adj_4255), 
            .CO(n46981));
    SB_LUT4 i47689_4_lut (.I0(n30), .I1(n10_adj_4245), .I2(n35_adj_4222), 
            .I3(n60223), .O(n62402));   // verilog/motorControl.v(56[14:36])
    defparam i47689_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 add_4578_3_lut (.I0(GND_net), .I1(n16059[0]), .I2(n171), .I3(n46979), 
            .O(n15611[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4578_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4578_3 (.CI(n46979), .I0(n16059[0]), .I1(n171), .CO(n46980));
    SB_LUT4 add_4578_2_lut (.I0(GND_net), .I1(n29_adj_4256), .I2(n98), 
            .I3(GND_net), .O(n15611[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4578_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i46408_3_lut (.I0(n61955), .I1(n233[15]), .I2(n31), .I3(GND_net), 
            .O(n61121));   // verilog/motorControl.v(56[14:36])
    defparam i46408_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i48089_4_lut (.I0(n61121), .I1(n62402), .I2(n35_adj_4222), 
            .I3(n60235), .O(n62802));   // verilog/motorControl.v(56[14:36])
    defparam i48089_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i48090_3_lut (.I0(n62802), .I1(n233[18]), .I2(n37), .I3(GND_net), 
            .O(n62803));   // verilog/motorControl.v(56[14:36])
    defparam i48090_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut (.I0(n17997[2]), .I1(n6_adj_4257), .I2(\Ki[4] ), 
            .I3(n341), .O(n17940[3]));   // verilog/motorControl.v(61[29:40])
    defparam i1_4_lut.LUT_INIT = 16'h9666;
    SB_LUT4 i48088_3_lut (.I0(n62803), .I1(n233[19]), .I2(n39), .I3(GND_net), 
            .O(n62801));   // verilog/motorControl.v(56[14:36])
    defparam i48088_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i45481_4_lut (.I0(n43), .I1(n41_adj_4219), .I2(n39), .I3(n62769), 
            .O(n60193));
    defparam i45481_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i47840_4_lut (.I0(n61119), .I1(n61877), .I2(n45_adj_4216), 
            .I3(n60182), .O(n62553));   // verilog/motorControl.v(56[14:36])
    defparam i47840_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i46414_3_lut (.I0(n62801), .I1(n233[20]), .I2(n41_adj_4219), 
            .I3(GND_net), .O(n61127));   // verilog/motorControl.v(56[14:36])
    defparam i46414_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i48040_4_lut (.I0(n61127), .I1(n62553), .I2(n45_adj_4216), 
            .I3(n60193), .O(n62753));   // verilog/motorControl.v(56[14:36])
    defparam i48040_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i48041_3_lut (.I0(n62753), .I1(IntegralLimit[23]), .I2(n233[23]), 
            .I3(GND_net), .O(n258));   // verilog/motorControl.v(56[14:36])
    defparam i48041_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 LessThan_19_i45_2_lut (.I0(n233[22]), .I1(n285[22]), .I2(GND_net), 
            .I3(GND_net), .O(n45_adj_4258));   // verilog/motorControl.v(58[23:46])
    defparam LessThan_19_i45_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_19_i41_2_lut (.I0(n233[20]), .I1(n285[20]), .I2(GND_net), 
            .I3(GND_net), .O(n41_adj_4259));   // verilog/motorControl.v(58[23:46])
    defparam LessThan_19_i41_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_4_lut_adj_928 (.I0(n18055[0]), .I1(n45772), .I2(\Ki[2] ), 
            .I3(n339), .O(n18034[1]));   // verilog/motorControl.v(61[29:40])
    defparam i1_4_lut_adj_928.LUT_INIT = 16'h9666;
    SB_LUT4 mux_21_i22_3_lut (.I0(n233[21]), .I1(n285[21]), .I2(n284), 
            .I3(GND_net), .O(n310[21]));   // verilog/motorControl.v(58[20] 60[14])
    defparam mux_21_i22_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_19_i43_2_lut (.I0(n233[21]), .I1(n285[21]), .I2(GND_net), 
            .I3(GND_net), .O(n43_adj_4260));   // verilog/motorControl.v(58[23:46])
    defparam LessThan_19_i43_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_19_i39_2_lut (.I0(n233[19]), .I1(n285[19]), .I2(GND_net), 
            .I3(GND_net), .O(n39_adj_4261));   // verilog/motorControl.v(58[23:46])
    defparam LessThan_19_i39_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mux_22_i22_3_lut (.I0(n310[21]), .I1(IntegralLimit[21]), .I2(n258), 
            .I3(GND_net), .O(n338));   // verilog/motorControl.v(58[20] 60[14])
    defparam mux_22_i22_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_21_i21_3_lut (.I0(n233[20]), .I1(n285[20]), .I2(n284), 
            .I3(GND_net), .O(n310[20]));   // verilog/motorControl.v(58[20] 60[14])
    defparam mux_21_i21_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_22_i21_3_lut (.I0(n310[20]), .I1(IntegralLimit[20]), .I2(n258), 
            .I3(GND_net), .O(n339));   // verilog/motorControl.v(58[20] 60[14])
    defparam mux_22_i21_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_19_i37_2_lut (.I0(n233[18]), .I1(n285[18]), .I2(GND_net), 
            .I3(GND_net), .O(n37_adj_4264));   // verilog/motorControl.v(58[23:46])
    defparam LessThan_19_i37_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mux_21_i24_3_lut (.I0(n233[23]), .I1(n285[23]), .I2(n284), 
            .I3(GND_net), .O(n310[23]));   // verilog/motorControl.v(58[20] 60[14])
    defparam mux_21_i24_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_22_i24_3_lut (.I0(n310[23]), .I1(IntegralLimit[23]), .I2(n258), 
            .I3(GND_net), .O(n336));   // verilog/motorControl.v(58[20] 60[14])
    defparam mux_22_i24_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_21_i23_3_lut (.I0(n233[22]), .I1(n285[22]), .I2(n284), 
            .I3(GND_net), .O(n310[22]));   // verilog/motorControl.v(58[20] 60[14])
    defparam mux_21_i23_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_22_i23_3_lut (.I0(n310[22]), .I1(IntegralLimit[22]), .I2(n258), 
            .I3(GND_net), .O(n337));   // verilog/motorControl.v(58[20] 60[14])
    defparam mux_22_i23_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_21_i20_3_lut (.I0(n233[19]), .I1(n285[19]), .I2(n284), 
            .I3(GND_net), .O(n310[19]));   // verilog/motorControl.v(58[20] 60[14])
    defparam mux_21_i20_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_4578_2 (.CI(GND_net), .I0(n29_adj_4256), .I1(n98), .CO(n46979));
    SB_LUT4 mux_22_i20_3_lut (.I0(n310[19]), .I1(IntegralLimit[19]), .I2(n258), 
            .I3(GND_net), .O(n340));   // verilog/motorControl.v(58[20] 60[14])
    defparam mux_22_i20_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_19_i31_2_lut (.I0(n233[15]), .I1(n285[15]), .I2(GND_net), 
            .I3(GND_net), .O(n31_adj_4266));   // verilog/motorControl.v(58[23:46])
    defparam LessThan_19_i31_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_19_i33_2_lut (.I0(n233[16]), .I1(n285[16]), .I2(GND_net), 
            .I3(GND_net), .O(n33_adj_4267));   // verilog/motorControl.v(58[23:46])
    defparam LessThan_19_i33_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_24_i365_2_lut (.I0(\Ki[7] ), .I1(n349), .I2(GND_net), 
            .I3(GND_net), .O(n542));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i365_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_21_i19_3_lut (.I0(n233[18]), .I1(n285[18]), .I2(n284), 
            .I3(GND_net), .O(n310[18]));   // verilog/motorControl.v(58[20] 60[14])
    defparam mux_21_i19_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_22_i19_3_lut (.I0(n310[18]), .I1(IntegralLimit[18]), .I2(n258), 
            .I3(GND_net), .O(n341));   // verilog/motorControl.v(58[20] 60[14])
    defparam mux_22_i19_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_23_i698_2_lut (.I0(\Kp[14] ), .I1(n207[9]), .I2(GND_net), 
            .I3(GND_net), .O(n1038));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i698_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_19_i29_2_lut (.I0(n233[14]), .I1(n285[14]), .I2(GND_net), 
            .I3(GND_net), .O(n29_adj_4268));   // verilog/motorControl.v(58[23:46])
    defparam LessThan_19_i29_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_4_lut_adj_929 (.I0(\Ki[1] ), .I1(\Ki[0] ), .I2(n337), .I3(n336), 
            .O(n56496));   // verilog/motorControl.v(61[29:40])
    defparam i1_4_lut_adj_929.LUT_INIT = 16'h93a0;
    SB_LUT4 i1_4_lut_adj_930 (.I0(\Ki[5] ), .I1(\Ki[4] ), .I2(n341), .I3(n340), 
            .O(n56500));   // verilog/motorControl.v(61[29:40])
    defparam i1_4_lut_adj_930.LUT_INIT = 16'h6ca0;
    SB_LUT4 i1_4_lut_adj_931 (.I0(\Ki[3] ), .I1(\Ki[2] ), .I2(n339), .I3(n338), 
            .O(n56498));   // verilog/motorControl.v(61[29:40])
    defparam i1_4_lut_adj_931.LUT_INIT = 16'h6ca0;
    SB_LUT4 n9440_bdd_4_lut_48718 (.I0(n9440), .I1(n59903), .I2(setpoint[17]), 
            .I3(n4357), .O(n63461));
    defparam n9440_bdd_4_lut_48718.LUT_INIT = 16'he4aa;
    SB_LUT4 LessThan_19_i27_2_lut (.I0(n233[13]), .I1(n285[13]), .I2(GND_net), 
            .I3(GND_net), .O(n27_adj_4269));   // verilog/motorControl.v(58[23:46])
    defparam LessThan_19_i27_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_4_lut_adj_932 (.I0(n56498), .I1(n45721), .I2(n56500), .I3(n56496), 
            .O(n56506));   // verilog/motorControl.v(61[29:40])
    defparam i1_4_lut_adj_932.LUT_INIT = 16'h6996;
    SB_LUT4 i32319_4_lut (.I0(n18055[0]), .I1(\Ki[2] ), .I2(n45772), .I3(n339), 
            .O(n4_adj_4270));   // verilog/motorControl.v(61[29:40])
    defparam i32319_4_lut.LUT_INIT = 16'he8a0;
    SB_LUT4 i45375_4_lut (.I0(n21_adj_4271), .I1(n19_adj_4272), .I2(n17_adj_4273), 
            .I3(n9_adj_4274), .O(n60087));
    defparam i45375_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i32436_4_lut (.I0(n17997[2]), .I1(\Ki[4] ), .I2(n6_adj_4257), 
            .I3(n341), .O(n8_adj_4275));   // verilog/motorControl.v(61[29:40])
    defparam i32436_4_lut.LUT_INIT = 16'he8a0;
    SB_LUT4 i1_4_lut_adj_933 (.I0(n6_adj_4276), .I1(n8_adj_4275), .I2(n4_adj_4270), 
            .I3(n56506), .O(n55441));   // verilog/motorControl.v(61[29:40])
    defparam i1_4_lut_adj_933.LUT_INIT = 16'h6996;
    SB_LUT4 i45339_4_lut (.I0(n27_adj_4269), .I1(n15_adj_4277), .I2(n13_adj_4278), 
            .I3(n11_adj_4279), .O(n60051));
    defparam i45339_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 LessThan_19_i12_3_lut (.I0(n285[7]), .I1(n285[16]), .I2(n33_adj_4267), 
            .I3(GND_net), .O(n12_adj_4280));   // verilog/motorControl.v(58[23:46])
    defparam LessThan_19_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_23_i67_2_lut (.I0(\Kp[1] ), .I1(n207[12]), .I2(GND_net), 
            .I3(GND_net), .O(n98));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i67_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i20_2_lut (.I0(\Kp[0] ), .I1(n207[13]), .I2(GND_net), 
            .I3(GND_net), .O(n29_adj_4256));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i20_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i116_2_lut (.I0(\Kp[2] ), .I1(n207[12]), .I2(GND_net), 
            .I3(GND_net), .O(n171));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i116_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i265_2_lut (.I0(\Kp[5] ), .I1(n207[13]), .I2(GND_net), 
            .I3(GND_net), .O(n393));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i265_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_4754_7_lut (.I0(GND_net), .I1(n55441), .I2(n490), .I3(n46978), 
            .O(n17859[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4754_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_19_i10_3_lut (.I0(n285[5]), .I1(n285[6]), .I2(n13_adj_4278), 
            .I3(GND_net), .O(n10_adj_4281));   // verilog/motorControl.v(58[23:46])
    defparam LessThan_19_i10_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_4754_6_lut (.I0(GND_net), .I1(n17940[3]), .I2(n417), .I3(n46977), 
            .O(n17859[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4754_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4754_6 (.CI(n46977), .I0(n17940[3]), .I1(n417), .CO(n46978));
    SB_LUT4 add_4754_5_lut (.I0(GND_net), .I1(n17940[2]), .I2(n344_adj_1), 
            .I3(n46976), .O(n17859[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4754_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4754_5 (.CI(n46976), .I0(n17940[2]), .I1(n344_adj_1), 
            .CO(n46977));
    SB_LUT4 add_4754_4_lut (.I0(GND_net), .I1(n17940[1]), .I2(n271), .I3(n46975), 
            .O(n17859[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4754_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_23_i314_2_lut (.I0(\Kp[6] ), .I1(n207[13]), .I2(GND_net), 
            .I3(GND_net), .O(n466));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i314_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_4754_4 (.CI(n46975), .I0(n17940[1]), .I1(n271), .CO(n46976));
    SB_LUT4 add_4754_3_lut (.I0(GND_net), .I1(n17940[0]), .I2(n198), .I3(n46974), 
            .O(n17859[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4754_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4754_3 (.CI(n46974), .I0(n17940[0]), .I1(n198), .CO(n46975));
    SB_LUT4 add_4754_2_lut (.I0(GND_net), .I1(n56), .I2(n125), .I3(GND_net), 
            .O(n17859[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4754_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 n9440_bdd_4_lut (.I0(n9440), .I1(n59930), .I2(setpoint[0]), 
            .I3(n4357), .O(n63677));
    defparam n9440_bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_LUT4 n63677_bdd_4_lut (.I0(n63677), .I1(n535[0]), .I2(n455[0]), 
            .I3(n4357), .O(n63680));
    defparam n63677_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_CARRY add_4754_2 (.CI(GND_net), .I0(n56), .I1(n125), .CO(n46974));
    SB_LUT4 add_4606_15_lut (.I0(GND_net), .I1(n16449[12]), .I2(n1050), 
            .I3(n46973), .O(n16059[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4606_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4606_14_lut (.I0(GND_net), .I1(n16449[11]), .I2(n977), 
            .I3(n46972), .O(n16059[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4606_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_23_i165_2_lut (.I0(\Kp[3] ), .I1(n207[12]), .I2(GND_net), 
            .I3(GND_net), .O(n244_adj_4255));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i165_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_4606_14 (.CI(n46972), .I0(n16449[11]), .I1(n977), .CO(n46973));
    SB_LUT4 add_4606_13_lut (.I0(GND_net), .I1(n16449[10]), .I2(n904), 
            .I3(n46971), .O(n16059[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4606_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4606_13 (.CI(n46971), .I0(n16449[10]), .I1(n904), .CO(n46972));
    SB_LUT4 add_4606_12_lut (.I0(GND_net), .I1(n16449[9]), .I2(n831), 
            .I3(n46970), .O(n16059[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4606_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4606_12 (.CI(n46970), .I0(n16449[9]), .I1(n831), .CO(n46971));
    SB_LUT4 add_4606_11_lut (.I0(GND_net), .I1(n16449[8]), .I2(n758), 
            .I3(n46969), .O(n16059[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4606_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 n63461_bdd_4_lut (.I0(n63461), .I1(n535[17]), .I2(n455[17]), 
            .I3(n4357), .O(n63464));
    defparam n63461_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n9440_bdd_4_lut_48713 (.I0(n9440), .I1(n59902), .I2(setpoint[16]), 
            .I3(n4357), .O(n63455));
    defparam n9440_bdd_4_lut_48713.LUT_INIT = 16'he4aa;
    SB_LUT4 n63455_bdd_4_lut (.I0(n63455), .I1(n535[16]), .I2(n455[16]), 
            .I3(n4357), .O(n63458));
    defparam n63455_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 mult_23_i214_2_lut (.I0(\Kp[4] ), .I1(n207[12]), .I2(GND_net), 
            .I3(GND_net), .O(n317));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i214_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_4606_11 (.CI(n46969), .I0(n16449[8]), .I1(n758), .CO(n46970));
    SB_LUT4 mult_23_i263_2_lut (.I0(\Kp[5] ), .I1(n207[12]), .I2(GND_net), 
            .I3(GND_net), .O(n390));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i263_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_4606_10_lut (.I0(GND_net), .I1(n16449[7]), .I2(n685), 
            .I3(n46968), .O(n16059[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4606_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4606_10 (.CI(n46968), .I0(n16449[7]), .I1(n685), .CO(n46969));
    SB_LUT4 add_4606_9_lut (.I0(GND_net), .I1(n16449[6]), .I2(n612), .I3(n46967), 
            .O(n16059[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4606_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 counter_1940_1941_add_4_15_lut (.I0(GND_net), .I1(GND_net), 
            .I2(counter[13]), .I3(n46625), .O(n61[13])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_1940_1941_add_4_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 n9440_bdd_4_lut_48708 (.I0(n9440), .I1(n59901), .I2(setpoint[15]), 
            .I3(n4357), .O(n63449));
    defparam n9440_bdd_4_lut_48708.LUT_INIT = 16'he4aa;
    SB_LUT4 counter_1940_1941_add_4_14_lut (.I0(GND_net), .I1(GND_net), 
            .I2(counter[12]), .I3(n46624), .O(n61[12])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_1940_1941_add_4_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4606_9 (.CI(n46967), .I0(n16449[6]), .I1(n612), .CO(n46968));
    SB_CARRY counter_1940_1941_add_4_14 (.CI(n46624), .I0(GND_net), .I1(counter[12]), 
            .CO(n46625));
    SB_LUT4 counter_1940_1941_add_4_13_lut (.I0(GND_net), .I1(GND_net), 
            .I2(counter[11]), .I3(n46623), .O(n61[11])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_1940_1941_add_4_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_1940_1941_add_4_13 (.CI(n46623), .I0(GND_net), .I1(counter[11]), 
            .CO(n46624));
    SB_LUT4 add_4606_8_lut (.I0(GND_net), .I1(n16449[5]), .I2(n539_adj_4285), 
            .I3(n46966), .O(n16059[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4606_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4606_8 (.CI(n46966), .I0(n16449[5]), .I1(n539_adj_4285), 
            .CO(n46967));
    SB_LUT4 LessThan_19_i30_3_lut (.I0(n12_adj_4280), .I1(n292), .I2(n35), 
            .I3(GND_net), .O(n30_adj_4287));   // verilog/motorControl.v(58[23:46])
    defparam LessThan_19_i30_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 counter_1940_1941_add_4_12_lut (.I0(GND_net), .I1(GND_net), 
            .I2(counter[10]), .I3(n46622), .O(n61[10])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_1940_1941_add_4_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_23_i312_2_lut (.I0(\Kp[6] ), .I1(n207[12]), .I2(GND_net), 
            .I3(GND_net), .O(n463));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i312_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_4606_7_lut (.I0(GND_net), .I1(n16449[4]), .I2(n466), .I3(n46965), 
            .O(n16059[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4606_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4606_7 (.CI(n46965), .I0(n16449[4]), .I1(n466), .CO(n46966));
    SB_CARRY counter_1940_1941_add_4_12 (.CI(n46622), .I0(GND_net), .I1(counter[10]), 
            .CO(n46623));
    SB_LUT4 add_4606_6_lut (.I0(GND_net), .I1(n16449[3]), .I2(n393), .I3(n46964), 
            .O(n16059[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4606_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 counter_1940_1941_add_4_11_lut (.I0(GND_net), .I1(GND_net), 
            .I2(counter[9]), .I3(n46621), .O(n61[9])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_1940_1941_add_4_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4606_6 (.CI(n46964), .I0(n16449[3]), .I1(n393), .CO(n46965));
    SB_LUT4 n63449_bdd_4_lut (.I0(n63449), .I1(n535[15]), .I2(n455[15]), 
            .I3(n4357), .O(n63452));
    defparam n63449_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 add_4606_5_lut (.I0(GND_net), .I1(n16449[2]), .I2(n320), .I3(n46963), 
            .O(n16059[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4606_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_1940_1941_add_4_11 (.CI(n46621), .I0(GND_net), .I1(counter[9]), 
            .CO(n46622));
    SB_LUT4 counter_1940_1941_add_4_10_lut (.I0(GND_net), .I1(GND_net), 
            .I2(counter[8]), .I3(n46620), .O(n61[8])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_1940_1941_add_4_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_1940_1941_add_4_10 (.CI(n46620), .I0(GND_net), .I1(counter[8]), 
            .CO(n46621));
    SB_CARRY add_4606_5 (.CI(n46963), .I0(n16449[2]), .I1(n320), .CO(n46964));
    SB_LUT4 add_4606_4_lut (.I0(GND_net), .I1(n16449[1]), .I2(n247_adj_4224), 
            .I3(n46962), .O(n16059[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4606_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 counter_1940_1941_add_4_9_lut (.I0(GND_net), .I1(GND_net), .I2(counter[7]), 
            .I3(n46619), .O(n61[7])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_1940_1941_add_4_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_1940_1941_add_4_9 (.CI(n46619), .I0(GND_net), .I1(counter[7]), 
            .CO(n46620));
    SB_LUT4 counter_1940_1941_add_4_8_lut (.I0(GND_net), .I1(GND_net), .I2(counter[6]), 
            .I3(n46618), .O(n61[6])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_1940_1941_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4606_4 (.CI(n46962), .I0(n16449[1]), .I1(n247_adj_4224), 
            .CO(n46963));
    SB_LUT4 add_4606_3_lut (.I0(GND_net), .I1(n16449[0]), .I2(n174), .I3(n46961), 
            .O(n16059[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4606_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_23_i361_2_lut (.I0(\Kp[7] ), .I1(n207[12]), .I2(GND_net), 
            .I3(GND_net), .O(n536));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i361_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY counter_1940_1941_add_4_8 (.CI(n46618), .I0(GND_net), .I1(counter[6]), 
            .CO(n46619));
    SB_LUT4 counter_1940_1941_add_4_7_lut (.I0(GND_net), .I1(GND_net), .I2(counter[5]), 
            .I3(n46617), .O(n61[5])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_1940_1941_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_1940_1941_add_4_7 (.CI(n46617), .I0(GND_net), .I1(counter[5]), 
            .CO(n46618));
    SB_CARRY add_4606_3 (.CI(n46961), .I0(n16449[0]), .I1(n174), .CO(n46962));
    SB_LUT4 counter_1940_1941_add_4_6_lut (.I0(GND_net), .I1(GND_net), .I2(counter[4]), 
            .I3(n46616), .O(n61[4])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_1940_1941_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_23_i410_2_lut (.I0(\Kp[8] ), .I1(n207[12]), .I2(GND_net), 
            .I3(GND_net), .O(n609));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i410_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_4606_2_lut (.I0(GND_net), .I1(n32), .I2(n101), .I3(GND_net), 
            .O(n16059[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4606_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i46364_4_lut (.I0(n13_adj_4278), .I1(n11_adj_4279), .I2(n9_adj_4274), 
            .I3(n60168), .O(n61076));
    defparam i46364_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 n9440_bdd_4_lut_48703 (.I0(n9440), .I1(n59900), .I2(setpoint[14]), 
            .I3(n4357), .O(n63443));
    defparam n9440_bdd_4_lut_48703.LUT_INIT = 16'he4aa;
    SB_LUT4 i46344_4_lut (.I0(n19_adj_4272), .I1(n17_adj_4273), .I2(n15_adj_4277), 
            .I3(n61076), .O(n61056));
    defparam i46344_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 n63443_bdd_4_lut (.I0(n63443), .I1(n535[14]), .I2(n455[14]), 
            .I3(n4357), .O(n63446));
    defparam n63443_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 mult_23_i459_2_lut (.I0(\Kp[9] ), .I1(n207[12]), .I2(GND_net), 
            .I3(GND_net), .O(n682));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i459_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY counter_1940_1941_add_4_6 (.CI(n46616), .I0(GND_net), .I1(counter[4]), 
            .CO(n46617));
    SB_LUT4 i47816_4_lut (.I0(n25_adj_4289), .I1(n23_adj_4290), .I2(n21_adj_4271), 
            .I3(n61056), .O(n62529));
    defparam i47816_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 n9440_bdd_4_lut_48698 (.I0(n9440), .I1(n59899), .I2(setpoint[13]), 
            .I3(n4357), .O(n63437));
    defparam n9440_bdd_4_lut_48698.LUT_INIT = 16'he4aa;
    SB_CARRY add_4606_2 (.CI(GND_net), .I0(n32), .I1(n101), .CO(n46961));
    SB_LUT4 add_4632_14_lut (.I0(GND_net), .I1(n16785[11]), .I2(n980), 
            .I3(n46960), .O(n16449[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4632_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 counter_1940_1941_add_4_5_lut (.I0(GND_net), .I1(GND_net), .I2(counter[3]), 
            .I3(n46615), .O(n61[3])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_1940_1941_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 n63437_bdd_4_lut (.I0(n63437), .I1(n535[13]), .I2(n455[13]), 
            .I3(n4357), .O(n63440));
    defparam n63437_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i47120_4_lut (.I0(n31_adj_4266), .I1(n29_adj_4268), .I2(n27_adj_4269), 
            .I3(n62529), .O(n61833));
    defparam i47120_4_lut.LUT_INIT = 16'hfeff;
    SB_CARRY counter_1940_1941_add_4_5 (.CI(n46615), .I0(GND_net), .I1(counter[3]), 
            .CO(n46616));
    SB_LUT4 i48024_4_lut (.I0(n37_adj_4264), .I1(n35), .I2(n33_adj_4267), 
            .I3(n61833), .O(n62737));
    defparam i48024_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 add_4632_13_lut (.I0(GND_net), .I1(n16785[10]), .I2(n907), 
            .I3(n46959), .O(n16449[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4632_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4632_13 (.CI(n46959), .I0(n16785[10]), .I1(n907), .CO(n46960));
    SB_LUT4 add_4632_12_lut (.I0(GND_net), .I1(n16785[9]), .I2(n834_adj_4292), 
            .I3(n46958), .O(n16449[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4632_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4632_12 (.CI(n46958), .I0(n16785[9]), .I1(n834_adj_4292), 
            .CO(n46959));
    SB_LUT4 add_4632_11_lut (.I0(GND_net), .I1(n16785[8]), .I2(n761_adj_4293), 
            .I3(n46957), .O(n16449[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4632_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 counter_1940_1941_add_4_4_lut (.I0(GND_net), .I1(GND_net), .I2(counter[2]), 
            .I3(n46614), .O(n61[2])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_1940_1941_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_1940_1941_add_4_4 (.CI(n46614), .I0(GND_net), .I1(counter[2]), 
            .CO(n46615));
    SB_CARRY add_4632_11 (.CI(n46957), .I0(n16785[8]), .I1(n761_adj_4293), 
            .CO(n46958));
    SB_LUT4 add_4632_10_lut (.I0(GND_net), .I1(n16785[7]), .I2(n688_adj_4294), 
            .I3(n46956), .O(n16449[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4632_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4632_10 (.CI(n46956), .I0(n16785[7]), .I1(n688_adj_4294), 
            .CO(n46957));
    SB_LUT4 counter_1940_1941_add_4_3_lut (.I0(GND_net), .I1(GND_net), .I2(counter[1]), 
            .I3(n46613), .O(n61[1])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_1940_1941_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 n9440_bdd_4_lut_48693 (.I0(n9440), .I1(n59898), .I2(setpoint[12]), 
            .I3(n4357), .O(n63431));
    defparam n9440_bdd_4_lut_48693.LUT_INIT = 16'he4aa;
    SB_LUT4 add_4632_9_lut (.I0(GND_net), .I1(n16785[6]), .I2(n615_adj_4295), 
            .I3(n46955), .O(n16449[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4632_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 n63431_bdd_4_lut (.I0(n63431), .I1(n535[12]), .I2(n455[12]), 
            .I3(n4357), .O(n63434));
    defparam n63431_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_CARRY add_4632_9 (.CI(n46955), .I0(n16785[6]), .I1(n615_adj_4295), 
            .CO(n46956));
    SB_LUT4 add_4632_8_lut (.I0(GND_net), .I1(n16785[5]), .I2(n542_adj_4296), 
            .I3(n46954), .O(n16449[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4632_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_19_i16_3_lut (.I0(n285[9]), .I1(n285[21]), .I2(n43_adj_4260), 
            .I3(GND_net), .O(n16_adj_4297));   // verilog/motorControl.v(58[23:46])
    defparam LessThan_19_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY counter_1940_1941_add_4_3 (.CI(n46613), .I0(GND_net), .I1(counter[1]), 
            .CO(n46614));
    SB_LUT4 counter_1940_1941_add_4_2_lut (.I0(GND_net), .I1(GND_net), .I2(counter[0]), 
            .I3(VCC_net), .O(n61[0])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_1940_1941_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_1940_1941_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(counter[0]), 
            .CO(n46613));
    SB_LUT4 n9440_bdd_4_lut_48688 (.I0(n9440), .I1(n59897), .I2(setpoint[11]), 
            .I3(n4357), .O(n63425));
    defparam n9440_bdd_4_lut_48688.LUT_INIT = 16'he4aa;
    SB_CARRY add_4632_8 (.CI(n46954), .I0(n16785[5]), .I1(n542_adj_4296), 
            .CO(n46955));
    SB_LUT4 add_4632_7_lut (.I0(GND_net), .I1(n16785[4]), .I2(n469_adj_4298), 
            .I3(n46953), .O(n16449[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4632_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4632_7 (.CI(n46953), .I0(n16785[4]), .I1(n469_adj_4298), 
            .CO(n46954));
    SB_LUT4 n63425_bdd_4_lut (.I0(n63425), .I1(n535[11]), .I2(n455[11]), 
            .I3(n4357), .O(n63428));
    defparam n63425_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 mult_23_i508_2_lut (.I0(\Kp[10] ), .I1(n207[12]), .I2(GND_net), 
            .I3(GND_net), .O(n755));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i508_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_4632_6_lut (.I0(GND_net), .I1(n16785[3]), .I2(n396_adj_4300), 
            .I3(n46952), .O(n16449[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4632_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_23_i363_2_lut (.I0(\Kp[7] ), .I1(n207[13]), .I2(GND_net), 
            .I3(GND_net), .O(n539_adj_4285));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i363_2_lut.LUT_INIT = 16'h8888;
    SB_DFFR \PID_CONTROLLER.integral_i0_i1  (.Q(\PID_CONTROLLER.integral [1]), 
            .C(clk16MHz), .D(n26870), .R(reset));   // verilog/motorControl.v(42[14] 73[8])
    SB_DFFR \PID_CONTROLLER.integral_i0_i2  (.Q(\PID_CONTROLLER.integral [2]), 
            .C(clk16MHz), .D(n26869), .R(reset));   // verilog/motorControl.v(42[14] 73[8])
    SB_DFFR \PID_CONTROLLER.integral_i0_i3  (.Q(\PID_CONTROLLER.integral [3]), 
            .C(clk16MHz), .D(n26868), .R(reset));   // verilog/motorControl.v(42[14] 73[8])
    SB_DFFR \PID_CONTROLLER.integral_i0_i4  (.Q(\PID_CONTROLLER.integral [4]), 
            .C(clk16MHz), .D(n26867), .R(reset));   // verilog/motorControl.v(42[14] 73[8])
    SB_DFFR \PID_CONTROLLER.integral_i0_i5  (.Q(\PID_CONTROLLER.integral [5]), 
            .C(clk16MHz), .D(n26866), .R(reset));   // verilog/motorControl.v(42[14] 73[8])
    SB_DFFR \PID_CONTROLLER.integral_i0_i6  (.Q(\PID_CONTROLLER.integral [6]), 
            .C(clk16MHz), .D(n26865), .R(reset));   // verilog/motorControl.v(42[14] 73[8])
    SB_DFFR \PID_CONTROLLER.integral_i0_i7  (.Q(\PID_CONTROLLER.integral [7]), 
            .C(clk16MHz), .D(n26864), .R(reset));   // verilog/motorControl.v(42[14] 73[8])
    SB_DFFR \PID_CONTROLLER.integral_i0_i8  (.Q(\PID_CONTROLLER.integral [8]), 
            .C(clk16MHz), .D(n26863), .R(reset));   // verilog/motorControl.v(42[14] 73[8])
    SB_DFFR \PID_CONTROLLER.integral_i0_i9  (.Q(\PID_CONTROLLER.integral [9]), 
            .C(clk16MHz), .D(n26862), .R(reset));   // verilog/motorControl.v(42[14] 73[8])
    SB_DFFR \PID_CONTROLLER.integral_i0_i10  (.Q(\PID_CONTROLLER.integral [10]), 
            .C(clk16MHz), .D(n26861), .R(reset));   // verilog/motorControl.v(42[14] 73[8])
    SB_DFFR \PID_CONTROLLER.integral_i0_i11  (.Q(\PID_CONTROLLER.integral [11]), 
            .C(clk16MHz), .D(n26860), .R(reset));   // verilog/motorControl.v(42[14] 73[8])
    SB_DFFR \PID_CONTROLLER.integral_i0_i12  (.Q(\PID_CONTROLLER.integral [12]), 
            .C(clk16MHz), .D(n26859), .R(reset));   // verilog/motorControl.v(42[14] 73[8])
    SB_LUT4 i47736_3_lut (.I0(n6_adj_4301), .I1(n285[10]), .I2(n21_adj_4271), 
            .I3(GND_net), .O(n62449));   // verilog/motorControl.v(58[23:46])
    defparam i47736_3_lut.LUT_INIT = 16'hcaca;
    SB_DFFR \PID_CONTROLLER.integral_i0_i13  (.Q(\PID_CONTROLLER.integral [13]), 
            .C(clk16MHz), .D(n26858), .R(reset));   // verilog/motorControl.v(42[14] 73[8])
    SB_DFFR \PID_CONTROLLER.integral_i0_i14  (.Q(\PID_CONTROLLER.integral [14]), 
            .C(clk16MHz), .D(n26857), .R(reset));   // verilog/motorControl.v(42[14] 73[8])
    SB_DFFR \PID_CONTROLLER.integral_i0_i15  (.Q(\PID_CONTROLLER.integral [15]), 
            .C(clk16MHz), .D(n26856), .R(reset));   // verilog/motorControl.v(42[14] 73[8])
    SB_DFFR \PID_CONTROLLER.integral_i0_i16  (.Q(\PID_CONTROLLER.integral [16]), 
            .C(clk16MHz), .D(n26855), .R(reset));   // verilog/motorControl.v(42[14] 73[8])
    SB_DFFR \PID_CONTROLLER.integral_i0_i17  (.Q(\PID_CONTROLLER.integral [17]), 
            .C(clk16MHz), .D(n26854), .R(reset));   // verilog/motorControl.v(42[14] 73[8])
    SB_DFFR \PID_CONTROLLER.integral_i0_i18  (.Q(\PID_CONTROLLER.integral [18]), 
            .C(clk16MHz), .D(n26853), .R(reset));   // verilog/motorControl.v(42[14] 73[8])
    SB_DFFR \PID_CONTROLLER.integral_i0_i19  (.Q(\PID_CONTROLLER.integral [19]), 
            .C(clk16MHz), .D(n26852), .R(reset));   // verilog/motorControl.v(42[14] 73[8])
    SB_DFFR \PID_CONTROLLER.integral_i0_i20  (.Q(\PID_CONTROLLER.integral [20]), 
            .C(clk16MHz), .D(n26851), .R(reset));   // verilog/motorControl.v(42[14] 73[8])
    SB_DFFR \PID_CONTROLLER.integral_i0_i21  (.Q(\PID_CONTROLLER.integral [21]), 
            .C(clk16MHz), .D(n26850), .R(reset));   // verilog/motorControl.v(42[14] 73[8])
    SB_DFFR \PID_CONTROLLER.integral_i0_i22  (.Q(\PID_CONTROLLER.integral [22]), 
            .C(clk16MHz), .D(n26849), .R(reset));   // verilog/motorControl.v(42[14] 73[8])
    SB_LUT4 i47737_3_lut (.I0(n62449), .I1(n285[11]), .I2(n23_adj_4290), 
            .I3(GND_net), .O(n62450));   // verilog/motorControl.v(58[23:46])
    defparam i47737_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_4632_6 (.CI(n46952), .I0(n16785[3]), .I1(n396_adj_4300), 
            .CO(n46953));
    SB_LUT4 mult_23_i412_2_lut (.I0(\Kp[8] ), .I1(n207[13]), .I2(GND_net), 
            .I3(GND_net), .O(n612));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i412_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i461_2_lut (.I0(\Kp[9] ), .I1(n207[13]), .I2(GND_net), 
            .I3(GND_net), .O(n685));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i461_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_4632_5_lut (.I0(GND_net), .I1(n16785[2]), .I2(n323_adj_4302), 
            .I3(n46951), .O(n16449[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4632_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 n9440_bdd_4_lut_48683 (.I0(n9440), .I1(n59896), .I2(setpoint[10]), 
            .I3(n4357), .O(n63419));
    defparam n9440_bdd_4_lut_48683.LUT_INIT = 16'he4aa;
    SB_LUT4 n63419_bdd_4_lut (.I0(n63419), .I1(n535[10]), .I2(n455[10]), 
            .I3(n4357), .O(n63422));
    defparam n63419_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 mult_23_i510_2_lut (.I0(\Kp[10] ), .I1(n207[13]), .I2(GND_net), 
            .I3(GND_net), .O(n758));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i510_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_4632_5 (.CI(n46951), .I0(n16785[2]), .I1(n323_adj_4302), 
            .CO(n46952));
    SB_LUT4 mult_23_i559_2_lut (.I0(\Kp[11] ), .I1(n207[13]), .I2(GND_net), 
            .I3(GND_net), .O(n831));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i559_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i608_2_lut (.I0(\Kp[12] ), .I1(n207[13]), .I2(GND_net), 
            .I3(GND_net), .O(n904));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i608_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_19_i8_3_lut (.I0(n285[4]), .I1(n285[8]), .I2(n17_adj_4273), 
            .I3(GND_net), .O(n8_adj_4304));   // verilog/motorControl.v(58[23:46])
    defparam LessThan_19_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_4632_4_lut (.I0(GND_net), .I1(n16785[1]), .I2(n250_adj_4305), 
            .I3(n46950), .O(n16449[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4632_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_23_i557_2_lut (.I0(\Kp[11] ), .I1(n207[12]), .I2(GND_net), 
            .I3(GND_net), .O(n828));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i557_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_19_i24_3_lut (.I0(n16_adj_4297), .I1(n285[22]), .I2(n45_adj_4258), 
            .I3(GND_net), .O(n24_adj_4306));   // verilog/motorControl.v(58[23:46])
    defparam LessThan_19_i24_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_23_i606_2_lut (.I0(\Kp[12] ), .I1(n207[12]), .I2(GND_net), 
            .I3(GND_net), .O(n901));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i606_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i45271_4_lut (.I0(n43_adj_4260), .I1(n25_adj_4289), .I2(n23_adj_4290), 
            .I3(n60087), .O(n59983));
    defparam i45271_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 mult_23_i655_2_lut (.I0(\Kp[13] ), .I1(n207[12]), .I2(GND_net), 
            .I3(GND_net), .O(n974));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i655_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i704_2_lut (.I0(\Kp[14] ), .I1(n207[12]), .I2(GND_net), 
            .I3(GND_net), .O(n1047));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i704_2_lut.LUT_INIT = 16'h8888;
    SB_DFFR \PID_CONTROLLER.integral_i0_i23  (.Q(\PID_CONTROLLER.integral [23]), 
            .C(clk16MHz), .D(n26780), .R(reset));   // verilog/motorControl.v(42[14] 73[8])
    SB_CARRY add_4632_4 (.CI(n46950), .I0(n16785[1]), .I1(n250_adj_4305), 
            .CO(n46951));
    SB_LUT4 add_4632_3_lut (.I0(GND_net), .I1(n16785[0]), .I2(n177_adj_4307), 
            .I3(n46949), .O(n16449[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4632_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_23_i657_2_lut (.I0(\Kp[13] ), .I1(n207[13]), .I2(GND_net), 
            .I3(GND_net), .O(n977));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i657_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i706_2_lut (.I0(\Kp[14] ), .I1(n207[13]), .I2(GND_net), 
            .I3(GND_net), .O(n1050));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i706_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i47166_4_lut (.I0(n24_adj_4306), .I1(n8_adj_4304), .I2(n45_adj_4258), 
            .I3(n59981), .O(n61879));   // verilog/motorControl.v(58[23:46])
    defparam i47166_4_lut.LUT_INIT = 16'haaac;
    SB_CARRY add_4632_3 (.CI(n46949), .I0(n16785[0]), .I1(n177_adj_4307), 
            .CO(n46950));
    SB_LUT4 mult_23_i753_2_lut (.I0(\Kp[15] ), .I1(n207[12]), .I2(GND_net), 
            .I3(GND_net), .O(n1120));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i753_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_4632_2_lut (.I0(GND_net), .I1(n35_adj_4308), .I2(n104_adj_4309), 
            .I3(GND_net), .O(n16449[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4632_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_23_i65_2_lut (.I0(\Kp[1] ), .I1(n207[11]), .I2(GND_net), 
            .I3(GND_net), .O(n95));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i65_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i47520_3_lut (.I0(n62450), .I1(n285[12]), .I2(n25_adj_4289), 
            .I3(GND_net), .O(n62233));   // verilog/motorControl.v(58[23:46])
    defparam i47520_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_23_i18_2_lut (.I0(\Kp[0] ), .I1(n207[12]), .I2(GND_net), 
            .I3(GND_net), .O(n26));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i18_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i114_2_lut (.I0(\Kp[2] ), .I1(n207[11]), .I2(GND_net), 
            .I3(GND_net), .O(n168));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i114_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i163_2_lut (.I0(\Kp[3] ), .I1(n207[11]), .I2(GND_net), 
            .I3(GND_net), .O(n241_adj_4253));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i163_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i212_2_lut (.I0(\Kp[4] ), .I1(n207[11]), .I2(GND_net), 
            .I3(GND_net), .O(n314));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i212_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i261_2_lut (.I0(\Kp[5] ), .I1(n207[11]), .I2(GND_net), 
            .I3(GND_net), .O(n387));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i261_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 n9440_bdd_4_lut_48678 (.I0(n9440), .I1(n59886), .I2(setpoint[9]), 
            .I3(n4357), .O(n63407));
    defparam n9440_bdd_4_lut_48678.LUT_INIT = 16'he4aa;
    SB_LUT4 n63407_bdd_4_lut (.I0(n63407), .I1(n535[9]), .I2(n455[9]), 
            .I3(n4357), .O(n63410));
    defparam n63407_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n9440_bdd_4_lut_48668 (.I0(n9440), .I1(n59885), .I2(setpoint[8]), 
            .I3(n4357), .O(n63401));
    defparam n9440_bdd_4_lut_48668.LUT_INIT = 16'he4aa;
    SB_LUT4 mult_23_i310_2_lut (.I0(\Kp[6] ), .I1(n207[11]), .I2(GND_net), 
            .I3(GND_net), .O(n460_adj_4249));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i310_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_4632_2 (.CI(GND_net), .I0(n35_adj_4308), .I1(n104_adj_4309), 
            .CO(n46949));
    SB_LUT4 add_4656_13_lut (.I0(GND_net), .I1(n17071[10]), .I2(n910_adj_4310), 
            .I3(n46948), .O(n16785[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4656_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_23_i359_2_lut (.I0(\Kp[7] ), .I1(n207[11]), .I2(GND_net), 
            .I3(GND_net), .O(n533));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i359_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_4656_12_lut (.I0(GND_net), .I1(n17071[9]), .I2(n837_adj_4311), 
            .I3(n46947), .O(n16785[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4656_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4656_12 (.CI(n46947), .I0(n17071[9]), .I1(n837_adj_4311), 
            .CO(n46948));
    SB_LUT4 add_4656_11_lut (.I0(GND_net), .I1(n17071[8]), .I2(n764_adj_4312), 
            .I3(n46946), .O(n16785[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4656_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4656_11 (.CI(n46946), .I0(n17071[8]), .I1(n764_adj_4312), 
            .CO(n46947));
    SB_LUT4 LessThan_19_i4_4_lut (.I0(n233[0]), .I1(n285[1]), .I2(n233[1]), 
            .I3(n285[0]), .O(n4_adj_4313));   // verilog/motorControl.v(58[23:46])
    defparam LessThan_19_i4_4_lut.LUT_INIT = 16'h4d0c;
    SB_LUT4 add_4656_10_lut (.I0(GND_net), .I1(n17071[7]), .I2(n691_adj_4314), 
            .I3(n46945), .O(n16785[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4656_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i47734_3_lut (.I0(n4_adj_4313), .I1(n285[13]), .I2(n27_adj_4269), 
            .I3(GND_net), .O(n62447));   // verilog/motorControl.v(58[23:46])
    defparam i47734_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 n63401_bdd_4_lut (.I0(n63401), .I1(n535[8]), .I2(n455[8]), 
            .I3(n4357), .O(n63404));
    defparam n63401_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFFSR counter_1940_1941__i1 (.Q(counter[0]), .C(clk16MHz), .D(n61[0]), 
            .R(counter_31__N_3487));   // verilog/motorControl.v(25[16:25])
    SB_LUT4 i47735_3_lut (.I0(n62447), .I1(n285[14]), .I2(n29_adj_4268), 
            .I3(GND_net), .O(n62448));   // verilog/motorControl.v(58[23:46])
    defparam i47735_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_4656_10 (.CI(n46945), .I0(n17071[7]), .I1(n691_adj_4314), 
            .CO(n46946));
    SB_LUT4 add_4656_9_lut (.I0(GND_net), .I1(n17071[6]), .I2(n618_adj_4315), 
            .I3(n46944), .O(n16785[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4656_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4656_9 (.CI(n46944), .I0(n17071[6]), .I1(n618_adj_4315), 
            .CO(n46945));
    SB_LUT4 n9440_bdd_4_lut_48663 (.I0(n9440), .I1(n59884), .I2(setpoint[7]), 
            .I3(n4357), .O(n63395));
    defparam n9440_bdd_4_lut_48663.LUT_INIT = 16'he4aa;
    SB_LUT4 mult_23_i408_2_lut (.I0(\Kp[8] ), .I1(n207[11]), .I2(GND_net), 
            .I3(GND_net), .O(n606));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i408_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_4656_8_lut (.I0(GND_net), .I1(n17071[5]), .I2(n545_adj_4316), 
            .I3(n46943), .O(n16785[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4656_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4656_8 (.CI(n46943), .I0(n17071[5]), .I1(n545_adj_4316), 
            .CO(n46944));
    SB_LUT4 add_4656_7_lut (.I0(GND_net), .I1(n17071[4]), .I2(n472_adj_4317), 
            .I3(n46942), .O(n16785[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4656_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4656_7 (.CI(n46942), .I0(n17071[4]), .I1(n472_adj_4317), 
            .CO(n46943));
    SB_LUT4 n63395_bdd_4_lut (.I0(n63395), .I1(n535[7]), .I2(n455[7]), 
            .I3(n4357), .O(n63398));
    defparam n63395_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 add_4656_6_lut (.I0(GND_net), .I1(n17071[3]), .I2(n399_adj_4319), 
            .I3(n46941), .O(n16785[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4656_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4656_6 (.CI(n46941), .I0(n17071[3]), .I1(n399_adj_4319), 
            .CO(n46942));
    SB_LUT4 add_4656_5_lut (.I0(GND_net), .I1(n17071[2]), .I2(n326_adj_4320), 
            .I3(n46940), .O(n16785[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4656_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4656_5 (.CI(n46940), .I0(n17071[2]), .I1(n326_adj_4320), 
            .CO(n46941));
    SB_LUT4 add_4656_4_lut (.I0(GND_net), .I1(n17071[1]), .I2(n253_adj_4321), 
            .I3(n46939), .O(n16785[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4656_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4656_4 (.CI(n46939), .I0(n17071[1]), .I1(n253_adj_4321), 
            .CO(n46940));
    SB_LUT4 add_4656_3_lut (.I0(GND_net), .I1(n17071[0]), .I2(n180_adj_4322), 
            .I3(n46938), .O(n16785[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4656_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4656_3 (.CI(n46938), .I0(n17071[0]), .I1(n180_adj_4322), 
            .CO(n46939));
    SB_LUT4 add_4656_2_lut (.I0(GND_net), .I1(n38_adj_4323), .I2(n107_adj_4324), 
            .I3(GND_net), .O(n16785[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4656_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4656_2 (.CI(GND_net), .I0(n38_adj_4323), .I1(n107_adj_4324), 
            .CO(n46938));
    SB_LUT4 mult_24_add_1225_24_lut (.I0(n336), .I1(n10031[21]), .I2(GND_net), 
            .I3(n46937), .O(n9524[0])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_24_add_1225_24_lut.LUT_INIT = 16'h6996;
    SB_LUT4 mult_24_add_1225_23_lut (.I0(GND_net), .I1(n10031[20]), .I2(GND_net), 
            .I3(n46936), .O(n42[22])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_24_add_1225_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i45307_4_lut (.I0(n33_adj_4267), .I1(n31_adj_4266), .I2(n29_adj_4268), 
            .I3(n60051), .O(n60019));
    defparam i45307_4_lut.LUT_INIT = 16'haaab;
    SB_CARRY mult_24_add_1225_23 (.CI(n46936), .I0(n10031[20]), .I1(GND_net), 
            .CO(n46937));
    SB_LUT4 mult_24_add_1225_22_lut (.I0(GND_net), .I1(n10031[19]), .I2(GND_net), 
            .I3(n46935), .O(n42[21])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_24_add_1225_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_23_i457_2_lut (.I0(\Kp[9] ), .I1(n207[11]), .I2(GND_net), 
            .I3(GND_net), .O(n679));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i457_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY mult_24_add_1225_22 (.CI(n46935), .I0(n10031[19]), .I1(GND_net), 
            .CO(n46936));
    SB_LUT4 mult_24_add_1225_21_lut (.I0(GND_net), .I1(n10031[18]), .I2(GND_net), 
            .I3(n46934), .O(n42[20])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_24_add_1225_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_24_add_1225_21 (.CI(n46934), .I0(n10031[18]), .I1(GND_net), 
            .CO(n46935));
    SB_LUT4 mult_24_add_1225_20_lut (.I0(GND_net), .I1(n10031[17]), .I2(GND_net), 
            .I3(n46933), .O(n42[19])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_24_add_1225_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_24_add_1225_20 (.CI(n46933), .I0(n10031[17]), .I1(GND_net), 
            .CO(n46934));
    SB_LUT4 i48062_4_lut (.I0(n30_adj_4287), .I1(n10_adj_4281), .I2(n35), 
            .I3(n60010), .O(n62775));   // verilog/motorControl.v(58[23:46])
    defparam i48062_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 mult_24_add_1225_19_lut (.I0(GND_net), .I1(n10031[16]), .I2(GND_net), 
            .I3(n46932), .O(n42[18])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_24_add_1225_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_24_add_1225_19 (.CI(n46932), .I0(n10031[16]), .I1(GND_net), 
            .CO(n46933));
    SB_LUT4 mult_24_add_1225_18_lut (.I0(GND_net), .I1(n10031[15]), .I2(GND_net), 
            .I3(n46931), .O(n42[17])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_24_add_1225_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_24_add_1225_18 (.CI(n46931), .I0(n10031[15]), .I1(GND_net), 
            .CO(n46932));
    SB_LUT4 mult_24_add_1225_17_lut (.I0(GND_net), .I1(n10031[14]), .I2(GND_net), 
            .I3(n46930), .O(n42[16])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_24_add_1225_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_24_add_1225_17 (.CI(n46930), .I0(n10031[14]), .I1(GND_net), 
            .CO(n46931));
    SB_LUT4 mult_24_add_1225_16_lut (.I0(GND_net), .I1(n10031[13]), .I2(n1096), 
            .I3(n46929), .O(n42[15])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_24_add_1225_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_24_add_1225_16 (.CI(n46929), .I0(n10031[13]), .I1(n1096), 
            .CO(n46930));
    SB_LUT4 mult_24_add_1225_15_lut (.I0(GND_net), .I1(n10031[12]), .I2(n1023), 
            .I3(n46928), .O(n42[14])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_24_add_1225_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i47522_3_lut (.I0(n62448), .I1(n285[15]), .I2(n31_adj_4266), 
            .I3(GND_net), .O(n62235));   // verilog/motorControl.v(58[23:46])
    defparam i47522_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY mult_24_add_1225_15 (.CI(n46928), .I0(n10031[12]), .I1(n1023), 
            .CO(n46929));
    SB_LUT4 mult_24_add_1225_14_lut (.I0(GND_net), .I1(n10031[11]), .I2(n950), 
            .I3(n46927), .O(n42[13])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_24_add_1225_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_24_add_1225_14 (.CI(n46927), .I0(n10031[11]), .I1(n950), 
            .CO(n46928));
    SB_LUT4 mult_24_add_1225_13_lut (.I0(GND_net), .I1(n10031[10]), .I2(n877), 
            .I3(n46926), .O(n42[12])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_24_add_1225_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_24_add_1225_13 (.CI(n46926), .I0(n10031[10]), .I1(n877), 
            .CO(n46927));
    SB_LUT4 mult_24_add_1225_12_lut (.I0(GND_net), .I1(n10031[9]), .I2(n804), 
            .I3(n46925), .O(n42[11])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_24_add_1225_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_24_add_1225_12 (.CI(n46925), .I0(n10031[9]), .I1(n804), 
            .CO(n46926));
    SB_LUT4 mult_24_add_1225_11_lut (.I0(GND_net), .I1(n10031[8]), .I2(n731), 
            .I3(n46924), .O(n42[10])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_24_add_1225_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_24_add_1225_11 (.CI(n46924), .I0(n10031[8]), .I1(n731), 
            .CO(n46925));
    SB_LUT4 mult_24_add_1225_10_lut (.I0(GND_net), .I1(n10031[7]), .I2(n658), 
            .I3(n46923), .O(n42[9])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_24_add_1225_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_24_add_1225_10 (.CI(n46923), .I0(n10031[7]), .I1(n658), 
            .CO(n46924));
    SB_LUT4 mult_24_add_1225_9_lut (.I0(GND_net), .I1(n10031[6]), .I2(n585), 
            .I3(n46922), .O(n42[8])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_24_add_1225_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_23_i506_2_lut (.I0(\Kp[10] ), .I1(n207[11]), .I2(GND_net), 
            .I3(GND_net), .O(n752));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i506_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY mult_24_add_1225_9 (.CI(n46922), .I0(n10031[6]), .I1(n585), 
            .CO(n46923));
    SB_LUT4 mult_24_add_1225_8_lut (.I0(GND_net), .I1(n10031[5]), .I2(n512), 
            .I3(n46921), .O(n42[7])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_24_add_1225_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_24_add_1225_8 (.CI(n46921), .I0(n10031[5]), .I1(n512), 
            .CO(n46922));
    SB_LUT4 mult_23_i555_2_lut (.I0(\Kp[11] ), .I1(n207[11]), .I2(GND_net), 
            .I3(GND_net), .O(n825));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i555_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 n9440_bdd_4_lut_48658 (.I0(n9440), .I1(n59883), .I2(setpoint[6]), 
            .I3(n4357), .O(n63389));
    defparam n9440_bdd_4_lut_48658.LUT_INIT = 16'he4aa;
    SB_LUT4 mult_24_add_1225_7_lut (.I0(GND_net), .I1(n10031[4]), .I2(n439_adj_4325), 
            .I3(n46920), .O(n42[6])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_24_add_1225_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_24_add_1225_7 (.CI(n46920), .I0(n10031[4]), .I1(n439_adj_4325), 
            .CO(n46921));
    SB_LUT4 mult_24_add_1225_6_lut (.I0(GND_net), .I1(n10031[3]), .I2(n366), 
            .I3(n46919), .O(n42[5])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_24_add_1225_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_24_add_1225_6 (.CI(n46919), .I0(n10031[3]), .I1(n366), 
            .CO(n46920));
    SB_LUT4 mult_24_add_1225_5_lut (.I0(GND_net), .I1(n10031[2]), .I2(n293_adj_4326), 
            .I3(n46918), .O(n42[4])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_24_add_1225_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_24_add_1225_5 (.CI(n46918), .I0(n10031[2]), .I1(n293_adj_4326), 
            .CO(n46919));
    SB_LUT4 mult_24_add_1225_4_lut (.I0(GND_net), .I1(n10031[1]), .I2(n220_adj_4327), 
            .I3(n46917), .O(n42[3])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_24_add_1225_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_24_add_1225_4 (.CI(n46917), .I0(n10031[1]), .I1(n220_adj_4327), 
            .CO(n46918));
    SB_LUT4 mult_24_add_1225_3_lut (.I0(GND_net), .I1(n10031[0]), .I2(n147), 
            .I3(n46916), .O(n42[2])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_24_add_1225_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_24_add_1225_3 (.CI(n46916), .I0(n10031[0]), .I1(n147), 
            .CO(n46917));
    SB_LUT4 mult_24_add_1225_2_lut (.I0(GND_net), .I1(n5_adj_4328), .I2(n74_adj_4329), 
            .I3(GND_net), .O(n42[1])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_24_add_1225_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_24_add_1225_2 (.CI(GND_net), .I0(n5_adj_4328), .I1(n74_adj_4329), 
            .CO(n46916));
    SB_LUT4 add_4304_23_lut (.I0(GND_net), .I1(n11044[20]), .I2(GND_net), 
            .I3(n46915), .O(n10031[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4304_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4304_22_lut (.I0(GND_net), .I1(n11044[19]), .I2(GND_net), 
            .I3(n46914), .O(n10031[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4304_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4304_22 (.CI(n46914), .I0(n11044[19]), .I1(GND_net), 
            .CO(n46915));
    SB_LUT4 add_4304_21_lut (.I0(GND_net), .I1(n11044[18]), .I2(GND_net), 
            .I3(n46913), .O(n10031[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4304_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4304_21 (.CI(n46913), .I0(n11044[18]), .I1(GND_net), 
            .CO(n46914));
    SB_LUT4 add_4304_20_lut (.I0(GND_net), .I1(n11044[17]), .I2(GND_net), 
            .I3(n46912), .O(n10031[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4304_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4304_20 (.CI(n46912), .I0(n11044[17]), .I1(GND_net), 
            .CO(n46913));
    SB_LUT4 add_4304_19_lut (.I0(GND_net), .I1(n11044[16]), .I2(GND_net), 
            .I3(n46911), .O(n10031[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4304_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4304_19 (.CI(n46911), .I0(n11044[16]), .I1(GND_net), 
            .CO(n46912));
    SB_LUT4 add_4304_18_lut (.I0(GND_net), .I1(n11044[15]), .I2(GND_net), 
            .I3(n46910), .O(n10031[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4304_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4304_18 (.CI(n46910), .I0(n11044[15]), .I1(GND_net), 
            .CO(n46911));
    SB_LUT4 add_4304_17_lut (.I0(GND_net), .I1(n11044[14]), .I2(GND_net), 
            .I3(n46909), .O(n10031[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4304_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4304_17 (.CI(n46909), .I0(n11044[14]), .I1(GND_net), 
            .CO(n46910));
    SB_LUT4 add_4304_16_lut (.I0(GND_net), .I1(n11044[13]), .I2(n1099), 
            .I3(n46908), .O(n10031[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4304_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4304_16 (.CI(n46908), .I0(n11044[13]), .I1(n1099), .CO(n46909));
    SB_LUT4 add_4304_15_lut (.I0(GND_net), .I1(n11044[12]), .I2(n1026), 
            .I3(n46907), .O(n10031[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4304_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4304_15 (.CI(n46907), .I0(n11044[12]), .I1(n1026), .CO(n46908));
    SB_LUT4 add_4304_14_lut (.I0(GND_net), .I1(n11044[11]), .I2(n953), 
            .I3(n46906), .O(n10031[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4304_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4304_14 (.CI(n46906), .I0(n11044[11]), .I1(n953), .CO(n46907));
    SB_LUT4 add_4304_13_lut (.I0(GND_net), .I1(n11044[10]), .I2(n880), 
            .I3(n46905), .O(n10031[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4304_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4304_13 (.CI(n46905), .I0(n11044[10]), .I1(n880), .CO(n46906));
    SB_LUT4 add_4304_12_lut (.I0(GND_net), .I1(n11044[9]), .I2(n807), 
            .I3(n46904), .O(n10031[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4304_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4304_12 (.CI(n46904), .I0(n11044[9]), .I1(n807), .CO(n46905));
    SB_LUT4 add_4304_11_lut (.I0(GND_net), .I1(n11044[8]), .I2(n734), 
            .I3(n46903), .O(n10031[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4304_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4304_11 (.CI(n46903), .I0(n11044[8]), .I1(n734), .CO(n46904));
    SB_LUT4 add_4304_10_lut (.I0(GND_net), .I1(n11044[7]), .I2(n661), 
            .I3(n46902), .O(n10031[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4304_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4304_10 (.CI(n46902), .I0(n11044[7]), .I1(n661), .CO(n46903));
    SB_LUT4 add_4304_9_lut (.I0(GND_net), .I1(n11044[6]), .I2(n588), .I3(n46901), 
            .O(n10031[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4304_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4304_9 (.CI(n46901), .I0(n11044[6]), .I1(n588), .CO(n46902));
    SB_LUT4 add_4304_8_lut (.I0(GND_net), .I1(n11044[5]), .I2(n515), .I3(n46900), 
            .O(n10031[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4304_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4304_8 (.CI(n46900), .I0(n11044[5]), .I1(n515), .CO(n46901));
    SB_LUT4 add_4304_7_lut (.I0(GND_net), .I1(n11044[4]), .I2(n442_adj_4330), 
            .I3(n46899), .O(n10031[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4304_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4304_7 (.CI(n46899), .I0(n11044[4]), .I1(n442_adj_4330), 
            .CO(n46900));
    SB_LUT4 add_4304_6_lut (.I0(GND_net), .I1(n11044[3]), .I2(n369), .I3(n46898), 
            .O(n10031[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4304_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4304_6 (.CI(n46898), .I0(n11044[3]), .I1(n369), .CO(n46899));
    SB_LUT4 i48250_4_lut (.I0(n62235), .I1(n62775), .I2(n35), .I3(n60019), 
            .O(n62963));   // verilog/motorControl.v(58[23:46])
    defparam i48250_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 add_4304_5_lut (.I0(GND_net), .I1(n11044[2]), .I2(n296_adj_4331), 
            .I3(n46897), .O(n10031[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4304_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i48251_3_lut (.I0(n62963), .I1(n285[18]), .I2(n37_adj_4264), 
            .I3(GND_net), .O(n62964));   // verilog/motorControl.v(58[23:46])
    defparam i48251_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_4304_5 (.CI(n46897), .I0(n11044[2]), .I1(n296_adj_4331), 
            .CO(n46898));
    SB_LUT4 add_4304_4_lut (.I0(GND_net), .I1(n11044[1]), .I2(n223_adj_4332), 
            .I3(n46896), .O(n10031[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4304_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4304_4 (.CI(n46896), .I0(n11044[1]), .I1(n223_adj_4332), 
            .CO(n46897));
    SB_LUT4 add_4304_3_lut (.I0(GND_net), .I1(n11044[0]), .I2(n150), .I3(n46895), 
            .O(n10031[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4304_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4304_3 (.CI(n46895), .I0(n11044[0]), .I1(n150), .CO(n46896));
    SB_LUT4 add_4304_2_lut (.I0(GND_net), .I1(n8_adj_4333), .I2(n77), 
            .I3(GND_net), .O(n10031[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4304_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4304_2 (.CI(GND_net), .I0(n8_adj_4333), .I1(n77), .CO(n46895));
    SB_LUT4 i48196_3_lut (.I0(n62964), .I1(n285[19]), .I2(n39_adj_4261), 
            .I3(GND_net), .O(n62909));   // verilog/motorControl.v(58[23:46])
    defparam i48196_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_4349_22_lut (.I0(GND_net), .I1(n11965[19]), .I2(GND_net), 
            .I3(n46894), .O(n11044[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4349_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4349_21_lut (.I0(GND_net), .I1(n11965[18]), .I2(GND_net), 
            .I3(n46893), .O(n11044[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4349_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4349_21 (.CI(n46893), .I0(n11965[18]), .I1(GND_net), 
            .CO(n46894));
    SB_LUT4 add_4349_20_lut (.I0(GND_net), .I1(n11965[17]), .I2(GND_net), 
            .I3(n46892), .O(n11044[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4349_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4349_20 (.CI(n46892), .I0(n11965[17]), .I1(GND_net), 
            .CO(n46893));
    SB_LUT4 add_4349_19_lut (.I0(GND_net), .I1(n11965[16]), .I2(GND_net), 
            .I3(n46891), .O(n11044[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4349_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4349_19 (.CI(n46891), .I0(n11965[16]), .I1(GND_net), 
            .CO(n46892));
    SB_LUT4 i45275_4_lut (.I0(n43_adj_4260), .I1(n41_adj_4259), .I2(n39_adj_4261), 
            .I3(n62737), .O(n59987));
    defparam i45275_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 add_4349_18_lut (.I0(GND_net), .I1(n11965[15]), .I2(GND_net), 
            .I3(n46890), .O(n11044[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4349_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4349_18 (.CI(n46890), .I0(n11965[15]), .I1(GND_net), 
            .CO(n46891));
    SB_LUT4 i47525_4_lut (.I0(n62233), .I1(n61879), .I2(n45_adj_4258), 
            .I3(n59983), .O(n62238));   // verilog/motorControl.v(58[23:46])
    defparam i47525_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 add_4349_17_lut (.I0(GND_net), .I1(n11965[14]), .I2(GND_net), 
            .I3(n46889), .O(n11044[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4349_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4349_17 (.CI(n46889), .I0(n11965[14]), .I1(GND_net), 
            .CO(n46890));
    SB_LUT4 i48151_3_lut (.I0(n62909), .I1(n285[20]), .I2(n41_adj_4259), 
            .I3(GND_net), .O(n40));   // verilog/motorControl.v(58[23:46])
    defparam i48151_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_4349_16_lut (.I0(GND_net), .I1(n11965[13]), .I2(n1102), 
            .I3(n46888), .O(n11044[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4349_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4349_16 (.CI(n46888), .I0(n11965[13]), .I1(n1102), .CO(n46889));
    SB_LUT4 add_4349_15_lut (.I0(GND_net), .I1(n11965[12]), .I2(n1029), 
            .I3(n46887), .O(n11044[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4349_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4349_15 (.CI(n46887), .I0(n11965[12]), .I1(n1029), .CO(n46888));
    SB_LUT4 i47844_4_lut (.I0(n40), .I1(n62238), .I2(n45_adj_4258), .I3(n59987), 
            .O(n62557));   // verilog/motorControl.v(58[23:46])
    defparam i47844_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i47845_3_lut (.I0(n62557), .I1(n233[23]), .I2(n285[23]), .I3(GND_net), 
            .O(n284));   // verilog/motorControl.v(58[23:46])
    defparam i47845_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 mult_23_i604_2_lut (.I0(\Kp[12] ), .I1(n207[11]), .I2(GND_net), 
            .I3(GND_net), .O(n898));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i604_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i653_2_lut (.I0(\Kp[13] ), .I1(n207[11]), .I2(GND_net), 
            .I3(GND_net), .O(n971));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i653_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_4349_14_lut (.I0(GND_net), .I1(n11965[11]), .I2(n956), 
            .I3(n46886), .O(n11044[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4349_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4349_14 (.CI(n46886), .I0(n11965[11]), .I1(n956), .CO(n46887));
    SB_LUT4 add_4349_13_lut (.I0(GND_net), .I1(n11965[10]), .I2(n883), 
            .I3(n46885), .O(n11044[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4349_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4349_13 (.CI(n46885), .I0(n11965[10]), .I1(n883), .CO(n46886));
    SB_LUT4 add_4349_12_lut (.I0(GND_net), .I1(n11965[9]), .I2(n810), 
            .I3(n46884), .O(n11044[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4349_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4349_12 (.CI(n46884), .I0(n11965[9]), .I1(n810), .CO(n46885));
    SB_LUT4 mux_21_i16_3_lut (.I0(n233[15]), .I1(n285[15]), .I2(n284), 
            .I3(GND_net), .O(n310[15]));   // verilog/motorControl.v(58[20] 60[14])
    defparam mux_21_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_22_i16_3_lut (.I0(n310[15]), .I1(IntegralLimit[15]), .I2(n258), 
            .I3(GND_net), .O(n344));   // verilog/motorControl.v(58[20] 60[14])
    defparam mux_22_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_24_i424_2_lut (.I0(\Ki[8] ), .I1(n344), .I2(GND_net), 
            .I3(GND_net), .O(n630));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i424_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_4349_11_lut (.I0(GND_net), .I1(n11965[8]), .I2(n737), 
            .I3(n46883), .O(n11044[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4349_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4349_11 (.CI(n46883), .I0(n11965[8]), .I1(n737), .CO(n46884));
    SB_LUT4 add_4349_10_lut (.I0(GND_net), .I1(n11965[7]), .I2(n664), 
            .I3(n46882), .O(n11044[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4349_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4349_10 (.CI(n46882), .I0(n11965[7]), .I1(n664), .CO(n46883));
    SB_LUT4 mult_23_i702_2_lut (.I0(\Kp[14] ), .I1(n207[11]), .I2(GND_net), 
            .I3(GND_net), .O(n1044));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i702_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i751_2_lut (.I0(\Kp[15] ), .I1(n207[11]), .I2(GND_net), 
            .I3(GND_net), .O(n1117));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i751_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_4349_9_lut (.I0(GND_net), .I1(n11965[6]), .I2(n591), .I3(n46881), 
            .O(n11044[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4349_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_24_i83_2_lut (.I0(\Ki[1] ), .I1(n343), .I2(GND_net), 
            .I3(GND_net), .O(n122_adj_4240));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i83_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_4349_9 (.CI(n46881), .I0(n11965[6]), .I1(n591), .CO(n46882));
    SB_LUT4 add_4349_8_lut (.I0(GND_net), .I1(n11965[5]), .I2(n518), .I3(n46880), 
            .O(n11044[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4349_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4349_8 (.CI(n46880), .I0(n11965[5]), .I1(n518), .CO(n46881));
    SB_LUT4 mult_24_i414_2_lut (.I0(\Ki[8] ), .I1(n349), .I2(GND_net), 
            .I3(GND_net), .O(n615));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i414_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_27_inv_0_i2_1_lut (.I0(\deadband[1] ), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n28[1]));   // verilog/motorControl.v(62[45:54])
    defparam unary_minus_27_inv_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_4349_7_lut (.I0(GND_net), .I1(n11965[4]), .I2(n445_adj_4334), 
            .I3(n46879), .O(n11044[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4349_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4349_7 (.CI(n46879), .I0(n11965[4]), .I1(n445_adj_4334), 
            .CO(n46880));
    SB_LUT4 mult_23_i747_2_lut (.I0(\Kp[15] ), .I1(n207[9]), .I2(GND_net), 
            .I3(GND_net), .O(n1111));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i747_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_4349_6_lut (.I0(GND_net), .I1(n11965[3]), .I2(n372), .I3(n46878), 
            .O(n11044[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4349_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4349_6 (.CI(n46878), .I0(n11965[3]), .I1(n372), .CO(n46879));
    SB_LUT4 n63389_bdd_4_lut (.I0(n63389), .I1(n535[6]), .I2(n455[6]), 
            .I3(n4357), .O(n63392));
    defparam n63389_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 add_4349_5_lut (.I0(GND_net), .I1(n11965[2]), .I2(n299_adj_4335), 
            .I3(n46877), .O(n11044[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4349_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4349_5 (.CI(n46877), .I0(n11965[2]), .I1(n299_adj_4335), 
            .CO(n46878));
    SB_LUT4 add_4349_4_lut (.I0(GND_net), .I1(n11965[1]), .I2(n226_adj_4336), 
            .I3(n46876), .O(n11044[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4349_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4349_4 (.CI(n46876), .I0(n11965[1]), .I1(n226_adj_4336), 
            .CO(n46877));
    SB_LUT4 add_4349_3_lut (.I0(GND_net), .I1(n11965[0]), .I2(n153), .I3(n46875), 
            .O(n11044[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4349_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4349_3 (.CI(n46875), .I0(n11965[0]), .I1(n153), .CO(n46876));
    SB_LUT4 add_4349_2_lut (.I0(GND_net), .I1(n11_adj_4337), .I2(n80), 
            .I3(GND_net), .O(n11044[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4349_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4349_2 (.CI(GND_net), .I0(n11_adj_4337), .I1(n80), .CO(n46875));
    SB_LUT4 add_4390_21_lut (.I0(GND_net), .I1(n12802[18]), .I2(GND_net), 
            .I3(n46874), .O(n11965[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4390_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4390_20_lut (.I0(GND_net), .I1(n12802[17]), .I2(GND_net), 
            .I3(n46873), .O(n11965[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4390_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4390_20 (.CI(n46873), .I0(n12802[17]), .I1(GND_net), 
            .CO(n46874));
    SB_LUT4 add_4390_19_lut (.I0(GND_net), .I1(n12802[16]), .I2(GND_net), 
            .I3(n46872), .O(n11965[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4390_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4390_19 (.CI(n46872), .I0(n12802[16]), .I1(GND_net), 
            .CO(n46873));
    SB_LUT4 add_4390_18_lut (.I0(GND_net), .I1(n12802[15]), .I2(GND_net), 
            .I3(n46871), .O(n11965[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4390_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4390_18 (.CI(n46871), .I0(n12802[15]), .I1(GND_net), 
            .CO(n46872));
    SB_LUT4 add_4390_17_lut (.I0(GND_net), .I1(n12802[14]), .I2(GND_net), 
            .I3(n46870), .O(n11965[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4390_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4390_17 (.CI(n46870), .I0(n12802[14]), .I1(GND_net), 
            .CO(n46871));
    SB_LUT4 add_4390_16_lut (.I0(GND_net), .I1(n12802[13]), .I2(n1105), 
            .I3(n46869), .O(n11965[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4390_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4390_16 (.CI(n46869), .I0(n12802[13]), .I1(n1105), .CO(n46870));
    SB_LUT4 add_4390_15_lut (.I0(GND_net), .I1(n12802[12]), .I2(n1032), 
            .I3(n46868), .O(n11965[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4390_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4390_15 (.CI(n46868), .I0(n12802[12]), .I1(n1032), .CO(n46869));
    SB_LUT4 add_4390_14_lut (.I0(GND_net), .I1(n12802[11]), .I2(n959), 
            .I3(n46867), .O(n11965[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4390_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4390_14 (.CI(n46867), .I0(n12802[11]), .I1(n959), .CO(n46868));
    SB_LUT4 add_4390_13_lut (.I0(GND_net), .I1(n12802[10]), .I2(n886), 
            .I3(n46866), .O(n11965[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4390_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4390_13 (.CI(n46866), .I0(n12802[10]), .I1(n886), .CO(n46867));
    SB_LUT4 add_4390_12_lut (.I0(GND_net), .I1(n12802[9]), .I2(n813), 
            .I3(n46865), .O(n11965[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4390_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4390_12 (.CI(n46865), .I0(n12802[9]), .I1(n813), .CO(n46866));
    SB_DFFER result_i0_i23 (.Q(duty[23]), .C(clk16MHz), .E(control_update), 
            .D(n63554), .R(reset));   // verilog/motorControl.v(42[14] 73[8])
    SB_DFFER result_i0_i22 (.Q(duty[22]), .C(clk16MHz), .E(control_update), 
            .D(n63512), .R(reset));   // verilog/motorControl.v(42[14] 73[8])
    SB_DFFER result_i0_i21 (.Q(duty[21]), .C(clk16MHz), .E(control_update), 
            .D(n63506), .R(reset));   // verilog/motorControl.v(42[14] 73[8])
    SB_DFFER result_i0_i20 (.Q(duty[20]), .C(clk16MHz), .E(control_update), 
            .D(n63488), .R(reset));   // verilog/motorControl.v(42[14] 73[8])
    SB_DFFER result_i0_i19 (.Q(duty[19]), .C(clk16MHz), .E(control_update), 
            .D(n63482), .R(reset));   // verilog/motorControl.v(42[14] 73[8])
    SB_DFFER result_i0_i18 (.Q(duty[18]), .C(clk16MHz), .E(control_update), 
            .D(n63470), .R(reset));   // verilog/motorControl.v(42[14] 73[8])
    SB_DFFER result_i0_i17 (.Q(duty[17]), .C(clk16MHz), .E(control_update), 
            .D(n63464), .R(reset));   // verilog/motorControl.v(42[14] 73[8])
    SB_DFFER result_i0_i16 (.Q(duty[16]), .C(clk16MHz), .E(control_update), 
            .D(n63458), .R(reset));   // verilog/motorControl.v(42[14] 73[8])
    SB_DFFER result_i0_i15 (.Q(duty[15]), .C(clk16MHz), .E(control_update), 
            .D(n63452), .R(reset));   // verilog/motorControl.v(42[14] 73[8])
    SB_DFFER result_i0_i14 (.Q(duty[14]), .C(clk16MHz), .E(control_update), 
            .D(n63446), .R(reset));   // verilog/motorControl.v(42[14] 73[8])
    SB_DFFER result_i0_i13 (.Q(duty[13]), .C(clk16MHz), .E(control_update), 
            .D(n63440), .R(reset));   // verilog/motorControl.v(42[14] 73[8])
    SB_DFFER result_i0_i12 (.Q(duty[12]), .C(clk16MHz), .E(control_update), 
            .D(n63434), .R(reset));   // verilog/motorControl.v(42[14] 73[8])
    SB_DFFER result_i0_i11 (.Q(duty[11]), .C(clk16MHz), .E(control_update), 
            .D(n63428), .R(reset));   // verilog/motorControl.v(42[14] 73[8])
    SB_DFFER result_i0_i10 (.Q(duty[10]), .C(clk16MHz), .E(control_update), 
            .D(n63422), .R(reset));   // verilog/motorControl.v(42[14] 73[8])
    SB_DFFER result_i0_i9 (.Q(duty[9]), .C(clk16MHz), .E(control_update), 
            .D(n63410), .R(reset));   // verilog/motorControl.v(42[14] 73[8])
    SB_DFFER result_i0_i8 (.Q(duty[8]), .C(clk16MHz), .E(control_update), 
            .D(n63404), .R(reset));   // verilog/motorControl.v(42[14] 73[8])
    SB_DFFER result_i0_i7 (.Q(duty[7]), .C(clk16MHz), .E(control_update), 
            .D(n63398), .R(reset));   // verilog/motorControl.v(42[14] 73[8])
    SB_DFFER result_i0_i6 (.Q(duty[6]), .C(clk16MHz), .E(control_update), 
            .D(n63392), .R(reset));   // verilog/motorControl.v(42[14] 73[8])
    SB_DFFER result_i0_i5 (.Q(duty[5]), .C(clk16MHz), .E(control_update), 
            .D(n63380), .R(reset));   // verilog/motorControl.v(42[14] 73[8])
    SB_DFFER result_i0_i4 (.Q(duty[4]), .C(clk16MHz), .E(control_update), 
            .D(n63368), .R(reset));   // verilog/motorControl.v(42[14] 73[8])
    SB_DFFER result_i0_i3 (.Q(duty[3]), .C(clk16MHz), .E(control_update), 
            .D(n63356), .R(reset));   // verilog/motorControl.v(42[14] 73[8])
    SB_DFFER result_i0_i2 (.Q(duty[2]), .C(clk16MHz), .E(control_update), 
            .D(n63344), .R(reset));   // verilog/motorControl.v(42[14] 73[8])
    SB_DFFER result_i0_i1 (.Q(duty[1]), .C(clk16MHz), .E(control_update), 
            .D(n63278), .R(reset));   // verilog/motorControl.v(42[14] 73[8])
    SB_LUT4 add_4390_11_lut (.I0(GND_net), .I1(n12802[8]), .I2(n740), 
            .I3(n46864), .O(n11965[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4390_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4390_11 (.CI(n46864), .I0(n12802[8]), .I1(n740), .CO(n46865));
    SB_LUT4 add_4390_10_lut (.I0(GND_net), .I1(n12802[7]), .I2(n667), 
            .I3(n46863), .O(n11965[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4390_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4390_10 (.CI(n46863), .I0(n12802[7]), .I1(n667), .CO(n46864));
    SB_LUT4 add_4390_9_lut (.I0(GND_net), .I1(n12802[6]), .I2(n594), .I3(n46862), 
            .O(n11965[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4390_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4390_9 (.CI(n46862), .I0(n12802[6]), .I1(n594), .CO(n46863));
    SB_LUT4 add_4390_8_lut (.I0(GND_net), .I1(n12802[5]), .I2(n521), .I3(n46861), 
            .O(n11965[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4390_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4390_8 (.CI(n46861), .I0(n12802[5]), .I1(n521), .CO(n46862));
    SB_LUT4 add_4390_7_lut (.I0(GND_net), .I1(n12802[4]), .I2(n448_adj_4338), 
            .I3(n46860), .O(n11965[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4390_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4390_7 (.CI(n46860), .I0(n12802[4]), .I1(n448_adj_4338), 
            .CO(n46861));
    SB_LUT4 add_4390_6_lut (.I0(GND_net), .I1(n12802[3]), .I2(n375), .I3(n46859), 
            .O(n11965[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4390_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4390_6 (.CI(n46859), .I0(n12802[3]), .I1(n375), .CO(n46860));
    SB_DFFSR counter_1940_1941__i2 (.Q(counter[1]), .C(clk16MHz), .D(n61[1]), 
            .R(counter_31__N_3487));   // verilog/motorControl.v(25[16:25])
    SB_DFFSR counter_1940_1941__i3 (.Q(counter[2]), .C(clk16MHz), .D(n61[2]), 
            .R(counter_31__N_3487));   // verilog/motorControl.v(25[16:25])
    SB_DFFSR counter_1940_1941__i4 (.Q(counter[3]), .C(clk16MHz), .D(n61[3]), 
            .R(counter_31__N_3487));   // verilog/motorControl.v(25[16:25])
    SB_DFFSR counter_1940_1941__i5 (.Q(counter[4]), .C(clk16MHz), .D(n61[4]), 
            .R(counter_31__N_3487));   // verilog/motorControl.v(25[16:25])
    SB_DFFSR counter_1940_1941__i6 (.Q(counter[5]), .C(clk16MHz), .D(n61[5]), 
            .R(counter_31__N_3487));   // verilog/motorControl.v(25[16:25])
    SB_DFFSR counter_1940_1941__i7 (.Q(counter[6]), .C(clk16MHz), .D(n61[6]), 
            .R(counter_31__N_3487));   // verilog/motorControl.v(25[16:25])
    SB_DFFSR counter_1940_1941__i8 (.Q(counter[7]), .C(clk16MHz), .D(n61[7]), 
            .R(counter_31__N_3487));   // verilog/motorControl.v(25[16:25])
    SB_DFFSR counter_1940_1941__i9 (.Q(counter[8]), .C(clk16MHz), .D(n61[8]), 
            .R(counter_31__N_3487));   // verilog/motorControl.v(25[16:25])
    SB_DFFSR counter_1940_1941__i10 (.Q(counter[9]), .C(clk16MHz), .D(n61[9]), 
            .R(counter_31__N_3487));   // verilog/motorControl.v(25[16:25])
    SB_DFFSR counter_1940_1941__i11 (.Q(counter[10]), .C(clk16MHz), .D(n61[10]), 
            .R(counter_31__N_3487));   // verilog/motorControl.v(25[16:25])
    SB_DFFSR counter_1940_1941__i12 (.Q(counter[11]), .C(clk16MHz), .D(n61[11]), 
            .R(counter_31__N_3487));   // verilog/motorControl.v(25[16:25])
    SB_DFFSR counter_1940_1941__i13 (.Q(counter[12]), .C(clk16MHz), .D(n61[12]), 
            .R(counter_31__N_3487));   // verilog/motorControl.v(25[16:25])
    SB_DFFSR counter_1940_1941__i14 (.Q(counter[13]), .C(clk16MHz), .D(n61[13]), 
            .R(counter_31__N_3487));   // verilog/motorControl.v(25[16:25])
    SB_LUT4 add_4390_5_lut (.I0(GND_net), .I1(n12802[2]), .I2(n302_adj_4339), 
            .I3(n46858), .O(n11965[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4390_5_lut.LUT_INIT = 16'hC33C;
    SB_DFFR \PID_CONTROLLER.integral_i0_i0  (.Q(\PID_CONTROLLER.integral [0]), 
            .C(clk16MHz), .D(n26085), .R(reset));   // verilog/motorControl.v(42[14] 73[8])
    SB_CARRY add_4390_5 (.CI(n46858), .I0(n12802[2]), .I1(n302_adj_4339), 
            .CO(n46859));
    SB_LUT4 add_4390_4_lut (.I0(GND_net), .I1(n12802[1]), .I2(n229), .I3(n46857), 
            .O(n11965[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4390_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4390_4 (.CI(n46857), .I0(n12802[1]), .I1(n229), .CO(n46858));
    SB_LUT4 add_4390_3_lut (.I0(GND_net), .I1(n12802[0]), .I2(n156), .I3(n46856), 
            .O(n11965[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4390_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4390_3 (.CI(n46856), .I0(n12802[0]), .I1(n156), .CO(n46857));
    SB_LUT4 add_4390_2_lut (.I0(GND_net), .I1(n14_adj_4340), .I2(n83), 
            .I3(GND_net), .O(n11965[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4390_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4390_2 (.CI(GND_net), .I0(n14_adj_4340), .I1(n83), .CO(n46856));
    SB_LUT4 add_4678_12_lut (.I0(GND_net), .I1(n17311[9]), .I2(n840_adj_4341), 
            .I3(n46855), .O(n17071[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4678_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4678_11_lut (.I0(GND_net), .I1(n17311[8]), .I2(n767_adj_4342), 
            .I3(n46854), .O(n17071[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4678_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4678_11 (.CI(n46854), .I0(n17311[8]), .I1(n767_adj_4342), 
            .CO(n46855));
    SB_LUT4 add_4678_10_lut (.I0(GND_net), .I1(n17311[7]), .I2(n694_adj_4343), 
            .I3(n46853), .O(n17071[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4678_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4678_10 (.CI(n46853), .I0(n17311[7]), .I1(n694_adj_4343), 
            .CO(n46854));
    SB_LUT4 add_4678_9_lut (.I0(GND_net), .I1(n17311[6]), .I2(n621_adj_4344), 
            .I3(n46852), .O(n17071[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4678_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4678_9 (.CI(n46852), .I0(n17311[6]), .I1(n621_adj_4344), 
            .CO(n46853));
    SB_LUT4 add_4678_8_lut (.I0(GND_net), .I1(n17311[5]), .I2(n548_adj_4345), 
            .I3(n46851), .O(n17071[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4678_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4678_8 (.CI(n46851), .I0(n17311[5]), .I1(n548_adj_4345), 
            .CO(n46852));
    SB_LUT4 add_4678_7_lut (.I0(GND_net), .I1(n17311[4]), .I2(n475_adj_4346), 
            .I3(n46850), .O(n17071[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4678_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4678_7 (.CI(n46850), .I0(n17311[4]), .I1(n475_adj_4346), 
            .CO(n46851));
    SB_LUT4 add_4678_6_lut (.I0(GND_net), .I1(n17311[3]), .I2(n402_adj_4347), 
            .I3(n46849), .O(n17071[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4678_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4678_6 (.CI(n46849), .I0(n17311[3]), .I1(n402_adj_4347), 
            .CO(n46850));
    SB_LUT4 add_4678_5_lut (.I0(GND_net), .I1(n17311[2]), .I2(n329_adj_4348), 
            .I3(n46848), .O(n17071[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4678_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_25_25_lut (.I0(GND_net), .I1(n10055[0]), .I2(n9524[0]), 
            .I3(n46095), .O(n455[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_25_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4678_5 (.CI(n46848), .I0(n17311[2]), .I1(n329_adj_4348), 
            .CO(n46849));
    SB_LUT4 add_4678_4_lut (.I0(GND_net), .I1(n17311[1]), .I2(n256_adj_4349), 
            .I3(n46847), .O(n17071[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4678_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4678_4 (.CI(n46847), .I0(n17311[1]), .I1(n256_adj_4349), 
            .CO(n46848));
    SB_LUT4 add_25_24_lut (.I0(GND_net), .I1(n360[22]), .I2(n42[22]), 
            .I3(n46094), .O(n455[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_25_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_25_24 (.CI(n46094), .I0(n360[22]), .I1(n42[22]), .CO(n46095));
    SB_LUT4 add_25_23_lut (.I0(GND_net), .I1(n360[21]), .I2(n42[21]), 
            .I3(n46093), .O(n455[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_25_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_25_23 (.CI(n46093), .I0(n360[21]), .I1(n42[21]), .CO(n46094));
    SB_LUT4 add_4678_3_lut (.I0(GND_net), .I1(n17311[0]), .I2(n183_adj_4351), 
            .I3(n46846), .O(n17071[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4678_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4678_3 (.CI(n46846), .I0(n17311[0]), .I1(n183_adj_4351), 
            .CO(n46847));
    SB_LUT4 add_4678_2_lut (.I0(GND_net), .I1(n41_adj_4352), .I2(n110_adj_4353), 
            .I3(GND_net), .O(n17071[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4678_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4678_2 (.CI(GND_net), .I0(n41_adj_4352), .I1(n110_adj_4353), 
            .CO(n46846));
    SB_LUT4 add_4429_20_lut (.I0(GND_net), .I1(n13559[17]), .I2(GND_net), 
            .I3(n46845), .O(n12802[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4429_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4429_19_lut (.I0(GND_net), .I1(n13559[16]), .I2(GND_net), 
            .I3(n46844), .O(n12802[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4429_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4429_19 (.CI(n46844), .I0(n13559[16]), .I1(GND_net), 
            .CO(n46845));
    SB_LUT4 add_25_22_lut (.I0(GND_net), .I1(n360[20]), .I2(n42[20]), 
            .I3(n46092), .O(n455[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_25_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_25_22 (.CI(n46092), .I0(n360[20]), .I1(n42[20]), .CO(n46093));
    SB_LUT4 add_25_21_lut (.I0(GND_net), .I1(n360[19]), .I2(n42[19]), 
            .I3(n46091), .O(n455[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_25_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4429_18_lut (.I0(GND_net), .I1(n13559[15]), .I2(GND_net), 
            .I3(n46843), .O(n12802[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4429_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4429_18 (.CI(n46843), .I0(n13559[15]), .I1(GND_net), 
            .CO(n46844));
    SB_LUT4 add_4429_17_lut (.I0(GND_net), .I1(n13559[14]), .I2(GND_net), 
            .I3(n46842), .O(n12802[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4429_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4429_17 (.CI(n46842), .I0(n13559[14]), .I1(GND_net), 
            .CO(n46843));
    SB_LUT4 add_4429_16_lut (.I0(GND_net), .I1(n13559[13]), .I2(n1108), 
            .I3(n46841), .O(n12802[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4429_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4429_16 (.CI(n46841), .I0(n13559[13]), .I1(n1108), .CO(n46842));
    SB_LUT4 add_4429_15_lut (.I0(GND_net), .I1(n13559[12]), .I2(n1035), 
            .I3(n46840), .O(n12802[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4429_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4429_15 (.CI(n46840), .I0(n13559[12]), .I1(n1035), .CO(n46841));
    SB_LUT4 add_4429_14_lut (.I0(GND_net), .I1(n13559[11]), .I2(n962), 
            .I3(n46839), .O(n12802[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4429_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4429_14 (.CI(n46839), .I0(n13559[11]), .I1(n962), .CO(n46840));
    SB_LUT4 add_4429_13_lut (.I0(GND_net), .I1(n13559[10]), .I2(n889), 
            .I3(n46838), .O(n12802[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4429_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_25_21 (.CI(n46091), .I0(n360[19]), .I1(n42[19]), .CO(n46092));
    SB_CARRY add_4429_13 (.CI(n46838), .I0(n13559[10]), .I1(n889), .CO(n46839));
    SB_LUT4 add_4429_12_lut (.I0(GND_net), .I1(n13559[9]), .I2(n816), 
            .I3(n46837), .O(n12802[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4429_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4429_12 (.CI(n46837), .I0(n13559[9]), .I1(n816), .CO(n46838));
    SB_LUT4 add_4429_11_lut (.I0(GND_net), .I1(n13559[8]), .I2(n743), 
            .I3(n46836), .O(n12802[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4429_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4429_11 (.CI(n46836), .I0(n13559[8]), .I1(n743), .CO(n46837));
    SB_LUT4 add_4429_10_lut (.I0(GND_net), .I1(n13559[7]), .I2(n670), 
            .I3(n46835), .O(n12802[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4429_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4429_10 (.CI(n46835), .I0(n13559[7]), .I1(n670), .CO(n46836));
    SB_LUT4 add_4429_9_lut (.I0(GND_net), .I1(n13559[6]), .I2(n597), .I3(n46834), 
            .O(n12802[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4429_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4429_9 (.CI(n46834), .I0(n13559[6]), .I1(n597), .CO(n46835));
    SB_LUT4 add_4429_8_lut (.I0(GND_net), .I1(n13559[5]), .I2(n524), .I3(n46833), 
            .O(n12802[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4429_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4429_8 (.CI(n46833), .I0(n13559[5]), .I1(n524), .CO(n46834));
    SB_LUT4 add_4429_7_lut (.I0(GND_net), .I1(n13559[4]), .I2(n451_adj_4355), 
            .I3(n46832), .O(n12802[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4429_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4429_7 (.CI(n46832), .I0(n13559[4]), .I1(n451_adj_4355), 
            .CO(n46833));
    SB_LUT4 add_4429_6_lut (.I0(GND_net), .I1(n13559[3]), .I2(n378), .I3(n46831), 
            .O(n12802[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4429_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4429_6 (.CI(n46831), .I0(n13559[3]), .I1(n378), .CO(n46832));
    SB_LUT4 add_4429_5_lut (.I0(GND_net), .I1(n13559[2]), .I2(n305_adj_4356), 
            .I3(n46830), .O(n12802[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4429_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4429_5 (.CI(n46830), .I0(n13559[2]), .I1(n305_adj_4356), 
            .CO(n46831));
    SB_LUT4 add_4429_4_lut (.I0(GND_net), .I1(n13559[1]), .I2(n232), .I3(n46829), 
            .O(n12802[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4429_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4429_4 (.CI(n46829), .I0(n13559[1]), .I1(n232), .CO(n46830));
    SB_LUT4 add_4429_3_lut (.I0(GND_net), .I1(n13559[0]), .I2(n159), .I3(n46828), 
            .O(n12802[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4429_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4429_3 (.CI(n46828), .I0(n13559[0]), .I1(n159), .CO(n46829));
    SB_LUT4 add_4429_2_lut (.I0(GND_net), .I1(n17_adj_4357), .I2(n86), 
            .I3(GND_net), .O(n12802[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4429_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4429_2 (.CI(GND_net), .I0(n17_adj_4357), .I1(n86), .CO(n46828));
    SB_LUT4 add_4466_19_lut (.I0(GND_net), .I1(n14240[16]), .I2(GND_net), 
            .I3(n46827), .O(n13559[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4466_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4466_18_lut (.I0(GND_net), .I1(n14240[15]), .I2(GND_net), 
            .I3(n46826), .O(n13559[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4466_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4466_18 (.CI(n46826), .I0(n14240[15]), .I1(GND_net), 
            .CO(n46827));
    SB_LUT4 add_4466_17_lut (.I0(GND_net), .I1(n14240[14]), .I2(GND_net), 
            .I3(n46825), .O(n13559[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4466_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4466_17 (.CI(n46825), .I0(n14240[14]), .I1(GND_net), 
            .CO(n46826));
    SB_LUT4 add_4466_16_lut (.I0(GND_net), .I1(n14240[13]), .I2(n1111_adj_4358), 
            .I3(n46824), .O(n13559[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4466_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4466_16 (.CI(n46824), .I0(n14240[13]), .I1(n1111_adj_4358), 
            .CO(n46825));
    SB_LUT4 add_4466_15_lut (.I0(GND_net), .I1(n14240[12]), .I2(n1038_adj_4359), 
            .I3(n46823), .O(n13559[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4466_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4466_15 (.CI(n46823), .I0(n14240[12]), .I1(n1038_adj_4359), 
            .CO(n46824));
    SB_LUT4 add_4466_14_lut (.I0(GND_net), .I1(n14240[11]), .I2(n965_adj_4360), 
            .I3(n46822), .O(n13559[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4466_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4466_14 (.CI(n46822), .I0(n14240[11]), .I1(n965_adj_4360), 
            .CO(n46823));
    SB_LUT4 add_4466_13_lut (.I0(GND_net), .I1(n14240[10]), .I2(n892_adj_4361), 
            .I3(n46821), .O(n13559[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4466_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_24_i463_2_lut (.I0(\Ki[9] ), .I1(n349), .I2(GND_net), 
            .I3(GND_net), .O(n688));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i463_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_4466_13 (.CI(n46821), .I0(n14240[10]), .I1(n892_adj_4361), 
            .CO(n46822));
    SB_LUT4 add_4466_12_lut (.I0(GND_net), .I1(n14240[9]), .I2(n819_adj_4362), 
            .I3(n46820), .O(n13559[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4466_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4466_12 (.CI(n46820), .I0(n14240[9]), .I1(n819_adj_4362), 
            .CO(n46821));
    SB_LUT4 add_4466_11_lut (.I0(GND_net), .I1(n14240[8]), .I2(n746_adj_4363), 
            .I3(n46819), .O(n13559[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4466_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4466_11 (.CI(n46819), .I0(n14240[8]), .I1(n746_adj_4363), 
            .CO(n46820));
    SB_LUT4 add_4466_10_lut (.I0(GND_net), .I1(n14240[7]), .I2(n673_adj_4364), 
            .I3(n46818), .O(n13559[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4466_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4466_10 (.CI(n46818), .I0(n14240[7]), .I1(n673_adj_4364), 
            .CO(n46819));
    SB_LUT4 add_4466_9_lut (.I0(GND_net), .I1(n14240[6]), .I2(n600_adj_4365), 
            .I3(n46817), .O(n13559[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4466_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_24_i512_2_lut (.I0(\Ki[10] ), .I1(n349), .I2(GND_net), 
            .I3(GND_net), .O(n761));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i512_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_4466_9 (.CI(n46817), .I0(n14240[6]), .I1(n600_adj_4365), 
            .CO(n46818));
    SB_LUT4 add_4466_8_lut (.I0(GND_net), .I1(n14240[5]), .I2(n527_adj_4366), 
            .I3(n46816), .O(n13559[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4466_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4466_8 (.CI(n46816), .I0(n14240[5]), .I1(n527_adj_4366), 
            .CO(n46817));
    SB_LUT4 add_4466_7_lut (.I0(GND_net), .I1(n14240[4]), .I2(n454_adj_4367), 
            .I3(n46815), .O(n13559[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4466_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4466_7 (.CI(n46815), .I0(n14240[4]), .I1(n454_adj_4367), 
            .CO(n46816));
    SB_LUT4 add_4466_6_lut (.I0(GND_net), .I1(n14240[3]), .I2(n381_adj_4368), 
            .I3(n46814), .O(n13559[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4466_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4466_6 (.CI(n46814), .I0(n14240[3]), .I1(n381_adj_4368), 
            .CO(n46815));
    SB_LUT4 add_4466_5_lut (.I0(GND_net), .I1(n14240[2]), .I2(n308_adj_4369), 
            .I3(n46813), .O(n13559[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4466_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4466_5 (.CI(n46813), .I0(n14240[2]), .I1(n308_adj_4369), 
            .CO(n46814));
    SB_LUT4 add_4466_4_lut (.I0(GND_net), .I1(n14240[1]), .I2(n235_adj_4370), 
            .I3(n46812), .O(n13559[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4466_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4466_4 (.CI(n46812), .I0(n14240[1]), .I1(n235_adj_4370), 
            .CO(n46813));
    SB_LUT4 add_4466_3_lut (.I0(GND_net), .I1(n14240[0]), .I2(n162_adj_4371), 
            .I3(n46811), .O(n13559[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4466_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4466_3 (.CI(n46811), .I0(n14240[0]), .I1(n162_adj_4371), 
            .CO(n46812));
    SB_LUT4 add_4466_2_lut (.I0(GND_net), .I1(n20_adj_4372), .I2(n89_adj_4373), 
            .I3(GND_net), .O(n13559[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4466_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4466_2 (.CI(GND_net), .I0(n20_adj_4372), .I1(n89_adj_4373), 
            .CO(n46811));
    SB_LUT4 add_4698_11_lut (.I0(GND_net), .I1(n17509[8]), .I2(n770), 
            .I3(n46810), .O(n17311[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4698_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4698_10_lut (.I0(GND_net), .I1(n17509[7]), .I2(n697), 
            .I3(n46809), .O(n17311[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4698_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_25_20_lut (.I0(GND_net), .I1(n360[18]), .I2(n42[18]), 
            .I3(n46090), .O(n455[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_25_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_25_20 (.CI(n46090), .I0(n360[18]), .I1(n42[18]), .CO(n46091));
    SB_LUT4 add_25_19_lut (.I0(GND_net), .I1(n360[17]), .I2(n42[17]), 
            .I3(n46089), .O(n455[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_25_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_25_19 (.CI(n46089), .I0(n360[17]), .I1(n42[17]), .CO(n46090));
    SB_LUT4 sub_15_add_2_25_lut (.I0(GND_net), .I1(setpoint[23]), .I2(\motor_state[23] ), 
            .I3(n46241), .O(n207[23])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_15_add_2_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_15_add_2_24_lut (.I0(GND_net), .I1(setpoint[22]), .I2(\motor_state[22] ), 
            .I3(n46240), .O(n207[22])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_15_add_2_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_15_add_2_24 (.CI(n46240), .I0(setpoint[22]), .I1(\motor_state[22] ), 
            .CO(n46241));
    SB_LUT4 add_25_18_lut (.I0(GND_net), .I1(n360[16]), .I2(n42[16]), 
            .I3(n46088), .O(n455[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_25_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4698_10 (.CI(n46809), .I0(n17509[7]), .I1(n697), .CO(n46810));
    SB_LUT4 add_4698_9_lut (.I0(GND_net), .I1(n17509[6]), .I2(n624), .I3(n46808), 
            .O(n17311[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4698_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4698_9 (.CI(n46808), .I0(n17509[6]), .I1(n624), .CO(n46809));
    SB_LUT4 add_4698_8_lut (.I0(GND_net), .I1(n17509[5]), .I2(n551_adj_4375), 
            .I3(n46807), .O(n17311[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4698_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_15_add_2_23_lut (.I0(GND_net), .I1(setpoint[21]), .I2(\motor_state[21] ), 
            .I3(n46239), .O(n207[21])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_15_add_2_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_15_add_2_23 (.CI(n46239), .I0(setpoint[21]), .I1(\motor_state[21] ), 
            .CO(n46240));
    SB_CARRY add_25_18 (.CI(n46088), .I0(n360[16]), .I1(n42[16]), .CO(n46089));
    SB_LUT4 add_4690_11_lut (.I0(GND_net), .I1(n17432[8]), .I2(n770_adj_4376), 
            .I3(n47175), .O(n17215[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4690_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4690_10_lut (.I0(GND_net), .I1(n17432[7]), .I2(n697_adj_4377), 
            .I3(n47174), .O(n17215[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4690_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4698_8 (.CI(n46807), .I0(n17509[5]), .I1(n551_adj_4375), 
            .CO(n46808));
    SB_LUT4 add_4698_7_lut (.I0(GND_net), .I1(n17509[4]), .I2(n478), .I3(n46806), 
            .O(n17311[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4698_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4690_10 (.CI(n47174), .I0(n17432[7]), .I1(n697_adj_4377), 
            .CO(n47175));
    SB_LUT4 add_4690_9_lut (.I0(GND_net), .I1(n17432[6]), .I2(n624_adj_4378), 
            .I3(n47173), .O(n17215[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4690_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4698_7 (.CI(n46806), .I0(n17509[4]), .I1(n478), .CO(n46807));
    SB_LUT4 sub_15_add_2_22_lut (.I0(GND_net), .I1(setpoint[20]), .I2(\motor_state[20] ), 
            .I3(n46238), .O(n207[20])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_15_add_2_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_15_add_2_22 (.CI(n46238), .I0(setpoint[20]), .I1(\motor_state[20] ), 
            .CO(n46239));
    SB_LUT4 sub_15_add_2_21_lut (.I0(GND_net), .I1(setpoint[19]), .I2(\motor_state[19] ), 
            .I3(n46237), .O(n207[19])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_15_add_2_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_15_add_2_21 (.CI(n46237), .I0(setpoint[19]), .I1(\motor_state[19] ), 
            .CO(n46238));
    SB_CARRY add_4690_9 (.CI(n47173), .I0(n17432[6]), .I1(n624_adj_4378), 
            .CO(n47174));
    SB_LUT4 add_25_17_lut (.I0(GND_net), .I1(n360[15]), .I2(n42[15]), 
            .I3(n46087), .O(n455[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_25_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_15_add_2_20_lut (.I0(GND_net), .I1(setpoint[18]), .I2(\motor_state[18] ), 
            .I3(n46236), .O(n207[18])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_15_add_2_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_15_add_2_20 (.CI(n46236), .I0(setpoint[18]), .I1(\motor_state[18] ), 
            .CO(n46237));
    SB_LUT4 add_4690_8_lut (.I0(GND_net), .I1(n17432[5]), .I2(n551_adj_4379), 
            .I3(n47172), .O(n17215[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4690_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_25_17 (.CI(n46087), .I0(n360[15]), .I1(n42[15]), .CO(n46088));
    SB_CARRY add_4690_8 (.CI(n47172), .I0(n17432[5]), .I1(n551_adj_4379), 
            .CO(n47173));
    SB_LUT4 add_4690_7_lut (.I0(GND_net), .I1(n17432[4]), .I2(n478_adj_4380), 
            .I3(n47171), .O(n17215[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4690_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4698_6_lut (.I0(GND_net), .I1(n17509[3]), .I2(n405), .I3(n46805), 
            .O(n17311[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4698_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4690_7 (.CI(n47171), .I0(n17432[4]), .I1(n478_adj_4380), 
            .CO(n47172));
    SB_LUT4 add_4690_6_lut (.I0(GND_net), .I1(n17432[3]), .I2(n405_adj_4381), 
            .I3(n47170), .O(n17215[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4690_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4698_6 (.CI(n46805), .I0(n17509[3]), .I1(n405), .CO(n46806));
    SB_LUT4 add_4698_5_lut (.I0(GND_net), .I1(n17509[2]), .I2(n332), .I3(n46804), 
            .O(n17311[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4698_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4690_6 (.CI(n47170), .I0(n17432[3]), .I1(n405_adj_4381), 
            .CO(n47171));
    SB_LUT4 add_4690_5_lut (.I0(GND_net), .I1(n17432[2]), .I2(n332_adj_4382), 
            .I3(n47169), .O(n17215[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4690_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4690_5 (.CI(n47169), .I0(n17432[2]), .I1(n332_adj_4382), 
            .CO(n47170));
    SB_CARRY add_4698_5 (.CI(n46804), .I0(n17509[2]), .I1(n332), .CO(n46805));
    SB_LUT4 add_4698_4_lut (.I0(GND_net), .I1(n17509[1]), .I2(n259), .I3(n46803), 
            .O(n17311[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4698_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4690_4_lut (.I0(GND_net), .I1(n17432[1]), .I2(n259_adj_4383), 
            .I3(n47168), .O(n17215[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4690_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4690_4 (.CI(n47168), .I0(n17432[1]), .I1(n259_adj_4383), 
            .CO(n47169));
    SB_CARRY add_4698_4 (.CI(n46803), .I0(n17509[1]), .I1(n259), .CO(n46804));
    SB_LUT4 add_4690_3_lut (.I0(GND_net), .I1(n17432[0]), .I2(n186), .I3(n47167), 
            .O(n17215[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4690_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_15_add_2_19_lut (.I0(GND_net), .I1(setpoint[17]), .I2(\motor_state[17] ), 
            .I3(n46235), .O(n207[17])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_15_add_2_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_15_add_2_19 (.CI(n46235), .I0(setpoint[17]), .I1(\motor_state[17] ), 
            .CO(n46236));
    SB_LUT4 sub_15_add_2_18_lut (.I0(GND_net), .I1(setpoint[16]), .I2(\motor_state[16] ), 
            .I3(n46234), .O(n207[16])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_15_add_2_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_15_add_2_18 (.CI(n46234), .I0(setpoint[16]), .I1(\motor_state[16] ), 
            .CO(n46235));
    SB_CARRY add_4690_3 (.CI(n47167), .I0(n17432[0]), .I1(n186), .CO(n47168));
    SB_LUT4 sub_15_add_2_17_lut (.I0(GND_net), .I1(setpoint[15]), .I2(\motor_state[15] ), 
            .I3(n46233), .O(n207[15])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_15_add_2_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_15_add_2_17 (.CI(n46233), .I0(setpoint[15]), .I1(\motor_state[15] ), 
            .CO(n46234));
    SB_LUT4 sub_15_add_2_16_lut (.I0(GND_net), .I1(setpoint[14]), .I2(\motor_state[14] ), 
            .I3(n46232), .O(n207[14])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_15_add_2_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_15_add_2_16 (.CI(n46232), .I0(setpoint[14]), .I1(\motor_state[14] ), 
            .CO(n46233));
    SB_LUT4 add_4698_3_lut (.I0(GND_net), .I1(n17509[0]), .I2(n186_adj_4384), 
            .I3(n46802), .O(n17311[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4698_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4690_2_lut (.I0(GND_net), .I1(n44), .I2(n113), .I3(GND_net), 
            .O(n17215[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4690_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4690_2 (.CI(GND_net), .I0(n44), .I1(n113), .CO(n47167));
    SB_CARRY add_4698_3 (.CI(n46802), .I0(n17509[0]), .I1(n186_adj_4384), 
            .CO(n46803));
    SB_LUT4 add_4698_2_lut (.I0(GND_net), .I1(n44_adj_4385), .I2(n113_adj_4386), 
            .I3(GND_net), .O(n17311[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4698_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_23_add_1221_24_lut (.I0(n207[23]), .I1(n10514[21]), .I2(GND_net), 
            .I3(n47166), .O(n10055[0])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_23_add_1221_24_lut.LUT_INIT = 16'h6996;
    SB_LUT4 mult_23_add_1221_23_lut (.I0(GND_net), .I1(n10514[20]), .I2(GND_net), 
            .I3(n47165), .O(n360[22])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_23_add_1221_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4698_2 (.CI(GND_net), .I0(n44_adj_4385), .I1(n113_adj_4386), 
            .CO(n46802));
    SB_LUT4 add_4501_18_lut (.I0(GND_net), .I1(n14849[15]), .I2(GND_net), 
            .I3(n46801), .O(n14240[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4501_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_23_add_1221_23 (.CI(n47165), .I0(n10514[20]), .I1(GND_net), 
            .CO(n47166));
    SB_LUT4 add_25_16_lut (.I0(GND_net), .I1(n360[14]), .I2(n42[14]), 
            .I3(n46086), .O(n455[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_25_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_23_add_1221_22_lut (.I0(GND_net), .I1(n10514[19]), .I2(GND_net), 
            .I3(n47164), .O(n360[21])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_23_add_1221_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_23_add_1221_22 (.CI(n47164), .I0(n10514[19]), .I1(GND_net), 
            .CO(n47165));
    SB_LUT4 add_4501_17_lut (.I0(GND_net), .I1(n14849[14]), .I2(GND_net), 
            .I3(n46800), .O(n14240[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4501_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_15_add_2_15_lut (.I0(GND_net), .I1(setpoint[13]), .I2(\motor_state[13] ), 
            .I3(n46231), .O(n207[13])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_15_add_2_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_15_add_2_15 (.CI(n46231), .I0(setpoint[13]), .I1(\motor_state[13] ), 
            .CO(n46232));
    SB_CARRY add_25_16 (.CI(n46086), .I0(n360[14]), .I1(n42[14]), .CO(n46087));
    SB_LUT4 sub_15_add_2_14_lut (.I0(GND_net), .I1(setpoint[12]), .I2(\motor_state[12] ), 
            .I3(n46230), .O(n207[12])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_15_add_2_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_25_15_lut (.I0(GND_net), .I1(n360[13]), .I2(n42[13]), 
            .I3(n46085), .O(n455[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_25_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_25_15 (.CI(n46085), .I0(n360[13]), .I1(n42[13]), .CO(n46086));
    SB_CARRY add_4501_17 (.CI(n46800), .I0(n14849[14]), .I1(GND_net), 
            .CO(n46801));
    SB_LUT4 add_4501_16_lut (.I0(GND_net), .I1(n14849[13]), .I2(n1114_adj_4388), 
            .I3(n46799), .O(n14240[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4501_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_23_add_1221_21_lut (.I0(GND_net), .I1(n10514[18]), .I2(GND_net), 
            .I3(n47163), .O(n360[20])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_23_add_1221_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_23_add_1221_21 (.CI(n47163), .I0(n10514[18]), .I1(GND_net), 
            .CO(n47164));
    SB_CARRY add_4501_16 (.CI(n46799), .I0(n14849[13]), .I1(n1114_adj_4388), 
            .CO(n46800));
    SB_LUT4 add_4501_15_lut (.I0(GND_net), .I1(n14849[12]), .I2(n1041_adj_4389), 
            .I3(n46798), .O(n14240[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4501_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_23_add_1221_20_lut (.I0(GND_net), .I1(n10514[17]), .I2(GND_net), 
            .I3(n47162), .O(n360[19])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_23_add_1221_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_23_add_1221_20 (.CI(n47162), .I0(n10514[17]), .I1(GND_net), 
            .CO(n47163));
    SB_CARRY add_4501_15 (.CI(n46798), .I0(n14849[12]), .I1(n1041_adj_4389), 
            .CO(n46799));
    SB_LUT4 add_4501_14_lut (.I0(GND_net), .I1(n14849[11]), .I2(n968_adj_4390), 
            .I3(n46797), .O(n14240[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4501_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_23_add_1221_19_lut (.I0(GND_net), .I1(n10514[16]), .I2(GND_net), 
            .I3(n47161), .O(n360[18])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_23_add_1221_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_15_add_2_14 (.CI(n46230), .I0(setpoint[12]), .I1(\motor_state[12] ), 
            .CO(n46231));
    SB_LUT4 sub_15_add_2_13_lut (.I0(GND_net), .I1(setpoint[11]), .I2(n35211), 
            .I3(n46229), .O(n207[11])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_15_add_2_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_23_add_1221_19 (.CI(n47161), .I0(n10514[16]), .I1(GND_net), 
            .CO(n47162));
    SB_LUT4 mult_23_add_1221_18_lut (.I0(GND_net), .I1(n10514[15]), .I2(GND_net), 
            .I3(n47160), .O(n360[17])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_23_add_1221_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_15_add_2_13 (.CI(n46229), .I0(setpoint[11]), .I1(n35211), 
            .CO(n46230));
    SB_LUT4 sub_15_add_2_12_lut (.I0(GND_net), .I1(setpoint[10]), .I2(\motor_state[10] ), 
            .I3(n46228), .O(n207[10])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_15_add_2_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_15_add_2_12 (.CI(n46228), .I0(setpoint[10]), .I1(\motor_state[10] ), 
            .CO(n46229));
    SB_LUT4 sub_15_add_2_11_lut (.I0(GND_net), .I1(setpoint[9]), .I2(\motor_state[9] ), 
            .I3(n46227), .O(n207[9])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_15_add_2_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_23_add_1221_18 (.CI(n47160), .I0(n10514[15]), .I1(GND_net), 
            .CO(n47161));
    SB_CARRY sub_15_add_2_11 (.CI(n46227), .I0(setpoint[9]), .I1(\motor_state[9] ), 
            .CO(n46228));
    SB_LUT4 sub_15_add_2_10_lut (.I0(GND_net), .I1(setpoint[8]), .I2(\motor_state[8] ), 
            .I3(n46226), .O(n207[8])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_15_add_2_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_23_add_1221_17_lut (.I0(GND_net), .I1(n10514[14]), .I2(GND_net), 
            .I3(n47159), .O(n360[16])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_23_add_1221_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_23_add_1221_17 (.CI(n47159), .I0(n10514[14]), .I1(GND_net), 
            .CO(n47160));
    SB_LUT4 mult_23_add_1221_16_lut (.I0(GND_net), .I1(n10514[13]), .I2(n1096_adj_4391), 
            .I3(n47158), .O(n360[15])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_23_add_1221_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4501_14 (.CI(n46797), .I0(n14849[11]), .I1(n968_adj_4390), 
            .CO(n46798));
    SB_LUT4 add_4501_13_lut (.I0(GND_net), .I1(n14849[10]), .I2(n895_adj_4392), 
            .I3(n46796), .O(n14240[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4501_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_23_add_1221_16 (.CI(n47158), .I0(n10514[13]), .I1(n1096_adj_4391), 
            .CO(n47159));
    SB_LUT4 mult_23_add_1221_15_lut (.I0(GND_net), .I1(n10514[12]), .I2(n1023_adj_4393), 
            .I3(n47157), .O(n360[14])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_23_add_1221_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4501_13 (.CI(n46796), .I0(n14849[10]), .I1(n895_adj_4392), 
            .CO(n46797));
    SB_LUT4 add_4501_12_lut (.I0(GND_net), .I1(n14849[9]), .I2(n822_adj_4394), 
            .I3(n46795), .O(n14240[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4501_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_23_add_1221_15 (.CI(n47157), .I0(n10514[12]), .I1(n1023_adj_4393), 
            .CO(n47158));
    SB_LUT4 mult_23_add_1221_14_lut (.I0(GND_net), .I1(n10514[11]), .I2(n950_adj_4395), 
            .I3(n47156), .O(n360[13])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_23_add_1221_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4501_12 (.CI(n46795), .I0(n14849[9]), .I1(n822_adj_4394), 
            .CO(n46796));
    SB_CARRY mult_23_add_1221_14 (.CI(n47156), .I0(n10514[11]), .I1(n950_adj_4395), 
            .CO(n47157));
    SB_LUT4 mult_23_add_1221_13_lut (.I0(GND_net), .I1(n10514[10]), .I2(n877_adj_4396), 
            .I3(n47155), .O(n360[12])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_23_add_1221_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4501_11_lut (.I0(GND_net), .I1(n14849[8]), .I2(n749_adj_4397), 
            .I3(n46794), .O(n14240[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4501_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_15_add_2_10 (.CI(n46226), .I0(setpoint[8]), .I1(\motor_state[8] ), 
            .CO(n46227));
    SB_CARRY mult_23_add_1221_13 (.CI(n47155), .I0(n10514[10]), .I1(n877_adj_4396), 
            .CO(n47156));
    SB_LUT4 sub_15_add_2_9_lut (.I0(GND_net), .I1(setpoint[7]), .I2(\motor_state[7] ), 
            .I3(n46225), .O(n207[7])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_15_add_2_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_23_add_1221_12_lut (.I0(GND_net), .I1(n10514[9]), .I2(n804_adj_4399), 
            .I3(n47154), .O(n360[11])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_23_add_1221_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_15_add_2_9 (.CI(n46225), .I0(setpoint[7]), .I1(\motor_state[7] ), 
            .CO(n46226));
    SB_CARRY mult_23_add_1221_12 (.CI(n47154), .I0(n10514[9]), .I1(n804_adj_4399), 
            .CO(n47155));
    SB_LUT4 sub_15_add_2_8_lut (.I0(GND_net), .I1(setpoint[6]), .I2(n33792), 
            .I3(n46224), .O(n207[6])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_15_add_2_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_23_add_1221_11_lut (.I0(GND_net), .I1(n10514[8]), .I2(n731_adj_4400), 
            .I3(n47153), .O(n360[10])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_23_add_1221_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_15_add_2_8 (.CI(n46224), .I0(setpoint[6]), .I1(n33792), 
            .CO(n46225));
    SB_LUT4 sub_15_add_2_7_lut (.I0(GND_net), .I1(setpoint[5]), .I2(\motor_state[5] ), 
            .I3(n46223), .O(n207[5])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_15_add_2_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_23_add_1221_11 (.CI(n47153), .I0(n10514[8]), .I1(n731_adj_4400), 
            .CO(n47154));
    SB_CARRY sub_15_add_2_7 (.CI(n46223), .I0(setpoint[5]), .I1(\motor_state[5] ), 
            .CO(n46224));
    SB_LUT4 sub_15_add_2_6_lut (.I0(GND_net), .I1(setpoint[4]), .I2(\motor_state[4] ), 
            .I3(n46222), .O(n207[4])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_15_add_2_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_15_add_2_6 (.CI(n46222), .I0(setpoint[4]), .I1(\motor_state[4] ), 
            .CO(n46223));
    SB_CARRY sub_15_add_2_5 (.CI(n46221), .I0(setpoint[3]), .I1(\motor_state[3] ), 
            .CO(n46222));
    SB_CARRY sub_15_add_2_4 (.CI(n46220), .I0(setpoint[2]), .I1(\motor_state[2] ), 
            .CO(n46221));
    SB_LUT4 mult_23_add_1221_10_lut (.I0(GND_net), .I1(n10514[7]), .I2(n658_adj_4401), 
            .I3(n47152), .O(n360[9])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_23_add_1221_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_23_add_1221_10 (.CI(n47152), .I0(n10514[7]), .I1(n658_adj_4401), 
            .CO(n47153));
    SB_LUT4 mult_23_add_1221_9_lut (.I0(GND_net), .I1(n10514[6]), .I2(n585_adj_4403), 
            .I3(n47151), .O(n360[8])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_23_add_1221_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4501_11 (.CI(n46794), .I0(n14849[8]), .I1(n749_adj_4397), 
            .CO(n46795));
    SB_LUT4 add_4501_10_lut (.I0(GND_net), .I1(n14849[7]), .I2(n676_adj_4404), 
            .I3(n46793), .O(n14240[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4501_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_23_add_1221_9 (.CI(n47151), .I0(n10514[6]), .I1(n585_adj_4403), 
            .CO(n47152));
    SB_LUT4 mult_23_add_1221_8_lut (.I0(GND_net), .I1(n10514[5]), .I2(n512_adj_4405), 
            .I3(n47150), .O(n360[7])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_23_add_1221_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_25_14_lut (.I0(GND_net), .I1(n360[12]), .I2(n42[12]), 
            .I3(n46084), .O(n455[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_25_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4501_10 (.CI(n46793), .I0(n14849[7]), .I1(n676_adj_4404), 
            .CO(n46794));
    SB_LUT4 add_4501_9_lut (.I0(GND_net), .I1(n14849[6]), .I2(n603_adj_4406), 
            .I3(n46792), .O(n14240[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4501_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_15_add_2_3 (.CI(n46219), .I0(setpoint[1]), .I1(n1), .CO(n46220));
    SB_CARRY sub_15_add_2_2 (.CI(VCC_net), .I0(setpoint[0]), .I1(\motor_state[0] ), 
            .CO(n46219));
    SB_CARRY mult_23_add_1221_8 (.CI(n47150), .I0(n10514[5]), .I1(n512_adj_4405), 
            .CO(n47151));
    SB_LUT4 unary_minus_33_add_3_25_lut (.I0(GND_net), .I1(GND_net), .I2(n46[23]), 
            .I3(n46218), .O(n535[23])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_33_add_3_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_23_add_1221_7_lut (.I0(GND_net), .I1(n10514[4]), .I2(n439_adj_4409), 
            .I3(n47149), .O(n360[6])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_23_add_1221_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_33_add_3_24_lut (.I0(GND_net), .I1(GND_net), .I2(n46[22]), 
            .I3(n46217), .O(n535[22])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_33_add_3_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_23_add_1221_7 (.CI(n47149), .I0(n10514[4]), .I1(n439_adj_4409), 
            .CO(n47150));
    SB_LUT4 mult_23_add_1221_6_lut (.I0(GND_net), .I1(n10514[3]), .I2(n366_adj_4412), 
            .I3(n47148), .O(n360[5])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_23_add_1221_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4501_9 (.CI(n46792), .I0(n14849[6]), .I1(n603_adj_4406), 
            .CO(n46793));
    SB_CARRY mult_23_add_1221_6 (.CI(n47148), .I0(n10514[3]), .I1(n366_adj_4412), 
            .CO(n47149));
    SB_LUT4 mult_23_add_1221_5_lut (.I0(GND_net), .I1(n10514[2]), .I2(n293_adj_4413), 
            .I3(n47147), .O(n360[4])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_23_add_1221_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4501_8_lut (.I0(GND_net), .I1(n14849[5]), .I2(n530_adj_4414), 
            .I3(n46791), .O(n14240[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4501_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_33_add_3_24 (.CI(n46217), .I0(GND_net), .I1(n46[22]), 
            .CO(n46218));
    SB_CARRY mult_23_add_1221_5 (.CI(n47147), .I0(n10514[2]), .I1(n293_adj_4413), 
            .CO(n47148));
    SB_LUT4 mult_23_add_1221_4_lut (.I0(GND_net), .I1(n10514[1]), .I2(n220_adj_4415), 
            .I3(n47146), .O(n360[3])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_23_add_1221_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_23_add_1221_4 (.CI(n47146), .I0(n10514[1]), .I1(n220_adj_4415), 
            .CO(n47147));
    SB_LUT4 unary_minus_33_add_3_23_lut (.I0(GND_net), .I1(GND_net), .I2(n46[21]), 
            .I3(n46216), .O(n535[21])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_33_add_3_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_23_add_1221_3_lut (.I0(GND_net), .I1(n10514[0]), .I2(n147_adj_4418), 
            .I3(n47145), .O(n360[2])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_23_add_1221_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4501_8 (.CI(n46791), .I0(n14849[5]), .I1(n530_adj_4414), 
            .CO(n46792));
    SB_LUT4 add_4501_7_lut (.I0(GND_net), .I1(n14849[4]), .I2(n457_adj_4419), 
            .I3(n46790), .O(n14240[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4501_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_23_add_1221_3 (.CI(n47145), .I0(n10514[0]), .I1(n147_adj_4418), 
            .CO(n47146));
    SB_LUT4 mult_23_add_1221_2_lut (.I0(GND_net), .I1(n5_adj_4420), .I2(n74_adj_4421), 
            .I3(GND_net), .O(n360[1])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_23_add_1221_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4501_7 (.CI(n46790), .I0(n14849[4]), .I1(n457_adj_4419), 
            .CO(n46791));
    SB_LUT4 add_4501_6_lut (.I0(GND_net), .I1(n14849[3]), .I2(n384_adj_4422), 
            .I3(n46789), .O(n14240[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4501_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_23_add_1221_2 (.CI(GND_net), .I0(n5_adj_4420), .I1(n74_adj_4421), 
            .CO(n47145));
    SB_CARRY unary_minus_33_add_3_23 (.CI(n46216), .I0(GND_net), .I1(n46[21]), 
            .CO(n46217));
    SB_LUT4 unary_minus_33_add_3_22_lut (.I0(GND_net), .I1(GND_net), .I2(n46[20]), 
            .I3(n46215), .O(n535[20])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_33_add_3_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_33_add_3_22 (.CI(n46215), .I0(GND_net), .I1(n46[20]), 
            .CO(n46216));
    SB_LUT4 unary_minus_33_add_3_21_lut (.I0(GND_net), .I1(GND_net), .I2(n46[19]), 
            .I3(n46214), .O(n535[19])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_33_add_3_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_33_add_3_21 (.CI(n46214), .I0(GND_net), .I1(n46[19]), 
            .CO(n46215));
    SB_LUT4 unary_minus_33_add_3_20_lut (.I0(GND_net), .I1(GND_net), .I2(n46[18]), 
            .I3(n46213), .O(n535[18])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_33_add_3_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_33_add_3_20 (.CI(n46213), .I0(GND_net), .I1(n46[18]), 
            .CO(n46214));
    SB_LUT4 unary_minus_33_add_3_19_lut (.I0(GND_net), .I1(GND_net), .I2(n46[17]), 
            .I3(n46212), .O(n535[17])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_33_add_3_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_25_14 (.CI(n46084), .I0(n360[12]), .I1(n42[12]), .CO(n46085));
    SB_LUT4 add_25_13_lut (.I0(GND_net), .I1(n360[11]), .I2(n42[11]), 
            .I3(n46083), .O(n455[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_25_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_25_13 (.CI(n46083), .I0(n360[11]), .I1(n42[11]), .CO(n46084));
    SB_CARRY unary_minus_33_add_3_19 (.CI(n46212), .I0(GND_net), .I1(n46[17]), 
            .CO(n46213));
    SB_LUT4 unary_minus_33_add_3_18_lut (.I0(GND_net), .I1(GND_net), .I2(n46[16]), 
            .I3(n46211), .O(n535[16])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_33_add_3_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_33_add_3_18 (.CI(n46211), .I0(GND_net), .I1(n46[16]), 
            .CO(n46212));
    SB_LUT4 add_25_12_lut (.I0(GND_net), .I1(n360[10]), .I2(n42[10]), 
            .I3(n46082), .O(n455[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_25_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4325_23_lut (.I0(GND_net), .I1(n11481[20]), .I2(GND_net), 
            .I3(n47144), .O(n10514[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4325_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_25_12 (.CI(n46082), .I0(n360[10]), .I1(n42[10]), .CO(n46083));
    SB_LUT4 add_25_11_lut (.I0(GND_net), .I1(n360[9]), .I2(n42[9]), .I3(n46081), 
            .O(n455[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_25_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_33_add_3_17_lut (.I0(GND_net), .I1(GND_net), .I2(n46[15]), 
            .I3(n46210), .O(n535[15])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_33_add_3_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4325_22_lut (.I0(GND_net), .I1(n11481[19]), .I2(GND_net), 
            .I3(n47143), .O(n10514[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4325_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4325_22 (.CI(n47143), .I0(n11481[19]), .I1(GND_net), 
            .CO(n47144));
    SB_CARRY add_4501_6 (.CI(n46789), .I0(n14849[3]), .I1(n384_adj_4422), 
            .CO(n46790));
    SB_LUT4 add_4501_5_lut (.I0(GND_net), .I1(n14849[2]), .I2(n311_adj_4429), 
            .I3(n46788), .O(n14240[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4501_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4325_21_lut (.I0(GND_net), .I1(n11481[18]), .I2(GND_net), 
            .I3(n47142), .O(n10514[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4325_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4325_21 (.CI(n47142), .I0(n11481[18]), .I1(GND_net), 
            .CO(n47143));
    SB_CARRY add_4501_5 (.CI(n46788), .I0(n14849[2]), .I1(n311_adj_4429), 
            .CO(n46789));
    SB_LUT4 add_4501_4_lut (.I0(GND_net), .I1(n14849[1]), .I2(n238_adj_4430), 
            .I3(n46787), .O(n14240[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4501_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4325_20_lut (.I0(GND_net), .I1(n11481[17]), .I2(GND_net), 
            .I3(n47141), .O(n10514[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4325_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4325_20 (.CI(n47141), .I0(n11481[17]), .I1(GND_net), 
            .CO(n47142));
    SB_CARRY add_4501_4 (.CI(n46787), .I0(n14849[1]), .I1(n238_adj_4430), 
            .CO(n46788));
    SB_LUT4 add_4501_3_lut (.I0(GND_net), .I1(n14849[0]), .I2(n165_adj_4431), 
            .I3(n46786), .O(n14240[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4501_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4325_19_lut (.I0(GND_net), .I1(n11481[16]), .I2(GND_net), 
            .I3(n47140), .O(n10514[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4325_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4325_19 (.CI(n47140), .I0(n11481[16]), .I1(GND_net), 
            .CO(n47141));
    SB_LUT4 add_4325_18_lut (.I0(GND_net), .I1(n11481[15]), .I2(GND_net), 
            .I3(n47139), .O(n10514[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4325_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4501_3 (.CI(n46786), .I0(n14849[0]), .I1(n165_adj_4431), 
            .CO(n46787));
    SB_LUT4 add_4501_2_lut (.I0(GND_net), .I1(n23_adj_4432), .I2(n92_adj_4433), 
            .I3(GND_net), .O(n14240[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4501_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4325_18 (.CI(n47139), .I0(n11481[15]), .I1(GND_net), 
            .CO(n47140));
    SB_LUT4 add_4325_17_lut (.I0(GND_net), .I1(n11481[14]), .I2(GND_net), 
            .I3(n47138), .O(n10514[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4325_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4501_2 (.CI(GND_net), .I0(n23_adj_4432), .I1(n92_adj_4433), 
            .CO(n46786));
    SB_LUT4 add_4534_17_lut (.I0(GND_net), .I1(n15390[14]), .I2(GND_net), 
            .I3(n46785), .O(n14849[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4534_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4325_17 (.CI(n47138), .I0(n11481[14]), .I1(GND_net), 
            .CO(n47139));
    SB_LUT4 add_4325_16_lut (.I0(GND_net), .I1(n11481[13]), .I2(n1099_adj_4434), 
            .I3(n47137), .O(n10514[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4325_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_33_add_3_17 (.CI(n46210), .I0(GND_net), .I1(n46[15]), 
            .CO(n46211));
    SB_LUT4 unary_minus_33_add_3_16_lut (.I0(GND_net), .I1(GND_net), .I2(n46[14]), 
            .I3(n46209), .O(n535[14])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_33_add_3_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_33_add_3_16 (.CI(n46209), .I0(GND_net), .I1(n46[14]), 
            .CO(n46210));
    SB_CARRY add_25_11 (.CI(n46081), .I0(n360[9]), .I1(n42[9]), .CO(n46082));
    SB_LUT4 unary_minus_33_add_3_15_lut (.I0(GND_net), .I1(GND_net), .I2(n46[13]), 
            .I3(n46208), .O(n535[13])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_33_add_3_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_33_add_3_15 (.CI(n46208), .I0(GND_net), .I1(n46[13]), 
            .CO(n46209));
    SB_LUT4 unary_minus_33_add_3_14_lut (.I0(GND_net), .I1(GND_net), .I2(n46[12]), 
            .I3(n46207), .O(n535[12])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_33_add_3_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_33_add_3_14 (.CI(n46207), .I0(GND_net), .I1(n46[12]), 
            .CO(n46208));
    SB_LUT4 unary_minus_33_add_3_13_lut (.I0(GND_net), .I1(GND_net), .I2(n46[11]), 
            .I3(n46206), .O(n535[11])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_33_add_3_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_25_10_lut (.I0(GND_net), .I1(n360[8]), .I2(n42[8]), .I3(n46080), 
            .O(n455[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_25_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_33_add_3_13 (.CI(n46206), .I0(GND_net), .I1(n46[11]), 
            .CO(n46207));
    SB_CARRY add_25_10 (.CI(n46080), .I0(n360[8]), .I1(n42[8]), .CO(n46081));
    SB_LUT4 add_25_9_lut (.I0(GND_net), .I1(n360[7]), .I2(n42[7]), .I3(n46079), 
            .O(n455[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_25_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4325_16 (.CI(n47137), .I0(n11481[13]), .I1(n1099_adj_4434), 
            .CO(n47138));
    SB_LUT4 add_4325_15_lut (.I0(GND_net), .I1(n11481[12]), .I2(n1026_adj_4439), 
            .I3(n47136), .O(n10514[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4325_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4534_16_lut (.I0(GND_net), .I1(n15390[13]), .I2(n1117_adj_4440), 
            .I3(n46784), .O(n14849[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4534_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4534_16 (.CI(n46784), .I0(n15390[13]), .I1(n1117_adj_4440), 
            .CO(n46785));
    SB_CARRY add_4325_15 (.CI(n47136), .I0(n11481[12]), .I1(n1026_adj_4439), 
            .CO(n47137));
    SB_LUT4 add_4325_14_lut (.I0(GND_net), .I1(n11481[11]), .I2(n953_adj_4441), 
            .I3(n47135), .O(n10514[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4325_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4534_15_lut (.I0(GND_net), .I1(n15390[12]), .I2(n1044_adj_4442), 
            .I3(n46783), .O(n14849[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4534_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4534_15 (.CI(n46783), .I0(n15390[12]), .I1(n1044_adj_4442), 
            .CO(n46784));
    SB_CARRY add_4325_14 (.CI(n47135), .I0(n11481[11]), .I1(n953_adj_4441), 
            .CO(n47136));
    SB_LUT4 add_4325_13_lut (.I0(GND_net), .I1(n11481[10]), .I2(n880_adj_4443), 
            .I3(n47134), .O(n10514[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4325_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_33_add_3_12_lut (.I0(GND_net), .I1(GND_net), .I2(n46[10]), 
            .I3(n46205), .O(n535[10])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_33_add_3_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4534_14_lut (.I0(GND_net), .I1(n15390[11]), .I2(n971_adj_4445), 
            .I3(n46782), .O(n14849[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4534_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4534_14 (.CI(n46782), .I0(n15390[11]), .I1(n971_adj_4445), 
            .CO(n46783));
    SB_CARRY add_4325_13 (.CI(n47134), .I0(n11481[10]), .I1(n880_adj_4443), 
            .CO(n47135));
    SB_LUT4 add_4325_12_lut (.I0(GND_net), .I1(n11481[9]), .I2(n807_adj_4446), 
            .I3(n47133), .O(n10514[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4325_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4534_13_lut (.I0(GND_net), .I1(n15390[10]), .I2(n898_adj_4447), 
            .I3(n46781), .O(n14849[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4534_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4534_13 (.CI(n46781), .I0(n15390[10]), .I1(n898_adj_4447), 
            .CO(n46782));
    SB_CARRY add_4325_12 (.CI(n47133), .I0(n11481[9]), .I1(n807_adj_4446), 
            .CO(n47134));
    SB_LUT4 add_4325_11_lut (.I0(GND_net), .I1(n11481[8]), .I2(n734_adj_4448), 
            .I3(n47132), .O(n10514[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4325_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_25_9 (.CI(n46079), .I0(n360[7]), .I1(n42[7]), .CO(n46080));
    SB_CARRY unary_minus_33_add_3_12 (.CI(n46205), .I0(GND_net), .I1(n46[10]), 
            .CO(n46206));
    SB_LUT4 unary_minus_33_add_3_11_lut (.I0(GND_net), .I1(GND_net), .I2(n46[9]), 
            .I3(n46204), .O(n535[9])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_33_add_3_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4325_11 (.CI(n47132), .I0(n11481[8]), .I1(n734_adj_4448), 
            .CO(n47133));
    SB_CARRY unary_minus_33_add_3_11 (.CI(n46204), .I0(GND_net), .I1(n46[9]), 
            .CO(n46205));
    SB_LUT4 add_4325_10_lut (.I0(GND_net), .I1(n11481[7]), .I2(n661_adj_4450), 
            .I3(n47131), .O(n10514[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4325_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4325_10 (.CI(n47131), .I0(n11481[7]), .I1(n661_adj_4450), 
            .CO(n47132));
    SB_LUT4 unary_minus_33_add_3_10_lut (.I0(GND_net), .I1(GND_net), .I2(n46[8]), 
            .I3(n46203), .O(n535[8])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_33_add_3_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_33_add_3_10 (.CI(n46203), .I0(GND_net), .I1(n46[8]), 
            .CO(n46204));
    SB_LUT4 unary_minus_33_add_3_9_lut (.I0(GND_net), .I1(GND_net), .I2(n46[7]), 
            .I3(n46202), .O(n535[7])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_33_add_3_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_25_8_lut (.I0(GND_net), .I1(n360[6]), .I2(n42[6]), .I3(n46078), 
            .O(n455[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_25_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4325_9_lut (.I0(GND_net), .I1(n11481[6]), .I2(n588_adj_4453), 
            .I3(n47130), .O(n10514[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4325_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4325_9 (.CI(n47130), .I0(n11481[6]), .I1(n588_adj_4453), 
            .CO(n47131));
    SB_LUT4 add_4325_8_lut (.I0(GND_net), .I1(n11481[5]), .I2(n515_adj_4454), 
            .I3(n47129), .O(n10514[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4325_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4325_8 (.CI(n47129), .I0(n11481[5]), .I1(n515_adj_4454), 
            .CO(n47130));
    SB_LUT4 add_4325_7_lut (.I0(GND_net), .I1(n11481[4]), .I2(n442_adj_4455), 
            .I3(n47128), .O(n10514[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4325_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4534_12_lut (.I0(GND_net), .I1(n15390[9]), .I2(n825_adj_4456), 
            .I3(n46780), .O(n14849[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4534_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4534_12 (.CI(n46780), .I0(n15390[9]), .I1(n825_adj_4456), 
            .CO(n46781));
    SB_CARRY add_4325_7 (.CI(n47128), .I0(n11481[4]), .I1(n442_adj_4455), 
            .CO(n47129));
    SB_LUT4 add_4325_6_lut (.I0(GND_net), .I1(n11481[3]), .I2(n369_adj_4457), 
            .I3(n47127), .O(n10514[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4325_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4534_11_lut (.I0(GND_net), .I1(n15390[8]), .I2(n752_adj_4458), 
            .I3(n46779), .O(n14849[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4534_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4534_11 (.CI(n46779), .I0(n15390[8]), .I1(n752_adj_4458), 
            .CO(n46780));
    SB_CARRY add_4325_6 (.CI(n47127), .I0(n11481[3]), .I1(n369_adj_4457), 
            .CO(n47128));
    SB_LUT4 add_4325_5_lut (.I0(GND_net), .I1(n11481[2]), .I2(n296_adj_4459), 
            .I3(n47126), .O(n10514[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4325_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4534_10_lut (.I0(GND_net), .I1(n15390[7]), .I2(n679_adj_4460), 
            .I3(n46778), .O(n14849[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4534_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4534_10 (.CI(n46778), .I0(n15390[7]), .I1(n679_adj_4460), 
            .CO(n46779));
    SB_CARRY add_4325_5 (.CI(n47126), .I0(n11481[2]), .I1(n296_adj_4459), 
            .CO(n47127));
    SB_LUT4 add_4325_4_lut (.I0(GND_net), .I1(n11481[1]), .I2(n223_adj_4461), 
            .I3(n47125), .O(n10514[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4325_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_33_add_3_9 (.CI(n46202), .I0(GND_net), .I1(n46[7]), 
            .CO(n46203));
    SB_CARRY add_25_8 (.CI(n46078), .I0(n360[6]), .I1(n42[6]), .CO(n46079));
    SB_LUT4 add_25_7_lut (.I0(GND_net), .I1(n360[5]), .I2(n42[5]), .I3(n46077), 
            .O(n455[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_25_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_33_add_3_8_lut (.I0(GND_net), .I1(GND_net), .I2(n46[6]), 
            .I3(n46201), .O(n535[6])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_33_add_3_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_33_add_3_8 (.CI(n46201), .I0(GND_net), .I1(n46[6]), 
            .CO(n46202));
    SB_LUT4 unary_minus_33_add_3_7_lut (.I0(GND_net), .I1(GND_net), .I2(n46[5]), 
            .I3(n46200), .O(n535[5])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_33_add_3_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_25_7 (.CI(n46077), .I0(n360[5]), .I1(n42[5]), .CO(n46078));
    SB_CARRY unary_minus_33_add_3_7 (.CI(n46200), .I0(GND_net), .I1(n46[5]), 
            .CO(n46201));
    SB_CARRY add_4325_4 (.CI(n47125), .I0(n11481[1]), .I1(n223_adj_4461), 
            .CO(n47126));
    SB_LUT4 unary_minus_33_add_3_6_lut (.I0(GND_net), .I1(GND_net), .I2(n46[4]), 
            .I3(n46199), .O(n535[4])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_33_add_3_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_33_add_3_6 (.CI(n46199), .I0(GND_net), .I1(n46[4]), 
            .CO(n46200));
    SB_LUT4 add_25_6_lut (.I0(GND_net), .I1(n360[4]), .I2(n42[4]), .I3(n46076), 
            .O(n455[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_25_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_33_add_3_5_lut (.I0(GND_net), .I1(GND_net), .I2(n46[3]), 
            .I3(n46198), .O(n535[3])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_33_add_3_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4325_3_lut (.I0(GND_net), .I1(n11481[0]), .I2(n150_adj_4467), 
            .I3(n47124), .O(n10514[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4325_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_25_6 (.CI(n46076), .I0(n360[4]), .I1(n42[4]), .CO(n46077));
    SB_LUT4 add_25_5_lut (.I0(GND_net), .I1(n360[3]), .I2(n42[3]), .I3(n46075), 
            .O(n455[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_25_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_25_5 (.CI(n46075), .I0(n360[3]), .I1(n42[3]), .CO(n46076));
    SB_LUT4 add_25_4_lut (.I0(GND_net), .I1(n360[2]), .I2(n42[2]), .I3(n46074), 
            .O(n455[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_25_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_25_4 (.CI(n46074), .I0(n360[2]), .I1(n42[2]), .CO(n46075));
    SB_CARRY unary_minus_33_add_3_5 (.CI(n46198), .I0(GND_net), .I1(n46[3]), 
            .CO(n46199));
    SB_LUT4 add_25_3_lut (.I0(GND_net), .I1(n360[1]), .I2(n42[1]), .I3(n46073), 
            .O(n455[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_25_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4325_3 (.CI(n47124), .I0(n11481[0]), .I1(n150_adj_4467), 
            .CO(n47125));
    SB_LUT4 add_4534_9_lut (.I0(GND_net), .I1(n15390[6]), .I2(n606_adj_4469), 
            .I3(n46777), .O(n14849[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4534_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4534_9 (.CI(n46777), .I0(n15390[6]), .I1(n606_adj_4469), 
            .CO(n46778));
    SB_LUT4 add_4534_8_lut (.I0(GND_net), .I1(n15390[5]), .I2(n533_adj_4470), 
            .I3(n46776), .O(n14849[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4534_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4325_2_lut (.I0(GND_net), .I1(n8_adj_4471), .I2(n77_adj_4472), 
            .I3(GND_net), .O(n10514[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4325_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4325_2 (.CI(GND_net), .I0(n8_adj_4471), .I1(n77_adj_4472), 
            .CO(n47124));
    SB_CARRY add_4534_8 (.CI(n46776), .I0(n15390[5]), .I1(n533_adj_4470), 
            .CO(n46777));
    SB_LUT4 add_4534_7_lut (.I0(GND_net), .I1(n15390[4]), .I2(n460_adj_4473), 
            .I3(n46775), .O(n14849[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4534_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4758_7_lut (.I0(GND_net), .I1(n54612), .I2(n490_adj_4474), 
            .I3(n47123), .O(n17891[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4758_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_33_add_3_4_lut (.I0(GND_net), .I1(GND_net), .I2(n46[2]), 
            .I3(n46197), .O(n535[2])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_33_add_3_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_25_3 (.CI(n46073), .I0(n360[1]), .I1(n42[1]), .CO(n46074));
    SB_LUT4 add_4758_6_lut (.I0(GND_net), .I1(n17961[3]), .I2(n417_adj_4477), 
            .I3(n47122), .O(n17891[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4758_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4758_6 (.CI(n47122), .I0(n17961[3]), .I1(n417_adj_4477), 
            .CO(n47123));
    SB_LUT4 add_4758_5_lut (.I0(GND_net), .I1(n17961[2]), .I2(n344_adj_4478), 
            .I3(n47121), .O(n17891[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4758_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4758_5 (.CI(n47121), .I0(n17961[2]), .I1(n344_adj_4478), 
            .CO(n47122));
    SB_LUT4 add_4758_4_lut (.I0(GND_net), .I1(n17961[1]), .I2(n271_adj_4479), 
            .I3(n47120), .O(n17891[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4758_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_33_add_3_4 (.CI(n46197), .I0(GND_net), .I1(n46[2]), 
            .CO(n46198));
    SB_LUT4 unary_minus_33_add_3_3_lut (.I0(GND_net), .I1(GND_net), .I2(n46[1]), 
            .I3(n46196), .O(n535[1])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_33_add_3_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4758_4 (.CI(n47120), .I0(n17961[1]), .I1(n271_adj_4479), 
            .CO(n47121));
    SB_CARRY unary_minus_33_add_3_3 (.CI(n46196), .I0(GND_net), .I1(n46[1]), 
            .CO(n46197));
    SB_LUT4 add_4758_3_lut (.I0(GND_net), .I1(n17961[0]), .I2(n198_adj_4481), 
            .I3(n47119), .O(n17891[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4758_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_33_add_3_2_lut (.I0(GND_net), .I1(GND_net), .I2(n46[0]), 
            .I3(VCC_net), .O(n535[0])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_33_add_3_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_25_2_lut (.I0(GND_net), .I1(n360[0]), .I2(n42[0]), .I3(GND_net), 
            .O(n455[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_25_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_25_2 (.CI(GND_net), .I0(n360[0]), .I1(n42[0]), .CO(n46073));
    SB_CARRY add_4758_3 (.CI(n47119), .I0(n17961[0]), .I1(n198_adj_4481), 
            .CO(n47120));
    SB_LUT4 add_16_25_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [23]), 
            .I2(n207[23]), .I3(n46072), .O(n233[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_16_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_33_add_3_2 (.CI(VCC_net), .I0(GND_net), .I1(n46[0]), 
            .CO(n46196));
    SB_LUT4 add_16_24_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [22]), 
            .I2(n207[23]), .I3(n46071), .O(n233[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_16_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_27_add_3_25_lut (.I0(n455[23]), .I1(GND_net), .I2(n28[23]), 
            .I3(n46195), .O(n47)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_27_add_3_25_lut.LUT_INIT = 16'h6996;
    SB_LUT4 add_4758_2_lut (.I0(GND_net), .I1(n56_adj_4484), .I2(n125_adj_4485), 
            .I3(GND_net), .O(n17891[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4758_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4758_2 (.CI(GND_net), .I0(n56_adj_4484), .I1(n125_adj_4485), 
            .CO(n47119));
    SB_LUT4 unary_minus_27_add_3_24_lut (.I0(GND_net), .I1(GND_net), .I2(n28[22]), 
            .I3(n46194), .O(n34[22])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_27_add_3_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_27_add_3_24 (.CI(n46194), .I0(GND_net), .I1(n28[22]), 
            .CO(n46195));
    SB_LUT4 add_4368_22_lut (.I0(GND_net), .I1(n12361[19]), .I2(GND_net), 
            .I3(n47118), .O(n11481[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4368_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_16_24 (.CI(n46071), .I0(\PID_CONTROLLER.integral [22]), 
            .I1(n207[23]), .CO(n46072));
    SB_LUT4 add_4368_21_lut (.I0(GND_net), .I1(n12361[18]), .I2(GND_net), 
            .I3(n47117), .O(n11481[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4368_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_16_23_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [21]), 
            .I2(n207[23]), .I3(n46070), .O(n233[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_16_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4368_21 (.CI(n47117), .I0(n12361[18]), .I1(GND_net), 
            .CO(n47118));
    SB_LUT4 unary_minus_27_add_3_23_lut (.I0(GND_net), .I1(GND_net), .I2(n28[21]), 
            .I3(n46193), .O(n34[21])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_27_add_3_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_16_23 (.CI(n46070), .I0(\PID_CONTROLLER.integral [21]), 
            .I1(n207[23]), .CO(n46071));
    SB_CARRY unary_minus_27_add_3_23 (.CI(n46193), .I0(GND_net), .I1(n28[21]), 
            .CO(n46194));
    SB_CARRY add_4534_7 (.CI(n46775), .I0(n15390[4]), .I1(n460_adj_4473), 
            .CO(n46776));
    SB_LUT4 add_4368_20_lut (.I0(GND_net), .I1(n12361[17]), .I2(GND_net), 
            .I3(n47116), .O(n11481[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4368_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4368_20 (.CI(n47116), .I0(n12361[17]), .I1(GND_net), 
            .CO(n47117));
    SB_LUT4 unary_minus_27_add_3_22_lut (.I0(GND_net), .I1(GND_net), .I2(n28[20]), 
            .I3(n46192), .O(n34[20])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_27_add_3_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_27_add_3_22 (.CI(n46192), .I0(GND_net), .I1(n28[20]), 
            .CO(n46193));
    SB_LUT4 add_4368_19_lut (.I0(GND_net), .I1(n12361[16]), .I2(GND_net), 
            .I3(n47115), .O(n11481[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4368_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_16_22_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [20]), 
            .I2(n207[23]), .I3(n46069), .O(n233[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_16_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_27_add_3_21_lut (.I0(GND_net), .I1(GND_net), .I2(n28[19]), 
            .I3(n46191), .O(n34[19])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_27_add_3_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_16_22 (.CI(n46069), .I0(\PID_CONTROLLER.integral [20]), 
            .I1(n207[23]), .CO(n46070));
    SB_CARRY add_4368_19 (.CI(n47115), .I0(n12361[16]), .I1(GND_net), 
            .CO(n47116));
    SB_LUT4 add_4534_6_lut (.I0(GND_net), .I1(n15390[3]), .I2(n387_adj_4491), 
            .I3(n46774), .O(n14849[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4534_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4368_18_lut (.I0(GND_net), .I1(n12361[15]), .I2(GND_net), 
            .I3(n47114), .O(n11481[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4368_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4368_18 (.CI(n47114), .I0(n12361[15]), .I1(GND_net), 
            .CO(n47115));
    SB_CARRY unary_minus_27_add_3_21 (.CI(n46191), .I0(GND_net), .I1(n28[19]), 
            .CO(n46192));
    SB_LUT4 add_4368_17_lut (.I0(GND_net), .I1(n12361[14]), .I2(GND_net), 
            .I3(n47113), .O(n11481[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4368_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_16_21_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [19]), 
            .I2(n207[23]), .I3(n46068), .O(n233[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_16_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_16_21 (.CI(n46068), .I0(\PID_CONTROLLER.integral [19]), 
            .I1(n207[23]), .CO(n46069));
    SB_CARRY add_4368_17 (.CI(n47113), .I0(n12361[14]), .I1(GND_net), 
            .CO(n47114));
    SB_LUT4 add_4368_16_lut (.I0(GND_net), .I1(n12361[13]), .I2(n1102_adj_4492), 
            .I3(n47112), .O(n11481[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4368_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4534_6 (.CI(n46774), .I0(n15390[3]), .I1(n387_adj_4491), 
            .CO(n46775));
    SB_LUT4 add_4534_5_lut (.I0(GND_net), .I1(n15390[2]), .I2(n314_adj_4493), 
            .I3(n46773), .O(n14849[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4534_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_27_add_3_20_lut (.I0(GND_net), .I1(GND_net), .I2(n28[18]), 
            .I3(n46190), .O(n34[18])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_27_add_3_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4368_16 (.CI(n47112), .I0(n12361[13]), .I1(n1102_adj_4492), 
            .CO(n47113));
    SB_LUT4 add_4368_15_lut (.I0(GND_net), .I1(n12361[12]), .I2(n1029_adj_4496), 
            .I3(n47111), .O(n11481[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4368_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_27_add_3_20 (.CI(n46190), .I0(GND_net), .I1(n28[18]), 
            .CO(n46191));
    SB_CARRY add_4534_5 (.CI(n46773), .I0(n15390[2]), .I1(n314_adj_4493), 
            .CO(n46774));
    SB_LUT4 add_16_20_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [18]), 
            .I2(n207[22]), .I3(n46067), .O(n233[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_16_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4534_4_lut (.I0(GND_net), .I1(n15390[1]), .I2(n241_adj_4497), 
            .I3(n46772), .O(n14849[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4534_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_27_add_3_19_lut (.I0(GND_net), .I1(GND_net), .I2(n28[17]), 
            .I3(n46189), .O(n34[17])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_27_add_3_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_16_20 (.CI(n46067), .I0(\PID_CONTROLLER.integral [18]), 
            .I1(n207[22]), .CO(n46068));
    SB_CARRY add_4368_15 (.CI(n47111), .I0(n12361[12]), .I1(n1029_adj_4496), 
            .CO(n47112));
    SB_LUT4 add_4368_14_lut (.I0(GND_net), .I1(n12361[11]), .I2(n956_adj_4499), 
            .I3(n47110), .O(n11481[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4368_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4534_4 (.CI(n46772), .I0(n15390[1]), .I1(n241_adj_4497), 
            .CO(n46773));
    SB_LUT4 add_4534_3_lut (.I0(GND_net), .I1(n15390[0]), .I2(n168_adj_4500), 
            .I3(n46771), .O(n14849[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4534_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4368_14 (.CI(n47110), .I0(n12361[11]), .I1(n956_adj_4499), 
            .CO(n47111));
    SB_LUT4 add_4368_13_lut (.I0(GND_net), .I1(n12361[10]), .I2(n883_adj_4501), 
            .I3(n47109), .O(n11481[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4368_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4534_3 (.CI(n46771), .I0(n15390[0]), .I1(n168_adj_4500), 
            .CO(n46772));
    SB_LUT4 add_4534_2_lut (.I0(GND_net), .I1(n26_adj_4502), .I2(n95_adj_4503), 
            .I3(GND_net), .O(n14849[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4534_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4368_13 (.CI(n47109), .I0(n12361[10]), .I1(n883_adj_4501), 
            .CO(n47110));
    SB_LUT4 add_4368_12_lut (.I0(GND_net), .I1(n12361[9]), .I2(n810_adj_4504), 
            .I3(n47108), .O(n11481[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4368_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4534_2 (.CI(GND_net), .I0(n26_adj_4502), .I1(n95_adj_4503), 
            .CO(n46771));
    SB_LUT4 add_4716_10_lut (.I0(GND_net), .I1(n17669[7]), .I2(n700), 
            .I3(n46770), .O(n17509[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4716_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_27_add_3_19 (.CI(n46189), .I0(GND_net), .I1(n28[17]), 
            .CO(n46190));
    SB_LUT4 unary_minus_27_add_3_18_lut (.I0(GND_net), .I1(GND_net), .I2(n28[16]), 
            .I3(n46188), .O(n34[16])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_27_add_3_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_16_19_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [17]), 
            .I2(n207[21]), .I3(n46066), .O(n240)) /* synthesis syn_instantiated=1 */ ;
    defparam add_16_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4368_12 (.CI(n47108), .I0(n12361[9]), .I1(n810_adj_4504), 
            .CO(n47109));
    SB_LUT4 add_4368_11_lut (.I0(GND_net), .I1(n12361[8]), .I2(n737_adj_4506), 
            .I3(n47107), .O(n11481[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4368_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_27_add_3_18 (.CI(n46188), .I0(GND_net), .I1(n28[16]), 
            .CO(n46189));
    SB_LUT4 unary_minus_27_add_3_17_lut (.I0(GND_net), .I1(GND_net), .I2(n28[15]), 
            .I3(n46187), .O(n34[15])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_27_add_3_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_27_add_3_17 (.CI(n46187), .I0(GND_net), .I1(n28[15]), 
            .CO(n46188));
    SB_CARRY add_16_19 (.CI(n46066), .I0(\PID_CONTROLLER.integral [17]), 
            .I1(n207[21]), .CO(n46067));
    SB_LUT4 add_16_18_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [16]), 
            .I2(n207[20]), .I3(n46065), .O(n233[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_16_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_27_add_3_16_lut (.I0(GND_net), .I1(GND_net), .I2(n28[14]), 
            .I3(n46186), .O(n34[14])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_27_add_3_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4368_11 (.CI(n47107), .I0(n12361[8]), .I1(n737_adj_4506), 
            .CO(n47108));
    SB_CARRY add_16_18 (.CI(n46065), .I0(\PID_CONTROLLER.integral [16]), 
            .I1(n207[20]), .CO(n46066));
    SB_CARRY unary_minus_27_add_3_16 (.CI(n46186), .I0(GND_net), .I1(n28[14]), 
            .CO(n46187));
    SB_LUT4 add_4368_10_lut (.I0(GND_net), .I1(n12361[7]), .I2(n664_adj_4510), 
            .I3(n47106), .O(n11481[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4368_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4368_10 (.CI(n47106), .I0(n12361[7]), .I1(n664_adj_4510), 
            .CO(n47107));
    SB_LUT4 add_4368_9_lut (.I0(GND_net), .I1(n12361[6]), .I2(n591_adj_4511), 
            .I3(n47105), .O(n11481[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4368_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4368_9 (.CI(n47105), .I0(n12361[6]), .I1(n591_adj_4511), 
            .CO(n47106));
    SB_LUT4 add_4716_9_lut (.I0(GND_net), .I1(n17669[6]), .I2(n627), .I3(n46769), 
            .O(n17509[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4716_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4716_9 (.CI(n46769), .I0(n17669[6]), .I1(n627), .CO(n46770));
    SB_LUT4 add_4368_8_lut (.I0(GND_net), .I1(n12361[5]), .I2(n518_adj_4512), 
            .I3(n47104), .O(n11481[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4368_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_27_add_3_15_lut (.I0(GND_net), .I1(GND_net), .I2(n28[13]), 
            .I3(n46185), .O(n34[13])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_27_add_3_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_27_add_3_15 (.CI(n46185), .I0(GND_net), .I1(n28[13]), 
            .CO(n46186));
    SB_CARRY add_4368_8 (.CI(n47104), .I0(n12361[5]), .I1(n518_adj_4512), 
            .CO(n47105));
    SB_LUT4 add_16_17_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [15]), 
            .I2(n207[19]), .I3(n46064), .O(n233[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_16_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4368_7_lut (.I0(GND_net), .I1(n12361[4]), .I2(n445_adj_4514), 
            .I3(n47103), .O(n11481[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4368_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4716_8_lut (.I0(GND_net), .I1(n17669[5]), .I2(n554_adj_4515), 
            .I3(n46768), .O(n17509[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4716_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4716_8 (.CI(n46768), .I0(n17669[5]), .I1(n554_adj_4515), 
            .CO(n46769));
    SB_CARRY add_4368_7 (.CI(n47103), .I0(n12361[4]), .I1(n445_adj_4514), 
            .CO(n47104));
    SB_LUT4 add_4368_6_lut (.I0(GND_net), .I1(n12361[3]), .I2(n372_adj_4516), 
            .I3(n47102), .O(n11481[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4368_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4716_7_lut (.I0(GND_net), .I1(n17669[4]), .I2(n481), .I3(n46767), 
            .O(n17509[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4716_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_16_17 (.CI(n46064), .I0(\PID_CONTROLLER.integral [15]), 
            .I1(n207[19]), .CO(n46065));
    SB_LUT4 unary_minus_27_add_3_14_lut (.I0(GND_net), .I1(GND_net), .I2(n28[12]), 
            .I3(n46184), .O(n34[12])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_27_add_3_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_16_16_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [14]), 
            .I2(n207[18]), .I3(n46063), .O(n233[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_16_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_27_add_3_14 (.CI(n46184), .I0(GND_net), .I1(n28[12]), 
            .CO(n46185));
    SB_CARRY add_4368_6 (.CI(n47102), .I0(n12361[3]), .I1(n372_adj_4516), 
            .CO(n47103));
    SB_LUT4 unary_minus_27_add_3_13_lut (.I0(GND_net), .I1(GND_net), .I2(n28[11]), 
            .I3(n46183), .O(n34[11])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_27_add_3_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4368_5_lut (.I0(GND_net), .I1(n12361[2]), .I2(n299_adj_4519), 
            .I3(n47101), .O(n11481[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4368_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4368_5 (.CI(n47101), .I0(n12361[2]), .I1(n299_adj_4519), 
            .CO(n47102));
    SB_LUT4 add_4368_4_lut (.I0(GND_net), .I1(n12361[1]), .I2(n226_adj_4520), 
            .I3(n47100), .O(n11481[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4368_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4716_7 (.CI(n46767), .I0(n17669[4]), .I1(n481), .CO(n46768));
    SB_CARRY add_4368_4 (.CI(n47100), .I0(n12361[1]), .I1(n226_adj_4520), 
            .CO(n47101));
    SB_LUT4 add_4368_3_lut (.I0(GND_net), .I1(n12361[0]), .I2(n153_adj_4521), 
            .I3(n47099), .O(n11481[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4368_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4716_6_lut (.I0(GND_net), .I1(n17669[3]), .I2(n408), .I3(n46766), 
            .O(n17509[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4716_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4716_6 (.CI(n46766), .I0(n17669[3]), .I1(n408), .CO(n46767));
    SB_CARRY add_4368_3 (.CI(n47099), .I0(n12361[0]), .I1(n153_adj_4521), 
            .CO(n47100));
    SB_CARRY unary_minus_27_add_3_13 (.CI(n46183), .I0(GND_net), .I1(n28[11]), 
            .CO(n46184));
    SB_LUT4 add_4368_2_lut (.I0(GND_net), .I1(n11_adj_4522), .I2(n80_adj_4523), 
            .I3(GND_net), .O(n11481[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4368_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4368_2 (.CI(GND_net), .I0(n11_adj_4522), .I1(n80_adj_4523), 
            .CO(n47099));
    SB_LUT4 add_4716_5_lut (.I0(GND_net), .I1(n17669[2]), .I2(n335), .I3(n46765), 
            .O(n17509[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4716_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_27_add_3_12_lut (.I0(GND_net), .I1(GND_net), .I2(n28[10]), 
            .I3(n46182), .O(n34[10])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_27_add_3_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_27_add_3_12 (.CI(n46182), .I0(GND_net), .I1(n28[10]), 
            .CO(n46183));
    SB_CARRY add_16_16 (.CI(n46063), .I0(\PID_CONTROLLER.integral [14]), 
            .I1(n207[18]), .CO(n46064));
    SB_LUT4 unary_minus_27_add_3_11_lut (.I0(GND_net), .I1(GND_net), .I2(n28[9]), 
            .I3(n46181), .O(n34[9])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_27_add_3_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_16_15_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [13]), 
            .I2(n207[17]), .I3(n46062), .O(n233[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_16_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_16_15 (.CI(n46062), .I0(\PID_CONTROLLER.integral [13]), 
            .I1(n207[17]), .CO(n46063));
    SB_CARRY add_4716_5 (.CI(n46765), .I0(n17669[2]), .I1(n335), .CO(n46766));
    SB_LUT4 add_4716_4_lut (.I0(GND_net), .I1(n17669[1]), .I2(n262), .I3(n46764), 
            .O(n17509[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4716_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_27_add_3_11 (.CI(n46181), .I0(GND_net), .I1(n28[9]), 
            .CO(n46182));
    SB_LUT4 add_4709_10_lut (.I0(GND_net), .I1(n17609[7]), .I2(n700_adj_4526), 
            .I3(n47098), .O(n17432[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4709_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4709_9_lut (.I0(GND_net), .I1(n17609[6]), .I2(n627_adj_4527), 
            .I3(n47097), .O(n17432[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4709_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4716_4 (.CI(n46764), .I0(n17669[1]), .I1(n262), .CO(n46765));
    SB_LUT4 add_4716_3_lut (.I0(GND_net), .I1(n17669[0]), .I2(n189), .I3(n46763), 
            .O(n17509[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4716_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_27_add_3_10_lut (.I0(GND_net), .I1(GND_net), .I2(n28[8]), 
            .I3(n46180), .O(n34[8])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_27_add_3_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_27_add_3_10 (.CI(n46180), .I0(GND_net), .I1(n28[8]), 
            .CO(n46181));
    SB_LUT4 add_16_14_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [12]), 
            .I2(n207[16]), .I3(n46061), .O(n233[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_16_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4709_9 (.CI(n47097), .I0(n17609[6]), .I1(n627_adj_4527), 
            .CO(n47098));
    SB_CARRY add_16_14 (.CI(n46061), .I0(\PID_CONTROLLER.integral [12]), 
            .I1(n207[16]), .CO(n46062));
    SB_LUT4 add_4709_8_lut (.I0(GND_net), .I1(n17609[5]), .I2(n554_adj_4529), 
            .I3(n47096), .O(n17432[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4709_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_27_add_3_9_lut (.I0(GND_net), .I1(GND_net), .I2(n28[7]), 
            .I3(n46179), .O(n34[7])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_27_add_3_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4709_8 (.CI(n47096), .I0(n17609[5]), .I1(n554_adj_4529), 
            .CO(n47097));
    SB_CARRY unary_minus_27_add_3_9 (.CI(n46179), .I0(GND_net), .I1(n28[7]), 
            .CO(n46180));
    SB_LUT4 unary_minus_27_add_3_8_lut (.I0(GND_net), .I1(GND_net), .I2(n28[6]), 
            .I3(n46178), .O(n34[6])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_27_add_3_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_27_add_3_8 (.CI(n46178), .I0(GND_net), .I1(n28[6]), 
            .CO(n46179));
    SB_LUT4 add_4709_7_lut (.I0(GND_net), .I1(n17609[4]), .I2(n481_adj_4532), 
            .I3(n47095), .O(n17432[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4709_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4709_7 (.CI(n47095), .I0(n17609[4]), .I1(n481_adj_4532), 
            .CO(n47096));
    SB_CARRY add_4716_3 (.CI(n46763), .I0(n17669[0]), .I1(n189), .CO(n46764));
    SB_LUT4 add_4716_2_lut (.I0(GND_net), .I1(n47_adj_4533), .I2(n116), 
            .I3(GND_net), .O(n17509[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4716_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4709_6_lut (.I0(GND_net), .I1(n17609[3]), .I2(n408_adj_4534), 
            .I3(n47094), .O(n17432[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4709_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4709_6 (.CI(n47094), .I0(n17609[3]), .I1(n408_adj_4534), 
            .CO(n47095));
    SB_LUT4 add_4709_5_lut (.I0(GND_net), .I1(n17609[2]), .I2(n335_adj_4535), 
            .I3(n47093), .O(n17432[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4709_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4716_2 (.CI(GND_net), .I0(n47_adj_4533), .I1(n116), .CO(n46763));
    SB_LUT4 add_4565_16_lut (.I0(GND_net), .I1(n15867[13]), .I2(n1120_adj_4536), 
            .I3(n46762), .O(n15390[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4565_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4709_5 (.CI(n47093), .I0(n17609[2]), .I1(n335_adj_4535), 
            .CO(n47094));
    SB_LUT4 add_4709_4_lut (.I0(GND_net), .I1(n17609[1]), .I2(n262_adj_4537), 
            .I3(n47092), .O(n17432[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4709_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4565_15_lut (.I0(GND_net), .I1(n15867[12]), .I2(n1047_adj_4538), 
            .I3(n46761), .O(n15390[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4565_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4565_15 (.CI(n46761), .I0(n15867[12]), .I1(n1047_adj_4538), 
            .CO(n46762));
    SB_CARRY add_4709_4 (.CI(n47092), .I0(n17609[1]), .I1(n262_adj_4537), 
            .CO(n47093));
    SB_LUT4 add_4709_3_lut (.I0(GND_net), .I1(n17609[0]), .I2(n189_adj_4539), 
            .I3(n47091), .O(n17432[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4709_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4565_14_lut (.I0(GND_net), .I1(n15867[11]), .I2(n974_adj_4540), 
            .I3(n46760), .O(n15390[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4565_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4565_14 (.CI(n46760), .I0(n15867[11]), .I1(n974_adj_4540), 
            .CO(n46761));
    SB_CARRY add_4709_3 (.CI(n47091), .I0(n17609[0]), .I1(n189_adj_4539), 
            .CO(n47092));
    SB_LUT4 add_4709_2_lut (.I0(GND_net), .I1(n47_adj_4541), .I2(n116_adj_4542), 
            .I3(GND_net), .O(n17432[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4709_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4565_13_lut (.I0(GND_net), .I1(n15867[10]), .I2(n901_adj_4543), 
            .I3(n46759), .O(n15390[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4565_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4565_13 (.CI(n46759), .I0(n15867[10]), .I1(n901_adj_4543), 
            .CO(n46760));
    SB_CARRY add_4709_2 (.CI(GND_net), .I0(n47_adj_4541), .I1(n116_adj_4542), 
            .CO(n47091));
    SB_LUT4 add_4408_21_lut (.I0(GND_net), .I1(n13159[18]), .I2(GND_net), 
            .I3(n47090), .O(n12361[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4408_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4408_20_lut (.I0(GND_net), .I1(n13159[17]), .I2(GND_net), 
            .I3(n47089), .O(n12361[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4408_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4565_12_lut (.I0(GND_net), .I1(n15867[9]), .I2(n828_adj_4544), 
            .I3(n46758), .O(n15390[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4565_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4565_12 (.CI(n46758), .I0(n15867[9]), .I1(n828_adj_4544), 
            .CO(n46759));
    SB_CARRY add_4408_20 (.CI(n47089), .I0(n13159[17]), .I1(GND_net), 
            .CO(n47090));
    SB_LUT4 add_4408_19_lut (.I0(GND_net), .I1(n13159[16]), .I2(GND_net), 
            .I3(n47088), .O(n12361[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4408_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4565_11_lut (.I0(GND_net), .I1(n15867[8]), .I2(n755_adj_4545), 
            .I3(n46757), .O(n15390[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4565_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4565_11 (.CI(n46757), .I0(n15867[8]), .I1(n755_adj_4545), 
            .CO(n46758));
    SB_LUT4 add_4565_10_lut (.I0(GND_net), .I1(n15867[7]), .I2(n682_adj_4546), 
            .I3(n46756), .O(n15390[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4565_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_27_add_3_7_lut (.I0(GND_net), .I1(GND_net), .I2(n28[5]), 
            .I3(n46177), .O(n34[5])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_27_add_3_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4565_10 (.CI(n46756), .I0(n15867[7]), .I1(n682_adj_4546), 
            .CO(n46757));
    SB_CARRY unary_minus_27_add_3_7 (.CI(n46177), .I0(GND_net), .I1(n28[5]), 
            .CO(n46178));
    SB_LUT4 unary_minus_27_add_3_6_lut (.I0(GND_net), .I1(GND_net), .I2(n28[4]), 
            .I3(n46176), .O(n34[4])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_27_add_3_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_16_13_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [11]), 
            .I2(n207[15]), .I3(n46060), .O(n233[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_16_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_16_13 (.CI(n46060), .I0(\PID_CONTROLLER.integral [11]), 
            .I1(n207[15]), .CO(n46061));
    SB_CARRY add_4408_19 (.CI(n47088), .I0(n13159[16]), .I1(GND_net), 
            .CO(n47089));
    SB_LUT4 add_4408_18_lut (.I0(GND_net), .I1(n13159[15]), .I2(GND_net), 
            .I3(n47087), .O(n12361[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4408_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4408_18 (.CI(n47087), .I0(n13159[15]), .I1(GND_net), 
            .CO(n47088));
    SB_LUT4 add_4565_9_lut (.I0(GND_net), .I1(n15867[6]), .I2(n609_adj_4548), 
            .I3(n46755), .O(n15390[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4565_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4565_9 (.CI(n46755), .I0(n15867[6]), .I1(n609_adj_4548), 
            .CO(n46756));
    SB_LUT4 add_4408_17_lut (.I0(GND_net), .I1(n13159[14]), .I2(GND_net), 
            .I3(n47086), .O(n12361[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4408_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4565_8_lut (.I0(GND_net), .I1(n15867[5]), .I2(n536_adj_4549), 
            .I3(n46754), .O(n15390[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4565_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4408_17 (.CI(n47086), .I0(n13159[14]), .I1(GND_net), 
            .CO(n47087));
    SB_CARRY add_4565_8 (.CI(n46754), .I0(n15867[5]), .I1(n536_adj_4549), 
            .CO(n46755));
    SB_LUT4 add_4408_16_lut (.I0(GND_net), .I1(n13159[13]), .I2(n1105_adj_4550), 
            .I3(n47085), .O(n12361[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4408_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4565_7_lut (.I0(GND_net), .I1(n15867[4]), .I2(n463_adj_4551), 
            .I3(n46753), .O(n15390[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4565_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4565_7 (.CI(n46753), .I0(n15867[4]), .I1(n463_adj_4551), 
            .CO(n46754));
    SB_CARRY add_4408_16 (.CI(n47085), .I0(n13159[13]), .I1(n1105_adj_4550), 
            .CO(n47086));
    SB_LUT4 add_4565_6_lut (.I0(GND_net), .I1(n15867[3]), .I2(n390_adj_4552), 
            .I3(n46752), .O(n15390[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4565_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4565_6 (.CI(n46752), .I0(n15867[3]), .I1(n390_adj_4552), 
            .CO(n46753));
    SB_LUT4 add_4408_15_lut (.I0(GND_net), .I1(n13159[12]), .I2(n1032_adj_4553), 
            .I3(n47084), .O(n12361[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4408_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4408_15 (.CI(n47084), .I0(n13159[12]), .I1(n1032_adj_4553), 
            .CO(n47085));
    SB_LUT4 add_4408_14_lut (.I0(GND_net), .I1(n13159[11]), .I2(n959_adj_4554), 
            .I3(n47083), .O(n12361[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4408_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4408_14 (.CI(n47083), .I0(n13159[11]), .I1(n959_adj_4554), 
            .CO(n47084));
    SB_LUT4 add_4408_13_lut (.I0(GND_net), .I1(n13159[10]), .I2(n886_adj_4555), 
            .I3(n47082), .O(n12361[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4408_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4408_13 (.CI(n47082), .I0(n13159[10]), .I1(n886_adj_4555), 
            .CO(n47083));
    SB_LUT4 add_4565_5_lut (.I0(GND_net), .I1(n15867[2]), .I2(n317_adj_4556), 
            .I3(n46751), .O(n15390[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4565_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4565_5 (.CI(n46751), .I0(n15867[2]), .I1(n317_adj_4556), 
            .CO(n46752));
    SB_LUT4 add_4408_12_lut (.I0(GND_net), .I1(n13159[9]), .I2(n813_adj_4557), 
            .I3(n47081), .O(n12361[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4408_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4408_12 (.CI(n47081), .I0(n13159[9]), .I1(n813_adj_4557), 
            .CO(n47082));
    SB_LUT4 add_4565_4_lut (.I0(GND_net), .I1(n15867[1]), .I2(n244_adj_4558), 
            .I3(n46750), .O(n15390[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4565_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4565_4 (.CI(n46750), .I0(n15867[1]), .I1(n244_adj_4558), 
            .CO(n46751));
    SB_LUT4 add_4408_11_lut (.I0(GND_net), .I1(n13159[8]), .I2(n740_adj_4559), 
            .I3(n47080), .O(n12361[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4408_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4408_11 (.CI(n47080), .I0(n13159[8]), .I1(n740_adj_4559), 
            .CO(n47081));
    SB_LUT4 add_4565_3_lut (.I0(GND_net), .I1(n15867[0]), .I2(n171_adj_4560), 
            .I3(n46749), .O(n15390[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4565_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4408_10_lut (.I0(GND_net), .I1(n13159[7]), .I2(n667_adj_4561), 
            .I3(n47079), .O(n12361[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4408_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4408_10 (.CI(n47079), .I0(n13159[7]), .I1(n667_adj_4561), 
            .CO(n47080));
    SB_CARRY add_4565_3 (.CI(n46749), .I0(n15867[0]), .I1(n171_adj_4560), 
            .CO(n46750));
    SB_LUT4 add_4408_9_lut (.I0(GND_net), .I1(n13159[6]), .I2(n594_adj_4562), 
            .I3(n47078), .O(n12361[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4408_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4565_2_lut (.I0(GND_net), .I1(n29_adj_4563), .I2(n98_adj_4564), 
            .I3(GND_net), .O(n15390[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4565_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4565_2 (.CI(GND_net), .I0(n29_adj_4563), .I1(n98_adj_4564), 
            .CO(n46749));
    SB_CARRY add_4408_9 (.CI(n47078), .I0(n13159[6]), .I1(n594_adj_4562), 
            .CO(n47079));
    SB_LUT4 add_4594_15_lut (.I0(GND_net), .I1(n16284[12]), .I2(n1050_adj_4565), 
            .I3(n46748), .O(n15867[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4594_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4594_14_lut (.I0(GND_net), .I1(n16284[11]), .I2(n977_adj_4566), 
            .I3(n46747), .O(n15867[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4594_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4408_8_lut (.I0(GND_net), .I1(n13159[5]), .I2(n521_adj_4567), 
            .I3(n47077), .O(n12361[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4408_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4594_14 (.CI(n46747), .I0(n16284[11]), .I1(n977_adj_4566), 
            .CO(n46748));
    SB_CARRY add_4408_8 (.CI(n47077), .I0(n13159[5]), .I1(n521_adj_4567), 
            .CO(n47078));
    SB_LUT4 add_4594_13_lut (.I0(GND_net), .I1(n16284[10]), .I2(n904_adj_4568), 
            .I3(n46746), .O(n15867[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4594_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4594_13 (.CI(n46746), .I0(n16284[10]), .I1(n904_adj_4568), 
            .CO(n46747));
    SB_LUT4 add_4408_7_lut (.I0(GND_net), .I1(n13159[4]), .I2(n448_adj_4569), 
            .I3(n47076), .O(n12361[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4408_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4408_7 (.CI(n47076), .I0(n13159[4]), .I1(n448_adj_4569), 
            .CO(n47077));
    SB_LUT4 add_4408_6_lut (.I0(GND_net), .I1(n13159[3]), .I2(n375_adj_4570), 
            .I3(n47075), .O(n12361[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4408_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4408_6 (.CI(n47075), .I0(n13159[3]), .I1(n375_adj_4570), 
            .CO(n47076));
    SB_LUT4 add_4408_5_lut (.I0(GND_net), .I1(n13159[2]), .I2(n302_adj_4571), 
            .I3(n47074), .O(n12361[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4408_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4594_12_lut (.I0(GND_net), .I1(n16284[9]), .I2(n831_adj_4572), 
            .I3(n46745), .O(n15867[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4594_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4408_5 (.CI(n47074), .I0(n13159[2]), .I1(n302_adj_4571), 
            .CO(n47075));
    SB_CARRY add_4594_12 (.CI(n46745), .I0(n16284[9]), .I1(n831_adj_4572), 
            .CO(n46746));
    SB_LUT4 add_4408_4_lut (.I0(GND_net), .I1(n13159[1]), .I2(n229_adj_4573), 
            .I3(n47073), .O(n12361[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4408_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4594_11_lut (.I0(GND_net), .I1(n16284[8]), .I2(n758_adj_4574), 
            .I3(n46744), .O(n15867[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4594_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4594_11 (.CI(n46744), .I0(n16284[8]), .I1(n758_adj_4574), 
            .CO(n46745));
    SB_CARRY add_4408_4 (.CI(n47073), .I0(n13159[1]), .I1(n229_adj_4573), 
            .CO(n47074));
    SB_LUT4 add_4594_10_lut (.I0(GND_net), .I1(n16284[7]), .I2(n685_adj_4575), 
            .I3(n46743), .O(n15867[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4594_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4594_10 (.CI(n46743), .I0(n16284[7]), .I1(n685_adj_4575), 
            .CO(n46744));
    SB_LUT4 add_4408_3_lut (.I0(GND_net), .I1(n13159[0]), .I2(n156_adj_4576), 
            .I3(n47072), .O(n12361[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4408_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4594_9_lut (.I0(GND_net), .I1(n16284[6]), .I2(n612_adj_4577), 
            .I3(n46742), .O(n15867[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4594_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4408_3 (.CI(n47072), .I0(n13159[0]), .I1(n156_adj_4576), 
            .CO(n47073));
    SB_LUT4 add_4408_2_lut (.I0(GND_net), .I1(n14_adj_4578), .I2(n83_adj_4579), 
            .I3(GND_net), .O(n12361[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4408_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4594_9 (.CI(n46742), .I0(n16284[6]), .I1(n612_adj_4577), 
            .CO(n46743));
    SB_CARRY add_4408_2 (.CI(GND_net), .I0(n14_adj_4578), .I1(n83_adj_4579), 
            .CO(n47072));
    SB_LUT4 add_4446_20_lut (.I0(GND_net), .I1(n13879[17]), .I2(GND_net), 
            .I3(n47071), .O(n13159[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4446_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4594_8_lut (.I0(GND_net), .I1(n16284[5]), .I2(n539_adj_4580), 
            .I3(n46741), .O(n15867[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4594_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4594_8 (.CI(n46741), .I0(n16284[5]), .I1(n539_adj_4580), 
            .CO(n46742));
    SB_LUT4 add_4446_19_lut (.I0(GND_net), .I1(n13879[16]), .I2(GND_net), 
            .I3(n47070), .O(n13159[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4446_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4446_19 (.CI(n47070), .I0(n13879[16]), .I1(GND_net), 
            .CO(n47071));
    SB_LUT4 add_4594_7_lut (.I0(GND_net), .I1(n16284[4]), .I2(n466_adj_4581), 
            .I3(n46740), .O(n15867[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4594_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4594_7 (.CI(n46740), .I0(n16284[4]), .I1(n466_adj_4581), 
            .CO(n46741));
    SB_LUT4 add_4446_18_lut (.I0(GND_net), .I1(n13879[15]), .I2(GND_net), 
            .I3(n47069), .O(n13159[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4446_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4446_18 (.CI(n47069), .I0(n13879[15]), .I1(GND_net), 
            .CO(n47070));
    SB_LUT4 add_4446_17_lut (.I0(GND_net), .I1(n13879[14]), .I2(GND_net), 
            .I3(n47068), .O(n13159[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4446_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4446_17 (.CI(n47068), .I0(n13879[14]), .I1(GND_net), 
            .CO(n47069));
    SB_LUT4 add_4446_16_lut (.I0(GND_net), .I1(n13879[13]), .I2(n1108_adj_4582), 
            .I3(n47067), .O(n13159[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4446_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4446_16 (.CI(n47067), .I0(n13879[13]), .I1(n1108_adj_4582), 
            .CO(n47068));
    SB_LUT4 add_4446_15_lut (.I0(GND_net), .I1(n13879[12]), .I2(n1035_adj_4583), 
            .I3(n47066), .O(n13159[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4446_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4446_15 (.CI(n47066), .I0(n13879[12]), .I1(n1035_adj_4583), 
            .CO(n47067));
    SB_LUT4 add_4446_14_lut (.I0(GND_net), .I1(n13879[11]), .I2(n962_adj_4584), 
            .I3(n47065), .O(n13159[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4446_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4446_14 (.CI(n47065), .I0(n13879[11]), .I1(n962_adj_4584), 
            .CO(n47066));
    SB_LUT4 add_4594_6_lut (.I0(GND_net), .I1(n16284[3]), .I2(n393_adj_4585), 
            .I3(n46739), .O(n15867[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4594_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4594_6 (.CI(n46739), .I0(n16284[3]), .I1(n393_adj_4585), 
            .CO(n46740));
    SB_LUT4 add_4446_13_lut (.I0(GND_net), .I1(n13879[10]), .I2(n889_adj_4586), 
            .I3(n47064), .O(n13159[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4446_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4594_5_lut (.I0(GND_net), .I1(n16284[2]), .I2(n320_adj_4587), 
            .I3(n46738), .O(n15867[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4594_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4594_5 (.CI(n46738), .I0(n16284[2]), .I1(n320_adj_4587), 
            .CO(n46739));
    SB_CARRY add_4446_13 (.CI(n47064), .I0(n13879[10]), .I1(n889_adj_4586), 
            .CO(n47065));
    SB_LUT4 add_4594_4_lut (.I0(GND_net), .I1(n16284[1]), .I2(n247_adj_4588), 
            .I3(n46737), .O(n15867[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4594_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4446_12_lut (.I0(GND_net), .I1(n13879[9]), .I2(n816_adj_4589), 
            .I3(n47063), .O(n13159[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4446_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4594_4 (.CI(n46737), .I0(n16284[1]), .I1(n247_adj_4588), 
            .CO(n46738));
    SB_LUT4 add_4594_3_lut (.I0(GND_net), .I1(n16284[0]), .I2(n174_adj_4590), 
            .I3(n46736), .O(n15867[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4594_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4446_12 (.CI(n47063), .I0(n13879[9]), .I1(n816_adj_4589), 
            .CO(n47064));
    SB_CARRY add_4594_3 (.CI(n46736), .I0(n16284[0]), .I1(n174_adj_4590), 
            .CO(n46737));
    SB_LUT4 add_4594_2_lut (.I0(GND_net), .I1(n32_adj_4591), .I2(n101_adj_4592), 
            .I3(GND_net), .O(n15867[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4594_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4446_11_lut (.I0(GND_net), .I1(n13879[8]), .I2(n743_adj_4593), 
            .I3(n47062), .O(n13159[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4446_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4446_11 (.CI(n47062), .I0(n13879[8]), .I1(n743_adj_4593), 
            .CO(n47063));
    SB_CARRY add_4594_2 (.CI(GND_net), .I0(n32_adj_4591), .I1(n101_adj_4592), 
            .CO(n46736));
    SB_LUT4 add_4732_9_lut (.I0(GND_net), .I1(n17795[6]), .I2(n630_adj_4594), 
            .I3(n46735), .O(n17669[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4732_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4446_10_lut (.I0(GND_net), .I1(n13879[7]), .I2(n670_adj_4595), 
            .I3(n47061), .O(n13159[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4446_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4446_10 (.CI(n47061), .I0(n13879[7]), .I1(n670_adj_4595), 
            .CO(n47062));
    SB_LUT4 add_4732_8_lut (.I0(GND_net), .I1(n17795[5]), .I2(n557_adj_4596), 
            .I3(n46734), .O(n17669[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4732_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4446_9_lut (.I0(GND_net), .I1(n13879[6]), .I2(n597_adj_4597), 
            .I3(n47060), .O(n13159[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4446_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4446_9 (.CI(n47060), .I0(n13879[6]), .I1(n597_adj_4597), 
            .CO(n47061));
    SB_CARRY add_4732_8 (.CI(n46734), .I0(n17795[5]), .I1(n557_adj_4596), 
            .CO(n46735));
    SB_LUT4 add_4446_8_lut (.I0(GND_net), .I1(n13879[5]), .I2(n524_adj_4598), 
            .I3(n47059), .O(n13159[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4446_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4446_8 (.CI(n47059), .I0(n13879[5]), .I1(n524_adj_4598), 
            .CO(n47060));
    SB_LUT4 add_4446_7_lut (.I0(GND_net), .I1(n13879[4]), .I2(n451_adj_4599), 
            .I3(n47058), .O(n13159[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4446_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4446_7 (.CI(n47058), .I0(n13879[4]), .I1(n451_adj_4599), 
            .CO(n47059));
    SB_LUT4 add_4446_6_lut (.I0(GND_net), .I1(n13879[3]), .I2(n378_adj_4600), 
            .I3(n47057), .O(n13159[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4446_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4446_6 (.CI(n47057), .I0(n13879[3]), .I1(n378_adj_4600), 
            .CO(n47058));
    SB_LUT4 add_4446_5_lut (.I0(GND_net), .I1(n13879[2]), .I2(n305_adj_4601), 
            .I3(n47056), .O(n13159[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4446_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4446_5 (.CI(n47056), .I0(n13879[2]), .I1(n305_adj_4601), 
            .CO(n47057));
    SB_LUT4 add_4446_4_lut (.I0(GND_net), .I1(n13879[1]), .I2(n232_adj_4602), 
            .I3(n47055), .O(n13159[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4446_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4446_4 (.CI(n47055), .I0(n13879[1]), .I1(n232_adj_4602), 
            .CO(n47056));
    SB_LUT4 n9440_bdd_4_lut_48653 (.I0(n9440), .I1(n59882), .I2(setpoint[5]), 
            .I3(n4357), .O(n63377));
    defparam n9440_bdd_4_lut_48653.LUT_INIT = 16'he4aa;
    SB_LUT4 add_4446_3_lut (.I0(GND_net), .I1(n13879[0]), .I2(n159_adj_4603), 
            .I3(n47054), .O(n13159[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4446_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4446_3 (.CI(n47054), .I0(n13879[0]), .I1(n159_adj_4603), 
            .CO(n47055));
    SB_LUT4 add_4446_2_lut (.I0(GND_net), .I1(n17_adj_4604), .I2(n86_adj_4605), 
            .I3(GND_net), .O(n13159[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4446_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4732_7_lut (.I0(GND_net), .I1(n17795[4]), .I2(n484_adj_4606), 
            .I3(n46733), .O(n17669[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4732_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 n63377_bdd_4_lut (.I0(n63377), .I1(n535[5]), .I2(n455[5]), 
            .I3(n4357), .O(n63380));
    defparam n63377_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_CARRY add_4446_2 (.CI(GND_net), .I0(n17_adj_4604), .I1(n86_adj_4605), 
            .CO(n47054));
    SB_CARRY add_4732_7 (.CI(n46733), .I0(n17795[4]), .I1(n484_adj_4606), 
            .CO(n46734));
    SB_LUT4 mult_24_i132_2_lut (.I0(\Ki[2] ), .I1(n343), .I2(GND_net), 
            .I3(GND_net), .O(n195_adj_4233));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i132_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_20_inv_0_i1_1_lut (.I0(IntegralLimit[0]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n36[0]));   // verilog/motorControl.v(59[24:38])
    defparam unary_minus_20_inv_0_i1_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_24_i561_2_lut (.I0(\Ki[11] ), .I1(n349), .I2(GND_net), 
            .I3(GND_net), .O(n834));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i561_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_20_inv_0_i2_1_lut (.I0(IntegralLimit[1]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n36[1]));   // verilog/motorControl.v(59[24:38])
    defparam unary_minus_20_inv_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_24_i181_2_lut (.I0(\Ki[3] ), .I1(n343), .I2(GND_net), 
            .I3(GND_net), .O(n268_adj_4229));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i181_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_17_i9_2_lut (.I0(IntegralLimit[4]), .I1(n233[4]), .I2(GND_net), 
            .I3(GND_net), .O(n9_adj_4238));   // verilog/motorControl.v(56[14:36])
    defparam LessThan_17_i9_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_17_i11_2_lut (.I0(IntegralLimit[5]), .I1(n233[5]), 
            .I2(GND_net), .I3(GND_net), .O(n11_adj_4243));   // verilog/motorControl.v(56[14:36])
    defparam LessThan_17_i11_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_17_i13_2_lut (.I0(IntegralLimit[6]), .I1(n233[6]), 
            .I2(GND_net), .I3(GND_net), .O(n13_adj_4242));   // verilog/motorControl.v(56[14:36])
    defparam LessThan_17_i13_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_17_i15_2_lut (.I0(IntegralLimit[7]), .I1(n233[7]), 
            .I2(GND_net), .I3(GND_net), .O(n15_adj_4241));   // verilog/motorControl.v(56[14:36])
    defparam LessThan_17_i15_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_17_i21_2_lut (.I0(IntegralLimit[10]), .I1(n233[10]), 
            .I2(GND_net), .I3(GND_net), .O(n21_adj_4235));   // verilog/motorControl.v(56[14:36])
    defparam LessThan_17_i21_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_17_i19_2_lut (.I0(IntegralLimit[9]), .I1(n233[9]), 
            .I2(GND_net), .I3(GND_net), .O(n19_adj_4236));   // verilog/motorControl.v(56[14:36])
    defparam LessThan_17_i19_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_17_i17_2_lut (.I0(IntegralLimit[8]), .I1(n233[8]), 
            .I2(GND_net), .I3(GND_net), .O(n17_adj_4237));   // verilog/motorControl.v(56[14:36])
    defparam LessThan_17_i17_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 unary_minus_20_inv_0_i3_1_lut (.I0(IntegralLimit[2]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n36[2]));   // verilog/motorControl.v(59[24:38])
    defparam unary_minus_20_inv_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 LessThan_17_i23_2_lut (.I0(IntegralLimit[11]), .I1(n233[11]), 
            .I2(GND_net), .I3(GND_net), .O(n23_adj_4247));   // verilog/motorControl.v(56[14:36])
    defparam LessThan_17_i23_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_17_i25_2_lut (.I0(IntegralLimit[12]), .I1(n233[12]), 
            .I2(GND_net), .I3(GND_net), .O(n25_adj_4246));   // verilog/motorControl.v(56[14:36])
    defparam LessThan_17_i25_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_19_i9_2_lut (.I0(n233[4]), .I1(n285[4]), .I2(GND_net), 
            .I3(GND_net), .O(n9_adj_4274));   // verilog/motorControl.v(58[23:46])
    defparam LessThan_19_i9_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_19_i11_2_lut (.I0(n233[5]), .I1(n285[5]), .I2(GND_net), 
            .I3(GND_net), .O(n11_adj_4279));   // verilog/motorControl.v(58[23:46])
    defparam LessThan_19_i11_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_19_i13_2_lut (.I0(n233[6]), .I1(n285[6]), .I2(GND_net), 
            .I3(GND_net), .O(n13_adj_4278));   // verilog/motorControl.v(58[23:46])
    defparam LessThan_19_i13_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_19_i15_2_lut (.I0(n233[7]), .I1(n285[7]), .I2(GND_net), 
            .I3(GND_net), .O(n15_adj_4277));   // verilog/motorControl.v(58[23:46])
    defparam LessThan_19_i15_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_19_i21_2_lut (.I0(n233[10]), .I1(n285[10]), .I2(GND_net), 
            .I3(GND_net), .O(n21_adj_4271));   // verilog/motorControl.v(58[23:46])
    defparam LessThan_19_i21_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_19_i19_2_lut (.I0(n233[9]), .I1(n285[9]), .I2(GND_net), 
            .I3(GND_net), .O(n19_adj_4272));   // verilog/motorControl.v(58[23:46])
    defparam LessThan_19_i19_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_19_i17_2_lut (.I0(n233[8]), .I1(n285[8]), .I2(GND_net), 
            .I3(GND_net), .O(n17_adj_4273));   // verilog/motorControl.v(58[23:46])
    defparam LessThan_19_i17_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_19_i23_2_lut (.I0(n233[11]), .I1(n285[11]), .I2(GND_net), 
            .I3(GND_net), .O(n23_adj_4290));   // verilog/motorControl.v(58[23:46])
    defparam LessThan_19_i23_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_19_i25_2_lut (.I0(n233[12]), .I1(n285[12]), .I2(GND_net), 
            .I3(GND_net), .O(n25_adj_4289));   // verilog/motorControl.v(58[23:46])
    defparam LessThan_19_i25_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_24_i230_2_lut (.I0(\Ki[4] ), .I1(n343), .I2(GND_net), 
            .I3(GND_net), .O(n341_adj_4226));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i230_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_20_inv_0_i4_1_lut (.I0(IntegralLimit[3]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n36[3]));   // verilog/motorControl.v(59[24:38])
    defparam unary_minus_20_inv_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 LessThan_32_i41_2_lut (.I0(n455[20]), .I1(n535[20]), .I2(GND_net), 
            .I3(GND_net), .O(n41_adj_4607));   // verilog/motorControl.v(65[25:41])
    defparam LessThan_32_i41_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_32_i39_2_lut (.I0(n455[19]), .I1(n535[19]), .I2(GND_net), 
            .I3(GND_net), .O(n39_adj_4608));   // verilog/motorControl.v(65[25:41])
    defparam LessThan_32_i39_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_32_i45_2_lut (.I0(n455[22]), .I1(n535[22]), .I2(GND_net), 
            .I3(GND_net), .O(n45_adj_4609));   // verilog/motorControl.v(65[25:41])
    defparam LessThan_32_i45_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_32_i43_2_lut (.I0(n455[21]), .I1(n535[21]), .I2(GND_net), 
            .I3(GND_net), .O(n43_adj_4610));   // verilog/motorControl.v(65[25:41])
    defparam LessThan_32_i43_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_32_i21_2_lut (.I0(n455[10]), .I1(n535[10]), .I2(GND_net), 
            .I3(GND_net), .O(n21_adj_4611));   // verilog/motorControl.v(65[25:41])
    defparam LessThan_32_i21_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_32_i23_2_lut (.I0(n455[11]), .I1(n535[11]), .I2(GND_net), 
            .I3(GND_net), .O(n23_adj_4612));   // verilog/motorControl.v(65[25:41])
    defparam LessThan_32_i23_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_32_i25_2_lut (.I0(n455[12]), .I1(n535[12]), .I2(GND_net), 
            .I3(GND_net), .O(n25_adj_4613));   // verilog/motorControl.v(65[25:41])
    defparam LessThan_32_i25_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_32_i17_2_lut (.I0(n455[8]), .I1(n535[8]), .I2(GND_net), 
            .I3(GND_net), .O(n17_adj_4614));   // verilog/motorControl.v(65[25:41])
    defparam LessThan_32_i17_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_32_i19_2_lut (.I0(n455[9]), .I1(n535[9]), .I2(GND_net), 
            .I3(GND_net), .O(n19_adj_4615));   // verilog/motorControl.v(65[25:41])
    defparam LessThan_32_i19_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_32_i37_2_lut (.I0(n455[18]), .I1(n535[18]), .I2(GND_net), 
            .I3(GND_net), .O(n37_adj_4616));   // verilog/motorControl.v(65[25:41])
    defparam LessThan_32_i37_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_32_i35_2_lut (.I0(n455[17]), .I1(n535[17]), .I2(GND_net), 
            .I3(GND_net), .O(n35_adj_4617));   // verilog/motorControl.v(65[25:41])
    defparam LessThan_32_i35_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_32_i27_2_lut (.I0(n455[13]), .I1(n535[13]), .I2(GND_net), 
            .I3(GND_net), .O(n27_adj_4618));   // verilog/motorControl.v(65[25:41])
    defparam LessThan_32_i27_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_32_i29_2_lut (.I0(n455[14]), .I1(n535[14]), .I2(GND_net), 
            .I3(GND_net), .O(n29_adj_4619));   // verilog/motorControl.v(65[25:41])
    defparam LessThan_32_i29_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_32_i31_2_lut (.I0(n455[15]), .I1(n535[15]), .I2(GND_net), 
            .I3(GND_net), .O(n31_adj_4620));   // verilog/motorControl.v(65[25:41])
    defparam LessThan_32_i31_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_32_i9_2_lut (.I0(n455[4]), .I1(n535[4]), .I2(GND_net), 
            .I3(GND_net), .O(n9_adj_4621));   // verilog/motorControl.v(65[25:41])
    defparam LessThan_32_i9_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_32_i11_2_lut (.I0(n455[5]), .I1(n535[5]), .I2(GND_net), 
            .I3(GND_net), .O(n11_adj_4622));   // verilog/motorControl.v(65[25:41])
    defparam LessThan_32_i11_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_32_i13_2_lut (.I0(n455[6]), .I1(n535[6]), .I2(GND_net), 
            .I3(GND_net), .O(n13_adj_4623));   // verilog/motorControl.v(65[25:41])
    defparam LessThan_32_i13_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_32_i15_2_lut (.I0(n455[7]), .I1(n535[7]), .I2(GND_net), 
            .I3(GND_net), .O(n15_adj_4624));   // verilog/motorControl.v(65[25:41])
    defparam LessThan_32_i15_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_11_i41_2_lut (.I0(setpoint[20]), .I1(n535[20]), .I2(GND_net), 
            .I3(GND_net), .O(n41_adj_4625));   // verilog/motorControl.v(47[25:43])
    defparam LessThan_11_i41_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_11_i39_2_lut (.I0(setpoint[19]), .I1(n535[19]), .I2(GND_net), 
            .I3(GND_net), .O(n39_adj_4626));   // verilog/motorControl.v(47[25:43])
    defparam LessThan_11_i39_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_11_i45_2_lut (.I0(setpoint[22]), .I1(n535[22]), .I2(GND_net), 
            .I3(GND_net), .O(n45_adj_4627));   // verilog/motorControl.v(47[25:43])
    defparam LessThan_11_i45_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_11_i43_2_lut (.I0(setpoint[21]), .I1(n535[21]), .I2(GND_net), 
            .I3(GND_net), .O(n43_adj_4628));   // verilog/motorControl.v(47[25:43])
    defparam LessThan_11_i43_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_11_i29_2_lut (.I0(setpoint[14]), .I1(n535[14]), .I2(GND_net), 
            .I3(GND_net), .O(n29_adj_4629));   // verilog/motorControl.v(47[25:43])
    defparam LessThan_11_i29_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_11_i31_2_lut (.I0(setpoint[15]), .I1(n535[15]), .I2(GND_net), 
            .I3(GND_net), .O(n31_adj_4630));   // verilog/motorControl.v(47[25:43])
    defparam LessThan_11_i31_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_11_i23_2_lut (.I0(setpoint[11]), .I1(n535[11]), .I2(GND_net), 
            .I3(GND_net), .O(n23_adj_4631));   // verilog/motorControl.v(47[25:43])
    defparam LessThan_11_i23_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_11_i25_2_lut (.I0(setpoint[12]), .I1(n535[12]), .I2(GND_net), 
            .I3(GND_net), .O(n25_adj_4632));   // verilog/motorControl.v(47[25:43])
    defparam LessThan_11_i25_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_11_i37_2_lut (.I0(setpoint[18]), .I1(n535[18]), .I2(GND_net), 
            .I3(GND_net), .O(n37_adj_4633));   // verilog/motorControl.v(47[25:43])
    defparam LessThan_11_i37_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_11_i35_2_lut (.I0(setpoint[17]), .I1(n535[17]), .I2(GND_net), 
            .I3(GND_net), .O(n35_adj_4634));   // verilog/motorControl.v(47[25:43])
    defparam LessThan_11_i35_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_11_i33_2_lut (.I0(setpoint[16]), .I1(n535[16]), .I2(GND_net), 
            .I3(GND_net), .O(n33_adj_4635));   // verilog/motorControl.v(47[25:43])
    defparam LessThan_11_i33_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_11_i11_2_lut (.I0(setpoint[5]), .I1(n535[5]), .I2(GND_net), 
            .I3(GND_net), .O(n11_adj_4636));   // verilog/motorControl.v(47[25:43])
    defparam LessThan_11_i11_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_11_i13_2_lut (.I0(setpoint[6]), .I1(n535[6]), .I2(GND_net), 
            .I3(GND_net), .O(n13_adj_4637));   // verilog/motorControl.v(47[25:43])
    defparam LessThan_11_i13_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_23_i326_2_lut (.I0(\Kp[6] ), .I1(n207[19]), .I2(GND_net), 
            .I3(GND_net), .O(n484_adj_4606));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i326_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_11_i15_2_lut (.I0(setpoint[7]), .I1(n535[7]), .I2(GND_net), 
            .I3(GND_net), .O(n15_adj_4638));   // verilog/motorControl.v(47[25:43])
    defparam LessThan_11_i15_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_23_i59_2_lut (.I0(\Kp[1] ), .I1(n207[8]), .I2(GND_net), 
            .I3(GND_net), .O(n86_adj_4605));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i59_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i12_2_lut (.I0(\Kp[0] ), .I1(n207[9]), .I2(GND_net), 
            .I3(GND_net), .O(n17_adj_4604));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i12_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_11_i27_2_lut (.I0(setpoint[13]), .I1(n535[13]), .I2(GND_net), 
            .I3(GND_net), .O(n27_adj_4639));   // verilog/motorControl.v(47[25:43])
    defparam LessThan_11_i27_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_23_i108_2_lut (.I0(\Kp[2] ), .I1(n207[8]), .I2(GND_net), 
            .I3(GND_net), .O(n159_adj_4603));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i108_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_11_i9_2_lut (.I0(setpoint[4]), .I1(n535[4]), .I2(GND_net), 
            .I3(GND_net), .O(n9_adj_4640));   // verilog/motorControl.v(47[25:43])
    defparam LessThan_11_i9_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_23_i157_2_lut (.I0(\Kp[3] ), .I1(n207[8]), .I2(GND_net), 
            .I3(GND_net), .O(n232_adj_4602));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i157_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i206_2_lut (.I0(\Kp[4] ), .I1(n207[8]), .I2(GND_net), 
            .I3(GND_net), .O(n305_adj_4601));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i206_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i255_2_lut (.I0(\Kp[5] ), .I1(n207[8]), .I2(GND_net), 
            .I3(GND_net), .O(n378_adj_4600));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i255_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_11_i17_2_lut (.I0(setpoint[8]), .I1(n535[8]), .I2(GND_net), 
            .I3(GND_net), .O(n17_adj_4641));   // verilog/motorControl.v(47[25:43])
    defparam LessThan_11_i17_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_23_i304_2_lut (.I0(\Kp[6] ), .I1(n207[8]), .I2(GND_net), 
            .I3(GND_net), .O(n451_adj_4599));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i304_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i353_2_lut (.I0(\Kp[7] ), .I1(n207[8]), .I2(GND_net), 
            .I3(GND_net), .O(n524_adj_4598));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i353_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_11_i19_2_lut (.I0(setpoint[9]), .I1(n535[9]), .I2(GND_net), 
            .I3(GND_net), .O(n19_adj_4642));   // verilog/motorControl.v(47[25:43])
    defparam LessThan_11_i19_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_23_i402_2_lut (.I0(\Kp[8] ), .I1(n207[8]), .I2(GND_net), 
            .I3(GND_net), .O(n597_adj_4597));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i402_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_11_i21_2_lut (.I0(setpoint[10]), .I1(n535[10]), .I2(GND_net), 
            .I3(GND_net), .O(n21_adj_4643));   // verilog/motorControl.v(47[25:43])
    defparam LessThan_11_i21_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_23_i375_2_lut (.I0(\Kp[7] ), .I1(n207[19]), .I2(GND_net), 
            .I3(GND_net), .O(n557_adj_4596));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i375_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i451_2_lut (.I0(\Kp[9] ), .I1(n207[8]), .I2(GND_net), 
            .I3(GND_net), .O(n670_adj_4595));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i451_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i424_2_lut (.I0(\Kp[8] ), .I1(n207[19]), .I2(GND_net), 
            .I3(GND_net), .O(n630_adj_4594));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i424_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i500_2_lut (.I0(\Kp[10] ), .I1(n207[8]), .I2(GND_net), 
            .I3(GND_net), .O(n743_adj_4593));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i500_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i69_2_lut (.I0(\Ki[1] ), .I1(n350), .I2(GND_net), 
            .I3(GND_net), .O(n101_adj_4592));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i69_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i45789_4_lut (.I0(n21_adj_4643), .I1(n19_adj_4642), .I2(n17_adj_4641), 
            .I3(n9_adj_4640), .O(n60501));
    defparam i45789_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 mult_24_i22_2_lut (.I0(\Ki[0] ), .I1(n349), .I2(GND_net), 
            .I3(GND_net), .O(n32_adj_4591));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i22_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i118_2_lut (.I0(\Ki[2] ), .I1(n350), .I2(GND_net), 
            .I3(GND_net), .O(n174_adj_4590));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i118_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i549_2_lut (.I0(\Kp[11] ), .I1(n207[8]), .I2(GND_net), 
            .I3(GND_net), .O(n816_adj_4589));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i549_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i167_2_lut (.I0(\Ki[3] ), .I1(n350), .I2(GND_net), 
            .I3(GND_net), .O(n247_adj_4588));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i167_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i216_2_lut (.I0(\Ki[4] ), .I1(n350), .I2(GND_net), 
            .I3(GND_net), .O(n320_adj_4587));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i216_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i45767_4_lut (.I0(n27_adj_4639), .I1(n15_adj_4638), .I2(n13_adj_4637), 
            .I3(n11_adj_4636), .O(n60479));
    defparam i45767_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 LessThan_11_i12_3_lut (.I0(n535[7]), .I1(n535[16]), .I2(n33_adj_4635), 
            .I3(GND_net), .O(n12_adj_4644));   // verilog/motorControl.v(47[25:43])
    defparam LessThan_11_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_23_i598_2_lut (.I0(\Kp[12] ), .I1(n207[8]), .I2(GND_net), 
            .I3(GND_net), .O(n889_adj_4586));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i598_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i265_2_lut (.I0(\Ki[5] ), .I1(n350), .I2(GND_net), 
            .I3(GND_net), .O(n393_adj_4585));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i265_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i647_2_lut (.I0(\Kp[13] ), .I1(n207[8]), .I2(GND_net), 
            .I3(GND_net), .O(n962_adj_4584));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i647_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i696_2_lut (.I0(\Kp[14] ), .I1(n207[8]), .I2(GND_net), 
            .I3(GND_net), .O(n1035_adj_4583));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i696_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i745_2_lut (.I0(\Kp[15] ), .I1(n207[8]), .I2(GND_net), 
            .I3(GND_net), .O(n1108_adj_4582));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i745_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_11_i10_3_lut (.I0(n535[5]), .I1(n535[6]), .I2(n13_adj_4637), 
            .I3(GND_net), .O(n10_adj_4645));   // verilog/motorControl.v(47[25:43])
    defparam LessThan_11_i10_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_24_i314_2_lut (.I0(\Ki[6] ), .I1(n350), .I2(GND_net), 
            .I3(GND_net), .O(n466_adj_4581));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i314_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i363_2_lut (.I0(\Ki[7] ), .I1(n350), .I2(GND_net), 
            .I3(GND_net), .O(n539_adj_4580));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i363_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_11_i30_3_lut (.I0(n12_adj_4644), .I1(n535[17]), .I2(n35_adj_4634), 
            .I3(GND_net), .O(n30_adj_4646));   // verilog/motorControl.v(47[25:43])
    defparam LessThan_11_i30_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_23_i57_2_lut (.I0(\Kp[1] ), .I1(n207[7]), .I2(GND_net), 
            .I3(GND_net), .O(n83_adj_4579));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i57_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i10_2_lut (.I0(\Kp[0] ), .I1(n207[8]), .I2(GND_net), 
            .I3(GND_net), .O(n14_adj_4578));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i10_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i412_2_lut (.I0(\Ki[8] ), .I1(n350), .I2(GND_net), 
            .I3(GND_net), .O(n612_adj_4577));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i412_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i106_2_lut (.I0(\Kp[2] ), .I1(n207[7]), .I2(GND_net), 
            .I3(GND_net), .O(n156_adj_4576));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i106_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i461_2_lut (.I0(\Ki[9] ), .I1(n350), .I2(GND_net), 
            .I3(GND_net), .O(n685_adj_4575));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i461_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i510_2_lut (.I0(\Ki[10] ), .I1(n350), .I2(GND_net), 
            .I3(GND_net), .O(n758_adj_4574));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i510_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i155_2_lut (.I0(\Kp[3] ), .I1(n207[7]), .I2(GND_net), 
            .I3(GND_net), .O(n229_adj_4573));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i155_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i46782_4_lut (.I0(n13_adj_4637), .I1(n11_adj_4636), .I2(n9_adj_4640), 
            .I3(n60553), .O(n61495));
    defparam i46782_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i46774_4_lut (.I0(n19_adj_4642), .I1(n17_adj_4641), .I2(n15_adj_4638), 
            .I3(n61495), .O(n61487));
    defparam i46774_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i47954_4_lut (.I0(n25_adj_4632), .I1(n23_adj_4631), .I2(n21_adj_4643), 
            .I3(n61487), .O(n62667));
    defparam i47954_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i47281_4_lut (.I0(n31_adj_4630), .I1(n29_adj_4629), .I2(n27_adj_4639), 
            .I3(n62667), .O(n61994));
    defparam i47281_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 mult_24_i559_2_lut (.I0(\Ki[11] ), .I1(n350), .I2(GND_net), 
            .I3(GND_net), .O(n831_adj_4572));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i559_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i204_2_lut (.I0(\Kp[4] ), .I1(n207[7]), .I2(GND_net), 
            .I3(GND_net), .O(n302_adj_4571));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i204_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i253_2_lut (.I0(\Kp[5] ), .I1(n207[7]), .I2(GND_net), 
            .I3(GND_net), .O(n375_adj_4570));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i253_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i302_2_lut (.I0(\Kp[6] ), .I1(n207[7]), .I2(GND_net), 
            .I3(GND_net), .O(n448_adj_4569));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i302_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i48097_4_lut (.I0(n37_adj_4633), .I1(n35_adj_4634), .I2(n33_adj_4635), 
            .I3(n61994), .O(n62810));
    defparam i48097_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 mult_24_i608_2_lut (.I0(\Ki[12] ), .I1(n350), .I2(GND_net), 
            .I3(GND_net), .O(n904_adj_4568));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i608_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i351_2_lut (.I0(\Kp[7] ), .I1(n207[7]), .I2(GND_net), 
            .I3(GND_net), .O(n521_adj_4567));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i351_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_11_i16_3_lut (.I0(n535[9]), .I1(n535[21]), .I2(n43_adj_4628), 
            .I3(GND_net), .O(n16_adj_4647));   // verilog/motorControl.v(47[25:43])
    defparam LessThan_11_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i47651_3_lut (.I0(n6_adj_4648), .I1(n535[10]), .I2(n21_adj_4643), 
            .I3(GND_net), .O(n62364));   // verilog/motorControl.v(47[25:43])
    defparam i47651_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_24_i657_2_lut (.I0(\Ki[13] ), .I1(n350), .I2(GND_net), 
            .I3(GND_net), .O(n977_adj_4566));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i657_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i706_2_lut (.I0(\Ki[14] ), .I1(n350), .I2(GND_net), 
            .I3(GND_net), .O(n1050_adj_4565));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i706_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i67_2_lut (.I0(\Ki[1] ), .I1(n351), .I2(GND_net), 
            .I3(GND_net), .O(n98_adj_4564));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i67_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i20_2_lut (.I0(\Ki[0] ), .I1(n350), .I2(GND_net), 
            .I3(GND_net), .O(n29_adj_4563));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i20_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i400_2_lut (.I0(\Kp[8] ), .I1(n207[7]), .I2(GND_net), 
            .I3(GND_net), .O(n594_adj_4562));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i400_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i449_2_lut (.I0(\Kp[9] ), .I1(n207[7]), .I2(GND_net), 
            .I3(GND_net), .O(n667_adj_4561));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i449_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i116_2_lut (.I0(\Ki[2] ), .I1(n351), .I2(GND_net), 
            .I3(GND_net), .O(n171_adj_4560));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i116_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i47652_3_lut (.I0(n62364), .I1(n535[11]), .I2(n23_adj_4631), 
            .I3(GND_net), .O(n62365));   // verilog/motorControl.v(47[25:43])
    defparam i47652_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_23_i498_2_lut (.I0(\Kp[10] ), .I1(n207[7]), .I2(GND_net), 
            .I3(GND_net), .O(n740_adj_4559));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i498_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i165_2_lut (.I0(\Ki[3] ), .I1(n351), .I2(GND_net), 
            .I3(GND_net), .O(n244_adj_4558));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i165_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i547_2_lut (.I0(\Kp[11] ), .I1(n207[7]), .I2(GND_net), 
            .I3(GND_net), .O(n813_adj_4557));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i547_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i214_2_lut (.I0(\Ki[4] ), .I1(n351), .I2(GND_net), 
            .I3(GND_net), .O(n317_adj_4556));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i214_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i596_2_lut (.I0(\Kp[12] ), .I1(n207[7]), .I2(GND_net), 
            .I3(GND_net), .O(n886_adj_4555));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i596_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i645_2_lut (.I0(\Kp[13] ), .I1(n207[7]), .I2(GND_net), 
            .I3(GND_net), .O(n959_adj_4554));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i645_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i694_2_lut (.I0(\Kp[14] ), .I1(n207[7]), .I2(GND_net), 
            .I3(GND_net), .O(n1032_adj_4553));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i694_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_11_i8_3_lut (.I0(n535[4]), .I1(n535[8]), .I2(n17_adj_4641), 
            .I3(GND_net), .O(n8_adj_4649));   // verilog/motorControl.v(47[25:43])
    defparam LessThan_11_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_24_i263_2_lut (.I0(\Ki[5] ), .I1(n351), .I2(GND_net), 
            .I3(GND_net), .O(n390_adj_4552));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i263_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i312_2_lut (.I0(\Ki[6] ), .I1(n351), .I2(GND_net), 
            .I3(GND_net), .O(n463_adj_4551));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i312_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i743_2_lut (.I0(\Kp[15] ), .I1(n207[7]), .I2(GND_net), 
            .I3(GND_net), .O(n1105_adj_4550));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i743_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i361_2_lut (.I0(\Ki[7] ), .I1(n351), .I2(GND_net), 
            .I3(GND_net), .O(n536_adj_4549));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i361_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i410_2_lut (.I0(\Ki[8] ), .I1(n351), .I2(GND_net), 
            .I3(GND_net), .O(n609_adj_4548));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i410_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_27_inv_0_i6_1_lut (.I0(\deadband[5] ), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n28[5]));   // verilog/motorControl.v(62[45:54])
    defparam unary_minus_27_inv_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_24_i459_2_lut (.I0(\Ki[9] ), .I1(n351), .I2(GND_net), 
            .I3(GND_net), .O(n682_adj_4546));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i459_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_11_i24_3_lut (.I0(n16_adj_4647), .I1(n535[22]), .I2(n45_adj_4627), 
            .I3(GND_net), .O(n24_adj_4650));   // verilog/motorControl.v(47[25:43])
    defparam LessThan_11_i24_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_24_i508_2_lut (.I0(\Ki[10] ), .I1(n351), .I2(GND_net), 
            .I3(GND_net), .O(n755_adj_4545));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i508_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i557_2_lut (.I0(\Ki[11] ), .I1(n351), .I2(GND_net), 
            .I3(GND_net), .O(n828_adj_4544));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i557_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i606_2_lut (.I0(\Ki[12] ), .I1(n351), .I2(GND_net), 
            .I3(GND_net), .O(n901_adj_4543));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i606_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i79_2_lut (.I0(\Ki[1] ), .I1(n345), .I2(GND_net), 
            .I3(GND_net), .O(n116_adj_4542));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i79_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i32_2_lut (.I0(\Ki[0] ), .I1(n344), .I2(GND_net), 
            .I3(GND_net), .O(n47_adj_4541));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i32_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i655_2_lut (.I0(\Ki[13] ), .I1(n351), .I2(GND_net), 
            .I3(GND_net), .O(n974_adj_4540));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i655_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i128_2_lut (.I0(\Ki[2] ), .I1(n345), .I2(GND_net), 
            .I3(GND_net), .O(n189_adj_4539));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i128_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i45693_4_lut (.I0(n43_adj_4628), .I1(n25_adj_4632), .I2(n23_adj_4631), 
            .I3(n60501), .O(n60405));
    defparam i45693_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 mult_24_i704_2_lut (.I0(\Ki[14] ), .I1(n351), .I2(GND_net), 
            .I3(GND_net), .O(n1047_adj_4538));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i704_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i177_2_lut (.I0(\Ki[3] ), .I1(n345), .I2(GND_net), 
            .I3(GND_net), .O(n262_adj_4537));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i177_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i753_2_lut (.I0(\Ki[15] ), .I1(n351), .I2(GND_net), 
            .I3(GND_net), .O(n1120_adj_4536));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i753_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i226_2_lut (.I0(\Ki[4] ), .I1(n345), .I2(GND_net), 
            .I3(GND_net), .O(n335_adj_4535));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i226_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i275_2_lut (.I0(\Ki[5] ), .I1(n345), .I2(GND_net), 
            .I3(GND_net), .O(n408_adj_4534));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i275_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i79_2_lut (.I0(\Kp[1] ), .I1(n207[18]), .I2(GND_net), 
            .I3(GND_net), .O(n116));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i79_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i32_2_lut (.I0(\Kp[0] ), .I1(n207[19]), .I2(GND_net), 
            .I3(GND_net), .O(n47_adj_4533));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i32_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i47162_4_lut (.I0(n24_adj_4650), .I1(n8_adj_4649), .I2(n45_adj_4627), 
            .I3(n60401), .O(n61875));   // verilog/motorControl.v(47[25:43])
    defparam i47162_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 mult_24_i324_2_lut (.I0(\Ki[6] ), .I1(n345), .I2(GND_net), 
            .I3(GND_net), .O(n481_adj_4532));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i324_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i46396_3_lut (.I0(n62365), .I1(n535[12]), .I2(n25_adj_4632), 
            .I3(GND_net), .O(n61109));   // verilog/motorControl.v(47[25:43])
    defparam i46396_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 unary_minus_27_inv_0_i7_1_lut (.I0(\deadband[6] ), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n28[6]));   // verilog/motorControl.v(62[45:54])
    defparam unary_minus_27_inv_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_27_inv_0_i8_1_lut (.I0(\deadband[7] ), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n28[7]));   // verilog/motorControl.v(62[45:54])
    defparam unary_minus_27_inv_0_i8_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_24_i373_2_lut (.I0(\Ki[7] ), .I1(n345), .I2(GND_net), 
            .I3(GND_net), .O(n554_adj_4529));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i373_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_27_inv_0_i9_1_lut (.I0(\deadband[8] ), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n28[8]));   // verilog/motorControl.v(62[45:54])
    defparam unary_minus_27_inv_0_i9_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_23_i128_2_lut (.I0(\Kp[2] ), .I1(n207[18]), .I2(GND_net), 
            .I3(GND_net), .O(n189));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i128_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i422_2_lut (.I0(\Ki[8] ), .I1(n345), .I2(GND_net), 
            .I3(GND_net), .O(n627_adj_4527));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i422_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_11_i4_4_lut (.I0(setpoint[0]), .I1(n535[1]), .I2(setpoint[1]), 
            .I3(n535[0]), .O(n4_adj_4651));   // verilog/motorControl.v(47[25:43])
    defparam LessThan_11_i4_4_lut.LUT_INIT = 16'h4d0c;
    SB_LUT4 i47647_3_lut (.I0(n4_adj_4651), .I1(n535[13]), .I2(n27_adj_4639), 
            .I3(GND_net), .O(n62360));   // verilog/motorControl.v(47[25:43])
    defparam i47647_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_24_i471_2_lut (.I0(\Ki[9] ), .I1(n345), .I2(GND_net), 
            .I3(GND_net), .O(n700_adj_4526));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i471_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i47648_3_lut (.I0(n62360), .I1(n535[14]), .I2(n29_adj_4629), 
            .I3(GND_net), .O(n62361));   // verilog/motorControl.v(47[25:43])
    defparam i47648_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_23_i177_2_lut (.I0(\Kp[3] ), .I1(n207[18]), .I2(GND_net), 
            .I3(GND_net), .O(n262));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i177_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_27_inv_0_i10_1_lut (.I0(\deadband[9] ), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n28[9]));   // verilog/motorControl.v(62[45:54])
    defparam unary_minus_27_inv_0_i10_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_27_inv_0_i11_1_lut (.I0(\deadband[10] ), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n28[10]));   // verilog/motorControl.v(62[45:54])
    defparam unary_minus_27_inv_0_i11_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_23_i226_2_lut (.I0(\Kp[4] ), .I1(n207[18]), .I2(GND_net), 
            .I3(GND_net), .O(n335));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i226_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i55_2_lut (.I0(\Kp[1] ), .I1(n207[6]), .I2(GND_net), 
            .I3(GND_net), .O(n80_adj_4523));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i55_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i45733_4_lut (.I0(n33_adj_4635), .I1(n31_adj_4630), .I2(n29_adj_4629), 
            .I3(n60479), .O(n60445));
    defparam i45733_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i48034_4_lut (.I0(n30_adj_4646), .I1(n10_adj_4645), .I2(n35_adj_4634), 
            .I3(n60441), .O(n62747));   // verilog/motorControl.v(47[25:43])
    defparam i48034_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 mult_23_i8_2_lut (.I0(\Kp[0] ), .I1(n207[7]), .I2(GND_net), 
            .I3(GND_net), .O(n11_adj_4522));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i8_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i46398_3_lut (.I0(n62361), .I1(n535[15]), .I2(n31_adj_4630), 
            .I3(GND_net), .O(n61111));   // verilog/motorControl.v(47[25:43])
    defparam i46398_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i48252_4_lut (.I0(n61111), .I1(n62747), .I2(n35_adj_4634), 
            .I3(n60445), .O(n62965));   // verilog/motorControl.v(47[25:43])
    defparam i48252_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 mult_23_i275_2_lut (.I0(\Kp[5] ), .I1(n207[18]), .I2(GND_net), 
            .I3(GND_net), .O(n408));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i275_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i48253_3_lut (.I0(n62965), .I1(n535[18]), .I2(n37_adj_4633), 
            .I3(GND_net), .O(n62966));   // verilog/motorControl.v(47[25:43])
    defparam i48253_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_23_i104_2_lut (.I0(\Kp[2] ), .I1(n207[6]), .I2(GND_net), 
            .I3(GND_net), .O(n153_adj_4521));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i104_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i153_2_lut (.I0(\Kp[3] ), .I1(n207[6]), .I2(GND_net), 
            .I3(GND_net), .O(n226_adj_4520));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i153_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i202_2_lut (.I0(\Kp[4] ), .I1(n207[6]), .I2(GND_net), 
            .I3(GND_net), .O(n299_adj_4519));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i202_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_27_inv_0_i12_1_lut (.I0(\deadband[11] ), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n28[11]));   // verilog/motorControl.v(62[45:54])
    defparam unary_minus_27_inv_0_i12_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_27_inv_0_i13_1_lut (.I0(\deadband[12] ), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n28[12]));   // verilog/motorControl.v(62[45:54])
    defparam unary_minus_27_inv_0_i13_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_23_i324_2_lut (.I0(\Kp[6] ), .I1(n207[18]), .I2(GND_net), 
            .I3(GND_net), .O(n481));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i324_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i251_2_lut (.I0(\Kp[5] ), .I1(n207[6]), .I2(GND_net), 
            .I3(GND_net), .O(n372_adj_4516));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i251_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i373_2_lut (.I0(\Kp[7] ), .I1(n207[18]), .I2(GND_net), 
            .I3(GND_net), .O(n554_adj_4515));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i373_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i48194_3_lut (.I0(n62966), .I1(n535[19]), .I2(n39_adj_4626), 
            .I3(GND_net), .O(n62907));   // verilog/motorControl.v(47[25:43])
    defparam i48194_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_23_i300_2_lut (.I0(\Kp[6] ), .I1(n207[6]), .I2(GND_net), 
            .I3(GND_net), .O(n445_adj_4514));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i300_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_27_inv_0_i14_1_lut (.I0(\deadband[13] ), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n28[13]));   // verilog/motorControl.v(62[45:54])
    defparam unary_minus_27_inv_0_i14_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_23_i349_2_lut (.I0(\Kp[7] ), .I1(n207[6]), .I2(GND_net), 
            .I3(GND_net), .O(n518_adj_4512));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i349_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i422_2_lut (.I0(\Kp[8] ), .I1(n207[18]), .I2(GND_net), 
            .I3(GND_net), .O(n627));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i422_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i398_2_lut (.I0(\Kp[8] ), .I1(n207[6]), .I2(GND_net), 
            .I3(GND_net), .O(n591_adj_4511));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i398_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i447_2_lut (.I0(\Kp[9] ), .I1(n207[6]), .I2(GND_net), 
            .I3(GND_net), .O(n664_adj_4510));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i447_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_27_inv_0_i15_1_lut (.I0(\deadband[14] ), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n28[14]));   // verilog/motorControl.v(62[45:54])
    defparam unary_minus_27_inv_0_i15_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i45700_4_lut (.I0(n43_adj_4628), .I1(n41_adj_4625), .I2(n39_adj_4626), 
            .I3(n62810), .O(n60412));
    defparam i45700_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 unary_minus_27_inv_0_i16_1_lut (.I0(\deadband[15] ), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n28[15]));   // verilog/motorControl.v(62[45:54])
    defparam unary_minus_27_inv_0_i16_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i47838_4_lut (.I0(n61109), .I1(n61875), .I2(n45_adj_4627), 
            .I3(n60405), .O(n62551));   // verilog/motorControl.v(47[25:43])
    defparam i47838_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 mult_23_i496_2_lut (.I0(\Kp[10] ), .I1(n207[6]), .I2(GND_net), 
            .I3(GND_net), .O(n737_adj_4506));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i496_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_27_inv_0_i17_1_lut (.I0(\deadband[16] ), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n28[16]));   // verilog/motorControl.v(62[45:54])
    defparam unary_minus_27_inv_0_i17_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_23_i471_2_lut (.I0(\Kp[9] ), .I1(n207[18]), .I2(GND_net), 
            .I3(GND_net), .O(n700));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i471_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i545_2_lut (.I0(\Kp[11] ), .I1(n207[6]), .I2(GND_net), 
            .I3(GND_net), .O(n810_adj_4504));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i545_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i65_2_lut (.I0(\Ki[1] ), .I1(n352), .I2(GND_net), 
            .I3(GND_net), .O(n95_adj_4503));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i65_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i18_2_lut (.I0(\Ki[0] ), .I1(n351), .I2(GND_net), 
            .I3(GND_net), .O(n26_adj_4502));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i18_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i46404_3_lut (.I0(n62907), .I1(n535[20]), .I2(n41_adj_4625), 
            .I3(GND_net), .O(n61117));   // verilog/motorControl.v(47[25:43])
    defparam i46404_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_23_i594_2_lut (.I0(\Kp[12] ), .I1(n207[6]), .I2(GND_net), 
            .I3(GND_net), .O(n883_adj_4501));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i594_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i48038_4_lut (.I0(n61117), .I1(n62551), .I2(n45_adj_4627), 
            .I3(n60412), .O(n62751));   // verilog/motorControl.v(47[25:43])
    defparam i48038_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 mult_24_i114_2_lut (.I0(\Ki[2] ), .I1(n352), .I2(GND_net), 
            .I3(GND_net), .O(n168_adj_4500));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i114_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i643_2_lut (.I0(\Kp[13] ), .I1(n207[6]), .I2(GND_net), 
            .I3(GND_net), .O(n956_adj_4499));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i643_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_27_inv_0_i18_1_lut (.I0(\deadband[17] ), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n28[17]));   // verilog/motorControl.v(62[45:54])
    defparam unary_minus_27_inv_0_i18_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_24_i163_2_lut (.I0(\Ki[3] ), .I1(n352), .I2(GND_net), 
            .I3(GND_net), .O(n241_adj_4497));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i163_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i48039_3_lut (.I0(n62751), .I1(setpoint[23]), .I2(n535[23]), 
            .I3(GND_net), .O(n131));   // verilog/motorControl.v(47[25:43])
    defparam i48039_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 mult_23_i692_2_lut (.I0(\Kp[14] ), .I1(n207[6]), .I2(GND_net), 
            .I3(GND_net), .O(n1029_adj_4496));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i692_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_27_inv_0_i19_1_lut (.I0(\deadband[18] ), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n28[18]));   // verilog/motorControl.v(62[45:54])
    defparam unary_minus_27_inv_0_i19_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 LessThan_30_i41_2_lut (.I0(PWMLimit[20]), .I1(n455[20]), .I2(GND_net), 
            .I3(GND_net), .O(n41_adj_4652));   // verilog/motorControl.v(63[16:31])
    defparam LessThan_30_i41_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_24_i212_2_lut (.I0(\Ki[4] ), .I1(n352), .I2(GND_net), 
            .I3(GND_net), .O(n314_adj_4493));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i212_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i741_2_lut (.I0(\Kp[15] ), .I1(n207[6]), .I2(GND_net), 
            .I3(GND_net), .O(n1102_adj_4492));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i741_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i261_2_lut (.I0(\Ki[5] ), .I1(n352), .I2(GND_net), 
            .I3(GND_net), .O(n387_adj_4491));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i261_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_27_inv_0_i20_1_lut (.I0(\deadband[19] ), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n28[19]));   // verilog/motorControl.v(62[45:54])
    defparam unary_minus_27_inv_0_i20_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_27_inv_0_i21_1_lut (.I0(\deadband[20] ), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n28[20]));   // verilog/motorControl.v(62[45:54])
    defparam unary_minus_27_inv_0_i21_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_27_inv_0_i22_1_lut (.I0(\deadband[21] ), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n28[21]));   // verilog/motorControl.v(62[45:54])
    defparam unary_minus_27_inv_0_i22_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_27_inv_0_i23_1_lut (.I0(\deadband[22] ), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n28[22]));   // verilog/motorControl.v(62[45:54])
    defparam unary_minus_27_inv_0_i23_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 LessThan_30_i39_2_lut (.I0(PWMLimit[19]), .I1(n455[19]), .I2(GND_net), 
            .I3(GND_net), .O(n39_adj_4653));   // verilog/motorControl.v(63[16:31])
    defparam LessThan_30_i39_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_30_i45_2_lut (.I0(PWMLimit[22]), .I1(n455[22]), .I2(GND_net), 
            .I3(GND_net), .O(n45_adj_4654));   // verilog/motorControl.v(63[16:31])
    defparam LessThan_30_i45_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_23_i85_2_lut (.I0(\Kp[1] ), .I1(n207[21]), .I2(GND_net), 
            .I3(GND_net), .O(n125_adj_4485));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i85_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i38_2_lut (.I0(\Kp[0] ), .I1(n207[22]), .I2(GND_net), 
            .I3(GND_net), .O(n56_adj_4484));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i38_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_27_inv_0_i24_1_lut (.I0(\deadband[23] ), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n28[23]));   // verilog/motorControl.v(62[45:54])
    defparam unary_minus_27_inv_0_i24_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_24_i2_2_lut (.I0(\Ki[0] ), .I1(n359), .I2(GND_net), .I3(GND_net), 
            .O(n42[0]));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i2_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i2_2_lut (.I0(\Kp[0] ), .I1(n207[4]), .I2(GND_net), 
            .I3(GND_net), .O(n360[0]));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i2_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_33_inv_0_i1_1_lut (.I0(PWMLimit[0]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n46[0]));   // verilog/motorControl.v(66[24:33])
    defparam unary_minus_33_inv_0_i1_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_23_i134_2_lut (.I0(\Kp[2] ), .I1(n207[21]), .I2(GND_net), 
            .I3(GND_net), .O(n198_adj_4481));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i134_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_30_i43_2_lut (.I0(PWMLimit[21]), .I1(n455[21]), .I2(GND_net), 
            .I3(GND_net), .O(n43_adj_4655));   // verilog/motorControl.v(63[16:31])
    defparam LessThan_30_i43_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_30_i37_2_lut (.I0(PWMLimit[18]), .I1(n455[18]), .I2(GND_net), 
            .I3(GND_net), .O(n37_adj_4656));   // verilog/motorControl.v(63[16:31])
    defparam LessThan_30_i37_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 unary_minus_33_inv_0_i2_1_lut (.I0(PWMLimit[1]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n46[1]));   // verilog/motorControl.v(66[24:33])
    defparam unary_minus_33_inv_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_23_i183_2_lut (.I0(\Kp[3] ), .I1(n207[21]), .I2(GND_net), 
            .I3(GND_net), .O(n271_adj_4479));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i183_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1_4_lut_adj_934 (.I0(n207[23]), .I1(\Kp[2] ), .I2(n45802), 
            .I3(n207[22]), .O(n56550));   // verilog/motorControl.v(61[20:26])
    defparam i1_4_lut_adj_934.LUT_INIT = 16'h6ca0;
    SB_LUT4 mult_23_i232_2_lut (.I0(\Kp[4] ), .I1(n207[21]), .I2(GND_net), 
            .I3(GND_net), .O(n344_adj_4478));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i232_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_30_i23_2_lut (.I0(PWMLimit[11]), .I1(n455[11]), .I2(GND_net), 
            .I3(GND_net), .O(n23_adj_4657));   // verilog/motorControl.v(63[16:31])
    defparam LessThan_30_i23_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_4_lut_adj_935 (.I0(n207[22]), .I1(n18009[1]), .I2(n4_adj_4658), 
            .I3(\Kp[3] ), .O(n17961[2]));   // verilog/motorControl.v(61[20:26])
    defparam i1_4_lut_adj_935.LUT_INIT = 16'hc66c;
    SB_LUT4 LessThan_30_i25_2_lut (.I0(PWMLimit[12]), .I1(n455[12]), .I2(GND_net), 
            .I3(GND_net), .O(n25_adj_4659));   // verilog/motorControl.v(63[16:31])
    defparam LessThan_30_i25_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_23_i281_2_lut (.I0(\Kp[5] ), .I1(n207[21]), .I2(GND_net), 
            .I3(GND_net), .O(n417_adj_4477));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i281_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i234_2_lut (.I0(\Kp[4] ), .I1(n207[22]), .I2(GND_net), 
            .I3(GND_net), .O(n347_c));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i234_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1_4_lut_adj_936 (.I0(n18009[1]), .I1(n6_adj_4660), .I2(n347_c), 
            .I3(n53040), .O(n17961[3]));   // verilog/motorControl.v(61[20:26])
    defparam i1_4_lut_adj_936.LUT_INIT = 16'h6996;
    SB_LUT4 unary_minus_33_inv_0_i3_1_lut (.I0(PWMLimit[2]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n46[2]));   // verilog/motorControl.v(66[24:33])
    defparam unary_minus_33_inv_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 LessThan_30_i29_2_lut (.I0(PWMLimit[14]), .I1(n455[14]), .I2(GND_net), 
            .I3(GND_net), .O(n29_adj_4661));   // verilog/motorControl.v(63[16:31])
    defparam LessThan_30_i29_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_3_lut (.I0(\Kp[0] ), .I1(\Kp[2] ), .I2(\Kp[1] ), .I3(GND_net), 
            .O(n56546));   // verilog/motorControl.v(61[20:26])
    defparam i1_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i1_2_lut (.I0(n56546), .I1(n207[23]), .I2(GND_net), .I3(GND_net), 
            .O(n4_adj_4658));   // verilog/motorControl.v(61[20:26])
    defparam i1_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i32508_4_lut (.I0(n18009[1]), .I1(\Kp[3] ), .I2(n4_adj_4658), 
            .I3(n207[22]), .O(n6_adj_4660));   // verilog/motorControl.v(61[20:26])
    defparam i32508_4_lut.LUT_INIT = 16'he800;
    SB_LUT4 mult_23_i46_2_lut (.I0(\Kp[0] ), .I1(n207[23]), .I2(GND_net), 
            .I3(GND_net), .O(n68_adj_4662));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i46_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i32446_2_lut (.I0(\Kp[0] ), .I1(\Kp[1] ), .I2(GND_net), .I3(GND_net), 
            .O(n45802));   // verilog/motorControl.v(61[20:26])
    defparam i32446_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_30_i31_2_lut (.I0(PWMLimit[15]), .I1(n455[15]), .I2(GND_net), 
            .I3(GND_net), .O(n31_adj_4663));   // verilog/motorControl.v(63[16:31])
    defparam LessThan_30_i31_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i41938_3_lut (.I0(n207[23]), .I1(n56546), .I2(\Kp[3] ), .I3(GND_net), 
            .O(n53040));   // verilog/motorControl.v(61[20:26])
    defparam i41938_3_lut.LUT_INIT = 16'h2828;
    SB_LUT4 i32455_3_lut (.I0(n207[23]), .I1(n45797), .I2(n47176), .I3(GND_net), 
            .O(n18009[1]));   // verilog/motorControl.v(61[20:26])
    defparam i32455_3_lut.LUT_INIT = 16'h6c6c;
    SB_LUT4 mult_23_i330_2_lut (.I0(\Kp[6] ), .I1(n207[21]), .I2(GND_net), 
            .I3(GND_net), .O(n490_adj_4474));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i330_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1_4_lut_adj_937 (.I0(n207[23]), .I1(\Kp[5] ), .I2(n47176), 
            .I3(n207[22]), .O(n56536));   // verilog/motorControl.v(61[20:26])
    defparam i1_4_lut_adj_937.LUT_INIT = 16'hc60a;
    SB_LUT4 i1_rep_584_2_lut (.I0(n18009[1]), .I1(n53040), .I2(GND_net), 
            .I3(GND_net), .O(n64292));   // verilog/motorControl.v(61[20:26])
    defparam i1_rep_584_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_4_lut_adj_938 (.I0(n45797), .I1(n56536), .I2(\Kp[4] ), 
            .I3(n207[23]), .O(n56540));   // verilog/motorControl.v(61[20:26])
    defparam i1_4_lut_adj_938.LUT_INIT = 16'h9666;
    SB_LUT4 i32516_4_lut (.I0(n64292), .I1(\Kp[4] ), .I2(n6_adj_4660), 
            .I3(n207[22]), .O(n8_adj_4664));   // verilog/motorControl.v(61[20:26])
    defparam i32516_4_lut.LUT_INIT = 16'he8a0;
    SB_LUT4 i32469_4_lut (.I0(n18009[1]), .I1(\Kp[3] ), .I2(n56546), .I3(n207[23]), 
            .O(n6_adj_4665));   // verilog/motorControl.v(61[20:26])
    defparam i32469_4_lut.LUT_INIT = 16'he800;
    SB_LUT4 i1_4_lut_adj_939 (.I0(n6_adj_4665), .I1(n8_adj_4664), .I2(n56540), 
            .I3(n53040), .O(n54612));   // verilog/motorControl.v(61[20:26])
    defparam i1_4_lut_adj_939.LUT_INIT = 16'h6996;
    SB_LUT4 LessThan_30_i35_2_lut (.I0(PWMLimit[17]), .I1(n455[17]), .I2(GND_net), 
            .I3(GND_net), .O(n35_adj_4666));   // verilog/motorControl.v(63[16:31])
    defparam LessThan_30_i35_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_24_i310_2_lut (.I0(\Ki[6] ), .I1(n352), .I2(GND_net), 
            .I3(GND_net), .O(n460_adj_4473));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i310_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i53_2_lut (.I0(\Kp[1] ), .I1(n207[5]), .I2(GND_net), 
            .I3(GND_net), .O(n77_adj_4472));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i53_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i6_2_lut (.I0(\Kp[0] ), .I1(n207[6]), .I2(GND_net), 
            .I3(GND_net), .O(n8_adj_4471));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i6_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i359_2_lut (.I0(\Ki[7] ), .I1(n352), .I2(GND_net), 
            .I3(GND_net), .O(n533_adj_4470));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i359_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i408_2_lut (.I0(\Ki[8] ), .I1(n352), .I2(GND_net), 
            .I3(GND_net), .O(n606_adj_4469));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i408_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i102_2_lut (.I0(\Kp[2] ), .I1(n207[5]), .I2(GND_net), 
            .I3(GND_net), .O(n150_adj_4467));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i102_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_33_inv_0_i4_1_lut (.I0(PWMLimit[3]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n46[3]));   // verilog/motorControl.v(66[24:33])
    defparam unary_minus_33_inv_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_33_inv_0_i5_1_lut (.I0(PWMLimit[4]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n46[4]));   // verilog/motorControl.v(66[24:33])
    defparam unary_minus_33_inv_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_33_inv_0_i6_1_lut (.I0(PWMLimit[5]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n46[5]));   // verilog/motorControl.v(66[24:33])
    defparam unary_minus_33_inv_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 LessThan_30_i33_2_lut (.I0(PWMLimit[16]), .I1(n455[16]), .I2(GND_net), 
            .I3(GND_net), .O(n33_adj_4667));   // verilog/motorControl.v(63[16:31])
    defparam LessThan_30_i33_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 unary_minus_33_inv_0_i7_1_lut (.I0(PWMLimit[6]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n46[6]));   // verilog/motorControl.v(66[24:33])
    defparam unary_minus_33_inv_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_23_i151_2_lut (.I0(\Kp[3] ), .I1(n207[5]), .I2(GND_net), 
            .I3(GND_net), .O(n223_adj_4461));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i151_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_30_i11_2_lut (.I0(PWMLimit[5]), .I1(n455[5]), .I2(GND_net), 
            .I3(GND_net), .O(n11_adj_4668));   // verilog/motorControl.v(63[16:31])
    defparam LessThan_30_i11_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_30_i13_2_lut (.I0(PWMLimit[6]), .I1(n455[6]), .I2(GND_net), 
            .I3(GND_net), .O(n13_adj_4669));   // verilog/motorControl.v(63[16:31])
    defparam LessThan_30_i13_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_24_i457_2_lut (.I0(\Ki[9] ), .I1(n352), .I2(GND_net), 
            .I3(GND_net), .O(n679_adj_4460));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i457_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_30_i15_2_lut (.I0(PWMLimit[7]), .I1(n455[7]), .I2(GND_net), 
            .I3(GND_net), .O(n15_adj_4670));   // verilog/motorControl.v(63[16:31])
    defparam LessThan_30_i15_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_23_i200_2_lut (.I0(\Kp[4] ), .I1(n207[5]), .I2(GND_net), 
            .I3(GND_net), .O(n296_adj_4459));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i200_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i506_2_lut (.I0(\Ki[10] ), .I1(n352), .I2(GND_net), 
            .I3(GND_net), .O(n752_adj_4458));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i506_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i249_2_lut (.I0(\Kp[5] ), .I1(n207[5]), .I2(GND_net), 
            .I3(GND_net), .O(n369_adj_4457));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i249_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i555_2_lut (.I0(\Ki[11] ), .I1(n352), .I2(GND_net), 
            .I3(GND_net), .O(n825_adj_4456));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i555_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i298_2_lut (.I0(\Kp[6] ), .I1(n207[5]), .I2(GND_net), 
            .I3(GND_net), .O(n442_adj_4455));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i298_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_30_i27_2_lut (.I0(PWMLimit[13]), .I1(n455[13]), .I2(GND_net), 
            .I3(GND_net), .O(n27_adj_4671));   // verilog/motorControl.v(63[16:31])
    defparam LessThan_30_i27_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_23_i347_2_lut (.I0(\Kp[7] ), .I1(n207[5]), .I2(GND_net), 
            .I3(GND_net), .O(n515_adj_4454));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i347_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i396_2_lut (.I0(\Kp[8] ), .I1(n207[5]), .I2(GND_net), 
            .I3(GND_net), .O(n588_adj_4453));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i396_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_33_inv_0_i8_1_lut (.I0(PWMLimit[7]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n46[7]));   // verilog/motorControl.v(66[24:33])
    defparam unary_minus_33_inv_0_i8_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 LessThan_30_i9_2_lut (.I0(PWMLimit[4]), .I1(n455[4]), .I2(GND_net), 
            .I3(GND_net), .O(n9_adj_4672));   // verilog/motorControl.v(63[16:31])
    defparam LessThan_30_i9_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_30_i17_2_lut (.I0(PWMLimit[8]), .I1(n455[8]), .I2(GND_net), 
            .I3(GND_net), .O(n17_adj_4673));   // verilog/motorControl.v(63[16:31])
    defparam LessThan_30_i17_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 unary_minus_33_inv_0_i9_1_lut (.I0(PWMLimit[8]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n46[8]));   // verilog/motorControl.v(66[24:33])
    defparam unary_minus_33_inv_0_i9_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_24_i610_2_lut (.I0(\Ki[12] ), .I1(n349), .I2(GND_net), 
            .I3(GND_net), .O(n907_adj_4210));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i610_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i445_2_lut (.I0(\Kp[9] ), .I1(n207[5]), .I2(GND_net), 
            .I3(GND_net), .O(n661_adj_4450));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i445_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_33_inv_0_i10_1_lut (.I0(PWMLimit[9]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n46[9]));   // verilog/motorControl.v(66[24:33])
    defparam unary_minus_33_inv_0_i10_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 LessThan_30_i19_2_lut (.I0(PWMLimit[9]), .I1(n455[9]), .I2(GND_net), 
            .I3(GND_net), .O(n19_adj_4674));   // verilog/motorControl.v(63[16:31])
    defparam LessThan_30_i19_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_23_i494_2_lut (.I0(\Kp[10] ), .I1(n207[5]), .I2(GND_net), 
            .I3(GND_net), .O(n734_adj_4448));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i494_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i604_2_lut (.I0(\Ki[12] ), .I1(n352), .I2(GND_net), 
            .I3(GND_net), .O(n898_adj_4447));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i604_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i543_2_lut (.I0(\Kp[11] ), .I1(n207[5]), .I2(GND_net), 
            .I3(GND_net), .O(n807_adj_4446));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i543_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i653_2_lut (.I0(\Ki[13] ), .I1(n352), .I2(GND_net), 
            .I3(GND_net), .O(n971_adj_4445));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i653_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_33_inv_0_i11_1_lut (.I0(PWMLimit[10]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n46[10]));   // verilog/motorControl.v(66[24:33])
    defparam unary_minus_33_inv_0_i11_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 LessThan_30_i21_2_lut (.I0(PWMLimit[10]), .I1(n455[10]), .I2(GND_net), 
            .I3(GND_net), .O(n21_adj_4675));   // verilog/motorControl.v(63[16:31])
    defparam LessThan_30_i21_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_23_i592_2_lut (.I0(\Kp[12] ), .I1(n207[5]), .I2(GND_net), 
            .I3(GND_net), .O(n880_adj_4443));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i592_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i702_2_lut (.I0(\Ki[14] ), .I1(n352), .I2(GND_net), 
            .I3(GND_net), .O(n1044_adj_4442));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i702_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i641_2_lut (.I0(\Kp[13] ), .I1(n207[5]), .I2(GND_net), 
            .I3(GND_net), .O(n953_adj_4441));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i641_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i751_2_lut (.I0(\Ki[15] ), .I1(n352), .I2(GND_net), 
            .I3(GND_net), .O(n1117_adj_4440));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i751_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i690_2_lut (.I0(\Kp[14] ), .I1(n207[5]), .I2(GND_net), 
            .I3(GND_net), .O(n1026_adj_4439));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i690_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_33_inv_0_i12_1_lut (.I0(PWMLimit[11]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n46[11]));   // verilog/motorControl.v(66[24:33])
    defparam unary_minus_33_inv_0_i12_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_33_inv_0_i13_1_lut (.I0(PWMLimit[12]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n46[12]));   // verilog/motorControl.v(66[24:33])
    defparam unary_minus_33_inv_0_i13_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i45998_4_lut (.I0(n21_adj_4675), .I1(n19_adj_4674), .I2(n17_adj_4673), 
            .I3(n9_adj_4672), .O(n60710));
    defparam i45998_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 unary_minus_33_inv_0_i14_1_lut (.I0(PWMLimit[13]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n46[13]));   // verilog/motorControl.v(66[24:33])
    defparam unary_minus_33_inv_0_i14_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_33_inv_0_i15_1_lut (.I0(PWMLimit[14]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n46[14]));   // verilog/motorControl.v(66[24:33])
    defparam unary_minus_33_inv_0_i15_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i45988_4_lut (.I0(n27_adj_4671), .I1(n15_adj_4670), .I2(n13_adj_4669), 
            .I3(n11_adj_4668), .O(n60700));
    defparam i45988_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 LessThan_30_i12_3_lut (.I0(n455[7]), .I1(n455[16]), .I2(n33_adj_4667), 
            .I3(GND_net), .O(n12_adj_4676));   // verilog/motorControl.v(63[16:31])
    defparam LessThan_30_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_23_i739_2_lut (.I0(\Kp[15] ), .I1(n207[5]), .I2(GND_net), 
            .I3(GND_net), .O(n1099_adj_4434));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i739_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_21_i17_3_lut (.I0(n233[16]), .I1(n285[16]), .I2(n284), 
            .I3(GND_net), .O(n310[16]));   // verilog/motorControl.v(58[20] 60[14])
    defparam mux_21_i17_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_24_i63_2_lut (.I0(\Ki[1] ), .I1(n353), .I2(GND_net), 
            .I3(GND_net), .O(n92_adj_4433));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i63_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i16_2_lut (.I0(\Ki[0] ), .I1(n352), .I2(GND_net), 
            .I3(GND_net), .O(n23_adj_4432));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i16_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i112_2_lut (.I0(\Ki[2] ), .I1(n353), .I2(GND_net), 
            .I3(GND_net), .O(n165_adj_4431));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i112_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_30_i10_3_lut (.I0(n455[5]), .I1(n455[6]), .I2(n13_adj_4669), 
            .I3(GND_net), .O(n10_adj_4677));   // verilog/motorControl.v(63[16:31])
    defparam LessThan_30_i10_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_24_i161_2_lut (.I0(\Ki[3] ), .I1(n353), .I2(GND_net), 
            .I3(GND_net), .O(n238_adj_4430));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i161_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i210_2_lut (.I0(\Ki[4] ), .I1(n353), .I2(GND_net), 
            .I3(GND_net), .O(n311_adj_4429));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i210_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_30_i30_3_lut (.I0(n12_adj_4676), .I1(n455[17]), .I2(n35_adj_4666), 
            .I3(GND_net), .O(n30_adj_4678));   // verilog/motorControl.v(63[16:31])
    defparam LessThan_30_i30_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 unary_minus_33_inv_0_i16_1_lut (.I0(PWMLimit[15]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n46[15]));   // verilog/motorControl.v(66[24:33])
    defparam unary_minus_33_inv_0_i16_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_33_inv_0_i17_1_lut (.I0(PWMLimit[16]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n46[16]));   // verilog/motorControl.v(66[24:33])
    defparam unary_minus_33_inv_0_i17_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_33_inv_0_i18_1_lut (.I0(PWMLimit[17]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n46[17]));   // verilog/motorControl.v(66[24:33])
    defparam unary_minus_33_inv_0_i18_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i46950_4_lut (.I0(n13_adj_4669), .I1(n11_adj_4668), .I2(n9_adj_4672), 
            .I3(n60732), .O(n61663));
    defparam i46950_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 unary_minus_33_inv_0_i19_1_lut (.I0(PWMLimit[18]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n46[18]));   // verilog/motorControl.v(66[24:33])
    defparam unary_minus_33_inv_0_i19_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_33_inv_0_i20_1_lut (.I0(PWMLimit[19]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n46[19]));   // verilog/motorControl.v(66[24:33])
    defparam unary_minus_33_inv_0_i20_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i46944_4_lut (.I0(n19_adj_4674), .I1(n17_adj_4673), .I2(n15_adj_4670), 
            .I3(n61663), .O(n61657));
    defparam i46944_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 unary_minus_33_inv_0_i21_1_lut (.I0(PWMLimit[20]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n46[20]));   // verilog/motorControl.v(66[24:33])
    defparam unary_minus_33_inv_0_i21_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i47996_4_lut (.I0(n25_adj_4659), .I1(n23_adj_4657), .I2(n21_adj_4675), 
            .I3(n61657), .O(n62709));
    defparam i47996_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 mux_22_i17_3_lut (.I0(n310[16]), .I1(IntegralLimit[16]), .I2(n258), 
            .I3(GND_net), .O(n343));   // verilog/motorControl.v(58[20] 60[14])
    defparam mux_22_i17_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_24_i259_2_lut (.I0(\Ki[5] ), .I1(n353), .I2(GND_net), 
            .I3(GND_net), .O(n384_adj_4422));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i259_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i51_2_lut (.I0(\Kp[1] ), .I1(n207[4]), .I2(GND_net), 
            .I3(GND_net), .O(n74_adj_4421));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i51_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i47377_4_lut (.I0(n31_adj_4663), .I1(n29_adj_4661), .I2(n27_adj_4671), 
            .I3(n62709), .O(n62090));
    defparam i47377_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i48113_4_lut (.I0(n37_adj_4656), .I1(n35_adj_4666), .I2(n33_adj_4667), 
            .I3(n62090), .O(n62826));
    defparam i48113_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 mult_24_i81_2_lut (.I0(\Ki[1] ), .I1(n344), .I2(GND_net), 
            .I3(GND_net), .O(n119_adj_4209));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i81_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i4_2_lut (.I0(\Kp[0] ), .I1(n207[5]), .I2(GND_net), 
            .I3(GND_net), .O(n5_adj_4420));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i4_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_30_i16_3_lut (.I0(n455[9]), .I1(n455[21]), .I2(n43_adj_4655), 
            .I3(GND_net), .O(n16_adj_4679));   // verilog/motorControl.v(63[16:31])
    defparam LessThan_30_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_24_i308_2_lut (.I0(\Ki[6] ), .I1(n353), .I2(GND_net), 
            .I3(GND_net), .O(n457_adj_4419));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i308_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i100_2_lut (.I0(\Kp[2] ), .I1(n207[4]), .I2(GND_net), 
            .I3(GND_net), .O(n147_adj_4418));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i100_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i47571_3_lut (.I0(n6_adj_4680), .I1(n455[10]), .I2(n21_adj_4675), 
            .I3(GND_net), .O(n62284));   // verilog/motorControl.v(63[16:31])
    defparam i47571_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 unary_minus_33_inv_0_i22_1_lut (.I0(PWMLimit[21]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n46[21]));   // verilog/motorControl.v(66[24:33])
    defparam unary_minus_33_inv_0_i22_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_23_i149_2_lut (.I0(\Kp[3] ), .I1(n207[4]), .I2(GND_net), 
            .I3(GND_net), .O(n220_adj_4415));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i149_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i47572_3_lut (.I0(n62284), .I1(n455[11]), .I2(n23_adj_4657), 
            .I3(GND_net), .O(n62285));   // verilog/motorControl.v(63[16:31])
    defparam i47572_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_24_i357_2_lut (.I0(\Ki[7] ), .I1(n353), .I2(GND_net), 
            .I3(GND_net), .O(n530_adj_4414));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i357_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_30_i8_3_lut (.I0(n455[4]), .I1(n455[8]), .I2(n17_adj_4673), 
            .I3(GND_net), .O(n8_adj_4681));   // verilog/motorControl.v(63[16:31])
    defparam LessThan_30_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_23_i198_2_lut (.I0(\Kp[4] ), .I1(n207[4]), .I2(GND_net), 
            .I3(GND_net), .O(n293_adj_4413));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i198_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i247_2_lut (.I0(\Kp[5] ), .I1(n207[4]), .I2(GND_net), 
            .I3(GND_net), .O(n366_adj_4412));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i247_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_33_inv_0_i23_1_lut (.I0(PWMLimit[22]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n46[22]));   // verilog/motorControl.v(66[24:33])
    defparam unary_minus_33_inv_0_i23_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_23_i296_2_lut (.I0(\Kp[6] ), .I1(n207[4]), .I2(GND_net), 
            .I3(GND_net), .O(n439_adj_4409));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i296_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_33_inv_0_i24_1_lut (.I0(PWMLimit[23]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n46[23]));   // verilog/motorControl.v(66[24:33])
    defparam unary_minus_33_inv_0_i24_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 LessThan_30_i24_3_lut (.I0(n16_adj_4679), .I1(n455[22]), .I2(n45_adj_4654), 
            .I3(GND_net), .O(n24_adj_4682));   // verilog/motorControl.v(63[16:31])
    defparam LessThan_30_i24_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i45942_4_lut (.I0(n43_adj_4655), .I1(n25_adj_4659), .I2(n23_adj_4657), 
            .I3(n60710), .O(n60654));
    defparam i45942_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 mult_24_i406_2_lut (.I0(\Ki[8] ), .I1(n353), .I2(GND_net), 
            .I3(GND_net), .O(n603_adj_4406));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i406_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i345_2_lut (.I0(\Kp[7] ), .I1(n207[4]), .I2(GND_net), 
            .I3(GND_net), .O(n512_adj_4405));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i345_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i455_2_lut (.I0(\Ki[9] ), .I1(n353), .I2(GND_net), 
            .I3(GND_net), .O(n676_adj_4404));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i455_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i47172_4_lut (.I0(n24_adj_4682), .I1(n8_adj_4681), .I2(n45_adj_4654), 
            .I3(n60650), .O(n61885));   // verilog/motorControl.v(63[16:31])
    defparam i47172_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 mult_23_i394_2_lut (.I0(\Kp[8] ), .I1(n207[4]), .I2(GND_net), 
            .I3(GND_net), .O(n585_adj_4403));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i394_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i443_2_lut (.I0(\Kp[9] ), .I1(n207[4]), .I2(GND_net), 
            .I3(GND_net), .O(n658_adj_4401));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i443_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i46434_3_lut (.I0(n62285), .I1(n455[12]), .I2(n25_adj_4659), 
            .I3(GND_net), .O(n61147));   // verilog/motorControl.v(63[16:31])
    defparam i46434_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_30_i4_4_lut (.I0(n455[0]), .I1(n455[1]), .I2(PWMLimit[1]), 
            .I3(PWMLimit[0]), .O(n4_adj_4683));   // verilog/motorControl.v(63[16:31])
    defparam LessThan_30_i4_4_lut.LUT_INIT = 16'h0c8e;
    SB_LUT4 i47569_3_lut (.I0(n4_adj_4683), .I1(n455[13]), .I2(n27_adj_4671), 
            .I3(GND_net), .O(n62282));   // verilog/motorControl.v(63[16:31])
    defparam i47569_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i47570_3_lut (.I0(n62282), .I1(n455[14]), .I2(n29_adj_4661), 
            .I3(GND_net), .O(n62283));   // verilog/motorControl.v(63[16:31])
    defparam i47570_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_23_i492_2_lut (.I0(\Kp[10] ), .I1(n207[4]), .I2(GND_net), 
            .I3(GND_net), .O(n731_adj_4400));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i492_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i541_2_lut (.I0(\Kp[11] ), .I1(n207[4]), .I2(GND_net), 
            .I3(GND_net), .O(n804_adj_4399));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i541_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i504_2_lut (.I0(\Ki[10] ), .I1(n353), .I2(GND_net), 
            .I3(GND_net), .O(n749_adj_4397));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i504_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i45975_4_lut (.I0(n33_adj_4667), .I1(n31_adj_4663), .I2(n29_adj_4661), 
            .I3(n60700), .O(n60687));
    defparam i45975_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 mult_23_i590_2_lut (.I0(\Kp[12] ), .I1(n207[4]), .I2(GND_net), 
            .I3(GND_net), .O(n877_adj_4396));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i590_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i34_2_lut (.I0(\Ki[0] ), .I1(n343), .I2(GND_net), 
            .I3(GND_net), .O(n50_adj_4208));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i34_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i639_2_lut (.I0(\Kp[13] ), .I1(n207[4]), .I2(GND_net), 
            .I3(GND_net), .O(n950_adj_4395));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i639_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i553_2_lut (.I0(\Ki[11] ), .I1(n353), .I2(GND_net), 
            .I3(GND_net), .O(n822_adj_4394));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i553_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i48077_4_lut (.I0(n30_adj_4678), .I1(n10_adj_4677), .I2(n35_adj_4666), 
            .I3(n60683), .O(n62790));   // verilog/motorControl.v(63[16:31])
    defparam i48077_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 mult_23_i688_2_lut (.I0(\Kp[14] ), .I1(n207[4]), .I2(GND_net), 
            .I3(GND_net), .O(n1023_adj_4393));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i688_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i602_2_lut (.I0(\Ki[12] ), .I1(n353), .I2(GND_net), 
            .I3(GND_net), .O(n895_adj_4392));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i602_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i737_2_lut (.I0(\Kp[15] ), .I1(n207[4]), .I2(GND_net), 
            .I3(GND_net), .O(n1096_adj_4391));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i737_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i46436_3_lut (.I0(n62283), .I1(n455[15]), .I2(n31_adj_4663), 
            .I3(GND_net), .O(n61149));   // verilog/motorControl.v(63[16:31])
    defparam i46436_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_21_i11_3_lut (.I0(n233[10]), .I1(n285[10]), .I2(n284), 
            .I3(GND_net), .O(n310[10]));   // verilog/motorControl.v(58[20] 60[14])
    defparam mux_21_i11_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i48187_4_lut (.I0(n61149), .I1(n62790), .I2(n35_adj_4666), 
            .I3(n60687), .O(n62900));   // verilog/motorControl.v(63[16:31])
    defparam i48187_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i48188_3_lut (.I0(n62900), .I1(n455[18]), .I2(n37_adj_4656), 
            .I3(GND_net), .O(n62901));   // verilog/motorControl.v(63[16:31])
    defparam i48188_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_24_i651_2_lut (.I0(\Ki[13] ), .I1(n353), .I2(GND_net), 
            .I3(GND_net), .O(n968_adj_4390));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i651_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i48163_3_lut (.I0(n62901), .I1(n455[19]), .I2(n39_adj_4653), 
            .I3(GND_net), .O(n62876));   // verilog/motorControl.v(63[16:31])
    defparam i48163_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i45944_4_lut (.I0(n43_adj_4655), .I1(n41_adj_4652), .I2(n39_adj_4653), 
            .I3(n62826), .O(n60656));
    defparam i45944_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 mux_22_i11_3_lut (.I0(n310[10]), .I1(IntegralLimit[10]), .I2(n258), 
            .I3(GND_net), .O(n349));   // verilog/motorControl.v(58[20] 60[14])
    defparam mux_22_i11_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_24_i700_2_lut (.I0(\Ki[14] ), .I1(n353), .I2(GND_net), 
            .I3(GND_net), .O(n1041_adj_4389));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i700_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i659_2_lut (.I0(\Ki[13] ), .I1(n349), .I2(GND_net), 
            .I3(GND_net), .O(n980_adj_4207));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i659_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i749_2_lut (.I0(\Ki[15] ), .I1(n353), .I2(GND_net), 
            .I3(GND_net), .O(n1114_adj_4388));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i749_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i77_2_lut (.I0(\Kp[1] ), .I1(n207[17]), .I2(GND_net), 
            .I3(GND_net), .O(n113_adj_4386));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i77_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i47850_4_lut (.I0(n61147), .I1(n61885), .I2(n45_adj_4654), 
            .I3(n60654), .O(n62563));   // verilog/motorControl.v(63[16:31])
    defparam i47850_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 mult_23_i30_2_lut (.I0(\Kp[0] ), .I1(n207[18]), .I2(GND_net), 
            .I3(GND_net), .O(n44_adj_4385));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i30_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i46442_3_lut (.I0(n62876), .I1(n455[20]), .I2(n41_adj_4652), 
            .I3(GND_net), .O(n61155));   // verilog/motorControl.v(63[16:31])
    defparam i46442_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_24_i77_2_lut (.I0(\Ki[1] ), .I1(n346), .I2(GND_net), 
            .I3(GND_net), .O(n113));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i77_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i30_2_lut (.I0(\Ki[0] ), .I1(n345), .I2(GND_net), 
            .I3(GND_net), .O(n44));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i30_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i126_2_lut (.I0(\Kp[2] ), .I1(n207[17]), .I2(GND_net), 
            .I3(GND_net), .O(n186_adj_4384));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i126_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i48042_4_lut (.I0(n61155), .I1(n62563), .I2(n45_adj_4654), 
            .I3(n60656), .O(n62755));   // verilog/motorControl.v(63[16:31])
    defparam i48042_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 LessThan_9_i41_2_lut (.I0(PWMLimit[20]), .I1(setpoint[20]), 
            .I2(GND_net), .I3(GND_net), .O(n41_adj_4684));   // verilog/motorControl.v(45[16:33])
    defparam LessThan_9_i41_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_9_i39_2_lut (.I0(PWMLimit[19]), .I1(setpoint[19]), 
            .I2(GND_net), .I3(GND_net), .O(n39_adj_4685));   // verilog/motorControl.v(45[16:33])
    defparam LessThan_9_i39_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_9_i45_2_lut (.I0(PWMLimit[22]), .I1(setpoint[22]), 
            .I2(GND_net), .I3(GND_net), .O(n45_adj_4686));   // verilog/motorControl.v(45[16:33])
    defparam LessThan_9_i45_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_9_i43_2_lut (.I0(PWMLimit[21]), .I1(setpoint[21]), 
            .I2(GND_net), .I3(GND_net), .O(n43_adj_4687));   // verilog/motorControl.v(45[16:33])
    defparam LessThan_9_i43_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_9_i37_2_lut (.I0(PWMLimit[18]), .I1(setpoint[18]), 
            .I2(GND_net), .I3(GND_net), .O(n37_adj_4688));   // verilog/motorControl.v(45[16:33])
    defparam LessThan_9_i37_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_24_i126_2_lut (.I0(\Ki[2] ), .I1(n346), .I2(GND_net), 
            .I3(GND_net), .O(n186));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i126_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_9_i29_2_lut (.I0(PWMLimit[14]), .I1(setpoint[14]), 
            .I2(GND_net), .I3(GND_net), .O(n29_adj_4689));   // verilog/motorControl.v(45[16:33])
    defparam LessThan_9_i29_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_24_i130_2_lut (.I0(\Ki[2] ), .I1(n344), .I2(GND_net), 
            .I3(GND_net), .O(n192_adj_4206));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i130_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_9_i31_2_lut (.I0(PWMLimit[15]), .I1(setpoint[15]), 
            .I2(GND_net), .I3(GND_net), .O(n31_adj_4690));   // verilog/motorControl.v(45[16:33])
    defparam LessThan_9_i31_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_24_i175_2_lut (.I0(\Ki[3] ), .I1(n346), .I2(GND_net), 
            .I3(GND_net), .O(n259_adj_4383));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i175_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i175_2_lut (.I0(\Kp[3] ), .I1(n207[17]), .I2(GND_net), 
            .I3(GND_net), .O(n259));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i175_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_9_i23_2_lut (.I0(PWMLimit[11]), .I1(setpoint[11]), 
            .I2(GND_net), .I3(GND_net), .O(n23_adj_4691));   // verilog/motorControl.v(45[16:33])
    defparam LessThan_9_i23_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_9_i25_2_lut (.I0(PWMLimit[12]), .I1(setpoint[12]), 
            .I2(GND_net), .I3(GND_net), .O(n25_adj_4692));   // verilog/motorControl.v(45[16:33])
    defparam LessThan_9_i25_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_24_i224_2_lut (.I0(\Ki[4] ), .I1(n346), .I2(GND_net), 
            .I3(GND_net), .O(n332_adj_4382));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i224_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i224_2_lut (.I0(\Kp[4] ), .I1(n207[17]), .I2(GND_net), 
            .I3(GND_net), .O(n332));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i224_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i273_2_lut (.I0(\Ki[5] ), .I1(n346), .I2(GND_net), 
            .I3(GND_net), .O(n405_adj_4381));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i273_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i273_2_lut (.I0(\Kp[5] ), .I1(n207[17]), .I2(GND_net), 
            .I3(GND_net), .O(n405));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i273_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i322_2_lut (.I0(\Ki[6] ), .I1(n346), .I2(GND_net), 
            .I3(GND_net), .O(n478_adj_4380));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i322_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i371_2_lut (.I0(\Ki[7] ), .I1(n346), .I2(GND_net), 
            .I3(GND_net), .O(n551_adj_4379));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i371_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_9_i35_2_lut (.I0(PWMLimit[17]), .I1(setpoint[17]), 
            .I2(GND_net), .I3(GND_net), .O(n35_adj_4693));   // verilog/motorControl.v(45[16:33])
    defparam LessThan_9_i35_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_9_i33_2_lut (.I0(PWMLimit[16]), .I1(setpoint[16]), 
            .I2(GND_net), .I3(GND_net), .O(n33_adj_4694));   // verilog/motorControl.v(45[16:33])
    defparam LessThan_9_i33_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_9_i11_2_lut (.I0(PWMLimit[5]), .I1(setpoint[5]), .I2(GND_net), 
            .I3(GND_net), .O(n11_adj_4695));   // verilog/motorControl.v(45[16:33])
    defparam LessThan_9_i11_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_9_i13_2_lut (.I0(PWMLimit[6]), .I1(setpoint[6]), .I2(GND_net), 
            .I3(GND_net), .O(n13_adj_4696));   // verilog/motorControl.v(45[16:33])
    defparam LessThan_9_i13_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_24_i420_2_lut (.I0(\Ki[8] ), .I1(n346), .I2(GND_net), 
            .I3(GND_net), .O(n624_adj_4378));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i420_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i322_2_lut (.I0(\Kp[6] ), .I1(n207[17]), .I2(GND_net), 
            .I3(GND_net), .O(n478));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i322_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i469_2_lut (.I0(\Ki[9] ), .I1(n346), .I2(GND_net), 
            .I3(GND_net), .O(n697_adj_4377));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i469_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i518_2_lut (.I0(\Ki[10] ), .I1(n346), .I2(GND_net), 
            .I3(GND_net), .O(n770_adj_4376));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i518_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i371_2_lut (.I0(\Kp[7] ), .I1(n207[17]), .I2(GND_net), 
            .I3(GND_net), .O(n551_adj_4375));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i371_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i420_2_lut (.I0(\Kp[8] ), .I1(n207[17]), .I2(GND_net), 
            .I3(GND_net), .O(n624));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i420_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_9_i27_2_lut (.I0(PWMLimit[13]), .I1(setpoint[13]), 
            .I2(GND_net), .I3(GND_net), .O(n27_adj_4697));   // verilog/motorControl.v(45[16:33])
    defparam LessThan_9_i27_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_9_i9_2_lut (.I0(PWMLimit[4]), .I1(setpoint[4]), .I2(GND_net), 
            .I3(GND_net), .O(n9_adj_4698));   // verilog/motorControl.v(45[16:33])
    defparam LessThan_9_i9_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i22198_1_lut (.I0(duty[0]), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n35713));   // verilog/motorControl.v(42[14] 73[8])
    defparam i22198_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 LessThan_9_i17_2_lut (.I0(PWMLimit[8]), .I1(setpoint[8]), .I2(GND_net), 
            .I3(GND_net), .O(n17_adj_4699));   // verilog/motorControl.v(45[16:33])
    defparam LessThan_9_i17_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_23_i469_2_lut (.I0(\Kp[9] ), .I1(n207[17]), .I2(GND_net), 
            .I3(GND_net), .O(n697));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i469_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i81_2_lut (.I0(\Kp[1] ), .I1(n207[19]), .I2(GND_net), 
            .I3(GND_net), .O(n119));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i81_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i518_2_lut (.I0(\Kp[10] ), .I1(n207[17]), .I2(GND_net), 
            .I3(GND_net), .O(n770));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i518_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i61_2_lut (.I0(\Ki[1] ), .I1(n354), .I2(GND_net), 
            .I3(GND_net), .O(n89_adj_4373));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i61_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i14_2_lut (.I0(\Ki[0] ), .I1(n353), .I2(GND_net), 
            .I3(GND_net), .O(n20_adj_4372));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i14_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_9_i21_2_lut (.I0(PWMLimit[10]), .I1(setpoint[10]), 
            .I2(GND_net), .I3(GND_net), .O(n21_adj_4700));   // verilog/motorControl.v(45[16:33])
    defparam LessThan_9_i21_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_24_i110_2_lut (.I0(\Ki[2] ), .I1(n354), .I2(GND_net), 
            .I3(GND_net), .O(n162_adj_4371));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i110_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i159_2_lut (.I0(\Ki[3] ), .I1(n354), .I2(GND_net), 
            .I3(GND_net), .O(n235_adj_4370));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i159_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i208_2_lut (.I0(\Ki[4] ), .I1(n354), .I2(GND_net), 
            .I3(GND_net), .O(n308_adj_4369));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i208_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i257_2_lut (.I0(\Ki[5] ), .I1(n354), .I2(GND_net), 
            .I3(GND_net), .O(n381_adj_4368));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i257_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i306_2_lut (.I0(\Ki[6] ), .I1(n354), .I2(GND_net), 
            .I3(GND_net), .O(n454_adj_4367));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i306_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i355_2_lut (.I0(\Ki[7] ), .I1(n354), .I2(GND_net), 
            .I3(GND_net), .O(n527_adj_4366));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i355_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i404_2_lut (.I0(\Ki[8] ), .I1(n354), .I2(GND_net), 
            .I3(GND_net), .O(n600_adj_4365));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i404_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i453_2_lut (.I0(\Ki[9] ), .I1(n354), .I2(GND_net), 
            .I3(GND_net), .O(n673_adj_4364));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i453_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i34_2_lut (.I0(\Kp[0] ), .I1(n207[20]), .I2(GND_net), 
            .I3(GND_net), .O(n50));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i34_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i502_2_lut (.I0(\Ki[10] ), .I1(n354), .I2(GND_net), 
            .I3(GND_net), .O(n746_adj_4363));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i502_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i551_2_lut (.I0(\Ki[11] ), .I1(n354), .I2(GND_net), 
            .I3(GND_net), .O(n819_adj_4362));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i551_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i600_2_lut (.I0(\Ki[12] ), .I1(n354), .I2(GND_net), 
            .I3(GND_net), .O(n892_adj_4361));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i600_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i649_2_lut (.I0(\Ki[13] ), .I1(n354), .I2(GND_net), 
            .I3(GND_net), .O(n965_adj_4360));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i649_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i698_2_lut (.I0(\Ki[14] ), .I1(n354), .I2(GND_net), 
            .I3(GND_net), .O(n1038_adj_4359));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i698_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i747_2_lut (.I0(\Ki[15] ), .I1(n354), .I2(GND_net), 
            .I3(GND_net), .O(n1111_adj_4358));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i747_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i5_4_lut (.I0(\control_mode[0] ), .I1(\control_mode[5] ), .I2(\control_mode[4] ), 
            .I3(n1_adj_2), .O(n12_adj_4702));
    defparam i5_4_lut.LUT_INIT = 16'h0002;
    SB_LUT4 mult_24_i59_2_lut (.I0(\Ki[1] ), .I1(n355), .I2(GND_net), 
            .I3(GND_net), .O(n86));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i59_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i12_2_lut (.I0(\Ki[0] ), .I1(n354), .I2(GND_net), 
            .I3(GND_net), .O(n17_adj_4357));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i12_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i6_4_lut (.I0(\control_mode[6] ), .I1(n12_adj_4702), .I2(\control_mode[7] ), 
            .I3(\control_mode[1] ), .O(n52622));
    defparam i6_4_lut.LUT_INIT = 16'h0400;
    SB_LUT4 i45940_4_lut (.I0(n21_adj_4700), .I1(n19), .I2(n17_adj_4699), 
            .I3(n9_adj_4698), .O(n60652));
    defparam i45940_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 mult_24_i108_2_lut (.I0(\Ki[2] ), .I1(n355), .I2(GND_net), 
            .I3(GND_net), .O(n159));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i108_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i45918_4_lut (.I0(n27_adj_4697), .I1(n15), .I2(n13_adj_4696), 
            .I3(n11_adj_4695), .O(n60630));
    defparam i45918_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 mult_24_i157_2_lut (.I0(\Ki[3] ), .I1(n355), .I2(GND_net), 
            .I3(GND_net), .O(n232));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i157_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i206_2_lut (.I0(\Ki[4] ), .I1(n355), .I2(GND_net), 
            .I3(GND_net), .O(n305_adj_4356));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i206_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i255_2_lut (.I0(\Ki[5] ), .I1(n355), .I2(GND_net), 
            .I3(GND_net), .O(n378));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i255_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i304_2_lut (.I0(\Ki[6] ), .I1(n355), .I2(GND_net), 
            .I3(GND_net), .O(n451_adj_4355));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i304_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i353_2_lut (.I0(\Ki[7] ), .I1(n355), .I2(GND_net), 
            .I3(GND_net), .O(n524));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i353_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_9_i30_3_lut (.I0(n12_adj_4705), .I1(setpoint[17]), 
            .I2(n35_adj_4693), .I3(GND_net), .O(n30_adj_4706));   // verilog/motorControl.v(45[16:33])
    defparam LessThan_9_i30_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_24_i402_2_lut (.I0(\Ki[8] ), .I1(n355), .I2(GND_net), 
            .I3(GND_net), .O(n597));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i402_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i451_2_lut (.I0(\Ki[9] ), .I1(n355), .I2(GND_net), 
            .I3(GND_net), .O(n670));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i451_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i500_2_lut (.I0(\Ki[10] ), .I1(n355), .I2(GND_net), 
            .I3(GND_net), .O(n743));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i500_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i549_2_lut (.I0(\Ki[11] ), .I1(n355), .I2(GND_net), 
            .I3(GND_net), .O(n816));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i549_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i598_2_lut (.I0(\Ki[12] ), .I1(n355), .I2(GND_net), 
            .I3(GND_net), .O(n889));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i598_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i647_2_lut (.I0(\Ki[13] ), .I1(n355), .I2(GND_net), 
            .I3(GND_net), .O(n962));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i647_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i696_2_lut (.I0(\Ki[14] ), .I1(n355), .I2(GND_net), 
            .I3(GND_net), .O(n1035));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i696_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i46900_4_lut (.I0(n13_adj_4696), .I1(n11_adj_4695), .I2(n9_adj_4698), 
            .I3(n60673), .O(n61613));
    defparam i46900_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 mult_24_i745_2_lut (.I0(\Ki[15] ), .I1(n355), .I2(GND_net), 
            .I3(GND_net), .O(n1108));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i745_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i46892_4_lut (.I0(n19), .I1(n17_adj_4699), .I2(n15), .I3(n61613), 
            .O(n61605));
    defparam i46892_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i47982_4_lut (.I0(n25_adj_4692), .I1(n23_adj_4691), .I2(n21_adj_4700), 
            .I3(n61605), .O(n62695));
    defparam i47982_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i47347_4_lut (.I0(n31_adj_4690), .I1(n29_adj_4689), .I2(n27_adj_4697), 
            .I3(n62695), .O(n62060));
    defparam i47347_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 mult_23_i75_2_lut (.I0(\Kp[1] ), .I1(n207[16]), .I2(GND_net), 
            .I3(GND_net), .O(n110_adj_4353));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i75_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i48107_4_lut (.I0(n37_adj_4688), .I1(n35_adj_4693), .I2(n33_adj_4694), 
            .I3(n62060), .O(n62820));
    defparam i48107_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 mult_23_i28_2_lut (.I0(\Kp[0] ), .I1(n207[17]), .I2(GND_net), 
            .I3(GND_net), .O(n41_adj_4352));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i28_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i124_2_lut (.I0(\Kp[2] ), .I1(n207[16]), .I2(GND_net), 
            .I3(GND_net), .O(n183_adj_4351));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i124_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i173_2_lut (.I0(\Kp[3] ), .I1(n207[16]), .I2(GND_net), 
            .I3(GND_net), .O(n256_adj_4349));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i173_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i222_2_lut (.I0(\Kp[4] ), .I1(n207[16]), .I2(GND_net), 
            .I3(GND_net), .O(n329_adj_4348));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i222_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i130_2_lut (.I0(\Kp[2] ), .I1(n207[19]), .I2(GND_net), 
            .I3(GND_net), .O(n192));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i130_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i271_2_lut (.I0(\Kp[5] ), .I1(n207[16]), .I2(GND_net), 
            .I3(GND_net), .O(n402_adj_4347));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i271_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i179_2_lut (.I0(\Ki[3] ), .I1(n344), .I2(GND_net), 
            .I3(GND_net), .O(n265_adj_4205));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i179_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i47657_3_lut (.I0(n6_adj_4707), .I1(setpoint[10]), .I2(n21_adj_4700), 
            .I3(GND_net), .O(n62370));   // verilog/motorControl.v(45[16:33])
    defparam i47657_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_23_i320_2_lut (.I0(\Kp[6] ), .I1(n207[16]), .I2(GND_net), 
            .I3(GND_net), .O(n475_adj_4346));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i320_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i47658_3_lut (.I0(n62370), .I1(setpoint[11]), .I2(n23_adj_4691), 
            .I3(GND_net), .O(n62371));   // verilog/motorControl.v(45[16:33])
    defparam i47658_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_23_i369_2_lut (.I0(\Kp[7] ), .I1(n207[16]), .I2(GND_net), 
            .I3(GND_net), .O(n548_adj_4345));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i369_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_9_i24_3_lut (.I0(n16_adj_4708), .I1(setpoint[22]), 
            .I2(n45_adj_4686), .I3(GND_net), .O(n24_adj_4709));   // verilog/motorControl.v(45[16:33])
    defparam LessThan_9_i24_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i45857_4_lut (.I0(n43_adj_4687), .I1(n25_adj_4692), .I2(n23_adj_4691), 
            .I3(n60652), .O(n60569));
    defparam i45857_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 mult_23_i418_2_lut (.I0(\Kp[8] ), .I1(n207[16]), .I2(GND_net), 
            .I3(GND_net), .O(n621_adj_4344));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i418_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i47160_4_lut (.I0(n24_adj_4709), .I1(n8_adj_4710), .I2(n45_adj_4686), 
            .I3(n60561), .O(n61873));   // verilog/motorControl.v(45[16:33])
    defparam i47160_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i46386_3_lut (.I0(n62371), .I1(setpoint[12]), .I2(n25_adj_4692), 
            .I3(GND_net), .O(n61099));   // verilog/motorControl.v(45[16:33])
    defparam i46386_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_9_i4_4_lut (.I0(PWMLimit[0]), .I1(setpoint[1]), .I2(PWMLimit[1]), 
            .I3(setpoint[0]), .O(n4_adj_4711));   // verilog/motorControl.v(45[16:33])
    defparam LessThan_9_i4_4_lut.LUT_INIT = 16'h4d0c;
    SB_LUT4 i47655_3_lut (.I0(n4_adj_4711), .I1(setpoint[13]), .I2(n27_adj_4697), 
            .I3(GND_net), .O(n62368));   // verilog/motorControl.v(45[16:33])
    defparam i47655_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i47656_3_lut (.I0(n62368), .I1(setpoint[14]), .I2(n29_adj_4689), 
            .I3(GND_net), .O(n62369));   // verilog/motorControl.v(45[16:33])
    defparam i47656_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i45899_4_lut (.I0(n33_adj_4694), .I1(n31_adj_4690), .I2(n29_adj_4689), 
            .I3(n60630), .O(n60611));
    defparam i45899_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 mult_23_i467_2_lut (.I0(\Kp[9] ), .I1(n207[16]), .I2(GND_net), 
            .I3(GND_net), .O(n694_adj_4343));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i467_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 n9440_bdd_4_lut_48892 (.I0(n9440), .I1(n59911), .I2(setpoint[23]), 
            .I3(n4357), .O(n63551));
    defparam n9440_bdd_4_lut_48892.LUT_INIT = 16'he4aa;
    SB_LUT4 i48032_4_lut (.I0(n30_adj_4706), .I1(n10_adj_4712), .I2(n35_adj_4693), 
            .I3(n60601), .O(n62745));   // verilog/motorControl.v(45[16:33])
    defparam i48032_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i46388_3_lut (.I0(n62369), .I1(setpoint[15]), .I2(n31_adj_4690), 
            .I3(GND_net), .O(n61101));   // verilog/motorControl.v(45[16:33])
    defparam i46388_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_23_i516_2_lut (.I0(\Kp[10] ), .I1(n207[16]), .I2(GND_net), 
            .I3(GND_net), .O(n767_adj_4342));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i516_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i565_2_lut (.I0(\Kp[11] ), .I1(n207[16]), .I2(GND_net), 
            .I3(GND_net), .O(n840_adj_4341));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i565_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i48248_4_lut (.I0(n61101), .I1(n62745), .I2(n35_adj_4693), 
            .I3(n60611), .O(n62961));   // verilog/motorControl.v(45[16:33])
    defparam i48248_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i48249_3_lut (.I0(n62961), .I1(setpoint[18]), .I2(n37_adj_4688), 
            .I3(GND_net), .O(n62962));   // verilog/motorControl.v(45[16:33])
    defparam i48249_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_24_i57_2_lut (.I0(\Ki[1] ), .I1(n356), .I2(GND_net), 
            .I3(GND_net), .O(n83));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i57_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i48200_3_lut (.I0(n62962), .I1(setpoint[19]), .I2(n39_adj_4685), 
            .I3(GND_net), .O(n62913));   // verilog/motorControl.v(45[16:33])
    defparam i48200_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_24_i10_2_lut (.I0(\Ki[0] ), .I1(n355), .I2(GND_net), 
            .I3(GND_net), .O(n14_adj_4340));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i10_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i45865_4_lut (.I0(n43_adj_4687), .I1(n41_adj_4684), .I2(n39_adj_4685), 
            .I3(n62820), .O(n60577));
    defparam i45865_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i47834_4_lut (.I0(n61099), .I1(n61873), .I2(n45_adj_4686), 
            .I3(n60569), .O(n62547));   // verilog/motorControl.v(45[16:33])
    defparam i47834_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i46394_3_lut (.I0(n62913), .I1(setpoint[20]), .I2(n41_adj_4684), 
            .I3(GND_net), .O(n61107));   // verilog/motorControl.v(45[16:33])
    defparam i46394_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i48036_4_lut (.I0(n61107), .I1(n62547), .I2(n45_adj_4686), 
            .I3(n60577), .O(n62749));   // verilog/motorControl.v(45[16:33])
    defparam i48036_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 mult_24_i106_2_lut (.I0(\Ki[2] ), .I1(n356), .I2(GND_net), 
            .I3(GND_net), .O(n156));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i106_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i48037_3_lut (.I0(n62749), .I1(PWMLimit[23]), .I2(setpoint[23]), 
            .I3(GND_net), .O(n105));   // verilog/motorControl.v(45[16:33])
    defparam i48037_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 mult_24_i155_2_lut (.I0(\Ki[3] ), .I1(n356), .I2(GND_net), 
            .I3(GND_net), .O(n229));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i155_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_32_i33_2_lut (.I0(n455[16]), .I1(n535[16]), .I2(GND_net), 
            .I3(GND_net), .O(n33_adj_4713));   // verilog/motorControl.v(65[25:41])
    defparam LessThan_32_i33_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_23_i179_2_lut (.I0(\Kp[3] ), .I1(n207[19]), .I2(GND_net), 
            .I3(GND_net), .O(n265));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i179_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i50_3_lut (.I0(n45), .I1(n455[1]), .I2(n34[1]), .I3(GND_net), 
            .O(n43_adj_4714));
    defparam i50_3_lut.LUT_INIT = 16'hb2b2;
    SB_LUT4 LessThan_26_i37_2_lut (.I0(\deadband[18] ), .I1(n455[18]), .I2(GND_net), 
            .I3(GND_net), .O(n37_adj_4715));   // verilog/motorControl.v(62[14:31])
    defparam LessThan_26_i37_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_24_i228_2_lut (.I0(\Ki[4] ), .I1(n344), .I2(GND_net), 
            .I3(GND_net), .O(n338_adj_4204));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i228_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_26_i33_2_lut (.I0(\deadband[16] ), .I1(n455[16]), .I2(GND_net), 
            .I3(GND_net), .O(n33_adj_4716));   // verilog/motorControl.v(62[14:31])
    defparam LessThan_26_i33_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_26_i31_2_lut (.I0(\deadband[15] ), .I1(n455[15]), .I2(GND_net), 
            .I3(GND_net), .O(n31_adj_4717));   // verilog/motorControl.v(62[14:31])
    defparam LessThan_26_i31_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_26_i4_4_lut (.I0(n28[0]), .I1(n455[1]), .I2(\deadband[1] ), 
            .I3(n455[0]), .O(n4_adj_4718));   // verilog/motorControl.v(62[14:31])
    defparam LessThan_26_i4_4_lut.LUT_INIT = 16'h8e0c;
    SB_LUT4 LessThan_26_i35_2_lut (.I0(\deadband[17] ), .I1(n455[17]), .I2(GND_net), 
            .I3(GND_net), .O(n35_adj_4719));   // verilog/motorControl.v(62[14:31])
    defparam LessThan_26_i35_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_26_i21_2_lut (.I0(\deadband[10] ), .I1(n455[10]), .I2(GND_net), 
            .I3(GND_net), .O(n21_adj_4720));   // verilog/motorControl.v(62[14:31])
    defparam LessThan_26_i21_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_24_i277_2_lut (.I0(\Ki[5] ), .I1(n344), .I2(GND_net), 
            .I3(GND_net), .O(n411_adj_4203));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i277_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_26_i23_2_lut (.I0(\deadband[11] ), .I1(n455[11]), .I2(GND_net), 
            .I3(GND_net), .O(n23_adj_4721));   // verilog/motorControl.v(62[14:31])
    defparam LessThan_26_i23_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_26_i25_2_lut (.I0(\deadband[12] ), .I1(n455[12]), .I2(GND_net), 
            .I3(GND_net), .O(n25_adj_4722));   // verilog/motorControl.v(62[14:31])
    defparam LessThan_26_i25_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_26_i27_2_lut (.I0(\deadband[13] ), .I1(n455[13]), .I2(GND_net), 
            .I3(GND_net), .O(n27_adj_4723));   // verilog/motorControl.v(62[14:31])
    defparam LessThan_26_i27_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_26_i29_2_lut (.I0(\deadband[14] ), .I1(n455[14]), .I2(GND_net), 
            .I3(GND_net), .O(n29_adj_4724));   // verilog/motorControl.v(62[14:31])
    defparam LessThan_26_i29_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_26_i13_2_lut (.I0(\deadband[6] ), .I1(n455[6]), .I2(GND_net), 
            .I3(GND_net), .O(n13_adj_4725));   // verilog/motorControl.v(62[14:31])
    defparam LessThan_26_i13_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_26_i15_2_lut (.I0(\deadband[7] ), .I1(n455[7]), .I2(GND_net), 
            .I3(GND_net), .O(n15_adj_4726));   // verilog/motorControl.v(62[14:31])
    defparam LessThan_26_i15_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_26_i17_2_lut (.I0(\deadband[8] ), .I1(n455[8]), .I2(GND_net), 
            .I3(GND_net), .O(n17_adj_4727));   // verilog/motorControl.v(62[14:31])
    defparam LessThan_26_i17_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 unary_minus_27_inv_0_i4_1_lut (.I0(\deadband[3] ), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n28[3]));   // verilog/motorControl.v(62[45:54])
    defparam unary_minus_27_inv_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 LessThan_26_i9_2_lut (.I0(\deadband[4] ), .I1(n455[4]), .I2(GND_net), 
            .I3(GND_net), .O(n9_adj_4728));   // verilog/motorControl.v(62[14:31])
    defparam LessThan_26_i9_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_26_i11_2_lut (.I0(\deadband[5] ), .I1(n455[5]), .I2(GND_net), 
            .I3(GND_net), .O(n11_adj_4729));   // verilog/motorControl.v(62[14:31])
    defparam LessThan_26_i11_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_26_i19_2_lut (.I0(\deadband[9] ), .I1(n455[9]), .I2(GND_net), 
            .I3(GND_net), .O(n19_adj_4730));   // verilog/motorControl.v(62[14:31])
    defparam LessThan_26_i19_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i46101_4_lut (.I0(n455[9]), .I1(n455[5]), .I2(n34[9]), .I3(n34[5]), 
            .O(n60813));
    defparam i46101_4_lut.LUT_INIT = 16'h7bde;
    SB_LUT4 i47016_3_lut (.I0(n455[10]), .I1(n60813), .I2(n34[10]), .I3(GND_net), 
            .O(n61729));
    defparam i47016_3_lut.LUT_INIT = 16'hdede;
    SB_LUT4 LessThan_28_i23_rep_131_2_lut (.I0(n455[11]), .I1(n34[11]), 
            .I2(GND_net), .I3(GND_net), .O(n63839));   // verilog/motorControl.v(62[35:55])
    defparam LessThan_28_i23_rep_131_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i46109_4_lut (.I0(n455[7]), .I1(n455[6]), .I2(n34[7]), .I3(n34[6]), 
            .O(n60821));
    defparam i46109_4_lut.LUT_INIT = 16'h7bde;
    SB_LUT4 i47026_3_lut (.I0(n455[8]), .I1(n60821), .I2(n34[8]), .I3(GND_net), 
            .O(n61739));
    defparam i47026_3_lut.LUT_INIT = 16'hdede;
    SB_LUT4 LessThan_28_i29_rep_145_2_lut (.I0(n455[14]), .I1(n34[14]), 
            .I2(GND_net), .I3(GND_net), .O(n63853));   // verilog/motorControl.v(62[35:55])
    defparam LessThan_28_i29_rep_145_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i47000_4_lut (.I0(n455[15]), .I1(n63853), .I2(n34[15]), .I3(n61739), 
            .O(n61713));
    defparam i47000_4_lut.LUT_INIT = 16'hdeff;
    SB_LUT4 LessThan_28_i33_rep_110_2_lut (.I0(n455[16]), .I1(n34[16]), 
            .I2(GND_net), .I3(GND_net), .O(n63818));   // verilog/motorControl.v(62[35:55])
    defparam LessThan_28_i33_rep_110_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_28_i14_3_lut (.I0(n34[8]), .I1(n34[17]), .I2(n455[17]), 
            .I3(GND_net), .O(n14_adj_4731));   // verilog/motorControl.v(62[35:55])
    defparam LessThan_28_i14_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i46051_4_lut (.I0(n455[17]), .I1(n455[8]), .I2(n34[17]), .I3(n34[8]), 
            .O(n60763));
    defparam i46051_4_lut.LUT_INIT = 16'h7bde;
    SB_LUT4 LessThan_28_i12_3_lut (.I0(n34[6]), .I1(n34[7]), .I2(n455[7]), 
            .I3(GND_net), .O(n12_adj_4732));   // verilog/motorControl.v(62[35:55])
    defparam LessThan_28_i12_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 LessThan_28_i32_3_lut (.I0(n14_adj_4731), .I1(n34[18]), .I2(n455[18]), 
            .I3(GND_net), .O(n32_adj_4733));   // verilog/motorControl.v(62[35:55])
    defparam LessThan_28_i32_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i46118_4_lut (.I0(n455[4]), .I1(n455[3]), .I2(n34[4]), .I3(n34[3]), 
            .O(n60830));
    defparam i46118_4_lut.LUT_INIT = 16'h7bde;
    SB_LUT4 n63551_bdd_4_lut (.I0(n63551), .I1(n535[23]), .I2(n455[23]), 
            .I3(n4357), .O(n63554));
    defparam n63551_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i47032_3_lut (.I0(n455[5]), .I1(n60830), .I2(n34[5]), .I3(GND_net), 
            .O(n61745));
    defparam i47032_3_lut.LUT_INIT = 16'hdede;
    SB_LUT4 LessThan_28_i13_rep_152_2_lut (.I0(n455[6]), .I1(n34[6]), .I2(GND_net), 
            .I3(GND_net), .O(n63860));   // verilog/motorControl.v(62[35:55])
    defparam LessThan_28_i13_rep_152_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i47030_4_lut (.I0(n455[7]), .I1(n63860), .I2(n34[7]), .I3(n61745), 
            .O(n61743));
    defparam i47030_4_lut.LUT_INIT = 16'hdeff;
    SB_LUT4 LessThan_28_i17_rep_141_2_lut (.I0(n455[8]), .I1(n34[8]), .I2(GND_net), 
            .I3(GND_net), .O(n63849));   // verilog/motorControl.v(62[35:55])
    defparam LessThan_28_i17_rep_141_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i46103_4_lut (.I0(n455[9]), .I1(n63849), .I2(n34[9]), .I3(n61743), 
            .O(n60815));
    defparam i46103_4_lut.LUT_INIT = 16'h5a7b;
    SB_LUT4 LessThan_28_i21_rep_121_2_lut (.I0(n455[10]), .I1(n34[10]), 
            .I2(GND_net), .I3(GND_net), .O(n63829));   // verilog/motorControl.v(62[35:55])
    defparam LessThan_28_i21_rep_121_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i47423_4_lut (.I0(n455[11]), .I1(n63829), .I2(n34[11]), .I3(n60815), 
            .O(n62136));
    defparam i47423_4_lut.LUT_INIT = 16'hffde;
    SB_LUT4 LessThan_28_i25_rep_130_2_lut (.I0(n455[12]), .I1(n34[12]), 
            .I2(GND_net), .I3(GND_net), .O(n63838));   // verilog/motorControl.v(62[35:55])
    defparam LessThan_28_i25_rep_130_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_24_i204_2_lut (.I0(\Ki[4] ), .I1(n356), .I2(GND_net), 
            .I3(GND_net), .O(n302_adj_4339));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i204_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i48014_4_lut (.I0(n455[13]), .I1(n63838), .I2(n34[13]), .I3(n62136), 
            .O(n62727));
    defparam i48014_4_lut.LUT_INIT = 16'hffde;
    SB_LUT4 i47006_4_lut (.I0(n455[15]), .I1(n63853), .I2(n34[15]), .I3(n62727), 
            .O(n61719));
    defparam i47006_4_lut.LUT_INIT = 16'hdeff;
    SB_LUT4 LessThan_26_i10_3_lut (.I0(n455[5]), .I1(n455[9]), .I2(n19_adj_4730), 
            .I3(GND_net), .O(n10_adj_4734));   // verilog/motorControl.v(62[14:31])
    defparam LessThan_26_i10_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i46255_4_lut (.I0(n11_adj_4729), .I1(n9_adj_4728), .I2(\deadband[3] ), 
            .I3(n455[3]), .O(n60967));
    defparam i46255_4_lut.LUT_INIT = 16'heffe;
    SB_LUT4 i47092_4_lut (.I0(n17_adj_4727), .I1(n15_adj_4726), .I2(n13_adj_4725), 
            .I3(n60967), .O(n61805));
    defparam i47092_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i47088_4_lut (.I0(n23_adj_4721), .I1(n21_adj_4720), .I2(n19_adj_4730), 
            .I3(n61805), .O(n61801));
    defparam i47088_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i45226_4_lut (.I0(n29_adj_4724), .I1(n27_adj_4723), .I2(n25_adj_4722), 
            .I3(n61801), .O(n59938));
    defparam i45226_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 LessThan_26_i14_3_lut (.I0(n455[8]), .I1(n455[17]), .I2(n35_adj_4719), 
            .I3(GND_net), .O(n14_adj_4735));   // verilog/motorControl.v(62[14:31])
    defparam LessThan_26_i14_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i18456_3_lut (.I0(n4_adj_4718), .I1(n455[2]), .I2(n32007), 
            .I3(GND_net), .O(n6_adj_4736));
    defparam i18456_3_lut.LUT_INIT = 16'he8e8;
    SB_LUT4 i47623_3_lut (.I0(n6_adj_4736), .I1(n455[14]), .I2(n29_adj_4724), 
            .I3(GND_net), .O(n62336));   // verilog/motorControl.v(62[14:31])
    defparam i47623_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i47624_3_lut (.I0(n62336), .I1(n455[15]), .I2(n31_adj_4717), 
            .I3(GND_net), .O(n62337));   // verilog/motorControl.v(62[14:31])
    defparam i47624_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i45220_4_lut (.I0(n29_adj_4724), .I1(n17_adj_4727), .I2(n15_adj_4726), 
            .I3(n13_adj_4725), .O(n59932));
    defparam i45220_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 LessThan_26_i12_3_lut (.I0(n455[6]), .I1(n455[7]), .I2(n15_adj_4726), 
            .I3(GND_net), .O(n12_adj_4737));   // verilog/motorControl.v(62[14:31])
    defparam LessThan_26_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_26_i32_3_lut (.I0(n14_adj_4735), .I1(n455[18]), .I2(n37_adj_4715), 
            .I3(GND_net), .O(n32_adj_4738));   // verilog/motorControl.v(62[14:31])
    defparam LessThan_26_i32_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i46186_4_lut (.I0(n35_adj_4719), .I1(n33_adj_4716), .I2(n31_adj_4717), 
            .I3(n59932), .O(n60898));
    defparam i46186_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i48068_4_lut (.I0(n32_adj_4738), .I1(n12_adj_4737), .I2(n37_adj_4715), 
            .I3(n60894), .O(n62781));   // verilog/motorControl.v(62[14:31])
    defparam i48068_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i46416_3_lut (.I0(n62337), .I1(n455[16]), .I2(n33_adj_4716), 
            .I3(GND_net), .O(n61129));   // verilog/motorControl.v(62[14:31])
    defparam i46416_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_28_i8_3_lut (.I0(n34[3]), .I1(n34[4]), .I2(n455[4]), 
            .I3(GND_net), .O(n8_adj_4739));   // verilog/motorControl.v(62[35:55])
    defparam LessThan_28_i8_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i47583_3_lut (.I0(n8_adj_4739), .I1(n34[11]), .I2(n455[11]), 
            .I3(GND_net), .O(n62296));   // verilog/motorControl.v(62[35:55])
    defparam i47583_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i47584_3_lut (.I0(n62296), .I1(n34[12]), .I2(n455[12]), .I3(GND_net), 
            .O(n62297));   // verilog/motorControl.v(62[35:55])
    defparam i47584_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 LessThan_28_i10_3_lut (.I0(n34[5]), .I1(n34[9]), .I2(n455[9]), 
            .I3(GND_net), .O(n10_adj_4740));   // verilog/motorControl.v(62[35:55])
    defparam LessThan_28_i10_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i47014_4_lut (.I0(n455[12]), .I1(n63839), .I2(n34[12]), .I3(n61729), 
            .O(n61727));
    defparam i47014_4_lut.LUT_INIT = 16'hdeff;
    SB_LUT4 LessThan_28_i27_rep_126_2_lut (.I0(n455[13]), .I1(n34[13]), 
            .I2(GND_net), .I3(GND_net), .O(n63834));   // verilog/motorControl.v(62[35:55])
    defparam LessThan_28_i27_rep_126_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i47170_3_lut (.I0(n10_adj_4740), .I1(n34[10]), .I2(n455[10]), 
            .I3(GND_net), .O(n61883));   // verilog/motorControl.v(62[35:55])
    defparam i47170_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i46424_3_lut (.I0(n62297), .I1(n34[13]), .I2(n455[13]), .I3(GND_net), 
            .O(n61137));   // verilog/motorControl.v(62[35:55])
    defparam i46424_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i18444_3_lut (.I0(n34[2]), .I1(n455[2]), .I2(n43_adj_4714), 
            .I3(GND_net), .O(n6_adj_4741));
    defparam i18444_3_lut.LUT_INIT = 16'hb2b2;
    SB_LUT4 i47577_3_lut (.I0(n6_adj_4741), .I1(n34[14]), .I2(n455[14]), 
            .I3(GND_net), .O(n62290));   // verilog/motorControl.v(62[35:55])
    defparam i47577_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i47578_3_lut (.I0(n62290), .I1(n34[15]), .I2(n455[15]), .I3(GND_net), 
            .O(n62291));   // verilog/motorControl.v(62[35:55])
    defparam i47578_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 mult_24_i253_2_lut (.I0(\Ki[5] ), .I1(n356), .I2(GND_net), 
            .I3(GND_net), .O(n375));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i253_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i46059_4_lut (.I0(n455[17]), .I1(n63818), .I2(n34[17]), .I3(n61713), 
            .O(n60771));
    defparam i46059_4_lut.LUT_INIT = 16'h5a7b;
    SB_LUT4 i48075_4_lut (.I0(n32_adj_4733), .I1(n12_adj_4732), .I2(n63827), 
            .I3(n60763), .O(n62788));   // verilog/motorControl.v(62[35:55])
    defparam i48075_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 mult_24_i302_2_lut (.I0(\Ki[6] ), .I1(n356), .I2(GND_net), 
            .I3(GND_net), .O(n448_adj_4338));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i302_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i351_2_lut (.I0(\Ki[7] ), .I1(n356), .I2(GND_net), 
            .I3(GND_net), .O(n521));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i351_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i46426_3_lut (.I0(n62291), .I1(n34[16]), .I2(n455[16]), .I3(GND_net), 
            .O(n61139));   // verilog/motorControl.v(62[35:55])
    defparam i46426_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i47774_4_lut (.I0(n455[17]), .I1(n63818), .I2(n34[17]), .I3(n61719), 
            .O(n62487));
    defparam i47774_4_lut.LUT_INIT = 16'hffde;
    SB_LUT4 LessThan_28_i37_rep_119_2_lut (.I0(n455[18]), .I1(n34[18]), 
            .I2(GND_net), .I3(GND_net), .O(n63827));   // verilog/motorControl.v(62[35:55])
    defparam LessThan_28_i37_rep_119_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_24_i400_2_lut (.I0(\Ki[8] ), .I1(n356), .I2(GND_net), 
            .I3(GND_net), .O(n594));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i400_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i449_2_lut (.I0(\Ki[9] ), .I1(n356), .I2(GND_net), 
            .I3(GND_net), .O(n667));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i449_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i48185_4_lut (.I0(n61139), .I1(n62788), .I2(n63827), .I3(n60771), 
            .O(n62898));   // verilog/motorControl.v(62[35:55])
    defparam i48185_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 mult_24_i498_2_lut (.I0(\Ki[10] ), .I1(n356), .I2(GND_net), 
            .I3(GND_net), .O(n740));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i498_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i47722_4_lut (.I0(n61137), .I1(n61883), .I2(n63834), .I3(n61727), 
            .O(n62435));   // verilog/motorControl.v(62[35:55])
    defparam i47722_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i48282_4_lut (.I0(n62435), .I1(n62898), .I2(n63827), .I3(n62487), 
            .O(n62995));   // verilog/motorControl.v(62[35:55])
    defparam i48282_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i48283_3_lut (.I0(n62995), .I1(n34[19]), .I2(n455[19]), .I3(GND_net), 
            .O(n62996));   // verilog/motorControl.v(62[35:55])
    defparam i48283_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i48074_3_lut (.I0(n62996), .I1(n34[20]), .I2(n455[20]), .I3(GND_net), 
            .O(n62787));   // verilog/motorControl.v(62[35:55])
    defparam i48074_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i47882_3_lut (.I0(n62787), .I1(n34[21]), .I2(n455[21]), .I3(GND_net), 
            .O(n62595));   // verilog/motorControl.v(62[35:55])
    defparam i47882_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i47883_3_lut (.I0(n62595), .I1(n34[22]), .I2(n455[22]), .I3(GND_net), 
            .O(n62596));   // verilog/motorControl.v(62[35:55])
    defparam i47883_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 mult_23_i228_2_lut (.I0(\Kp[4] ), .I1(n207[19]), .I2(GND_net), 
            .I3(GND_net), .O(n338_c));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i228_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_26_i8_3_lut (.I0(n455[3]), .I1(n455[4]), .I2(n9_adj_4728), 
            .I3(GND_net), .O(n8_adj_4742));   // verilog/motorControl.v(62[14:31])
    defparam LessThan_26_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i47730_3_lut (.I0(n8_adj_4742), .I1(n455[11]), .I2(n23_adj_4721), 
            .I3(GND_net), .O(n62443));   // verilog/motorControl.v(62[14:31])
    defparam i47730_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i47731_3_lut (.I0(n62443), .I1(n455[12]), .I2(n25_adj_4722), 
            .I3(GND_net), .O(n62444));   // verilog/motorControl.v(62[14:31])
    defparam i47731_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i46229_4_lut (.I0(n25_adj_4722), .I1(n23_adj_4721), .I2(n21_adj_4720), 
            .I3(n59961), .O(n60941));
    defparam i46229_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i47168_3_lut (.I0(n10_adj_4734), .I1(n455[10]), .I2(n21_adj_4720), 
            .I3(GND_net), .O(n61881));   // verilog/motorControl.v(62[14:31])
    defparam i47168_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i47528_3_lut (.I0(n62444), .I1(n455[13]), .I2(n27_adj_4723), 
            .I3(GND_net), .O(n62241));   // verilog/motorControl.v(62[14:31])
    defparam i47528_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i47447_4_lut (.I0(n35_adj_4719), .I1(n33_adj_4716), .I2(n31_adj_4717), 
            .I3(n59938), .O(n62160));
    defparam i47447_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i48183_4_lut (.I0(n61129), .I1(n62781), .I2(n37_adj_4715), 
            .I3(n60898), .O(n62896));   // verilog/motorControl.v(62[14:31])
    defparam i48183_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i47726_4_lut (.I0(n62241), .I1(n61881), .I2(n27_adj_4723), 
            .I3(n60941), .O(n62439));   // verilog/motorControl.v(62[14:31])
    defparam i47726_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i48294_4_lut (.I0(n62439), .I1(n62896), .I2(n37_adj_4715), 
            .I3(n62160), .O(n63007));   // verilog/motorControl.v(62[14:31])
    defparam i48294_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i48295_3_lut (.I0(n63007), .I1(n455[19]), .I2(\deadband[19] ), 
            .I3(GND_net), .O(n63008));   // verilog/motorControl.v(62[14:31])
    defparam i48295_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i48289_3_lut (.I0(n63008), .I1(n455[20]), .I2(\deadband[20] ), 
            .I3(GND_net), .O(n63002));   // verilog/motorControl.v(62[14:31])
    defparam i48289_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i47886_3_lut (.I0(n63002), .I1(n455[21]), .I2(\deadband[21] ), 
            .I3(GND_net), .O(n62599));   // verilog/motorControl.v(62[14:31])
    defparam i47886_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i47849_3_lut (.I0(n62596), .I1(n455[23]), .I2(n47), .I3(GND_net), 
            .O(n62562));   // verilog/motorControl.v(62[35:55])
    defparam i47849_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i47887_3_lut (.I0(n62599), .I1(n455[22]), .I2(\deadband[22] ), 
            .I3(GND_net), .O(n62600));   // verilog/motorControl.v(62[14:31])
    defparam i47887_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 mult_24_i326_2_lut (.I0(\Ki[6] ), .I1(n344), .I2(GND_net), 
            .I3(GND_net), .O(n484));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i326_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i21888_4_lut (.I0(n62600), .I1(n62562), .I2(\deadband[23] ), 
            .I3(n455[23]), .O(n35399));
    defparam i21888_4_lut.LUT_INIT = 16'hecfe;
    SB_LUT4 mult_24_i547_2_lut (.I0(\Ki[11] ), .I1(n356), .I2(GND_net), 
            .I3(GND_net), .O(n813));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i547_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i596_2_lut (.I0(\Ki[12] ), .I1(n356), .I2(GND_net), 
            .I3(GND_net), .O(n886));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i596_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i645_2_lut (.I0(\Ki[13] ), .I1(n356), .I2(GND_net), 
            .I3(GND_net), .O(n959));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i645_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i694_2_lut (.I0(\Ki[14] ), .I1(n356), .I2(GND_net), 
            .I3(GND_net), .O(n1032));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i694_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i743_2_lut (.I0(\Ki[15] ), .I1(n356), .I2(GND_net), 
            .I3(GND_net), .O(n1105));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i743_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i55_2_lut (.I0(\Ki[1] ), .I1(n357), .I2(GND_net), 
            .I3(GND_net), .O(n80));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i55_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i8_2_lut (.I0(\Ki[0] ), .I1(n356), .I2(GND_net), .I3(GND_net), 
            .O(n11_adj_4337));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i8_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i104_2_lut (.I0(\Ki[2] ), .I1(n357), .I2(GND_net), 
            .I3(GND_net), .O(n153));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i104_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i153_2_lut (.I0(\Ki[3] ), .I1(n357), .I2(GND_net), 
            .I3(GND_net), .O(n226_adj_4336));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i153_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i202_2_lut (.I0(\Ki[4] ), .I1(n357), .I2(GND_net), 
            .I3(GND_net), .O(n299_adj_4335));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i202_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i251_2_lut (.I0(\Ki[5] ), .I1(n357), .I2(GND_net), 
            .I3(GND_net), .O(n372));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i251_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i300_2_lut (.I0(\Ki[6] ), .I1(n357), .I2(GND_net), 
            .I3(GND_net), .O(n445_adj_4334));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i300_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i349_2_lut (.I0(\Ki[7] ), .I1(n357), .I2(GND_net), 
            .I3(GND_net), .O(n518));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i349_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i398_2_lut (.I0(\Ki[8] ), .I1(n357), .I2(GND_net), 
            .I3(GND_net), .O(n591));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i398_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i447_2_lut (.I0(\Ki[9] ), .I1(n357), .I2(GND_net), 
            .I3(GND_net), .O(n664));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i447_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i496_2_lut (.I0(\Ki[10] ), .I1(n357), .I2(GND_net), 
            .I3(GND_net), .O(n737));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i496_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i545_2_lut (.I0(\Ki[11] ), .I1(n357), .I2(GND_net), 
            .I3(GND_net), .O(n810));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i545_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i594_2_lut (.I0(\Ki[12] ), .I1(n357), .I2(GND_net), 
            .I3(GND_net), .O(n883));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i594_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i643_2_lut (.I0(\Ki[13] ), .I1(n357), .I2(GND_net), 
            .I3(GND_net), .O(n956));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i643_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i3_4_lut (.I0(n6646), .I1(n6648), .I2(n22268), .I3(n35687), 
            .O(n4357));
    defparam i3_4_lut.LUT_INIT = 16'hefff;
    SB_LUT4 i45891_4_lut (.I0(n27_adj_4618), .I1(n15_adj_4624), .I2(n13_adj_4623), 
            .I3(n11_adj_4622), .O(n60603));
    defparam i45891_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 LessThan_32_i12_3_lut (.I0(n535[7]), .I1(n535[16]), .I2(n33_adj_4713), 
            .I3(GND_net), .O(n12_adj_4743));   // verilog/motorControl.v(65[25:41])
    defparam LessThan_32_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_24_i692_2_lut (.I0(\Ki[14] ), .I1(n357), .I2(GND_net), 
            .I3(GND_net), .O(n1029));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i692_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i741_2_lut (.I0(\Ki[15] ), .I1(n357), .I2(GND_net), 
            .I3(GND_net), .O(n1102));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i741_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_32_i10_3_lut (.I0(n535[5]), .I1(n535[6]), .I2(n13_adj_4623), 
            .I3(GND_net), .O(n10_adj_4744));   // verilog/motorControl.v(65[25:41])
    defparam LessThan_32_i10_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_32_i30_3_lut (.I0(n12_adj_4743), .I1(n535[17]), .I2(n35_adj_4617), 
            .I3(GND_net), .O(n30_adj_4745));   // verilog/motorControl.v(65[25:41])
    defparam LessThan_32_i30_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i46868_4_lut (.I0(n13_adj_4623), .I1(n11_adj_4622), .I2(n9_adj_4621), 
            .I3(n60648), .O(n61581));
    defparam i46868_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i46858_4_lut (.I0(n19_adj_4615), .I1(n17_adj_4614), .I2(n15_adj_4624), 
            .I3(n61581), .O(n61571));
    defparam i46858_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i47978_4_lut (.I0(n25_adj_4613), .I1(n23_adj_4612), .I2(n21_adj_4611), 
            .I3(n61571), .O(n62691));
    defparam i47978_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i47333_4_lut (.I0(n31_adj_4620), .I1(n29_adj_4619), .I2(n27_adj_4618), 
            .I3(n62691), .O(n62046));
    defparam i47333_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i48105_4_lut (.I0(n37_adj_4616), .I1(n35_adj_4617), .I2(n33_adj_4713), 
            .I3(n62046), .O(n62818));
    defparam i48105_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i47563_3_lut (.I0(n6_adj_4746), .I1(n535[10]), .I2(n21_adj_4611), 
            .I3(GND_net), .O(n62276));   // verilog/motorControl.v(65[25:41])
    defparam i47563_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i47564_3_lut (.I0(n62276), .I1(n535[11]), .I2(n23_adj_4612), 
            .I3(GND_net), .O(n62277));   // verilog/motorControl.v(65[25:41])
    defparam i47564_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_32_i16_3_lut (.I0(n535[9]), .I1(n535[21]), .I2(n43_adj_4610), 
            .I3(GND_net), .O(n16_adj_4747));   // verilog/motorControl.v(65[25:41])
    defparam LessThan_32_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_32_i8_3_lut (.I0(n535[4]), .I1(n535[8]), .I2(n17_adj_4614), 
            .I3(GND_net), .O(n8_adj_4748));   // verilog/motorControl.v(65[25:41])
    defparam LessThan_32_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_32_i24_3_lut (.I0(n16_adj_4747), .I1(n535[22]), .I2(n45_adj_4609), 
            .I3(GND_net), .O(n24_adj_4749));   // verilog/motorControl.v(65[25:41])
    defparam LessThan_32_i24_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i45901_4_lut (.I0(n21_adj_4611), .I1(n19_adj_4615), .I2(n17_adj_4614), 
            .I3(n9_adj_4621), .O(n60613));
    defparam i45901_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i45847_4_lut (.I0(n43_adj_4610), .I1(n25_adj_4613), .I2(n23_adj_4612), 
            .I3(n60613), .O(n60559));
    defparam i45847_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i47174_4_lut (.I0(n24_adj_4749), .I1(n8_adj_4748), .I2(n45_adj_4609), 
            .I3(n60555), .O(n61887));   // verilog/motorControl.v(65[25:41])
    defparam i47174_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 mult_24_i53_2_lut (.I0(\Ki[1] ), .I1(n358), .I2(GND_net), 
            .I3(GND_net), .O(n77));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i53_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i6_2_lut (.I0(\Ki[0] ), .I1(n357), .I2(GND_net), .I3(GND_net), 
            .O(n8_adj_4333));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i6_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i46444_3_lut (.I0(n62277), .I1(n535[12]), .I2(n25_adj_4613), 
            .I3(GND_net), .O(n61157));   // verilog/motorControl.v(65[25:41])
    defparam i46444_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_24_i102_2_lut (.I0(\Ki[2] ), .I1(n358), .I2(GND_net), 
            .I3(GND_net), .O(n150));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i102_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i151_2_lut (.I0(\Ki[3] ), .I1(n358), .I2(GND_net), 
            .I3(GND_net), .O(n223_adj_4332));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i151_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i200_2_lut (.I0(\Ki[4] ), .I1(n358), .I2(GND_net), 
            .I3(GND_net), .O(n296_adj_4331));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i200_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i47559_3_lut (.I0(n4_adj_4750), .I1(n535[13]), .I2(n27_adj_4618), 
            .I3(GND_net), .O(n62272));   // verilog/motorControl.v(65[25:41])
    defparam i47559_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i47560_3_lut (.I0(n62272), .I1(n535[14]), .I2(n29_adj_4619), 
            .I3(GND_net), .O(n62273));   // verilog/motorControl.v(65[25:41])
    defparam i47560_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 n9440_bdd_4_lut_48643 (.I0(n9440), .I1(n59851), .I2(setpoint[4]), 
            .I3(n4357), .O(n63365));
    defparam n9440_bdd_4_lut_48643.LUT_INIT = 16'he4aa;
    SB_LUT4 i45877_4_lut (.I0(n33_adj_4713), .I1(n31_adj_4620), .I2(n29_adj_4619), 
            .I3(n60603), .O(n60589));
    defparam i45877_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 mult_24_i249_2_lut (.I0(\Ki[5] ), .I1(n358), .I2(GND_net), 
            .I3(GND_net), .O(n369));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i249_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i298_2_lut (.I0(\Ki[6] ), .I1(n358), .I2(GND_net), 
            .I3(GND_net), .O(n442_adj_4330));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i298_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i47870_4_lut (.I0(n30_adj_4745), .I1(n10_adj_4744), .I2(n35_adj_4617), 
            .I3(n60585), .O(n62583));   // verilog/motorControl.v(65[25:41])
    defparam i47870_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i46446_3_lut (.I0(n62273), .I1(n535[15]), .I2(n31_adj_4620), 
            .I3(GND_net), .O(n61159));   // verilog/motorControl.v(65[25:41])
    defparam i46446_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_24_i347_2_lut (.I0(\Ki[7] ), .I1(n358), .I2(GND_net), 
            .I3(GND_net), .O(n515));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i347_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i48189_4_lut (.I0(n61159), .I1(n62583), .I2(n35_adj_4617), 
            .I3(n60589), .O(n62902));   // verilog/motorControl.v(65[25:41])
    defparam i48189_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 mult_24_i396_2_lut (.I0(\Ki[8] ), .I1(n358), .I2(GND_net), 
            .I3(GND_net), .O(n588));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i396_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i48190_3_lut (.I0(n62902), .I1(n535[18]), .I2(n37_adj_4616), 
            .I3(GND_net), .O(n62903));   // verilog/motorControl.v(65[25:41])
    defparam i48190_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i48161_3_lut (.I0(n62903), .I1(n535[19]), .I2(n39_adj_4608), 
            .I3(GND_net), .O(n62874));   // verilog/motorControl.v(65[25:41])
    defparam i48161_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i45853_4_lut (.I0(n43_adj_4610), .I1(n41_adj_4607), .I2(n39_adj_4608), 
            .I3(n62818), .O(n60565));
    defparam i45853_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 mult_24_i445_2_lut (.I0(\Ki[9] ), .I1(n358), .I2(GND_net), 
            .I3(GND_net), .O(n661));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i445_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i47852_4_lut (.I0(n61157), .I1(n61887), .I2(n45_adj_4609), 
            .I3(n60559), .O(n62565));   // verilog/motorControl.v(65[25:41])
    defparam i47852_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 mult_24_i494_2_lut (.I0(\Ki[10] ), .I1(n358), .I2(GND_net), 
            .I3(GND_net), .O(n734));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i494_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i543_2_lut (.I0(\Ki[11] ), .I1(n358), .I2(GND_net), 
            .I3(GND_net), .O(n807));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i543_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i592_2_lut (.I0(\Ki[12] ), .I1(n358), .I2(GND_net), 
            .I3(GND_net), .O(n880));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i592_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i641_2_lut (.I0(\Ki[13] ), .I1(n358), .I2(GND_net), 
            .I3(GND_net), .O(n953));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i641_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 n63365_bdd_4_lut (.I0(n63365), .I1(n535[4]), .I2(n455[4]), 
            .I3(n4357), .O(n63368));
    defparam n63365_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i46452_3_lut (.I0(n62874), .I1(n535[20]), .I2(n41_adj_4607), 
            .I3(GND_net), .O(n61165));   // verilog/motorControl.v(65[25:41])
    defparam i46452_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_24_i690_2_lut (.I0(\Ki[14] ), .I1(n358), .I2(GND_net), 
            .I3(GND_net), .O(n1026));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i690_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i739_2_lut (.I0(\Ki[15] ), .I1(n358), .I2(GND_net), 
            .I3(GND_net), .O(n1099));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i739_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i51_2_lut (.I0(\Ki[1] ), .I1(n359), .I2(GND_net), 
            .I3(GND_net), .O(n74_adj_4329));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i51_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i4_2_lut (.I0(\Ki[0] ), .I1(n358), .I2(GND_net), .I3(GND_net), 
            .O(n5_adj_4328));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i4_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i100_2_lut (.I0(\Ki[2] ), .I1(n359), .I2(GND_net), 
            .I3(GND_net), .O(n147));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i100_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i149_2_lut (.I0(\Ki[3] ), .I1(n359), .I2(GND_net), 
            .I3(GND_net), .O(n220_adj_4327));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i149_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i198_2_lut (.I0(\Ki[4] ), .I1(n359), .I2(GND_net), 
            .I3(GND_net), .O(n293_adj_4326));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i198_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i247_2_lut (.I0(\Ki[5] ), .I1(n359), .I2(GND_net), 
            .I3(GND_net), .O(n366));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i247_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i296_2_lut (.I0(\Ki[6] ), .I1(n359), .I2(GND_net), 
            .I3(GND_net), .O(n439_adj_4325));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i296_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i32256_3_lut_4_lut (.I0(\Ki[0] ), .I1(n337), .I2(n338), .I3(\Ki[1] ), 
            .O(n18055[0]));   // verilog/motorControl.v(61[29:40])
    defparam i32256_3_lut_4_lut.LUT_INIT = 16'h7888;
    SB_LUT4 i48044_4_lut (.I0(n61165), .I1(n62565), .I2(n45_adj_4609), 
            .I3(n60565), .O(n62757));   // verilog/motorControl.v(65[25:41])
    defparam i48044_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 mult_24_i345_2_lut (.I0(\Ki[7] ), .I1(n359), .I2(GND_net), 
            .I3(GND_net), .O(n512));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i345_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i2_4_lut (.I0(n62757), .I1(n4_adj_4751), .I2(n455[23]), .I3(n535[23]), 
            .O(n54971));
    defparam i2_4_lut.LUT_INIT = 16'hdfcd;
    SB_LUT4 mult_24_i394_2_lut (.I0(\Ki[8] ), .I1(n359), .I2(GND_net), 
            .I3(GND_net), .O(n585));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i394_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i443_2_lut (.I0(\Ki[9] ), .I1(n359), .I2(GND_net), 
            .I3(GND_net), .O(n658));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i443_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i4200_4_lut (.I0(n6646), .I1(n4357), .I2(n54971), .I3(n22302), 
            .O(n9440));
    defparam i4200_4_lut.LUT_INIT = 16'hbbab;
    SB_LUT4 i32258_3_lut_4_lut (.I0(\Ki[0] ), .I1(n337), .I2(n338), .I3(\Ki[1] ), 
            .O(n45721));   // verilog/motorControl.v(61[29:40])
    defparam i32258_3_lut_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 mult_24_i492_2_lut (.I0(\Ki[10] ), .I1(n359), .I2(GND_net), 
            .I3(GND_net), .O(n731));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i492_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i541_2_lut (.I0(\Ki[11] ), .I1(n359), .I2(GND_net), 
            .I3(GND_net), .O(n804));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i541_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i590_2_lut (.I0(\Ki[12] ), .I1(n359), .I2(GND_net), 
            .I3(GND_net), .O(n877));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i590_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i279_2_lut (.I0(\Ki[5] ), .I1(n343), .I2(GND_net), 
            .I3(GND_net), .O(n414_adj_4223));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i279_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i639_2_lut (.I0(\Ki[13] ), .I1(n359), .I2(GND_net), 
            .I3(GND_net), .O(n950));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i639_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i41909_2_lut (.I0(counter[13]), .I1(counter[11]), .I2(GND_net), 
            .I3(GND_net), .O(n56609));
    defparam i41909_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i9_4_lut (.I0(counter[8]), .I1(counter[0]), .I2(counter[2]), 
            .I3(counter[4]), .O(n23_adj_4752));
    defparam i9_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i8_4_lut (.I0(counter[1]), .I1(counter[6]), .I2(counter[10]), 
            .I3(counter[5]), .O(n22_adj_4753));
    defparam i8_4_lut.LUT_INIT = 16'hffef;
    SB_LUT4 mult_24_i688_2_lut (.I0(\Ki[14] ), .I1(n359), .I2(GND_net), 
            .I3(GND_net), .O(n1023));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i688_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i12_4_lut (.I0(n23_adj_4752), .I1(counter[3]), .I2(n56609), 
            .I3(counter[9]), .O(n26_adj_4754));
    defparam i12_4_lut.LUT_INIT = 16'hefff;
    SB_LUT4 mux_21_i1_3_lut (.I0(n233[0]), .I1(n285[0]), .I2(n284), .I3(GND_net), 
            .O(n310[0]));   // verilog/motorControl.v(58[20] 60[14])
    defparam mux_21_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_22_i1_3_lut (.I0(n310[0]), .I1(IntegralLimit[0]), .I2(n258), 
            .I3(GND_net), .O(n359));   // verilog/motorControl.v(58[20] 60[14])
    defparam mux_22_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_24_i737_2_lut (.I0(\Ki[15] ), .I1(n359), .I2(GND_net), 
            .I3(GND_net), .O(n1096));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i737_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i48346_4_lut (.I0(counter[12]), .I1(n26_adj_4754), .I2(n22_adj_4753), 
            .I3(counter[7]), .O(counter_31__N_3487));   // verilog/motorControl.v(27[8:42])
    defparam i48346_4_lut.LUT_INIT = 16'h0200;
    SB_LUT4 unary_minus_20_inv_0_i5_1_lut (.I0(IntegralLimit[4]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n36[4]));   // verilog/motorControl.v(59[24:38])
    defparam unary_minus_20_inv_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_24_i328_2_lut (.I0(\Ki[6] ), .I1(n343), .I2(GND_net), 
            .I3(GND_net), .O(n487_adj_4220));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i328_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i73_2_lut (.I0(\Kp[1] ), .I1(n207[15]), .I2(GND_net), 
            .I3(GND_net), .O(n107_adj_4324));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i73_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i26_2_lut (.I0(\Kp[0] ), .I1(n207[16]), .I2(GND_net), 
            .I3(GND_net), .O(n38_adj_4323));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i26_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i122_2_lut (.I0(\Kp[2] ), .I1(n207[15]), .I2(GND_net), 
            .I3(GND_net), .O(n180_adj_4322));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i122_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i171_2_lut (.I0(\Kp[3] ), .I1(n207[15]), .I2(GND_net), 
            .I3(GND_net), .O(n253_adj_4321));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i171_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i220_2_lut (.I0(\Kp[4] ), .I1(n207[15]), .I2(GND_net), 
            .I3(GND_net), .O(n326_adj_4320));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i220_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i269_2_lut (.I0(\Kp[5] ), .I1(n207[15]), .I2(GND_net), 
            .I3(GND_net), .O(n399_adj_4319));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i269_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i318_2_lut (.I0(\Kp[6] ), .I1(n207[15]), .I2(GND_net), 
            .I3(GND_net), .O(n472_adj_4317));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i318_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i32306_2_lut_3_lut_4_lut (.I0(\Ki[0] ), .I1(n338), .I2(n339), 
            .I3(\Ki[1] ), .O(n18034[0]));   // verilog/motorControl.v(61[29:40])
    defparam i32306_2_lut_3_lut_4_lut.LUT_INIT = 16'h7888;
    SB_LUT4 mult_23_i367_2_lut (.I0(\Kp[7] ), .I1(n207[15]), .I2(GND_net), 
            .I3(GND_net), .O(n545_adj_4316));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i367_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i32308_2_lut_3_lut_4_lut (.I0(\Ki[0] ), .I1(n338), .I2(n339), 
            .I3(\Ki[1] ), .O(n45772));   // verilog/motorControl.v(61[29:40])
    defparam i32308_2_lut_3_lut_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i45843_2_lut_4_lut (.I0(n455[21]), .I1(n535[21]), .I2(n455[9]), 
            .I3(n535[9]), .O(n60555));
    defparam i45843_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 i1_3_lut_4_lut (.I0(\Ki[3] ), .I1(n340), .I2(n4_adj_4755), 
            .I3(n18034[1]), .O(n17997[2]));   // verilog/motorControl.v(61[29:40])
    defparam i1_3_lut_4_lut.LUT_INIT = 16'h8778;
    SB_LUT4 mult_23_i416_2_lut (.I0(\Kp[8] ), .I1(n207[15]), .I2(GND_net), 
            .I3(GND_net), .O(n618_adj_4315));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i416_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i45873_2_lut_4_lut (.I0(n455[16]), .I1(n535[16]), .I2(n455[7]), 
            .I3(n535[7]), .O(n60585));
    defparam i45873_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 i32374_3_lut_4_lut (.I0(\Ki[3] ), .I1(n340), .I2(n4_adj_4755), 
            .I3(n18034[1]), .O(n6_adj_4276));   // verilog/motorControl.v(61[29:40])
    defparam i32374_3_lut_4_lut.LUT_INIT = 16'hf880;
    SB_LUT4 i32366_3_lut_4_lut (.I0(\Ki[2] ), .I1(n340), .I2(n45825), 
            .I3(n18034[0]), .O(n4_adj_4755));   // verilog/motorControl.v(61[29:40])
    defparam i32366_3_lut_4_lut.LUT_INIT = 16'hf880;
    SB_LUT4 i1_3_lut_4_lut_adj_940 (.I0(\Ki[2] ), .I1(n340), .I2(n45825), 
            .I3(n18034[0]), .O(n17997[1]));   // verilog/motorControl.v(61[29:40])
    defparam i1_3_lut_4_lut_adj_940.LUT_INIT = 16'h8778;
    SB_LUT4 n9440_bdd_4_lut_48633 (.I0(n9440), .I1(n59843), .I2(setpoint[3]), 
            .I3(n4357), .O(n63353));
    defparam n9440_bdd_4_lut_48633.LUT_INIT = 16'he4aa;
    SB_LUT4 i1_2_lut_3_lut (.I0(n52622), .I1(control_update), .I2(n35399), 
            .I3(GND_net), .O(n22266));
    defparam i1_2_lut_3_lut.LUT_INIT = 16'hbfbf;
    SB_LUT4 i32353_2_lut_3_lut_4_lut (.I0(\Ki[0] ), .I1(n339), .I2(n340), 
            .I3(\Ki[1] ), .O(n17997[0]));   // verilog/motorControl.v(61[29:40])
    defparam i32353_2_lut_3_lut_4_lut.LUT_INIT = 16'h7888;
    SB_LUT4 i22175_2_lut_3_lut (.I0(n52622), .I1(control_update), .I2(n35399), 
            .I3(GND_net), .O(n35687));
    defparam i22175_2_lut_3_lut.LUT_INIT = 16'hfbfb;
    SB_LUT4 i32355_2_lut_3_lut_4_lut (.I0(\Ki[0] ), .I1(n339), .I2(n340), 
            .I3(\Ki[1] ), .O(n45825));   // verilog/motorControl.v(61[29:40])
    defparam i32355_2_lut_3_lut_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i32428_3_lut_4_lut (.I0(\Ki[3] ), .I1(n341), .I2(n4_adj_4756), 
            .I3(n17997[1]), .O(n6_adj_4257));   // verilog/motorControl.v(61[29:40])
    defparam i32428_3_lut_4_lut.LUT_INIT = 16'hf880;
    SB_LUT4 n63353_bdd_4_lut (.I0(n63353), .I1(n535[3]), .I2(n455[3]), 
            .I3(n4357), .O(n63356));
    defparam n63353_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 unary_minus_20_inv_0_i6_1_lut (.I0(IntegralLimit[5]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n36[5]));   // verilog/motorControl.v(59[24:38])
    defparam unary_minus_20_inv_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_24_i377_2_lut (.I0(\Ki[7] ), .I1(n343), .I2(GND_net), 
            .I3(GND_net), .O(n560_adj_4214));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i377_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i277_2_lut (.I0(\Kp[5] ), .I1(n207[19]), .I2(GND_net), 
            .I3(GND_net), .O(n411));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i277_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1_3_lut_4_lut_adj_941 (.I0(\Ki[3] ), .I1(n341), .I2(n4_adj_4756), 
            .I3(n17997[1]), .O(n17940[2]));   // verilog/motorControl.v(61[29:40])
    defparam i1_3_lut_4_lut_adj_941.LUT_INIT = 16'h8778;
    SB_LUT4 i1_3_lut_4_lut_adj_942 (.I0(\Ki[2] ), .I1(n341), .I2(n45885), 
            .I3(n17997[0]), .O(n17940[1]));   // verilog/motorControl.v(61[29:40])
    defparam i1_3_lut_4_lut_adj_942.LUT_INIT = 16'h8778;
    SB_LUT4 i32420_3_lut_4_lut (.I0(\Ki[2] ), .I1(n341), .I2(n45885), 
            .I3(n17997[0]), .O(n4_adj_4756));   // verilog/motorControl.v(61[29:40])
    defparam i32420_3_lut_4_lut.LUT_INIT = 16'hf880;
    SB_LUT4 i32407_2_lut_3_lut_4_lut (.I0(\Ki[0] ), .I1(n340), .I2(n341), 
            .I3(\Ki[1] ), .O(n17940[0]));   // verilog/motorControl.v(61[29:40])
    defparam i32407_2_lut_3_lut_4_lut.LUT_INIT = 16'h7888;
    SB_LUT4 mult_23_i63_2_lut (.I0(\Kp[1] ), .I1(n207[10]), .I2(GND_net), 
            .I3(GND_net), .O(n92));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i63_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i16_2_lut (.I0(\Kp[0] ), .I1(n207[11]), .I2(GND_net), 
            .I3(GND_net), .O(n23));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i16_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i46182_2_lut_4_lut (.I0(\deadband[17] ), .I1(n455[17]), .I2(\deadband[8] ), 
            .I3(n455[8]), .O(n60894));
    defparam i46182_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 mult_23_i112_2_lut (.I0(\Kp[2] ), .I1(n207[10]), .I2(GND_net), 
            .I3(GND_net), .O(n165));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i112_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i45249_2_lut_4_lut (.I0(\deadband[9] ), .I1(n455[9]), .I2(\deadband[5] ), 
            .I3(n455[5]), .O(n59961));
    defparam i45249_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 mult_23_i465_2_lut (.I0(\Kp[9] ), .I1(n207[15]), .I2(GND_net), 
            .I3(GND_net), .O(n691_adj_4314));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i465_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i32409_2_lut_3_lut_4_lut (.I0(\Ki[0] ), .I1(n340), .I2(n341), 
            .I3(\Ki[1] ), .O(n45885));   // verilog/motorControl.v(61[29:40])
    defparam i32409_2_lut_3_lut_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 LessThan_9_i8_3_lut_3_lut (.I0(setpoint[4]), .I1(setpoint[8]), 
            .I2(PWMLimit[8]), .I3(GND_net), .O(n8_adj_4710));   // verilog/motorControl.v(45[16:33])
    defparam LessThan_9_i8_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i45849_2_lut_4_lut (.I0(PWMLimit[21]), .I1(setpoint[21]), .I2(PWMLimit[9]), 
            .I3(setpoint[9]), .O(n60561));
    defparam i45849_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 LessThan_9_i16_3_lut_3_lut (.I0(setpoint[9]), .I1(setpoint[21]), 
            .I2(PWMLimit[21]), .I3(GND_net), .O(n16_adj_4708));   // verilog/motorControl.v(45[16:33])
    defparam LessThan_9_i16_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 mult_23_i514_2_lut (.I0(\Kp[10] ), .I1(n207[15]), .I2(GND_net), 
            .I3(GND_net), .O(n764_adj_4312));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i514_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_9_i10_3_lut_3_lut (.I0(setpoint[5]), .I1(setpoint[6]), 
            .I2(PWMLimit[6]), .I3(GND_net), .O(n10_adj_4712));   // verilog/motorControl.v(45[16:33])
    defparam LessThan_9_i10_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i45889_2_lut_4_lut (.I0(PWMLimit[16]), .I1(setpoint[16]), .I2(PWMLimit[7]), 
            .I3(setpoint[7]), .O(n60601));
    defparam i45889_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 LessThan_9_i12_3_lut_3_lut (.I0(setpoint[7]), .I1(setpoint[16]), 
            .I2(PWMLimit[16]), .I3(GND_net), .O(n12_adj_4705));   // verilog/motorControl.v(45[16:33])
    defparam LessThan_9_i12_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 mult_23_i563_2_lut (.I0(\Kp[11] ), .I1(n207[15]), .I2(GND_net), 
            .I3(GND_net), .O(n837_adj_4311));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i563_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_20_inv_0_i7_1_lut (.I0(IntegralLimit[6]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n36[6]));   // verilog/motorControl.v(59[24:38])
    defparam unary_minus_20_inv_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_20_inv_0_i8_1_lut (.I0(IntegralLimit[7]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n36[7]));   // verilog/motorControl.v(59[24:38])
    defparam unary_minus_20_inv_0_i8_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_23_i161_2_lut (.I0(\Kp[3] ), .I1(n207[10]), .I2(GND_net), 
            .I3(GND_net), .O(n238));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i161_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_20_inv_0_i9_1_lut (.I0(IntegralLimit[8]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n36[8]));   // verilog/motorControl.v(59[24:38])
    defparam unary_minus_20_inv_0_i9_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1_2_lut_3_lut_adj_943 (.I0(control_update), .I1(n52622), .I2(n105), 
            .I3(GND_net), .O(n6648));
    defparam i1_2_lut_3_lut_adj_943.LUT_INIT = 16'h8080;
    SB_LUT4 i1_2_lut_3_lut_4_lut (.I0(control_update), .I1(n52622), .I2(n131), 
            .I3(n105), .O(n22302));
    defparam i1_2_lut_3_lut_4_lut.LUT_INIT = 16'h0080;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_944 (.I0(control_update), .I1(n52622), 
            .I2(n131), .I3(n105), .O(n6646));
    defparam i1_2_lut_3_lut_4_lut_adj_944.LUT_INIT = 16'h0008;
    SB_LUT4 mult_23_i210_2_lut (.I0(\Kp[4] ), .I1(n207[10]), .I2(GND_net), 
            .I3(GND_net), .O(n311));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i210_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i259_2_lut (.I0(\Kp[5] ), .I1(n207[10]), .I2(GND_net), 
            .I3(GND_net), .O(n384));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i259_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_20_inv_0_i10_1_lut (.I0(IntegralLimit[9]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n36[9]));   // verilog/motorControl.v(59[24:38])
    defparam unary_minus_20_inv_0_i10_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 LessThan_9_i6_3_lut_3_lut (.I0(PWMLimit[3]), .I1(setpoint[3]), 
            .I2(setpoint[2]), .I3(GND_net), .O(n6_adj_4707));   // verilog/motorControl.v(45[16:33])
    defparam LessThan_9_i6_3_lut_3_lut.LUT_INIT = 16'hd4d4;
    SB_LUT4 i45961_3_lut_4_lut (.I0(PWMLimit[3]), .I1(setpoint[3]), .I2(setpoint[2]), 
            .I3(PWMLimit[2]), .O(n60673));   // verilog/motorControl.v(45[16:33])
    defparam i45961_3_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 mult_23_i308_2_lut (.I0(\Kp[6] ), .I1(n207[10]), .I2(GND_net), 
            .I3(GND_net), .O(n457));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i308_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_4_lut (.I0(n62755), .I1(PWMLimit[23]), .I2(n455[23]), 
            .I3(n22266), .O(n4_adj_4751));   // verilog/motorControl.v(63[16:31])
    defparam i1_2_lut_4_lut.LUT_INIT = 16'hff8e;
    SB_LUT4 i1_2_lut_4_lut_adj_945 (.I0(n62755), .I1(PWMLimit[23]), .I2(n455[23]), 
            .I3(n22266), .O(n22268));   // verilog/motorControl.v(63[16:31])
    defparam i1_2_lut_4_lut_adj_945.LUT_INIT = 16'hff71;
    SB_LUT4 LessThan_30_i6_3_lut_3_lut (.I0(PWMLimit[3]), .I1(n455[3]), 
            .I2(n455[2]), .I3(GND_net), .O(n6_adj_4680));   // verilog/motorControl.v(63[16:31])
    defparam LessThan_30_i6_3_lut_3_lut.LUT_INIT = 16'hd4d4;
    SB_LUT4 i46020_3_lut_4_lut (.I0(PWMLimit[3]), .I1(n455[3]), .I2(n455[2]), 
            .I3(PWMLimit[2]), .O(n60732));   // verilog/motorControl.v(63[16:31])
    defparam i46020_3_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 i32487_2_lut_3_lut (.I0(\Kp[1] ), .I1(n207[22]), .I2(n68_adj_4662), 
            .I3(GND_net), .O(n17961[0]));   // verilog/motorControl.v(61[20:26])
    defparam i32487_2_lut_3_lut.LUT_INIT = 16'h7878;
    SB_LUT4 i1_3_lut_4_lut_adj_946 (.I0(\Kp[1] ), .I1(n207[22]), .I2(n68_adj_4662), 
            .I3(n56550), .O(n17961[1]));   // verilog/motorControl.v(61[20:26])
    defparam i1_3_lut_4_lut_adj_946.LUT_INIT = 16'h7f80;
    SB_LUT4 n9440_bdd_4_lut_48624 (.I0(n9440), .I1(n59737), .I2(setpoint[2]), 
            .I3(n4357), .O(n63341));
    defparam n9440_bdd_4_lut_48624.LUT_INIT = 16'he4aa;
    SB_LUT4 n9440_bdd_4_lut_48787 (.I0(n9440), .I1(n59908), .I2(setpoint[22]), 
            .I3(n4357), .O(n63509));
    defparam n9440_bdd_4_lut_48787.LUT_INIT = 16'he4aa;
    SB_LUT4 unary_minus_20_inv_0_i11_1_lut (.I0(IntegralLimit[10]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n36[10]));   // verilog/motorControl.v(59[24:38])
    defparam unary_minus_20_inv_0_i11_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_23_i357_2_lut (.I0(\Kp[7] ), .I1(n207[10]), .I2(GND_net), 
            .I3(GND_net), .O(n530));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i357_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i45841_3_lut_4_lut (.I0(setpoint[3]), .I1(n535[3]), .I2(n535[2]), 
            .I3(setpoint[2]), .O(n60553));   // verilog/motorControl.v(47[25:43])
    defparam i45841_3_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 mult_23_i406_2_lut (.I0(\Kp[8] ), .I1(n207[10]), .I2(GND_net), 
            .I3(GND_net), .O(n603));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i406_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i45938_2_lut_4_lut (.I0(PWMLimit[21]), .I1(n455[21]), .I2(PWMLimit[9]), 
            .I3(n455[9]), .O(n60650));
    defparam i45938_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 LessThan_11_i6_3_lut_3_lut (.I0(setpoint[3]), .I1(n535[3]), 
            .I2(n535[2]), .I3(GND_net), .O(n6_adj_4648));   // verilog/motorControl.v(47[25:43])
    defparam LessThan_11_i6_3_lut_3_lut.LUT_INIT = 16'hd4d4;
    SB_LUT4 i45971_2_lut_4_lut (.I0(PWMLimit[16]), .I1(n455[16]), .I2(PWMLimit[7]), 
            .I3(n455[7]), .O(n60683));
    defparam i45971_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 mult_23_i612_2_lut (.I0(\Kp[12] ), .I1(n207[15]), .I2(GND_net), 
            .I3(GND_net), .O(n910_adj_4310));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i612_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i46188_2_lut_3_lut (.I0(n6648), .I1(n22268), .I2(PWMLimit[1]), 
            .I3(GND_net), .O(n59723));
    defparam i46188_2_lut_3_lut.LUT_INIT = 16'hb0b0;
    SB_LUT4 n63509_bdd_4_lut (.I0(n63509), .I1(n535[22]), .I2(n455[22]), 
            .I3(n4357), .O(n63512));
    defparam n63509_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i45558_2_lut_3_lut (.I0(n6648), .I1(n22268), .I2(PWMLimit[21]), 
            .I3(GND_net), .O(n59907));
    defparam i45558_2_lut_3_lut.LUT_INIT = 16'hb0b0;
    SB_LUT4 i32331_2_lut_3_lut (.I0(\Kp[0] ), .I1(n207[23]), .I2(\Kp[1] ), 
            .I3(GND_net), .O(n45797));   // verilog/motorControl.v(61[20:26])
    defparam i32331_2_lut_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 i45557_2_lut_3_lut (.I0(n6648), .I1(n22268), .I2(PWMLimit[22]), 
            .I3(GND_net), .O(n59908));
    defparam i45557_2_lut_3_lut.LUT_INIT = 16'hb0b0;
    SB_LUT4 i45426_2_lut_3_lut (.I0(n6648), .I1(n22268), .I2(PWMLimit[2]), 
            .I3(GND_net), .O(n59737));
    defparam i45426_2_lut_3_lut.LUT_INIT = 16'hb0b0;
    SB_LUT4 i32337_2_lut_3_lut (.I0(\Kp[0] ), .I1(\Kp[1] ), .I2(\Kp[2] ), 
            .I3(GND_net), .O(n47176));   // verilog/motorControl.v(61[20:26])
    defparam i32337_2_lut_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 i45548_2_lut_3_lut (.I0(n6648), .I1(n22268), .I2(PWMLimit[3]), 
            .I3(GND_net), .O(n59843));
    defparam i45548_2_lut_3_lut.LUT_INIT = 16'hb0b0;
    SB_LUT4 i45591_2_lut_3_lut (.I0(n6648), .I1(n22268), .I2(PWMLimit[4]), 
            .I3(GND_net), .O(n59851));
    defparam i45591_2_lut_3_lut.LUT_INIT = 16'hb0b0;
    SB_LUT4 LessThan_32_i4_4_lut_4_lut (.I0(n455[0]), .I1(n535[0]), .I2(n455[1]), 
            .I3(n535[1]), .O(n4_adj_4750));   // verilog/motorControl.v(61[20:40])
    defparam LessThan_32_i4_4_lut_4_lut.LUT_INIT = 16'h4f04;
    SB_LUT4 i45520_2_lut_3_lut (.I0(n6648), .I1(n22268), .I2(PWMLimit[23]), 
            .I3(GND_net), .O(n59911));
    defparam i45520_2_lut_3_lut.LUT_INIT = 16'hb0b0;
    SB_LUT4 n63341_bdd_4_lut (.I0(n63341), .I1(n535[2]), .I2(n455[2]), 
            .I3(n4357), .O(n63344));
    defparam n63341_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i45595_2_lut_3_lut (.I0(n6648), .I1(n22268), .I2(PWMLimit[5]), 
            .I3(GND_net), .O(n59882));
    defparam i45595_2_lut_3_lut.LUT_INIT = 16'hb0b0;
    SB_LUT4 i45571_2_lut_3_lut (.I0(n6648), .I1(n22268), .I2(PWMLimit[6]), 
            .I3(GND_net), .O(n59883));
    defparam i45571_2_lut_3_lut.LUT_INIT = 16'hb0b0;
    SB_LUT4 i45570_2_lut_3_lut (.I0(n6648), .I1(n22268), .I2(PWMLimit[7]), 
            .I3(GND_net), .O(n59884));
    defparam i45570_2_lut_3_lut.LUT_INIT = 16'hb0b0;
    SB_LUT4 i45689_2_lut_4_lut (.I0(setpoint[21]), .I1(n535[21]), .I2(setpoint[9]), 
            .I3(n535[9]), .O(n60401));
    defparam i45689_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 i45559_2_lut_3_lut (.I0(n6648), .I1(n22268), .I2(PWMLimit[20]), 
            .I3(GND_net), .O(n59906));
    defparam i45559_2_lut_3_lut.LUT_INIT = 16'hb0b0;
    SB_LUT4 i45729_2_lut_4_lut (.I0(setpoint[16]), .I1(n535[16]), .I2(setpoint[7]), 
            .I3(n535[7]), .O(n60441));
    defparam i45729_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 i45566_2_lut_3_lut (.I0(n6648), .I1(n22268), .I2(PWMLimit[13]), 
            .I3(GND_net), .O(n59899));
    defparam i45566_2_lut_3_lut.LUT_INIT = 16'hb0b0;
    SB_LUT4 mult_23_i71_2_lut (.I0(\Kp[1] ), .I1(n207[14]), .I2(GND_net), 
            .I3(GND_net), .O(n104_adj_4309));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i71_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i24_2_lut (.I0(\Kp[0] ), .I1(n207[15]), .I2(GND_net), 
            .I3(GND_net), .O(n35_adj_4308));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i24_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i45567_2_lut_3_lut (.I0(n6648), .I1(n22268), .I2(PWMLimit[12]), 
            .I3(GND_net), .O(n59898));
    defparam i45567_2_lut_3_lut.LUT_INIT = 16'hb0b0;
    SB_LUT4 i45561_2_lut_3_lut (.I0(n6648), .I1(n22268), .I2(PWMLimit[18]), 
            .I3(GND_net), .O(n59904));
    defparam i45561_2_lut_3_lut.LUT_INIT = 16'hb0b0;
    SB_LUT4 i45560_2_lut_3_lut (.I0(n6648), .I1(n22268), .I2(PWMLimit[19]), 
            .I3(GND_net), .O(n59905));
    defparam i45560_2_lut_3_lut.LUT_INIT = 16'hb0b0;
    SB_LUT4 unary_minus_20_inv_0_i12_1_lut (.I0(IntegralLimit[11]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n36[11]));   // verilog/motorControl.v(59[24:38])
    defparam unary_minus_20_inv_0_i12_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i46208_2_lut_3_lut (.I0(n6648), .I1(n22268), .I2(PWMLimit[0]), 
            .I3(GND_net), .O(n59930));
    defparam i46208_2_lut_3_lut.LUT_INIT = 16'hb0b0;
    SB_LUT4 i45563_2_lut_3_lut (.I0(n6648), .I1(n22268), .I2(PWMLimit[16]), 
            .I3(GND_net), .O(n59902));
    defparam i45563_2_lut_3_lut.LUT_INIT = 16'hb0b0;
    SB_LUT4 mux_21_i14_3_lut (.I0(n233[13]), .I1(n285[13]), .I2(n284), 
            .I3(GND_net), .O(n310[13]));   // verilog/motorControl.v(58[20] 60[14])
    defparam mux_21_i14_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_22_i14_3_lut (.I0(n310[13]), .I1(IntegralLimit[13]), .I2(n258), 
            .I3(GND_net), .O(n346));   // verilog/motorControl.v(58[20] 60[14])
    defparam mux_22_i14_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_24_i75_2_lut (.I0(\Ki[1] ), .I1(n347), .I2(GND_net), 
            .I3(GND_net), .O(n110));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i75_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i45564_2_lut_3_lut (.I0(n6648), .I1(n22268), .I2(PWMLimit[15]), 
            .I3(GND_net), .O(n59901));
    defparam i45564_2_lut_3_lut.LUT_INIT = 16'hb0b0;
    SB_LUT4 mult_24_i28_2_lut (.I0(\Ki[0] ), .I1(n346), .I2(GND_net), 
            .I3(GND_net), .O(n41));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i28_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i124_2_lut (.I0(\Ki[2] ), .I1(n347), .I2(GND_net), 
            .I3(GND_net), .O(n183));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i124_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i45565_2_lut_3_lut (.I0(n6648), .I1(n22268), .I2(PWMLimit[14]), 
            .I3(GND_net), .O(n59900));
    defparam i45565_2_lut_3_lut.LUT_INIT = 16'hb0b0;
    SB_LUT4 mult_23_i120_2_lut (.I0(\Kp[2] ), .I1(n207[14]), .I2(GND_net), 
            .I3(GND_net), .O(n177_adj_4307));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i120_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i45569_2_lut_3_lut (.I0(n6648), .I1(n22268), .I2(PWMLimit[9]), 
            .I3(GND_net), .O(n59886));
    defparam i45569_2_lut_3_lut.LUT_INIT = 16'hb0b0;
    SB_LUT4 i45402_2_lut_3_lut (.I0(n6648), .I1(n22268), .I2(PWMLimit[10]), 
            .I3(GND_net), .O(n59896));
    defparam i45402_2_lut_3_lut.LUT_INIT = 16'hb0b0;
    SB_LUT4 i45568_2_lut_3_lut (.I0(n6648), .I1(n22268), .I2(PWMLimit[11]), 
            .I3(GND_net), .O(n59897));
    defparam i45568_2_lut_3_lut.LUT_INIT = 16'hb0b0;
    SB_LUT4 mult_23_i455_2_lut (.I0(\Kp[9] ), .I1(n207[10]), .I2(GND_net), 
            .I3(GND_net), .O(n676));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i455_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i173_2_lut (.I0(\Ki[3] ), .I1(n347), .I2(GND_net), 
            .I3(GND_net), .O(n256));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i173_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i45562_2_lut_3_lut (.I0(n6648), .I1(n22268), .I2(PWMLimit[17]), 
            .I3(GND_net), .O(n59903));
    defparam i45562_2_lut_3_lut.LUT_INIT = 16'hb0b0;
    SB_LUT4 i45304_2_lut_3_lut (.I0(n6648), .I1(n22268), .I2(PWMLimit[8]), 
            .I3(GND_net), .O(n59885));
    defparam i45304_2_lut_3_lut.LUT_INIT = 16'hb0b0;
    SB_LUT4 n9440_bdd_4_lut_48753 (.I0(n9440), .I1(n59907), .I2(setpoint[21]), 
            .I3(n4357), .O(n63503));
    defparam n9440_bdd_4_lut_48753.LUT_INIT = 16'he4aa;
    SB_LUT4 i45936_3_lut_4_lut (.I0(n455[3]), .I1(n535[3]), .I2(n535[2]), 
            .I3(n455[2]), .O(n60648));   // verilog/motorControl.v(65[25:41])
    defparam i45936_3_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 mult_23_i504_2_lut (.I0(\Kp[10] ), .I1(n207[10]), .I2(GND_net), 
            .I3(GND_net), .O(n749));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i504_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_32_i6_3_lut_3_lut (.I0(n455[3]), .I1(n535[3]), .I2(n535[2]), 
            .I3(GND_net), .O(n6_adj_4746));   // verilog/motorControl.v(65[25:41])
    defparam LessThan_32_i6_3_lut_3_lut.LUT_INIT = 16'hd4d4;
    SB_LUT4 n63503_bdd_4_lut (.I0(n63503), .I1(n535[21]), .I2(n455[21]), 
            .I3(n4357), .O(n63506));
    defparam n63503_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 mult_23_i169_2_lut (.I0(\Kp[3] ), .I1(n207[14]), .I2(GND_net), 
            .I3(GND_net), .O(n250_adj_4305));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i169_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i218_2_lut (.I0(\Kp[4] ), .I1(n207[14]), .I2(GND_net), 
            .I3(GND_net), .O(n323_adj_4302));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i218_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_20_inv_0_i13_1_lut (.I0(IntegralLimit[12]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n36[12]));   // verilog/motorControl.v(59[24:38])
    defparam unary_minus_20_inv_0_i13_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_24_i222_2_lut (.I0(\Ki[4] ), .I1(n347), .I2(GND_net), 
            .I3(GND_net), .O(n329));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i222_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i553_2_lut (.I0(\Kp[11] ), .I1(n207[10]), .I2(GND_net), 
            .I3(GND_net), .O(n822));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i553_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i271_2_lut (.I0(\Ki[5] ), .I1(n347), .I2(GND_net), 
            .I3(GND_net), .O(n402));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i271_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i602_2_lut (.I0(\Kp[12] ), .I1(n207[10]), .I2(GND_net), 
            .I3(GND_net), .O(n895));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i602_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i45456_3_lut_4_lut (.I0(n233[3]), .I1(n285[3]), .I2(n285[2]), 
            .I3(n233[2]), .O(n60168));   // verilog/motorControl.v(58[23:46])
    defparam i45456_3_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 unary_minus_20_inv_0_i14_1_lut (.I0(IntegralLimit[13]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n36[13]));   // verilog/motorControl.v(59[24:38])
    defparam unary_minus_20_inv_0_i14_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 LessThan_19_i6_3_lut_3_lut (.I0(n233[3]), .I1(n285[3]), .I2(n285[2]), 
            .I3(GND_net), .O(n6_adj_4301));   // verilog/motorControl.v(58[23:46])
    defparam LessThan_19_i6_3_lut_3_lut.LUT_INIT = 16'hd4d4;
    SB_LUT4 mult_24_i320_2_lut (.I0(\Ki[6] ), .I1(n347), .I2(GND_net), 
            .I3(GND_net), .O(n475));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i320_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i651_2_lut (.I0(\Kp[13] ), .I1(n207[10]), .I2(GND_net), 
            .I3(GND_net), .O(n968));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i651_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i369_2_lut (.I0(\Ki[7] ), .I1(n347), .I2(GND_net), 
            .I3(GND_net), .O(n548));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i369_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i45687_3_lut_4_lut (.I0(IntegralLimit[3]), .I1(n233[3]), .I2(n233[2]), 
            .I3(IntegralLimit[2]), .O(n60399));   // verilog/motorControl.v(56[14:36])
    defparam i45687_3_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 mult_23_i700_2_lut (.I0(\Kp[14] ), .I1(n207[10]), .I2(GND_net), 
            .I3(GND_net), .O(n1041));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i700_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_17_i6_3_lut_3_lut (.I0(IntegralLimit[3]), .I1(n233[3]), 
            .I2(n233[2]), .I3(GND_net), .O(n6_adj_4250));   // verilog/motorControl.v(56[14:36])
    defparam LessThan_17_i6_3_lut_3_lut.LUT_INIT = 16'hd4d4;
    SB_LUT4 mult_23_i749_2_lut (.I0(\Kp[15] ), .I1(n207[10]), .I2(GND_net), 
            .I3(GND_net), .O(n1114));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i749_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i418_2_lut (.I0(\Ki[8] ), .I1(n347), .I2(GND_net), 
            .I3(GND_net), .O(n621));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i418_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i467_2_lut (.I0(\Ki[9] ), .I1(n347), .I2(GND_net), 
            .I3(GND_net), .O(n694));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i467_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i516_2_lut (.I0(\Ki[10] ), .I1(n347), .I2(GND_net), 
            .I3(GND_net), .O(n767));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i516_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i61_2_lut (.I0(\Kp[1] ), .I1(n207[9]), .I2(GND_net), 
            .I3(GND_net), .O(n89));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i61_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i14_2_lut (.I0(\Kp[0] ), .I1(n207[10]), .I2(GND_net), 
            .I3(GND_net), .O(n20));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i14_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_21_i15_3_lut (.I0(n233[14]), .I1(n285[14]), .I2(n284), 
            .I3(GND_net), .O(n310[14]));   // verilog/motorControl.v(58[20] 60[14])
    defparam mux_21_i15_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_22_i15_3_lut (.I0(n310[14]), .I1(IntegralLimit[14]), .I2(n258), 
            .I3(GND_net), .O(n345));   // verilog/motorControl.v(58[20] 60[14])
    defparam mux_22_i15_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_21_i10_3_lut (.I0(n233[9]), .I1(n285[9]), .I2(n284), .I3(GND_net), 
            .O(n310[9]));   // verilog/motorControl.v(58[20] 60[14])
    defparam mux_21_i10_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_22_i10_3_lut (.I0(n310[9]), .I1(IntegralLimit[9]), .I2(n258), 
            .I3(GND_net), .O(n350));   // verilog/motorControl.v(58[20] 60[14])
    defparam mux_22_i10_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_21_i9_3_lut (.I0(n233[8]), .I1(n285[8]), .I2(n284), .I3(GND_net), 
            .O(n310[8]));   // verilog/motorControl.v(58[20] 60[14])
    defparam mux_21_i9_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_22_i9_3_lut (.I0(n310[8]), .I1(IntegralLimit[8]), .I2(n258), 
            .I3(GND_net), .O(n351));   // verilog/motorControl.v(58[20] 60[14])
    defparam mux_22_i9_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_21_i8_3_lut (.I0(n233[7]), .I1(n285[7]), .I2(n284), .I3(GND_net), 
            .O(n310[7]));   // verilog/motorControl.v(58[20] 60[14])
    defparam mux_21_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_22_i8_3_lut (.I0(n310[7]), .I1(IntegralLimit[7]), .I2(n258), 
            .I3(GND_net), .O(n352));   // verilog/motorControl.v(58[20] 60[14])
    defparam mux_22_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_21_i7_3_lut (.I0(n233[6]), .I1(n285[6]), .I2(n284), .I3(GND_net), 
            .O(n310[6]));   // verilog/motorControl.v(58[20] 60[14])
    defparam mux_21_i7_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_22_i7_3_lut (.I0(n310[6]), .I1(IntegralLimit[6]), .I2(n258), 
            .I3(GND_net), .O(n353));   // verilog/motorControl.v(58[20] 60[14])
    defparam mux_22_i7_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_21_i6_3_lut (.I0(n233[5]), .I1(n285[5]), .I2(n284), .I3(GND_net), 
            .O(n310[5]));   // verilog/motorControl.v(58[20] 60[14])
    defparam mux_21_i6_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_24_i565_2_lut (.I0(\Ki[11] ), .I1(n347), .I2(GND_net), 
            .I3(GND_net), .O(n840));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i565_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_22_i6_3_lut (.I0(n310[5]), .I1(IntegralLimit[5]), .I2(n258), 
            .I3(GND_net), .O(n354));   // verilog/motorControl.v(58[20] 60[14])
    defparam mux_22_i6_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_23_i110_2_lut (.I0(\Kp[2] ), .I1(n207[9]), .I2(GND_net), 
            .I3(GND_net), .O(n162));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i110_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_21_i5_3_lut (.I0(n233[4]), .I1(n285[4]), .I2(n284), .I3(GND_net), 
            .O(n310[4]));   // verilog/motorControl.v(58[20] 60[14])
    defparam mux_21_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_22_i5_3_lut (.I0(n310[4]), .I1(IntegralLimit[4]), .I2(n258), 
            .I3(GND_net), .O(n355));   // verilog/motorControl.v(58[20] 60[14])
    defparam mux_22_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_21_i4_3_lut (.I0(n233[3]), .I1(n285[3]), .I2(n284), .I3(GND_net), 
            .O(n310[3]));   // verilog/motorControl.v(58[20] 60[14])
    defparam mux_21_i4_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_22_i4_3_lut (.I0(n310[3]), .I1(IntegralLimit[3]), .I2(n258), 
            .I3(GND_net), .O(n356));   // verilog/motorControl.v(58[20] 60[14])
    defparam mux_22_i4_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_21_i3_3_lut (.I0(n233[2]), .I1(n285[2]), .I2(n284), .I3(GND_net), 
            .O(n310[2]));   // verilog/motorControl.v(58[20] 60[14])
    defparam mux_21_i3_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_22_i3_3_lut (.I0(n310[2]), .I1(IntegralLimit[2]), .I2(n258), 
            .I3(GND_net), .O(n357));   // verilog/motorControl.v(58[20] 60[14])
    defparam mux_22_i3_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_21_i2_3_lut (.I0(n233[1]), .I1(n285[1]), .I2(n284), .I3(GND_net), 
            .O(n310[1]));   // verilog/motorControl.v(58[20] 60[14])
    defparam mux_21_i2_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_22_i2_3_lut (.I0(n310[1]), .I1(IntegralLimit[1]), .I2(n258), 
            .I3(GND_net), .O(n358));   // verilog/motorControl.v(58[20] 60[14])
    defparam mux_22_i2_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_23_i267_2_lut (.I0(\Kp[5] ), .I1(n207[14]), .I2(GND_net), 
            .I3(GND_net), .O(n396_adj_4300));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i267_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i45269_2_lut_4_lut (.I0(n233[21]), .I1(n285[21]), .I2(n233[9]), 
            .I3(n285[9]), .O(n59981));
    defparam i45269_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 mult_23_i83_2_lut (.I0(\Kp[1] ), .I1(n207[20]), .I2(GND_net), 
            .I3(GND_net), .O(n122));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i83_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i36_2_lut (.I0(\Kp[0] ), .I1(n207[21]), .I2(GND_net), 
            .I3(GND_net), .O(n53_c));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i36_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_20_inv_0_i15_1_lut (.I0(IntegralLimit[14]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n36[14]));   // verilog/motorControl.v(59[24:38])
    defparam unary_minus_20_inv_0_i15_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_23_i132_2_lut (.I0(\Kp[2] ), .I1(n207[20]), .I2(GND_net), 
            .I3(GND_net), .O(n195));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i132_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i159_2_lut (.I0(\Kp[3] ), .I1(n207[9]), .I2(GND_net), 
            .I3(GND_net), .O(n235));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i159_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i181_2_lut (.I0(\Kp[3] ), .I1(n207[20]), .I2(GND_net), 
            .I3(GND_net), .O(n268));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i181_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i45298_2_lut_4_lut (.I0(n233[16]), .I1(n285[16]), .I2(n233[7]), 
            .I3(n285[7]), .O(n60010));
    defparam i45298_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 mult_23_i316_2_lut (.I0(\Kp[6] ), .I1(n207[14]), .I2(GND_net), 
            .I3(GND_net), .O(n469_adj_4298));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i316_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 n9440_bdd_4_lut_48614 (.I0(n9440), .I1(n59723), .I2(setpoint[1]), 
            .I3(n4357), .O(n63275));
    defparam n9440_bdd_4_lut_48614.LUT_INIT = 16'he4aa;
    SB_LUT4 mult_23_i230_2_lut (.I0(\Kp[4] ), .I1(n207[20]), .I2(GND_net), 
            .I3(GND_net), .O(n341_c));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i230_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i279_2_lut (.I0(\Kp[5] ), .I1(n207[20]), .I2(GND_net), 
            .I3(GND_net), .O(n414));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i279_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 n63275_bdd_4_lut (.I0(n63275), .I1(n535[1]), .I2(n455[1]), 
            .I3(n4357), .O(n63278));
    defparam n63275_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 mult_23_i328_2_lut (.I0(\Kp[6] ), .I1(n207[20]), .I2(GND_net), 
            .I3(GND_net), .O(n487));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i328_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i208_2_lut (.I0(\Kp[4] ), .I1(n207[9]), .I2(GND_net), 
            .I3(GND_net), .O(n308));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i208_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i377_2_lut (.I0(\Kp[7] ), .I1(n207[20]), .I2(GND_net), 
            .I3(GND_net), .O(n560));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i377_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i45465_2_lut_4_lut (.I0(IntegralLimit[21]), .I1(n233[21]), .I2(IntegralLimit[9]), 
            .I3(n233[9]), .O(n60177));
    defparam i45465_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 unary_minus_20_inv_0_i16_1_lut (.I0(IntegralLimit[15]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n36[15]));   // verilog/motorControl.v(59[24:38])
    defparam unary_minus_20_inv_0_i16_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mux_21_i13_3_lut (.I0(n233[12]), .I1(n285[12]), .I2(n284), 
            .I3(GND_net), .O(n310[12]));   // verilog/motorControl.v(58[20] 60[14])
    defparam mux_21_i13_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_22_i13_3_lut (.I0(n310[12]), .I1(IntegralLimit[12]), .I2(n258), 
            .I3(GND_net), .O(n347));   // verilog/motorControl.v(58[20] 60[14])
    defparam mux_22_i13_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_23_i365_2_lut (.I0(\Kp[7] ), .I1(n207[14]), .I2(GND_net), 
            .I3(GND_net), .O(n542_adj_4296));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i365_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i73_2_lut (.I0(\Ki[1] ), .I1(n348), .I2(GND_net), 
            .I3(GND_net), .O(n107));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i73_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i414_2_lut (.I0(\Kp[8] ), .I1(n207[14]), .I2(GND_net), 
            .I3(GND_net), .O(n615_adj_4295));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i414_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i26_2_lut (.I0(\Ki[0] ), .I1(n347), .I2(GND_net), 
            .I3(GND_net), .O(n38));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i26_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i45511_2_lut_4_lut (.I0(IntegralLimit[16]), .I1(n233[16]), .I2(IntegralLimit[7]), 
            .I3(n233[7]), .O(n60223));
    defparam i45511_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 mult_23_i257_2_lut (.I0(\Kp[5] ), .I1(n207[9]), .I2(GND_net), 
            .I3(GND_net), .O(n381));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i257_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i122_2_lut (.I0(\Ki[2] ), .I1(n348), .I2(GND_net), 
            .I3(GND_net), .O(n180));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i122_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i463_2_lut (.I0(\Kp[9] ), .I1(n207[14]), .I2(GND_net), 
            .I3(GND_net), .O(n688_adj_4294));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i463_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i512_2_lut (.I0(\Kp[10] ), .I1(n207[14]), .I2(GND_net), 
            .I3(GND_net), .O(n761_adj_4293));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i512_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i561_2_lut (.I0(\Kp[11] ), .I1(n207[14]), .I2(GND_net), 
            .I3(GND_net), .O(n834_adj_4292));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i561_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_27_inv_0_i5_1_lut (.I0(\deadband[4] ), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n28[4]));   // verilog/motorControl.v(62[45:54])
    defparam unary_minus_27_inv_0_i5_1_lut.LUT_INIT = 16'h5555;
    
endmodule
