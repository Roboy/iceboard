// ******************************************************************************

// iCEcube Netlister

// Version:            2017.08.27940

// Build Date:         Sep 12 2017 08:25:46

// File Generated:     Mar 24 2020 18:54:39

// Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

// Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

// ******************************************************************************

// Verilog file for cell "TinyFPGA_B" view "INTERFACE"

module TinyFPGA_B (
    USBPU,
    SPI_IO2,
    PIN_9,
    PIN_8,
    PIN_7,
    PIN_6,
    PIN_5,
    PIN_4,
    PIN_3,
    PIN_24,
    PIN_23,
    PIN_22,
    PIN_21,
    PIN_20,
    PIN_2,
    PIN_19,
    PIN_18,
    PIN_17,
    PIN_16,
    PIN_15,
    PIN_14,
    PIN_13,
    PIN_12,
    PIN_11,
    PIN_10,
    PIN_1,
    LED,
    CLK);

    input USBPU;
    input SPI_IO2;
    input PIN_9;
    input PIN_8;
    input PIN_7;
    input PIN_6;
    input PIN_5;
    input PIN_4;
    input PIN_3;
    input PIN_24;
    input PIN_23;
    input PIN_22;
    input PIN_21;
    input PIN_20;
    output PIN_2;
    input PIN_19;
    output PIN_18;
    input PIN_17;
    input PIN_16;
    input PIN_15;
    input PIN_14;
    inout PIN_13;
    input PIN_12;
    input PIN_11;
    input PIN_10;
    input PIN_1;
    output LED;
    input CLK;

    wire N__5970;
    wire N__5969;
    wire N__5968;
    wire N__5961;
    wire N__5960;
    wire N__5959;
    wire N__5952;
    wire N__5951;
    wire N__5950;
    wire N__5943;
    wire N__5942;
    wire N__5941;
    wire N__5934;
    wire N__5933;
    wire N__5932;
    wire N__5915;
    wire N__5914;
    wire N__5911;
    wire N__5908;
    wire N__5903;
    wire N__5900;
    wire N__5899;
    wire N__5896;
    wire N__5893;
    wire N__5888;
    wire N__5885;
    wire N__5884;
    wire N__5881;
    wire N__5878;
    wire N__5873;
    wire N__5870;
    wire N__5869;
    wire N__5866;
    wire N__5863;
    wire N__5858;
    wire N__5855;
    wire N__5854;
    wire N__5851;
    wire N__5848;
    wire N__5843;
    wire N__5840;
    wire N__5837;
    wire N__5836;
    wire N__5833;
    wire N__5830;
    wire N__5825;
    wire N__5822;
    wire N__5819;
    wire N__5816;
    wire N__5815;
    wire N__5814;
    wire N__5813;
    wire N__5812;
    wire N__5809;
    wire N__5806;
    wire N__5805;
    wire N__5804;
    wire N__5801;
    wire N__5798;
    wire N__5795;
    wire N__5792;
    wire N__5789;
    wire N__5786;
    wire N__5783;
    wire N__5780;
    wire N__5775;
    wire N__5774;
    wire N__5771;
    wire N__5766;
    wire N__5763;
    wire N__5758;
    wire N__5755;
    wire N__5754;
    wire N__5751;
    wire N__5748;
    wire N__5745;
    wire N__5740;
    wire N__5737;
    wire N__5734;
    wire N__5731;
    wire N__5724;
    wire N__5717;
    wire N__5714;
    wire N__5711;
    wire N__5710;
    wire N__5709;
    wire N__5708;
    wire N__5707;
    wire N__5706;
    wire N__5705;
    wire N__5704;
    wire N__5703;
    wire N__5702;
    wire N__5701;
    wire N__5700;
    wire N__5697;
    wire N__5694;
    wire N__5691;
    wire N__5688;
    wire N__5685;
    wire N__5682;
    wire N__5675;
    wire N__5668;
    wire N__5651;
    wire N__5650;
    wire N__5647;
    wire N__5644;
    wire N__5639;
    wire N__5638;
    wire N__5635;
    wire N__5632;
    wire N__5627;
    wire N__5626;
    wire N__5623;
    wire N__5620;
    wire N__5617;
    wire N__5612;
    wire N__5611;
    wire N__5608;
    wire N__5605;
    wire N__5600;
    wire N__5599;
    wire N__5594;
    wire N__5591;
    wire N__5590;
    wire N__5587;
    wire N__5584;
    wire N__5579;
    wire N__5578;
    wire N__5575;
    wire N__5572;
    wire N__5567;
    wire N__5566;
    wire N__5563;
    wire N__5560;
    wire N__5557;
    wire N__5552;
    wire N__5551;
    wire N__5548;
    wire N__5545;
    wire N__5540;
    wire N__5537;
    wire N__5534;
    wire N__5533;
    wire N__5530;
    wire N__5527;
    wire N__5522;
    wire N__5521;
    wire N__5518;
    wire N__5515;
    wire N__5510;
    wire N__5509;
    wire N__5506;
    wire N__5503;
    wire N__5498;
    wire N__5495;
    wire N__5492;
    wire N__5489;
    wire N__5488;
    wire N__5485;
    wire N__5482;
    wire N__5477;
    wire N__5476;
    wire N__5475;
    wire N__5474;
    wire N__5473;
    wire N__5472;
    wire N__5469;
    wire N__5466;
    wire N__5461;
    wire N__5456;
    wire N__5447;
    wire N__5444;
    wire N__5443;
    wire N__5442;
    wire N__5439;
    wire N__5438;
    wire N__5437;
    wire N__5436;
    wire N__5433;
    wire N__5432;
    wire N__5429;
    wire N__5426;
    wire N__5423;
    wire N__5420;
    wire N__5415;
    wire N__5410;
    wire N__5399;
    wire N__5398;
    wire N__5397;
    wire N__5396;
    wire N__5395;
    wire N__5394;
    wire N__5393;
    wire N__5392;
    wire N__5391;
    wire N__5390;
    wire N__5389;
    wire N__5388;
    wire N__5387;
    wire N__5386;
    wire N__5385;
    wire N__5384;
    wire N__5383;
    wire N__5382;
    wire N__5381;
    wire N__5380;
    wire N__5379;
    wire N__5336;
    wire N__5333;
    wire N__5330;
    wire N__5329;
    wire N__5326;
    wire N__5323;
    wire N__5320;
    wire N__5319;
    wire N__5316;
    wire N__5313;
    wire N__5310;
    wire N__5303;
    wire N__5302;
    wire N__5299;
    wire N__5296;
    wire N__5293;
    wire N__5290;
    wire N__5287;
    wire N__5284;
    wire N__5281;
    wire N__5276;
    wire N__5275;
    wire N__5272;
    wire N__5269;
    wire N__5266;
    wire N__5263;
    wire N__5260;
    wire N__5257;
    wire N__5254;
    wire N__5251;
    wire N__5248;
    wire N__5245;
    wire N__5242;
    wire N__5239;
    wire N__5234;
    wire N__5231;
    wire N__5230;
    wire N__5227;
    wire N__5224;
    wire N__5219;
    wire N__5218;
    wire N__5215;
    wire N__5212;
    wire N__5207;
    wire N__5204;
    wire N__5203;
    wire N__5200;
    wire N__5197;
    wire N__5194;
    wire N__5189;
    wire N__5188;
    wire N__5185;
    wire N__5182;
    wire N__5177;
    wire N__5176;
    wire N__5173;
    wire N__5170;
    wire N__5167;
    wire N__5162;
    wire N__5161;
    wire N__5158;
    wire N__5155;
    wire N__5150;
    wire N__5147;
    wire N__5144;
    wire N__5141;
    wire N__5138;
    wire N__5137;
    wire N__5134;
    wire N__5131;
    wire N__5126;
    wire N__5125;
    wire N__5120;
    wire N__5119;
    wire N__5116;
    wire N__5113;
    wire N__5110;
    wire N__5105;
    wire N__5102;
    wire N__5099;
    wire N__5096;
    wire N__5093;
    wire N__5092;
    wire N__5089;
    wire N__5086;
    wire N__5083;
    wire N__5080;
    wire N__5075;
    wire N__5072;
    wire N__5069;
    wire N__5068;
    wire N__5065;
    wire N__5062;
    wire N__5057;
    wire N__5056;
    wire N__5053;
    wire N__5050;
    wire N__5045;
    wire N__5044;
    wire N__5041;
    wire N__5038;
    wire N__5033;
    wire N__5032;
    wire N__5029;
    wire N__5026;
    wire N__5023;
    wire N__5018;
    wire N__5017;
    wire N__5014;
    wire N__5011;
    wire N__5006;
    wire N__5003;
    wire N__5000;
    wire N__4999;
    wire N__4996;
    wire N__4993;
    wire N__4988;
    wire N__4987;
    wire N__4984;
    wire N__4981;
    wire N__4976;
    wire N__4975;
    wire N__4972;
    wire N__4969;
    wire N__4966;
    wire N__4961;
    wire N__4960;
    wire N__4957;
    wire N__4954;
    wire N__4949;
    wire N__4946;
    wire N__4945;
    wire N__4942;
    wire N__4939;
    wire N__4934;
    wire N__4931;
    wire N__4930;
    wire N__4927;
    wire N__4924;
    wire N__4919;
    wire N__4918;
    wire N__4915;
    wire N__4912;
    wire N__4907;
    wire N__4906;
    wire N__4903;
    wire N__4900;
    wire N__4895;
    wire N__4894;
    wire N__4893;
    wire N__4892;
    wire N__4891;
    wire N__4890;
    wire N__4889;
    wire N__4888;
    wire N__4877;
    wire N__4870;
    wire N__4865;
    wire N__4864;
    wire N__4861;
    wire N__4858;
    wire N__4853;
    wire N__4850;
    wire N__4849;
    wire N__4846;
    wire N__4843;
    wire N__4838;
    wire N__4835;
    wire N__4834;
    wire N__4831;
    wire N__4828;
    wire N__4823;
    wire N__4822;
    wire N__4819;
    wire N__4816;
    wire N__4811;
    wire N__4808;
    wire N__4807;
    wire N__4804;
    wire N__4801;
    wire N__4796;
    wire N__4793;
    wire N__4792;
    wire N__4789;
    wire N__4786;
    wire N__4781;
    wire N__4778;
    wire N__4775;
    wire N__4772;
    wire N__4771;
    wire N__4766;
    wire N__4763;
    wire N__4762;
    wire N__4757;
    wire N__4754;
    wire N__4751;
    wire N__4748;
    wire N__4745;
    wire N__4744;
    wire N__4739;
    wire N__4736;
    wire N__4733;
    wire N__4732;
    wire N__4731;
    wire N__4730;
    wire N__4729;
    wire N__4726;
    wire N__4725;
    wire N__4722;
    wire N__4721;
    wire N__4720;
    wire N__4719;
    wire N__4716;
    wire N__4713;
    wire N__4710;
    wire N__4707;
    wire N__4704;
    wire N__4697;
    wire N__4692;
    wire N__4679;
    wire N__4678;
    wire N__4677;
    wire N__4674;
    wire N__4673;
    wire N__4672;
    wire N__4667;
    wire N__4664;
    wire N__4663;
    wire N__4662;
    wire N__4657;
    wire N__4652;
    wire N__4649;
    wire N__4646;
    wire N__4637;
    wire N__4636;
    wire N__4633;
    wire N__4632;
    wire N__4631;
    wire N__4630;
    wire N__4629;
    wire N__4626;
    wire N__4623;
    wire N__4620;
    wire N__4617;
    wire N__4612;
    wire N__4605;
    wire N__4598;
    wire N__4597;
    wire N__4594;
    wire N__4591;
    wire N__4586;
    wire N__4583;
    wire N__4580;
    wire N__4577;
    wire N__4574;
    wire N__4571;
    wire N__4570;
    wire N__4569;
    wire N__4566;
    wire N__4563;
    wire N__4560;
    wire N__4553;
    wire N__4550;
    wire N__4549;
    wire N__4548;
    wire N__4547;
    wire N__4546;
    wire N__4543;
    wire N__4538;
    wire N__4533;
    wire N__4530;
    wire N__4523;
    wire N__4520;
    wire N__4519;
    wire N__4516;
    wire N__4513;
    wire N__4510;
    wire N__4505;
    wire N__4502;
    wire N__4499;
    wire N__4496;
    wire N__4493;
    wire N__4490;
    wire N__4487;
    wire N__4484;
    wire N__4481;
    wire N__4478;
    wire N__4475;
    wire N__4472;
    wire N__4469;
    wire N__4466;
    wire N__4463;
    wire N__4460;
    wire N__4457;
    wire N__4454;
    wire N__4451;
    wire N__4448;
    wire N__4445;
    wire N__4442;
    wire N__4439;
    wire N__4436;
    wire N__4433;
    wire N__4430;
    wire N__4427;
    wire N__4424;
    wire N__4421;
    wire N__4418;
    wire N__4415;
    wire N__4412;
    wire N__4409;
    wire N__4406;
    wire N__4403;
    wire N__4400;
    wire N__4397;
    wire N__4394;
    wire N__4391;
    wire N__4388;
    wire N__4385;
    wire N__4382;
    wire N__4379;
    wire N__4376;
    wire N__4373;
    wire N__4372;
    wire N__4369;
    wire N__4366;
    wire N__4361;
    wire N__4358;
    wire N__4355;
    wire N__4352;
    wire N__4349;
    wire N__4346;
    wire N__4343;
    wire N__4342;
    wire N__4337;
    wire N__4336;
    wire N__4333;
    wire N__4330;
    wire N__4325;
    wire N__4324;
    wire N__4323;
    wire N__4318;
    wire N__4315;
    wire N__4310;
    wire N__4309;
    wire N__4306;
    wire N__4303;
    wire N__4298;
    wire N__4297;
    wire N__4294;
    wire N__4291;
    wire N__4286;
    wire N__4285;
    wire N__4280;
    wire N__4279;
    wire N__4276;
    wire N__4273;
    wire N__4268;
    wire N__4265;
    wire N__4262;
    wire N__4259;
    wire N__4256;
    wire N__4253;
    wire N__4250;
    wire N__4247;
    wire N__4246;
    wire N__4243;
    wire N__4240;
    wire N__4237;
    wire N__4232;
    wire N__4229;
    wire N__4226;
    wire N__4223;
    wire N__4220;
    wire N__4219;
    wire N__4216;
    wire N__4213;
    wire N__4210;
    wire N__4205;
    wire N__4202;
    wire N__4199;
    wire N__4198;
    wire N__4193;
    wire N__4190;
    wire N__4187;
    wire N__4184;
    wire N__4181;
    wire N__4178;
    wire N__4175;
    wire N__4172;
    wire N__4169;
    wire N__4166;
    wire N__4163;
    wire N__4160;
    wire N__4157;
    wire N__4154;
    wire N__4151;
    wire N__4148;
    wire N__4145;
    wire N__4142;
    wire N__4139;
    wire N__4136;
    wire N__4133;
    wire N__4130;
    wire N__4127;
    wire N__4124;
    wire N__4121;
    wire N__4118;
    wire N__4115;
    wire N__4112;
    wire N__4109;
    wire N__4106;
    wire N__4103;
    wire N__4100;
    wire N__4097;
    wire N__4094;
    wire N__4091;
    wire N__4088;
    wire N__4085;
    wire N__4082;
    wire N__4079;
    wire N__4076;
    wire N__4073;
    wire N__4070;
    wire N__4067;
    wire N__4064;
    wire N__4061;
    wire N__4058;
    wire N__4055;
    wire N__4052;
    wire N__4049;
    wire N__4046;
    wire N__4043;
    wire N__4040;
    wire N__4037;
    wire N__4034;
    wire N__4031;
    wire N__4028;
    wire N__4025;
    wire N__4022;
    wire N__4019;
    wire N__4016;
    wire N__4013;
    wire N__4010;
    wire N__4007;
    wire N__4004;
    wire N__4001;
    wire N__3998;
    wire N__3995;
    wire N__3992;
    wire N__3989;
    wire N__3988;
    wire N__3985;
    wire N__3982;
    wire N__3979;
    wire N__3974;
    wire N__3973;
    wire N__3970;
    wire N__3967;
    wire N__3962;
    wire N__3961;
    wire N__3958;
    wire N__3955;
    wire N__3952;
    wire N__3947;
    wire N__3946;
    wire N__3943;
    wire N__3942;
    wire N__3939;
    wire N__3938;
    wire N__3935;
    wire N__3932;
    wire N__3929;
    wire N__3926;
    wire N__3921;
    wire N__3916;
    wire N__3911;
    wire N__3908;
    wire N__3905;
    wire N__3902;
    wire N__3899;
    wire N__3898;
    wire N__3895;
    wire N__3892;
    wire N__3887;
    wire N__3886;
    wire N__3883;
    wire N__3880;
    wire N__3875;
    wire N__3872;
    wire N__3869;
    wire N__3868;
    wire N__3865;
    wire N__3862;
    wire N__3857;
    wire N__3856;
    wire N__3853;
    wire N__3850;
    wire N__3845;
    wire N__3842;
    wire N__3841;
    wire N__3838;
    wire N__3835;
    wire N__3832;
    wire N__3827;
    wire N__3826;
    wire N__3823;
    wire N__3820;
    wire N__3815;
    wire N__3814;
    wire N__3811;
    wire N__3808;
    wire N__3803;
    wire N__3802;
    wire N__3799;
    wire N__3796;
    wire N__3791;
    wire N__3790;
    wire N__3787;
    wire N__3784;
    wire N__3781;
    wire N__3776;
    wire N__3775;
    wire N__3772;
    wire N__3769;
    wire N__3766;
    wire N__3761;
    wire N__3760;
    wire N__3757;
    wire N__3754;
    wire N__3749;
    wire N__3748;
    wire N__3745;
    wire N__3742;
    wire N__3739;
    wire N__3734;
    wire N__3731;
    wire N__3728;
    wire N__3727;
    wire N__3724;
    wire N__3721;
    wire N__3718;
    wire N__3713;
    wire N__3712;
    wire N__3709;
    wire N__3706;
    wire N__3703;
    wire N__3698;
    wire N__3695;
    wire N__3692;
    wire N__3691;
    wire N__3688;
    wire N__3683;
    wire N__3682;
    wire N__3679;
    wire N__3676;
    wire N__3673;
    wire N__3668;
    wire N__3665;
    wire N__3664;
    wire N__3659;
    wire N__3656;
    wire N__3655;
    wire N__3650;
    wire N__3647;
    wire N__3644;
    wire N__3643;
    wire N__3640;
    wire N__3637;
    wire N__3632;
    wire N__3631;
    wire N__3628;
    wire N__3625;
    wire N__3620;
    wire N__3619;
    wire N__3616;
    wire N__3613;
    wire N__3610;
    wire N__3605;
    wire N__3604;
    wire N__3601;
    wire N__3598;
    wire N__3593;
    wire N__3592;
    wire N__3589;
    wire N__3586;
    wire N__3583;
    wire N__3578;
    wire N__3577;
    wire N__3574;
    wire N__3571;
    wire N__3566;
    wire N__3565;
    wire N__3562;
    wire N__3559;
    wire N__3556;
    wire N__3551;
    wire N__3550;
    wire N__3547;
    wire N__3544;
    wire N__3539;
    wire N__3536;
    wire N__3533;
    wire N__3530;
    wire N__3527;
    wire N__3524;
    wire N__3521;
    wire N__3518;
    wire N__3515;
    wire N__3512;
    wire N__3509;
    wire N__3506;
    wire N__3505;
    wire N__3502;
    wire N__3499;
    wire N__3496;
    wire N__3491;
    wire N__3490;
    wire N__3487;
    wire N__3484;
    wire N__3481;
    wire N__3476;
    wire N__3473;
    wire N__3472;
    wire N__3469;
    wire N__3466;
    wire N__3463;
    wire N__3458;
    wire N__3455;
    wire N__3454;
    wire N__3451;
    wire N__3448;
    wire N__3445;
    wire N__3440;
    wire N__3439;
    wire N__3436;
    wire N__3433;
    wire N__3430;
    wire N__3425;
    wire N__3422;
    wire N__3421;
    wire N__3418;
    wire N__3415;
    wire N__3412;
    wire N__3407;
    wire N__3404;
    wire N__3401;
    wire N__3400;
    wire N__3397;
    wire N__3394;
    wire N__3391;
    wire N__3386;
    wire N__3385;
    wire N__3382;
    wire N__3379;
    wire N__3374;
    wire N__3371;
    wire N__3370;
    wire N__3367;
    wire N__3364;
    wire N__3361;
    wire N__3356;
    wire N__3353;
    wire N__3352;
    wire N__3349;
    wire N__3346;
    wire N__3343;
    wire N__3338;
    wire N__3335;
    wire N__3334;
    wire N__3331;
    wire N__3328;
    wire N__3325;
    wire N__3320;
    wire N__3319;
    wire N__3316;
    wire N__3313;
    wire N__3310;
    wire N__3305;
    wire N__3302;
    wire N__3299;
    wire N__3296;
    wire N__3293;
    wire N__3290;
    wire N__3289;
    wire N__3286;
    wire N__3283;
    wire N__3278;
    wire N__3277;
    wire N__3274;
    wire N__3271;
    wire N__3266;
    wire N__3265;
    wire N__3262;
    wire N__3259;
    wire N__3256;
    wire N__3251;
    wire N__3248;
    wire N__3247;
    wire N__3244;
    wire N__3241;
    wire N__3236;
    wire N__3233;
    wire N__3230;
    wire N__3227;
    wire N__3224;
    wire N__3221;
    wire N__3218;
    wire N__3217;
    wire N__3216;
    wire N__3215;
    wire N__3212;
    wire N__3209;
    wire N__3206;
    wire N__3203;
    wire N__3194;
    wire N__3193;
    wire N__3190;
    wire N__3187;
    wire N__3184;
    wire N__3179;
    wire N__3178;
    wire N__3175;
    wire N__3172;
    wire N__3167;
    wire N__3164;
    wire N__3161;
    wire N__3160;
    wire N__3157;
    wire N__3154;
    wire N__3149;
    wire N__3148;
    wire N__3145;
    wire N__3142;
    wire N__3137;
    wire N__3134;
    wire N__3133;
    wire N__3130;
    wire N__3127;
    wire N__3124;
    wire N__3119;
    wire N__3118;
    wire N__3115;
    wire N__3112;
    wire N__3107;
    wire N__3106;
    wire N__3103;
    wire N__3100;
    wire N__3097;
    wire N__3096;
    wire N__3095;
    wire N__3094;
    wire N__3091;
    wire N__3088;
    wire N__3085;
    wire N__3082;
    wire N__3079;
    wire N__3074;
    wire N__3065;
    wire N__3064;
    wire N__3061;
    wire N__3058;
    wire N__3053;
    wire N__3052;
    wire N__3049;
    wire N__3046;
    wire N__3041;
    wire N__3040;
    wire N__3037;
    wire N__3034;
    wire N__3031;
    wire N__3026;
    wire N__3025;
    wire N__3022;
    wire N__3019;
    wire N__3014;
    wire N__3011;
    wire N__3008;
    wire N__3005;
    wire N__3002;
    wire N__2999;
    wire N__2998;
    wire N__2995;
    wire N__2992;
    wire N__2987;
    wire N__2986;
    wire N__2983;
    wire N__2980;
    wire N__2975;
    wire N__2974;
    wire N__2971;
    wire N__2968;
    wire N__2965;
    wire N__2960;
    wire N__2959;
    wire N__2956;
    wire N__2953;
    wire N__2948;
    wire N__2947;
    wire N__2944;
    wire N__2941;
    wire N__2936;
    wire N__2935;
    wire N__2932;
    wire N__2929;
    wire N__2924;
    wire N__2921;
    wire N__2920;
    wire N__2917;
    wire N__2914;
    wire N__2909;
    wire N__2908;
    wire N__2905;
    wire N__2902;
    wire N__2897;
    wire N__2896;
    wire N__2893;
    wire N__2890;
    wire N__2885;
    wire N__2882;
    wire N__2879;
    wire N__2878;
    wire N__2875;
    wire N__2872;
    wire N__2869;
    wire N__2864;
    wire N__2861;
    wire N__2858;
    wire N__2855;
    wire N__2852;
    wire N__2849;
    wire N__2846;
    wire N__2843;
    wire N__2840;
    wire N__2837;
    wire N__2834;
    wire N__2831;
    wire N__2828;
    wire N__2825;
    wire N__2822;
    wire N__2819;
    wire N__2816;
    wire N__2813;
    wire N__2810;
    wire N__2807;
    wire N__2804;
    wire N__2801;
    wire N__2798;
    wire N__2795;
    wire N__2792;
    wire N__2789;
    wire N__2786;
    wire N__2783;
    wire N__2780;
    wire N__2777;
    wire N__2774;
    wire N__2771;
    wire N__2768;
    wire N__2765;
    wire N__2762;
    wire N__2759;
    wire N__2756;
    wire N__2753;
    wire N__2750;
    wire N__2747;
    wire N__2744;
    wire N__2741;
    wire N__2738;
    wire N__2735;
    wire N__2732;
    wire N__2729;
    wire N__2726;
    wire N__2723;
    wire N__2720;
    wire N__2717;
    wire N__2714;
    wire N__2711;
    wire N__2708;
    wire N__2705;
    wire N__2702;
    wire N__2699;
    wire N__2696;
    wire N__2693;
    wire N__2690;
    wire N__2687;
    wire N__2684;
    wire N__2681;
    wire N__2678;
    wire N__2675;
    wire N__2672;
    wire CLK_pad_gb_input;
    wire GNDG0;
    wire VCCG0;
    wire bfn_1_18_0_;
    wire \uart.n2132 ;
    wire \uart.n2133 ;
    wire \uart.n2134 ;
    wire \uart.n2135 ;
    wire \uart.n2136 ;
    wire \uart.n2137 ;
    wire \uart.n2138 ;
    wire \uart.n2139 ;
    wire bfn_1_19_0_;
    wire \uart.n2140 ;
    wire \uart.n2141 ;
    wire \uart.n2142 ;
    wire \uart.n2143 ;
    wire \uart.n2144 ;
    wire \uart.n2145 ;
    wire \uart.n2146 ;
    wire \uart.n2147 ;
    wire bfn_1_20_0_;
    wire \uart.n2148 ;
    wire \uart.n2149 ;
    wire \uart.n2150 ;
    wire \uart.n2151 ;
    wire \uart.n2152 ;
    wire \uart.n2153 ;
    wire \uart.n2154 ;
    wire \uart.n2155 ;
    wire bfn_1_21_0_;
    wire \uart.n2156 ;
    wire \uart.n2157 ;
    wire \uart.n2158 ;
    wire \uart.n2159 ;
    wire \uart.n2160 ;
    wire \uart.n2161 ;
    wire \uart.n2162 ;
    wire bfn_1_22_0_;
    wire n2226;
    wire n2227;
    wire n2228;
    wire n2229;
    wire n2230;
    wire n2231;
    wire n2232;
    wire n2233;
    wire bfn_1_23_0_;
    wire n2234;
    wire n2235;
    wire n2236;
    wire n2237;
    wire n2238;
    wire n2239;
    wire n2240;
    wire n2241;
    wire bfn_1_24_0_;
    wire n2242;
    wire n2243;
    wire n2244;
    wire n2245;
    wire n2246;
    wire n2247;
    wire n2248;
    wire n2249;
    wire bfn_1_25_0_;
    wire n2250;
    wire n2251;
    wire n2252;
    wire n2253;
    wire n2254;
    wire n2255;
    wire n2256;
    wire \uart.r_Clock_Count_2 ;
    wire \uart.r_Clock_Count_0 ;
    wire \uart.r_Clock_Count_1 ;
    wire \uart.r_Clock_Count_3 ;
    wire \uart.r_Clock_Count_5 ;
    wire \uart.r_Clock_Count_4 ;
    wire \uart.n2006_cascade_ ;
    wire \uart.r_Clock_Count_6 ;
    wire \uart.r_Clock_Count_10 ;
    wire \uart.r_Clock_Count_22 ;
    wire \uart.r_Clock_Count_26 ;
    wire \uart.r_Clock_Count_13 ;
    wire \uart.r_Clock_Count_12 ;
    wire \uart.r_Clock_Count_29 ;
    wire \uart.n42_cascade_ ;
    wire \uart.r_Clock_Count_7 ;
    wire \uart.n45_cascade_ ;
    wire \uart.n2385 ;
    wire r_SM_Main_2_N_233_1_cascade_;
    wire \uart.n1796 ;
    wire \uart.r_Clock_Count_8 ;
    wire \uart.r_Clock_Count_14 ;
    wire \uart.n34 ;
    wire \uart.r_Clock_Count_30 ;
    wire \uart.r_Clock_Count_28 ;
    wire \uart.r_Clock_Count_24 ;
    wire \uart.r_Clock_Count_23 ;
    wire \uart.n1 ;
    wire \uart.r_Clock_Count_11 ;
    wire \uart.r_Clock_Count_21 ;
    wire \uart.r_Clock_Count_17 ;
    wire \uart.r_Clock_Count_18 ;
    wire \uart.r_Clock_Count_20 ;
    wire \uart.r_Clock_Count_15 ;
    wire \uart.r_Clock_Count_25 ;
    wire \uart.r_Clock_Count_9 ;
    wire \uart.r_Clock_Count_27 ;
    wire \uart.r_Clock_Count_19 ;
    wire \uart.r_Clock_Count_16 ;
    wire \uart.r_Clock_Count_31 ;
    wire \uart.n39 ;
    wire \uart.n40 ;
    wire \uart.n37_cascade_ ;
    wire \uart.n38 ;
    wire \uart.n46 ;
    wire clk_divider_26;
    wire clk_divider_9;
    wire clk_divider_14;
    wire clk_divider_17;
    wire clk_divider_21;
    wire clk_divider_22;
    wire clk_divider_28;
    wire clk_divider_6;
    wire clk_divider_30;
    wire clk_divider_27;
    wire clk_divider_20;
    wire clk_divider_19;
    wire n44_adj_358;
    wire n42_adj_360_cascade_;
    wire n41_adj_361;
    wire clk_divider_4;
    wire clk_divider_0;
    wire clk_divider_3;
    wire clk_divider_31__N_139;
    wire \uart.n3 ;
    wire clk_divider_1;
    wire clk_divider_2;
    wire n6_adj_324;
    wire clk_divider_8;
    wire clk_divider_15;
    wire clk_divider_24;
    wire clk_divider_11;
    wire clk_divider_5;
    wire clk_divider_10;
    wire clk_divider_12;
    wire clk_divider_18;
    wire clk_divider_13;
    wire clk_divider_29;
    wire clk_divider_23;
    wire clk_divider_16;
    wire n43_adj_359;
    wire clk_divider_31;
    wire n50;
    wire n10;
    wire n26;
    wire bfn_2_23_0_;
    wire n25;
    wire n2163;
    wire n24;
    wire n2164;
    wire n23;
    wire n2165;
    wire n22;
    wire n2166;
    wire n21;
    wire n2167;
    wire n20;
    wire n2168;
    wire n19;
    wire n2169;
    wire n2170;
    wire n18;
    wire bfn_2_24_0_;
    wire n17;
    wire n2171;
    wire n16;
    wire n2172;
    wire n15;
    wire n2173;
    wire n14;
    wire n2174;
    wire n13;
    wire n2175;
    wire n12;
    wire n2176;
    wire n11;
    wire n2177;
    wire n2178;
    wire n10_adj_317;
    wire bfn_2_25_0_;
    wire n9;
    wire n2179;
    wire n8;
    wire n2180;
    wire n7;
    wire n2181;
    wire n6;
    wire n2182;
    wire n2183;
    wire n2184;
    wire n2185;
    wire n2186;
    wire bfn_2_26_0_;
    wire n2187;
    wire blink_counter_25;
    wire n2395_cascade_;
    wire LED_c;
    wire blink_counter_21;
    wire blink_counter_24;
    wire blink_counter_23;
    wire blink_counter_22;
    wire n2394;
    wire \uart.n1711 ;
    wire \uart.o_Tx_Serial_N_312 ;
    wire clk_divider_7;
    wire n40_adj_362;
    wire clk_divider_25;
    wire n45_adj_357;
    wire n49;
    wire counter_0;
    wire bfn_3_22_0_;
    wire counter_1;
    wire n2195;
    wire counter_2;
    wire n2196;
    wire counter_3;
    wire n2197;
    wire counter_4;
    wire n2198;
    wire counter_5;
    wire n2199;
    wire counter_6;
    wire n2200;
    wire counter_7;
    wire n2201;
    wire n2202;
    wire bfn_3_23_0_;
    wire n2203;
    wire n2204;
    wire n2205;
    wire n2206;
    wire n2207;
    wire n2208;
    wire n2209;
    wire n2210;
    wire bfn_3_24_0_;
    wire n2211;
    wire n2212;
    wire n2213;
    wire n2214;
    wire n2215;
    wire n2216;
    wire n2217;
    wire n2218;
    wire bfn_3_25_0_;
    wire n2219;
    wire n2220;
    wire n2221;
    wire n2222;
    wire n2223;
    wire n2224;
    wire n2225;
    wire \uart.r_Bit_Index_2 ;
    wire n2002_cascade_;
    wire r_SM_Main_2_N_233_1;
    wire n2308_cascade_;
    wire n2002;
    wire \uart.n2428_cascade_ ;
    wire \uart.n2431 ;
    wire r_Tx_Data_4;
    wire r_Tx_Data_5;
    wire \uart.n2422_cascade_ ;
    wire \uart.n2425 ;
    wire r_Tx_Data_6;
    wire r_SM_Main_1;
    wire r_SM_Main_0;
    wire r_SM_Main_2;
    wire r_Tx_Data_1;
    wire r_Tx_Data_3;
    wire r_Tx_Data_7;
    wire r_Tx_Data_0;
    wire n1757;
    wire r_Tx_Data_2;
    wire data_out_5;
    wire data_out_0;
    wire data_out_3;
    wire data_out_1;
    wire data_out_2;
    wire counter_13;
    wire counter_23;
    wire counter_11;
    wire counter_14;
    wire n38_cascade_;
    wire n44_cascade_;
    wire counter_31__N_172_cascade_;
    wire data_out_4;
    wire counter_31;
    wire n44;
    wire r_SM_Main_2_N_236_0;
    wire data_out_6;
    wire counter_22;
    wire counter_30;
    wire counter_19;
    wire counter_26;
    wire n36;
    wire counter_12;
    wire counter_8;
    wire counter_15;
    wire counter_25;
    wire n40;
    wire counter_17;
    wire counter_24;
    wire counter_21;
    wire counter_16;
    wire n39;
    wire counter_20;
    wire counter_10;
    wire counter_29;
    wire counter_28;
    wire n37;
    wire counter_18;
    wire counter_27;
    wire counter_9;
    wire n35;
    wire data_out_7;
    wire r_Bit_Index_0;
    wire \uart.r_Bit_Index_1 ;
    wire CLK_c;
    wire n2308;
    wire \uart.n2310 ;
    wire diff_input;
    wire integrator_0;
    wire bfn_5_23_0_;
    wire integrator_1;
    wire n2188;
    wire integrator_2;
    wire n2189;
    wire integrator_3;
    wire n2190;
    wire integrator_4;
    wire n2191;
    wire integrator_5;
    wire n2192;
    wire integrator_6;
    wire n2193;
    wire n2194;
    wire integrator_7;
    wire _gnd_net_;
    wire clk_slow;
    wire counter_31__N_172;

    defparam LED_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam LED_pad_iopad.PULLUP=1'b0;
    IO_PAD LED_pad_iopad (
            .OE(N__5970),
            .DIN(N__5969),
            .DOUT(N__5968),
            .PACKAGEPIN(LED));
    defparam LED_pad_preio.PIN_TYPE=6'b011001;
    defparam LED_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO LED_pad_preio (
            .PADOEN(N__5970),
            .PADOUT(N__5969),
            .PADIN(N__5968),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__4358),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    defparam PIN_18_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam PIN_18_pad_iopad.PULLUP=1'b0;
    IO_PAD PIN_18_pad_iopad (
            .OE(N__5961),
            .DIN(N__5960),
            .DOUT(N__5959),
            .PACKAGEPIN(PIN_18));
    defparam PIN_18_pad_preio.PIN_TYPE=6'b010101;
    defparam PIN_18_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO PIN_18_pad_preio (
            .PADOEN(N__5961),
            .PADOUT(N__5960),
            .PADIN(N__5959),
            .CLOCKENABLE(VCCG0),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__5276),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(N__5825),
            .OUTPUTENABLE());
    defparam PIN_2_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam PIN_2_pad_iopad.PULLUP=1'b0;
    IO_PAD PIN_2_pad_iopad (
            .OE(N__5952),
            .DIN(N__5951),
            .DOUT(N__5950),
            .PACKAGEPIN(PIN_2));
    defparam PIN_2_pad_preio.PIN_TYPE=6'b010101;
    defparam PIN_2_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO PIN_2_pad_preio (
            .PADOEN(N__5952),
            .PADOUT(N__5951),
            .PADIN(N__5950),
            .CLOCKENABLE(N__3107),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__3911),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(N__5399),
            .OUTPUTENABLE());
    defparam differential_input_iopad.IO_STANDARD="SB_LVDS_INPUT";
    defparam differential_input_iopad.PULLUP=1'b0;
    IO_PAD differential_input_iopad (
            .OE(N__5943),
            .DIN(N__5942),
            .DOUT(N__5941),
            .PACKAGEPIN(PIN_13));
    defparam differential_input_preio.PIN_TYPE=6'b000001;
    defparam differential_input_preio.NEG_TRIGGER=1'b0;
    PRE_IO differential_input_preio (
            .PADOEN(N__5943),
            .PADOUT(N__5942),
            .PADIN(N__5941),
            .CLOCKENABLE(),
            .DIN0(diff_input),
            .DIN1(),
            .DOUT0(GNDG0),
            .DOUT1(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    defparam CLK_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam CLK_pad_iopad.PULLUP=1'b0;
    IO_PAD CLK_pad_iopad (
            .OE(N__5934),
            .DIN(N__5933),
            .DOUT(N__5932),
            .PACKAGEPIN(CLK));
    defparam CLK_pad_preio.PIN_TYPE=6'b000001;
    defparam CLK_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO CLK_pad_preio (
            .PADOEN(N__5934),
            .PADOUT(N__5933),
            .PADIN(N__5932),
            .CLOCKENABLE(),
            .DIN0(CLK_pad_gb_input),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    InMux I__1307 (
            .O(N__5915),
            .I(N__5911));
    InMux I__1306 (
            .O(N__5914),
            .I(N__5908));
    LocalMux I__1305 (
            .O(N__5911),
            .I(integrator_2));
    LocalMux I__1304 (
            .O(N__5908),
            .I(integrator_2));
    InMux I__1303 (
            .O(N__5903),
            .I(n2189));
    InMux I__1302 (
            .O(N__5900),
            .I(N__5896));
    InMux I__1301 (
            .O(N__5899),
            .I(N__5893));
    LocalMux I__1300 (
            .O(N__5896),
            .I(integrator_3));
    LocalMux I__1299 (
            .O(N__5893),
            .I(integrator_3));
    InMux I__1298 (
            .O(N__5888),
            .I(n2190));
    InMux I__1297 (
            .O(N__5885),
            .I(N__5881));
    InMux I__1296 (
            .O(N__5884),
            .I(N__5878));
    LocalMux I__1295 (
            .O(N__5881),
            .I(integrator_4));
    LocalMux I__1294 (
            .O(N__5878),
            .I(integrator_4));
    InMux I__1293 (
            .O(N__5873),
            .I(n2191));
    InMux I__1292 (
            .O(N__5870),
            .I(N__5866));
    InMux I__1291 (
            .O(N__5869),
            .I(N__5863));
    LocalMux I__1290 (
            .O(N__5866),
            .I(integrator_5));
    LocalMux I__1289 (
            .O(N__5863),
            .I(integrator_5));
    InMux I__1288 (
            .O(N__5858),
            .I(n2192));
    InMux I__1287 (
            .O(N__5855),
            .I(N__5851));
    InMux I__1286 (
            .O(N__5854),
            .I(N__5848));
    LocalMux I__1285 (
            .O(N__5851),
            .I(integrator_6));
    LocalMux I__1284 (
            .O(N__5848),
            .I(integrator_6));
    InMux I__1283 (
            .O(N__5843),
            .I(n2193));
    InMux I__1282 (
            .O(N__5840),
            .I(n2194));
    InMux I__1281 (
            .O(N__5837),
            .I(N__5833));
    InMux I__1280 (
            .O(N__5836),
            .I(N__5830));
    LocalMux I__1279 (
            .O(N__5833),
            .I(integrator_7));
    LocalMux I__1278 (
            .O(N__5830),
            .I(integrator_7));
    ClkMux I__1277 (
            .O(N__5825),
            .I(N__5822));
    LocalMux I__1276 (
            .O(N__5822),
            .I(N__5819));
    Span4Mux_s2_h I__1275 (
            .O(N__5819),
            .I(N__5816));
    Span4Mux_h I__1274 (
            .O(N__5816),
            .I(N__5809));
    ClkMux I__1273 (
            .O(N__5815),
            .I(N__5806));
    ClkMux I__1272 (
            .O(N__5814),
            .I(N__5801));
    ClkMux I__1271 (
            .O(N__5813),
            .I(N__5798));
    ClkMux I__1270 (
            .O(N__5812),
            .I(N__5795));
    Sp12to4 I__1269 (
            .O(N__5809),
            .I(N__5792));
    LocalMux I__1268 (
            .O(N__5806),
            .I(N__5789));
    ClkMux I__1267 (
            .O(N__5805),
            .I(N__5786));
    ClkMux I__1266 (
            .O(N__5804),
            .I(N__5783));
    LocalMux I__1265 (
            .O(N__5801),
            .I(N__5780));
    LocalMux I__1264 (
            .O(N__5798),
            .I(N__5775));
    LocalMux I__1263 (
            .O(N__5795),
            .I(N__5775));
    Span12Mux_v I__1262 (
            .O(N__5792),
            .I(N__5771));
    Span4Mux_v I__1261 (
            .O(N__5789),
            .I(N__5766));
    LocalMux I__1260 (
            .O(N__5786),
            .I(N__5766));
    LocalMux I__1259 (
            .O(N__5783),
            .I(N__5763));
    Span4Mux_v I__1258 (
            .O(N__5780),
            .I(N__5758));
    Span4Mux_v I__1257 (
            .O(N__5775),
            .I(N__5758));
    ClkMux I__1256 (
            .O(N__5774),
            .I(N__5755));
    Span12Mux_h I__1255 (
            .O(N__5771),
            .I(N__5751));
    Span4Mux_h I__1254 (
            .O(N__5766),
            .I(N__5748));
    Span4Mux_v I__1253 (
            .O(N__5763),
            .I(N__5745));
    Span4Mux_s2_h I__1252 (
            .O(N__5758),
            .I(N__5740));
    LocalMux I__1251 (
            .O(N__5755),
            .I(N__5740));
    ClkMux I__1250 (
            .O(N__5754),
            .I(N__5737));
    Span12Mux_h I__1249 (
            .O(N__5751),
            .I(N__5734));
    Span4Mux_v I__1248 (
            .O(N__5748),
            .I(N__5731));
    Sp12to4 I__1247 (
            .O(N__5745),
            .I(N__5724));
    Sp12to4 I__1246 (
            .O(N__5740),
            .I(N__5724));
    LocalMux I__1245 (
            .O(N__5737),
            .I(N__5724));
    Odrv12 I__1244 (
            .O(N__5734),
            .I(clk_slow));
    Odrv4 I__1243 (
            .O(N__5731),
            .I(clk_slow));
    Odrv12 I__1242 (
            .O(N__5724),
            .I(clk_slow));
    SRMux I__1241 (
            .O(N__5717),
            .I(N__5714));
    LocalMux I__1240 (
            .O(N__5714),
            .I(N__5711));
    Span4Mux_s3_h I__1239 (
            .O(N__5711),
            .I(N__5697));
    SRMux I__1238 (
            .O(N__5710),
            .I(N__5694));
    SRMux I__1237 (
            .O(N__5709),
            .I(N__5691));
    SRMux I__1236 (
            .O(N__5708),
            .I(N__5688));
    SRMux I__1235 (
            .O(N__5707),
            .I(N__5685));
    InMux I__1234 (
            .O(N__5706),
            .I(N__5682));
    InMux I__1233 (
            .O(N__5705),
            .I(N__5675));
    InMux I__1232 (
            .O(N__5704),
            .I(N__5675));
    InMux I__1231 (
            .O(N__5703),
            .I(N__5675));
    InMux I__1230 (
            .O(N__5702),
            .I(N__5668));
    InMux I__1229 (
            .O(N__5701),
            .I(N__5668));
    InMux I__1228 (
            .O(N__5700),
            .I(N__5668));
    Odrv4 I__1227 (
            .O(N__5697),
            .I(counter_31__N_172));
    LocalMux I__1226 (
            .O(N__5694),
            .I(counter_31__N_172));
    LocalMux I__1225 (
            .O(N__5691),
            .I(counter_31__N_172));
    LocalMux I__1224 (
            .O(N__5688),
            .I(counter_31__N_172));
    LocalMux I__1223 (
            .O(N__5685),
            .I(counter_31__N_172));
    LocalMux I__1222 (
            .O(N__5682),
            .I(counter_31__N_172));
    LocalMux I__1221 (
            .O(N__5675),
            .I(counter_31__N_172));
    LocalMux I__1220 (
            .O(N__5668),
            .I(counter_31__N_172));
    InMux I__1219 (
            .O(N__5651),
            .I(N__5647));
    InMux I__1218 (
            .O(N__5650),
            .I(N__5644));
    LocalMux I__1217 (
            .O(N__5647),
            .I(counter_17));
    LocalMux I__1216 (
            .O(N__5644),
            .I(counter_17));
    InMux I__1215 (
            .O(N__5639),
            .I(N__5635));
    InMux I__1214 (
            .O(N__5638),
            .I(N__5632));
    LocalMux I__1213 (
            .O(N__5635),
            .I(counter_24));
    LocalMux I__1212 (
            .O(N__5632),
            .I(counter_24));
    CascadeMux I__1211 (
            .O(N__5627),
            .I(N__5623));
    InMux I__1210 (
            .O(N__5626),
            .I(N__5620));
    InMux I__1209 (
            .O(N__5623),
            .I(N__5617));
    LocalMux I__1208 (
            .O(N__5620),
            .I(counter_21));
    LocalMux I__1207 (
            .O(N__5617),
            .I(counter_21));
    InMux I__1206 (
            .O(N__5612),
            .I(N__5608));
    InMux I__1205 (
            .O(N__5611),
            .I(N__5605));
    LocalMux I__1204 (
            .O(N__5608),
            .I(counter_16));
    LocalMux I__1203 (
            .O(N__5605),
            .I(counter_16));
    InMux I__1202 (
            .O(N__5600),
            .I(N__5594));
    InMux I__1201 (
            .O(N__5599),
            .I(N__5594));
    LocalMux I__1200 (
            .O(N__5594),
            .I(n39));
    InMux I__1199 (
            .O(N__5591),
            .I(N__5587));
    InMux I__1198 (
            .O(N__5590),
            .I(N__5584));
    LocalMux I__1197 (
            .O(N__5587),
            .I(counter_20));
    LocalMux I__1196 (
            .O(N__5584),
            .I(counter_20));
    InMux I__1195 (
            .O(N__5579),
            .I(N__5575));
    InMux I__1194 (
            .O(N__5578),
            .I(N__5572));
    LocalMux I__1193 (
            .O(N__5575),
            .I(counter_10));
    LocalMux I__1192 (
            .O(N__5572),
            .I(counter_10));
    CascadeMux I__1191 (
            .O(N__5567),
            .I(N__5563));
    InMux I__1190 (
            .O(N__5566),
            .I(N__5560));
    InMux I__1189 (
            .O(N__5563),
            .I(N__5557));
    LocalMux I__1188 (
            .O(N__5560),
            .I(counter_29));
    LocalMux I__1187 (
            .O(N__5557),
            .I(counter_29));
    InMux I__1186 (
            .O(N__5552),
            .I(N__5548));
    InMux I__1185 (
            .O(N__5551),
            .I(N__5545));
    LocalMux I__1184 (
            .O(N__5548),
            .I(counter_28));
    LocalMux I__1183 (
            .O(N__5545),
            .I(counter_28));
    InMux I__1182 (
            .O(N__5540),
            .I(N__5537));
    LocalMux I__1181 (
            .O(N__5537),
            .I(n37));
    InMux I__1180 (
            .O(N__5534),
            .I(N__5530));
    InMux I__1179 (
            .O(N__5533),
            .I(N__5527));
    LocalMux I__1178 (
            .O(N__5530),
            .I(counter_18));
    LocalMux I__1177 (
            .O(N__5527),
            .I(counter_18));
    InMux I__1176 (
            .O(N__5522),
            .I(N__5518));
    InMux I__1175 (
            .O(N__5521),
            .I(N__5515));
    LocalMux I__1174 (
            .O(N__5518),
            .I(counter_27));
    LocalMux I__1173 (
            .O(N__5515),
            .I(counter_27));
    InMux I__1172 (
            .O(N__5510),
            .I(N__5506));
    InMux I__1171 (
            .O(N__5509),
            .I(N__5503));
    LocalMux I__1170 (
            .O(N__5506),
            .I(counter_9));
    LocalMux I__1169 (
            .O(N__5503),
            .I(counter_9));
    InMux I__1168 (
            .O(N__5498),
            .I(N__5495));
    LocalMux I__1167 (
            .O(N__5495),
            .I(n35));
    InMux I__1166 (
            .O(N__5492),
            .I(N__5489));
    LocalMux I__1165 (
            .O(N__5489),
            .I(N__5485));
    InMux I__1164 (
            .O(N__5488),
            .I(N__5482));
    Odrv12 I__1163 (
            .O(N__5485),
            .I(data_out_7));
    LocalMux I__1162 (
            .O(N__5482),
            .I(data_out_7));
    InMux I__1161 (
            .O(N__5477),
            .I(N__5469));
    InMux I__1160 (
            .O(N__5476),
            .I(N__5466));
    InMux I__1159 (
            .O(N__5475),
            .I(N__5461));
    InMux I__1158 (
            .O(N__5474),
            .I(N__5461));
    InMux I__1157 (
            .O(N__5473),
            .I(N__5456));
    InMux I__1156 (
            .O(N__5472),
            .I(N__5456));
    LocalMux I__1155 (
            .O(N__5469),
            .I(r_Bit_Index_0));
    LocalMux I__1154 (
            .O(N__5466),
            .I(r_Bit_Index_0));
    LocalMux I__1153 (
            .O(N__5461),
            .I(r_Bit_Index_0));
    LocalMux I__1152 (
            .O(N__5456),
            .I(r_Bit_Index_0));
    InMux I__1151 (
            .O(N__5447),
            .I(N__5444));
    LocalMux I__1150 (
            .O(N__5444),
            .I(N__5439));
    CascadeMux I__1149 (
            .O(N__5443),
            .I(N__5433));
    CascadeMux I__1148 (
            .O(N__5442),
            .I(N__5429));
    Span4Mux_h I__1147 (
            .O(N__5439),
            .I(N__5426));
    InMux I__1146 (
            .O(N__5438),
            .I(N__5423));
    InMux I__1145 (
            .O(N__5437),
            .I(N__5420));
    InMux I__1144 (
            .O(N__5436),
            .I(N__5415));
    InMux I__1143 (
            .O(N__5433),
            .I(N__5415));
    InMux I__1142 (
            .O(N__5432),
            .I(N__5410));
    InMux I__1141 (
            .O(N__5429),
            .I(N__5410));
    Odrv4 I__1140 (
            .O(N__5426),
            .I(\uart.r_Bit_Index_1 ));
    LocalMux I__1139 (
            .O(N__5423),
            .I(\uart.r_Bit_Index_1 ));
    LocalMux I__1138 (
            .O(N__5420),
            .I(\uart.r_Bit_Index_1 ));
    LocalMux I__1137 (
            .O(N__5415),
            .I(\uart.r_Bit_Index_1 ));
    LocalMux I__1136 (
            .O(N__5410),
            .I(\uart.r_Bit_Index_1 ));
    ClkMux I__1135 (
            .O(N__5399),
            .I(N__5336));
    ClkMux I__1134 (
            .O(N__5398),
            .I(N__5336));
    ClkMux I__1133 (
            .O(N__5397),
            .I(N__5336));
    ClkMux I__1132 (
            .O(N__5396),
            .I(N__5336));
    ClkMux I__1131 (
            .O(N__5395),
            .I(N__5336));
    ClkMux I__1130 (
            .O(N__5394),
            .I(N__5336));
    ClkMux I__1129 (
            .O(N__5393),
            .I(N__5336));
    ClkMux I__1128 (
            .O(N__5392),
            .I(N__5336));
    ClkMux I__1127 (
            .O(N__5391),
            .I(N__5336));
    ClkMux I__1126 (
            .O(N__5390),
            .I(N__5336));
    ClkMux I__1125 (
            .O(N__5389),
            .I(N__5336));
    ClkMux I__1124 (
            .O(N__5388),
            .I(N__5336));
    ClkMux I__1123 (
            .O(N__5387),
            .I(N__5336));
    ClkMux I__1122 (
            .O(N__5386),
            .I(N__5336));
    ClkMux I__1121 (
            .O(N__5385),
            .I(N__5336));
    ClkMux I__1120 (
            .O(N__5384),
            .I(N__5336));
    ClkMux I__1119 (
            .O(N__5383),
            .I(N__5336));
    ClkMux I__1118 (
            .O(N__5382),
            .I(N__5336));
    ClkMux I__1117 (
            .O(N__5381),
            .I(N__5336));
    ClkMux I__1116 (
            .O(N__5380),
            .I(N__5336));
    ClkMux I__1115 (
            .O(N__5379),
            .I(N__5336));
    GlobalMux I__1114 (
            .O(N__5336),
            .I(N__5333));
    gio2CtrlBuf I__1113 (
            .O(N__5333),
            .I(CLK_c));
    CEMux I__1112 (
            .O(N__5330),
            .I(N__5326));
    CEMux I__1111 (
            .O(N__5329),
            .I(N__5323));
    LocalMux I__1110 (
            .O(N__5326),
            .I(N__5320));
    LocalMux I__1109 (
            .O(N__5323),
            .I(N__5316));
    Span4Mux_v I__1108 (
            .O(N__5320),
            .I(N__5313));
    InMux I__1107 (
            .O(N__5319),
            .I(N__5310));
    Odrv4 I__1106 (
            .O(N__5316),
            .I(n2308));
    Odrv4 I__1105 (
            .O(N__5313),
            .I(n2308));
    LocalMux I__1104 (
            .O(N__5310),
            .I(n2308));
    SRMux I__1103 (
            .O(N__5303),
            .I(N__5299));
    SRMux I__1102 (
            .O(N__5302),
            .I(N__5296));
    LocalMux I__1101 (
            .O(N__5299),
            .I(N__5293));
    LocalMux I__1100 (
            .O(N__5296),
            .I(N__5290));
    Span4Mux_h I__1099 (
            .O(N__5293),
            .I(N__5287));
    Span4Mux_s3_h I__1098 (
            .O(N__5290),
            .I(N__5284));
    Span4Mux_s1_h I__1097 (
            .O(N__5287),
            .I(N__5281));
    Odrv4 I__1096 (
            .O(N__5284),
            .I(\uart.n2310 ));
    Odrv4 I__1095 (
            .O(N__5281),
            .I(\uart.n2310 ));
    IoInMux I__1094 (
            .O(N__5276),
            .I(N__5272));
    CascadeMux I__1093 (
            .O(N__5275),
            .I(N__5269));
    LocalMux I__1092 (
            .O(N__5272),
            .I(N__5266));
    InMux I__1091 (
            .O(N__5269),
            .I(N__5263));
    IoSpan4Mux I__1090 (
            .O(N__5266),
            .I(N__5260));
    LocalMux I__1089 (
            .O(N__5263),
            .I(N__5257));
    Span4Mux_s2_v I__1088 (
            .O(N__5260),
            .I(N__5254));
    Span4Mux_h I__1087 (
            .O(N__5257),
            .I(N__5251));
    Sp12to4 I__1086 (
            .O(N__5254),
            .I(N__5248));
    Sp12to4 I__1085 (
            .O(N__5251),
            .I(N__5245));
    Span12Mux_h I__1084 (
            .O(N__5248),
            .I(N__5242));
    Span12Mux_v I__1083 (
            .O(N__5245),
            .I(N__5239));
    Span12Mux_h I__1082 (
            .O(N__5242),
            .I(N__5234));
    Span12Mux_v I__1081 (
            .O(N__5239),
            .I(N__5234));
    Odrv12 I__1080 (
            .O(N__5234),
            .I(diff_input));
    InMux I__1079 (
            .O(N__5231),
            .I(N__5227));
    InMux I__1078 (
            .O(N__5230),
            .I(N__5224));
    LocalMux I__1077 (
            .O(N__5227),
            .I(integrator_0));
    LocalMux I__1076 (
            .O(N__5224),
            .I(integrator_0));
    InMux I__1075 (
            .O(N__5219),
            .I(N__5215));
    InMux I__1074 (
            .O(N__5218),
            .I(N__5212));
    LocalMux I__1073 (
            .O(N__5215),
            .I(integrator_1));
    LocalMux I__1072 (
            .O(N__5212),
            .I(integrator_1));
    InMux I__1071 (
            .O(N__5207),
            .I(n2188));
    InMux I__1070 (
            .O(N__5204),
            .I(N__5200));
    InMux I__1069 (
            .O(N__5203),
            .I(N__5197));
    LocalMux I__1068 (
            .O(N__5200),
            .I(N__5194));
    LocalMux I__1067 (
            .O(N__5197),
            .I(counter_13));
    Odrv4 I__1066 (
            .O(N__5194),
            .I(counter_13));
    InMux I__1065 (
            .O(N__5189),
            .I(N__5185));
    InMux I__1064 (
            .O(N__5188),
            .I(N__5182));
    LocalMux I__1063 (
            .O(N__5185),
            .I(counter_23));
    LocalMux I__1062 (
            .O(N__5182),
            .I(counter_23));
    CascadeMux I__1061 (
            .O(N__5177),
            .I(N__5173));
    InMux I__1060 (
            .O(N__5176),
            .I(N__5170));
    InMux I__1059 (
            .O(N__5173),
            .I(N__5167));
    LocalMux I__1058 (
            .O(N__5170),
            .I(counter_11));
    LocalMux I__1057 (
            .O(N__5167),
            .I(counter_11));
    InMux I__1056 (
            .O(N__5162),
            .I(N__5158));
    InMux I__1055 (
            .O(N__5161),
            .I(N__5155));
    LocalMux I__1054 (
            .O(N__5158),
            .I(counter_14));
    LocalMux I__1053 (
            .O(N__5155),
            .I(counter_14));
    CascadeMux I__1052 (
            .O(N__5150),
            .I(n38_cascade_));
    CascadeMux I__1051 (
            .O(N__5147),
            .I(n44_cascade_));
    CascadeMux I__1050 (
            .O(N__5144),
            .I(counter_31__N_172_cascade_));
    InMux I__1049 (
            .O(N__5141),
            .I(N__5138));
    LocalMux I__1048 (
            .O(N__5138),
            .I(N__5134));
    InMux I__1047 (
            .O(N__5137),
            .I(N__5131));
    Odrv12 I__1046 (
            .O(N__5134),
            .I(data_out_4));
    LocalMux I__1045 (
            .O(N__5131),
            .I(data_out_4));
    InMux I__1044 (
            .O(N__5126),
            .I(N__5120));
    InMux I__1043 (
            .O(N__5125),
            .I(N__5120));
    LocalMux I__1042 (
            .O(N__5120),
            .I(N__5116));
    InMux I__1041 (
            .O(N__5119),
            .I(N__5113));
    Span4Mux_h I__1040 (
            .O(N__5116),
            .I(N__5110));
    LocalMux I__1039 (
            .O(N__5113),
            .I(counter_31));
    Odrv4 I__1038 (
            .O(N__5110),
            .I(counter_31));
    InMux I__1037 (
            .O(N__5105),
            .I(N__5102));
    LocalMux I__1036 (
            .O(N__5102),
            .I(n44));
    CascadeMux I__1035 (
            .O(N__5099),
            .I(N__5096));
    InMux I__1034 (
            .O(N__5096),
            .I(N__5093));
    LocalMux I__1033 (
            .O(N__5093),
            .I(N__5089));
    CascadeMux I__1032 (
            .O(N__5092),
            .I(N__5086));
    Span4Mux_s3_h I__1031 (
            .O(N__5089),
            .I(N__5083));
    InMux I__1030 (
            .O(N__5086),
            .I(N__5080));
    Sp12to4 I__1029 (
            .O(N__5083),
            .I(N__5075));
    LocalMux I__1028 (
            .O(N__5080),
            .I(N__5075));
    Odrv12 I__1027 (
            .O(N__5075),
            .I(r_SM_Main_2_N_236_0));
    InMux I__1026 (
            .O(N__5072),
            .I(N__5069));
    LocalMux I__1025 (
            .O(N__5069),
            .I(N__5065));
    InMux I__1024 (
            .O(N__5068),
            .I(N__5062));
    Odrv12 I__1023 (
            .O(N__5065),
            .I(data_out_6));
    LocalMux I__1022 (
            .O(N__5062),
            .I(data_out_6));
    InMux I__1021 (
            .O(N__5057),
            .I(N__5053));
    InMux I__1020 (
            .O(N__5056),
            .I(N__5050));
    LocalMux I__1019 (
            .O(N__5053),
            .I(counter_22));
    LocalMux I__1018 (
            .O(N__5050),
            .I(counter_22));
    InMux I__1017 (
            .O(N__5045),
            .I(N__5041));
    InMux I__1016 (
            .O(N__5044),
            .I(N__5038));
    LocalMux I__1015 (
            .O(N__5041),
            .I(counter_30));
    LocalMux I__1014 (
            .O(N__5038),
            .I(counter_30));
    CascadeMux I__1013 (
            .O(N__5033),
            .I(N__5029));
    InMux I__1012 (
            .O(N__5032),
            .I(N__5026));
    InMux I__1011 (
            .O(N__5029),
            .I(N__5023));
    LocalMux I__1010 (
            .O(N__5026),
            .I(counter_19));
    LocalMux I__1009 (
            .O(N__5023),
            .I(counter_19));
    InMux I__1008 (
            .O(N__5018),
            .I(N__5014));
    InMux I__1007 (
            .O(N__5017),
            .I(N__5011));
    LocalMux I__1006 (
            .O(N__5014),
            .I(counter_26));
    LocalMux I__1005 (
            .O(N__5011),
            .I(counter_26));
    InMux I__1004 (
            .O(N__5006),
            .I(N__5003));
    LocalMux I__1003 (
            .O(N__5003),
            .I(n36));
    InMux I__1002 (
            .O(N__5000),
            .I(N__4996));
    InMux I__1001 (
            .O(N__4999),
            .I(N__4993));
    LocalMux I__1000 (
            .O(N__4996),
            .I(counter_12));
    LocalMux I__999 (
            .O(N__4993),
            .I(counter_12));
    InMux I__998 (
            .O(N__4988),
            .I(N__4984));
    InMux I__997 (
            .O(N__4987),
            .I(N__4981));
    LocalMux I__996 (
            .O(N__4984),
            .I(counter_8));
    LocalMux I__995 (
            .O(N__4981),
            .I(counter_8));
    CascadeMux I__994 (
            .O(N__4976),
            .I(N__4972));
    InMux I__993 (
            .O(N__4975),
            .I(N__4969));
    InMux I__992 (
            .O(N__4972),
            .I(N__4966));
    LocalMux I__991 (
            .O(N__4969),
            .I(counter_15));
    LocalMux I__990 (
            .O(N__4966),
            .I(counter_15));
    InMux I__989 (
            .O(N__4961),
            .I(N__4957));
    InMux I__988 (
            .O(N__4960),
            .I(N__4954));
    LocalMux I__987 (
            .O(N__4957),
            .I(counter_25));
    LocalMux I__986 (
            .O(N__4954),
            .I(counter_25));
    CascadeMux I__985 (
            .O(N__4949),
            .I(N__4946));
    InMux I__984 (
            .O(N__4946),
            .I(N__4942));
    InMux I__983 (
            .O(N__4945),
            .I(N__4939));
    LocalMux I__982 (
            .O(N__4942),
            .I(N__4934));
    LocalMux I__981 (
            .O(N__4939),
            .I(N__4934));
    Odrv4 I__980 (
            .O(N__4934),
            .I(n40));
    InMux I__979 (
            .O(N__4931),
            .I(N__4927));
    InMux I__978 (
            .O(N__4930),
            .I(N__4924));
    LocalMux I__977 (
            .O(N__4927),
            .I(r_Tx_Data_3));
    LocalMux I__976 (
            .O(N__4924),
            .I(r_Tx_Data_3));
    InMux I__975 (
            .O(N__4919),
            .I(N__4915));
    InMux I__974 (
            .O(N__4918),
            .I(N__4912));
    LocalMux I__973 (
            .O(N__4915),
            .I(r_Tx_Data_7));
    LocalMux I__972 (
            .O(N__4912),
            .I(r_Tx_Data_7));
    InMux I__971 (
            .O(N__4907),
            .I(N__4903));
    InMux I__970 (
            .O(N__4906),
            .I(N__4900));
    LocalMux I__969 (
            .O(N__4903),
            .I(r_Tx_Data_0));
    LocalMux I__968 (
            .O(N__4900),
            .I(r_Tx_Data_0));
    InMux I__967 (
            .O(N__4895),
            .I(N__4877));
    InMux I__966 (
            .O(N__4894),
            .I(N__4877));
    InMux I__965 (
            .O(N__4893),
            .I(N__4877));
    InMux I__964 (
            .O(N__4892),
            .I(N__4877));
    InMux I__963 (
            .O(N__4891),
            .I(N__4877));
    InMux I__962 (
            .O(N__4890),
            .I(N__4870));
    InMux I__961 (
            .O(N__4889),
            .I(N__4870));
    InMux I__960 (
            .O(N__4888),
            .I(N__4870));
    LocalMux I__959 (
            .O(N__4877),
            .I(n1757));
    LocalMux I__958 (
            .O(N__4870),
            .I(n1757));
    InMux I__957 (
            .O(N__4865),
            .I(N__4861));
    InMux I__956 (
            .O(N__4864),
            .I(N__4858));
    LocalMux I__955 (
            .O(N__4861),
            .I(r_Tx_Data_2));
    LocalMux I__954 (
            .O(N__4858),
            .I(r_Tx_Data_2));
    InMux I__953 (
            .O(N__4853),
            .I(N__4850));
    LocalMux I__952 (
            .O(N__4850),
            .I(N__4846));
    InMux I__951 (
            .O(N__4849),
            .I(N__4843));
    Odrv12 I__950 (
            .O(N__4846),
            .I(data_out_5));
    LocalMux I__949 (
            .O(N__4843),
            .I(data_out_5));
    InMux I__948 (
            .O(N__4838),
            .I(N__4835));
    LocalMux I__947 (
            .O(N__4835),
            .I(N__4831));
    InMux I__946 (
            .O(N__4834),
            .I(N__4828));
    Odrv4 I__945 (
            .O(N__4831),
            .I(data_out_0));
    LocalMux I__944 (
            .O(N__4828),
            .I(data_out_0));
    InMux I__943 (
            .O(N__4823),
            .I(N__4819));
    InMux I__942 (
            .O(N__4822),
            .I(N__4816));
    LocalMux I__941 (
            .O(N__4819),
            .I(data_out_3));
    LocalMux I__940 (
            .O(N__4816),
            .I(data_out_3));
    InMux I__939 (
            .O(N__4811),
            .I(N__4808));
    LocalMux I__938 (
            .O(N__4808),
            .I(N__4804));
    InMux I__937 (
            .O(N__4807),
            .I(N__4801));
    Odrv4 I__936 (
            .O(N__4804),
            .I(data_out_1));
    LocalMux I__935 (
            .O(N__4801),
            .I(data_out_1));
    InMux I__934 (
            .O(N__4796),
            .I(N__4793));
    LocalMux I__933 (
            .O(N__4793),
            .I(N__4789));
    InMux I__932 (
            .O(N__4792),
            .I(N__4786));
    Odrv12 I__931 (
            .O(N__4789),
            .I(data_out_2));
    LocalMux I__930 (
            .O(N__4786),
            .I(data_out_2));
    CascadeMux I__929 (
            .O(N__4781),
            .I(\uart.n2428_cascade_ ));
    InMux I__928 (
            .O(N__4778),
            .I(N__4775));
    LocalMux I__927 (
            .O(N__4775),
            .I(\uart.n2431 ));
    InMux I__926 (
            .O(N__4772),
            .I(N__4766));
    InMux I__925 (
            .O(N__4771),
            .I(N__4766));
    LocalMux I__924 (
            .O(N__4766),
            .I(r_Tx_Data_4));
    InMux I__923 (
            .O(N__4763),
            .I(N__4757));
    InMux I__922 (
            .O(N__4762),
            .I(N__4757));
    LocalMux I__921 (
            .O(N__4757),
            .I(r_Tx_Data_5));
    CascadeMux I__920 (
            .O(N__4754),
            .I(\uart.n2422_cascade_ ));
    InMux I__919 (
            .O(N__4751),
            .I(N__4748));
    LocalMux I__918 (
            .O(N__4748),
            .I(\uart.n2425 ));
    InMux I__917 (
            .O(N__4745),
            .I(N__4739));
    InMux I__916 (
            .O(N__4744),
            .I(N__4739));
    LocalMux I__915 (
            .O(N__4739),
            .I(r_Tx_Data_6));
    InMux I__914 (
            .O(N__4736),
            .I(N__4733));
    LocalMux I__913 (
            .O(N__4733),
            .I(N__4726));
    CascadeMux I__912 (
            .O(N__4732),
            .I(N__4722));
    CascadeMux I__911 (
            .O(N__4731),
            .I(N__4716));
    InMux I__910 (
            .O(N__4730),
            .I(N__4713));
    InMux I__909 (
            .O(N__4729),
            .I(N__4710));
    Span4Mux_v I__908 (
            .O(N__4726),
            .I(N__4707));
    InMux I__907 (
            .O(N__4725),
            .I(N__4704));
    InMux I__906 (
            .O(N__4722),
            .I(N__4697));
    InMux I__905 (
            .O(N__4721),
            .I(N__4697));
    InMux I__904 (
            .O(N__4720),
            .I(N__4697));
    InMux I__903 (
            .O(N__4719),
            .I(N__4692));
    InMux I__902 (
            .O(N__4716),
            .I(N__4692));
    LocalMux I__901 (
            .O(N__4713),
            .I(r_SM_Main_1));
    LocalMux I__900 (
            .O(N__4710),
            .I(r_SM_Main_1));
    Odrv4 I__899 (
            .O(N__4707),
            .I(r_SM_Main_1));
    LocalMux I__898 (
            .O(N__4704),
            .I(r_SM_Main_1));
    LocalMux I__897 (
            .O(N__4697),
            .I(r_SM_Main_1));
    LocalMux I__896 (
            .O(N__4692),
            .I(r_SM_Main_1));
    InMux I__895 (
            .O(N__4679),
            .I(N__4674));
    InMux I__894 (
            .O(N__4678),
            .I(N__4667));
    InMux I__893 (
            .O(N__4677),
            .I(N__4667));
    LocalMux I__892 (
            .O(N__4674),
            .I(N__4664));
    InMux I__891 (
            .O(N__4673),
            .I(N__4657));
    InMux I__890 (
            .O(N__4672),
            .I(N__4657));
    LocalMux I__889 (
            .O(N__4667),
            .I(N__4652));
    Span4Mux_v I__888 (
            .O(N__4664),
            .I(N__4652));
    InMux I__887 (
            .O(N__4663),
            .I(N__4649));
    InMux I__886 (
            .O(N__4662),
            .I(N__4646));
    LocalMux I__885 (
            .O(N__4657),
            .I(r_SM_Main_0));
    Odrv4 I__884 (
            .O(N__4652),
            .I(r_SM_Main_0));
    LocalMux I__883 (
            .O(N__4649),
            .I(r_SM_Main_0));
    LocalMux I__882 (
            .O(N__4646),
            .I(r_SM_Main_0));
    InMux I__881 (
            .O(N__4637),
            .I(N__4633));
    SRMux I__880 (
            .O(N__4636),
            .I(N__4626));
    LocalMux I__879 (
            .O(N__4633),
            .I(N__4623));
    InMux I__878 (
            .O(N__4632),
            .I(N__4620));
    InMux I__877 (
            .O(N__4631),
            .I(N__4617));
    InMux I__876 (
            .O(N__4630),
            .I(N__4612));
    InMux I__875 (
            .O(N__4629),
            .I(N__4612));
    LocalMux I__874 (
            .O(N__4626),
            .I(N__4605));
    Span4Mux_v I__873 (
            .O(N__4623),
            .I(N__4605));
    LocalMux I__872 (
            .O(N__4620),
            .I(N__4605));
    LocalMux I__871 (
            .O(N__4617),
            .I(r_SM_Main_2));
    LocalMux I__870 (
            .O(N__4612),
            .I(r_SM_Main_2));
    Odrv4 I__869 (
            .O(N__4605),
            .I(r_SM_Main_2));
    InMux I__868 (
            .O(N__4598),
            .I(N__4594));
    InMux I__867 (
            .O(N__4597),
            .I(N__4591));
    LocalMux I__866 (
            .O(N__4594),
            .I(r_Tx_Data_1));
    LocalMux I__865 (
            .O(N__4591),
            .I(r_Tx_Data_1));
    InMux I__864 (
            .O(N__4586),
            .I(n2221));
    InMux I__863 (
            .O(N__4583),
            .I(n2222));
    InMux I__862 (
            .O(N__4580),
            .I(n2223));
    InMux I__861 (
            .O(N__4577),
            .I(n2224));
    InMux I__860 (
            .O(N__4574),
            .I(n2225));
    InMux I__859 (
            .O(N__4571),
            .I(N__4566));
    InMux I__858 (
            .O(N__4570),
            .I(N__4563));
    InMux I__857 (
            .O(N__4569),
            .I(N__4560));
    LocalMux I__856 (
            .O(N__4566),
            .I(\uart.r_Bit_Index_2 ));
    LocalMux I__855 (
            .O(N__4563),
            .I(\uart.r_Bit_Index_2 ));
    LocalMux I__854 (
            .O(N__4560),
            .I(\uart.r_Bit_Index_2 ));
    CascadeMux I__853 (
            .O(N__4553),
            .I(n2002_cascade_));
    InMux I__852 (
            .O(N__4550),
            .I(N__4543));
    InMux I__851 (
            .O(N__4549),
            .I(N__4538));
    InMux I__850 (
            .O(N__4548),
            .I(N__4538));
    InMux I__849 (
            .O(N__4547),
            .I(N__4533));
    InMux I__848 (
            .O(N__4546),
            .I(N__4533));
    LocalMux I__847 (
            .O(N__4543),
            .I(N__4530));
    LocalMux I__846 (
            .O(N__4538),
            .I(r_SM_Main_2_N_233_1));
    LocalMux I__845 (
            .O(N__4533),
            .I(r_SM_Main_2_N_233_1));
    Odrv4 I__844 (
            .O(N__4530),
            .I(r_SM_Main_2_N_233_1));
    CascadeMux I__843 (
            .O(N__4523),
            .I(n2308_cascade_));
    InMux I__842 (
            .O(N__4520),
            .I(N__4516));
    InMux I__841 (
            .O(N__4519),
            .I(N__4513));
    LocalMux I__840 (
            .O(N__4516),
            .I(N__4510));
    LocalMux I__839 (
            .O(N__4513),
            .I(n2002));
    Odrv4 I__838 (
            .O(N__4510),
            .I(n2002));
    InMux I__837 (
            .O(N__4505),
            .I(n2211));
    InMux I__836 (
            .O(N__4502),
            .I(n2212));
    InMux I__835 (
            .O(N__4499),
            .I(n2213));
    InMux I__834 (
            .O(N__4496),
            .I(n2214));
    InMux I__833 (
            .O(N__4493),
            .I(n2215));
    InMux I__832 (
            .O(N__4490),
            .I(n2216));
    InMux I__831 (
            .O(N__4487),
            .I(n2217));
    InMux I__830 (
            .O(N__4484),
            .I(bfn_3_25_0_));
    InMux I__829 (
            .O(N__4481),
            .I(n2219));
    InMux I__828 (
            .O(N__4478),
            .I(n2220));
    InMux I__827 (
            .O(N__4475),
            .I(bfn_3_23_0_));
    InMux I__826 (
            .O(N__4472),
            .I(n2203));
    InMux I__825 (
            .O(N__4469),
            .I(n2204));
    InMux I__824 (
            .O(N__4466),
            .I(n2205));
    InMux I__823 (
            .O(N__4463),
            .I(n2206));
    InMux I__822 (
            .O(N__4460),
            .I(n2207));
    InMux I__821 (
            .O(N__4457),
            .I(n2208));
    InMux I__820 (
            .O(N__4454),
            .I(n2209));
    InMux I__819 (
            .O(N__4451),
            .I(bfn_3_24_0_));
    InMux I__818 (
            .O(N__4448),
            .I(N__4445));
    LocalMux I__817 (
            .O(N__4445),
            .I(counter_0));
    InMux I__816 (
            .O(N__4442),
            .I(bfn_3_22_0_));
    InMux I__815 (
            .O(N__4439),
            .I(N__4436));
    LocalMux I__814 (
            .O(N__4436),
            .I(counter_1));
    InMux I__813 (
            .O(N__4433),
            .I(n2195));
    InMux I__812 (
            .O(N__4430),
            .I(N__4427));
    LocalMux I__811 (
            .O(N__4427),
            .I(counter_2));
    InMux I__810 (
            .O(N__4424),
            .I(n2196));
    InMux I__809 (
            .O(N__4421),
            .I(N__4418));
    LocalMux I__808 (
            .O(N__4418),
            .I(counter_3));
    InMux I__807 (
            .O(N__4415),
            .I(n2197));
    InMux I__806 (
            .O(N__4412),
            .I(N__4409));
    LocalMux I__805 (
            .O(N__4409),
            .I(counter_4));
    InMux I__804 (
            .O(N__4406),
            .I(n2198));
    InMux I__803 (
            .O(N__4403),
            .I(N__4400));
    LocalMux I__802 (
            .O(N__4400),
            .I(counter_5));
    InMux I__801 (
            .O(N__4397),
            .I(n2199));
    InMux I__800 (
            .O(N__4394),
            .I(N__4391));
    LocalMux I__799 (
            .O(N__4391),
            .I(counter_6));
    InMux I__798 (
            .O(N__4388),
            .I(n2200));
    InMux I__797 (
            .O(N__4385),
            .I(N__4382));
    LocalMux I__796 (
            .O(N__4382),
            .I(counter_7));
    InMux I__795 (
            .O(N__4379),
            .I(n2201));
    InMux I__794 (
            .O(N__4376),
            .I(n2187));
    InMux I__793 (
            .O(N__4373),
            .I(N__4369));
    InMux I__792 (
            .O(N__4372),
            .I(N__4366));
    LocalMux I__791 (
            .O(N__4369),
            .I(blink_counter_25));
    LocalMux I__790 (
            .O(N__4366),
            .I(blink_counter_25));
    CascadeMux I__789 (
            .O(N__4361),
            .I(n2395_cascade_));
    IoInMux I__788 (
            .O(N__4358),
            .I(N__4355));
    LocalMux I__787 (
            .O(N__4355),
            .I(N__4352));
    Span4Mux_s1_v I__786 (
            .O(N__4352),
            .I(N__4349));
    Span4Mux_v I__785 (
            .O(N__4349),
            .I(N__4346));
    Odrv4 I__784 (
            .O(N__4346),
            .I(LED_c));
    InMux I__783 (
            .O(N__4343),
            .I(N__4337));
    InMux I__782 (
            .O(N__4342),
            .I(N__4337));
    LocalMux I__781 (
            .O(N__4337),
            .I(N__4333));
    InMux I__780 (
            .O(N__4336),
            .I(N__4330));
    Odrv4 I__779 (
            .O(N__4333),
            .I(blink_counter_21));
    LocalMux I__778 (
            .O(N__4330),
            .I(blink_counter_21));
    InMux I__777 (
            .O(N__4325),
            .I(N__4318));
    InMux I__776 (
            .O(N__4324),
            .I(N__4318));
    InMux I__775 (
            .O(N__4323),
            .I(N__4315));
    LocalMux I__774 (
            .O(N__4318),
            .I(blink_counter_24));
    LocalMux I__773 (
            .O(N__4315),
            .I(blink_counter_24));
    CascadeMux I__772 (
            .O(N__4310),
            .I(N__4306));
    CascadeMux I__771 (
            .O(N__4309),
            .I(N__4303));
    InMux I__770 (
            .O(N__4306),
            .I(N__4298));
    InMux I__769 (
            .O(N__4303),
            .I(N__4298));
    LocalMux I__768 (
            .O(N__4298),
            .I(N__4294));
    InMux I__767 (
            .O(N__4297),
            .I(N__4291));
    Odrv4 I__766 (
            .O(N__4294),
            .I(blink_counter_23));
    LocalMux I__765 (
            .O(N__4291),
            .I(blink_counter_23));
    InMux I__764 (
            .O(N__4286),
            .I(N__4280));
    InMux I__763 (
            .O(N__4285),
            .I(N__4280));
    LocalMux I__762 (
            .O(N__4280),
            .I(N__4276));
    InMux I__761 (
            .O(N__4279),
            .I(N__4273));
    Odrv4 I__760 (
            .O(N__4276),
            .I(blink_counter_22));
    LocalMux I__759 (
            .O(N__4273),
            .I(blink_counter_22));
    InMux I__758 (
            .O(N__4268),
            .I(N__4265));
    LocalMux I__757 (
            .O(N__4265),
            .I(n2394));
    InMux I__756 (
            .O(N__4262),
            .I(N__4259));
    LocalMux I__755 (
            .O(N__4259),
            .I(\uart.n1711 ));
    InMux I__754 (
            .O(N__4256),
            .I(N__4253));
    LocalMux I__753 (
            .O(N__4253),
            .I(\uart.o_Tx_Serial_N_312 ));
    InMux I__752 (
            .O(N__4250),
            .I(N__4247));
    LocalMux I__751 (
            .O(N__4247),
            .I(N__4243));
    InMux I__750 (
            .O(N__4246),
            .I(N__4240));
    Span4Mux_h I__749 (
            .O(N__4243),
            .I(N__4237));
    LocalMux I__748 (
            .O(N__4240),
            .I(clk_divider_7));
    Odrv4 I__747 (
            .O(N__4237),
            .I(clk_divider_7));
    InMux I__746 (
            .O(N__4232),
            .I(N__4229));
    LocalMux I__745 (
            .O(N__4229),
            .I(n40_adj_362));
    CascadeMux I__744 (
            .O(N__4226),
            .I(N__4223));
    InMux I__743 (
            .O(N__4223),
            .I(N__4220));
    LocalMux I__742 (
            .O(N__4220),
            .I(N__4216));
    InMux I__741 (
            .O(N__4219),
            .I(N__4213));
    Span4Mux_h I__740 (
            .O(N__4216),
            .I(N__4210));
    LocalMux I__739 (
            .O(N__4213),
            .I(clk_divider_25));
    Odrv4 I__738 (
            .O(N__4210),
            .I(clk_divider_25));
    InMux I__737 (
            .O(N__4205),
            .I(N__4202));
    LocalMux I__736 (
            .O(N__4202),
            .I(n45_adj_357));
    InMux I__735 (
            .O(N__4199),
            .I(N__4193));
    InMux I__734 (
            .O(N__4198),
            .I(N__4193));
    LocalMux I__733 (
            .O(N__4193),
            .I(n49));
    InMux I__732 (
            .O(N__4190),
            .I(N__4187));
    LocalMux I__731 (
            .O(N__4187),
            .I(n9));
    InMux I__730 (
            .O(N__4184),
            .I(n2179));
    InMux I__729 (
            .O(N__4181),
            .I(N__4178));
    LocalMux I__728 (
            .O(N__4178),
            .I(n8));
    InMux I__727 (
            .O(N__4175),
            .I(n2180));
    InMux I__726 (
            .O(N__4172),
            .I(N__4169));
    LocalMux I__725 (
            .O(N__4169),
            .I(n7));
    InMux I__724 (
            .O(N__4166),
            .I(n2181));
    InMux I__723 (
            .O(N__4163),
            .I(N__4160));
    LocalMux I__722 (
            .O(N__4160),
            .I(n6));
    InMux I__721 (
            .O(N__4157),
            .I(n2182));
    InMux I__720 (
            .O(N__4154),
            .I(n2183));
    InMux I__719 (
            .O(N__4151),
            .I(n2184));
    InMux I__718 (
            .O(N__4148),
            .I(n2185));
    InMux I__717 (
            .O(N__4145),
            .I(bfn_2_26_0_));
    InMux I__716 (
            .O(N__4142),
            .I(N__4139));
    LocalMux I__715 (
            .O(N__4139),
            .I(n18));
    InMux I__714 (
            .O(N__4136),
            .I(bfn_2_24_0_));
    InMux I__713 (
            .O(N__4133),
            .I(N__4130));
    LocalMux I__712 (
            .O(N__4130),
            .I(n17));
    InMux I__711 (
            .O(N__4127),
            .I(n2171));
    InMux I__710 (
            .O(N__4124),
            .I(N__4121));
    LocalMux I__709 (
            .O(N__4121),
            .I(n16));
    InMux I__708 (
            .O(N__4118),
            .I(n2172));
    InMux I__707 (
            .O(N__4115),
            .I(N__4112));
    LocalMux I__706 (
            .O(N__4112),
            .I(n15));
    InMux I__705 (
            .O(N__4109),
            .I(n2173));
    InMux I__704 (
            .O(N__4106),
            .I(N__4103));
    LocalMux I__703 (
            .O(N__4103),
            .I(n14));
    InMux I__702 (
            .O(N__4100),
            .I(n2174));
    InMux I__701 (
            .O(N__4097),
            .I(N__4094));
    LocalMux I__700 (
            .O(N__4094),
            .I(n13));
    InMux I__699 (
            .O(N__4091),
            .I(n2175));
    InMux I__698 (
            .O(N__4088),
            .I(N__4085));
    LocalMux I__697 (
            .O(N__4085),
            .I(n12));
    InMux I__696 (
            .O(N__4082),
            .I(n2176));
    InMux I__695 (
            .O(N__4079),
            .I(N__4076));
    LocalMux I__694 (
            .O(N__4076),
            .I(n11));
    InMux I__693 (
            .O(N__4073),
            .I(n2177));
    InMux I__692 (
            .O(N__4070),
            .I(N__4067));
    LocalMux I__691 (
            .O(N__4067),
            .I(n10_adj_317));
    InMux I__690 (
            .O(N__4064),
            .I(bfn_2_25_0_));
    InMux I__689 (
            .O(N__4061),
            .I(N__4058));
    LocalMux I__688 (
            .O(N__4058),
            .I(n26));
    InMux I__687 (
            .O(N__4055),
            .I(bfn_2_23_0_));
    InMux I__686 (
            .O(N__4052),
            .I(N__4049));
    LocalMux I__685 (
            .O(N__4049),
            .I(n25));
    InMux I__684 (
            .O(N__4046),
            .I(n2163));
    InMux I__683 (
            .O(N__4043),
            .I(N__4040));
    LocalMux I__682 (
            .O(N__4040),
            .I(n24));
    InMux I__681 (
            .O(N__4037),
            .I(n2164));
    InMux I__680 (
            .O(N__4034),
            .I(N__4031));
    LocalMux I__679 (
            .O(N__4031),
            .I(n23));
    InMux I__678 (
            .O(N__4028),
            .I(n2165));
    InMux I__677 (
            .O(N__4025),
            .I(N__4022));
    LocalMux I__676 (
            .O(N__4022),
            .I(n22));
    InMux I__675 (
            .O(N__4019),
            .I(n2166));
    InMux I__674 (
            .O(N__4016),
            .I(N__4013));
    LocalMux I__673 (
            .O(N__4013),
            .I(n21));
    InMux I__672 (
            .O(N__4010),
            .I(n2167));
    InMux I__671 (
            .O(N__4007),
            .I(N__4004));
    LocalMux I__670 (
            .O(N__4004),
            .I(n20));
    InMux I__669 (
            .O(N__4001),
            .I(n2168));
    InMux I__668 (
            .O(N__3998),
            .I(N__3995));
    LocalMux I__667 (
            .O(N__3995),
            .I(n19));
    InMux I__666 (
            .O(N__3992),
            .I(n2169));
    InMux I__665 (
            .O(N__3989),
            .I(N__3985));
    InMux I__664 (
            .O(N__3988),
            .I(N__3982));
    LocalMux I__663 (
            .O(N__3985),
            .I(N__3979));
    LocalMux I__662 (
            .O(N__3982),
            .I(clk_divider_4));
    Odrv4 I__661 (
            .O(N__3979),
            .I(clk_divider_4));
    InMux I__660 (
            .O(N__3974),
            .I(N__3970));
    InMux I__659 (
            .O(N__3973),
            .I(N__3967));
    LocalMux I__658 (
            .O(N__3970),
            .I(clk_divider_0));
    LocalMux I__657 (
            .O(N__3967),
            .I(clk_divider_0));
    CascadeMux I__656 (
            .O(N__3962),
            .I(N__3958));
    InMux I__655 (
            .O(N__3961),
            .I(N__3955));
    InMux I__654 (
            .O(N__3958),
            .I(N__3952));
    LocalMux I__653 (
            .O(N__3955),
            .I(clk_divider_3));
    LocalMux I__652 (
            .O(N__3952),
            .I(clk_divider_3));
    SRMux I__651 (
            .O(N__3947),
            .I(N__3943));
    SRMux I__650 (
            .O(N__3946),
            .I(N__3939));
    LocalMux I__649 (
            .O(N__3943),
            .I(N__3935));
    SRMux I__648 (
            .O(N__3942),
            .I(N__3932));
    LocalMux I__647 (
            .O(N__3939),
            .I(N__3929));
    SRMux I__646 (
            .O(N__3938),
            .I(N__3926));
    Span4Mux_v I__645 (
            .O(N__3935),
            .I(N__3921));
    LocalMux I__644 (
            .O(N__3932),
            .I(N__3921));
    Span4Mux_v I__643 (
            .O(N__3929),
            .I(N__3916));
    LocalMux I__642 (
            .O(N__3926),
            .I(N__3916));
    Odrv4 I__641 (
            .O(N__3921),
            .I(clk_divider_31__N_139));
    Odrv4 I__640 (
            .O(N__3916),
            .I(clk_divider_31__N_139));
    IoInMux I__639 (
            .O(N__3911),
            .I(N__3908));
    LocalMux I__638 (
            .O(N__3908),
            .I(N__3905));
    Span12Mux_s1_v I__637 (
            .O(N__3905),
            .I(N__3902));
    Odrv12 I__636 (
            .O(N__3902),
            .I(\uart.n3 ));
    InMux I__635 (
            .O(N__3899),
            .I(N__3895));
    InMux I__634 (
            .O(N__3898),
            .I(N__3892));
    LocalMux I__633 (
            .O(N__3895),
            .I(clk_divider_1));
    LocalMux I__632 (
            .O(N__3892),
            .I(clk_divider_1));
    InMux I__631 (
            .O(N__3887),
            .I(N__3883));
    InMux I__630 (
            .O(N__3886),
            .I(N__3880));
    LocalMux I__629 (
            .O(N__3883),
            .I(clk_divider_2));
    LocalMux I__628 (
            .O(N__3880),
            .I(clk_divider_2));
    InMux I__627 (
            .O(N__3875),
            .I(N__3872));
    LocalMux I__626 (
            .O(N__3872),
            .I(n6_adj_324));
    InMux I__625 (
            .O(N__3869),
            .I(N__3865));
    InMux I__624 (
            .O(N__3868),
            .I(N__3862));
    LocalMux I__623 (
            .O(N__3865),
            .I(clk_divider_8));
    LocalMux I__622 (
            .O(N__3862),
            .I(clk_divider_8));
    InMux I__621 (
            .O(N__3857),
            .I(N__3853));
    InMux I__620 (
            .O(N__3856),
            .I(N__3850));
    LocalMux I__619 (
            .O(N__3853),
            .I(clk_divider_15));
    LocalMux I__618 (
            .O(N__3850),
            .I(clk_divider_15));
    CascadeMux I__617 (
            .O(N__3845),
            .I(N__3842));
    InMux I__616 (
            .O(N__3842),
            .I(N__3838));
    InMux I__615 (
            .O(N__3841),
            .I(N__3835));
    LocalMux I__614 (
            .O(N__3838),
            .I(N__3832));
    LocalMux I__613 (
            .O(N__3835),
            .I(clk_divider_24));
    Odrv4 I__612 (
            .O(N__3832),
            .I(clk_divider_24));
    InMux I__611 (
            .O(N__3827),
            .I(N__3823));
    InMux I__610 (
            .O(N__3826),
            .I(N__3820));
    LocalMux I__609 (
            .O(N__3823),
            .I(clk_divider_11));
    LocalMux I__608 (
            .O(N__3820),
            .I(clk_divider_11));
    InMux I__607 (
            .O(N__3815),
            .I(N__3811));
    InMux I__606 (
            .O(N__3814),
            .I(N__3808));
    LocalMux I__605 (
            .O(N__3811),
            .I(clk_divider_5));
    LocalMux I__604 (
            .O(N__3808),
            .I(clk_divider_5));
    InMux I__603 (
            .O(N__3803),
            .I(N__3799));
    InMux I__602 (
            .O(N__3802),
            .I(N__3796));
    LocalMux I__601 (
            .O(N__3799),
            .I(clk_divider_10));
    LocalMux I__600 (
            .O(N__3796),
            .I(clk_divider_10));
    CascadeMux I__599 (
            .O(N__3791),
            .I(N__3787));
    InMux I__598 (
            .O(N__3790),
            .I(N__3784));
    InMux I__597 (
            .O(N__3787),
            .I(N__3781));
    LocalMux I__596 (
            .O(N__3784),
            .I(clk_divider_12));
    LocalMux I__595 (
            .O(N__3781),
            .I(clk_divider_12));
    InMux I__594 (
            .O(N__3776),
            .I(N__3772));
    InMux I__593 (
            .O(N__3775),
            .I(N__3769));
    LocalMux I__592 (
            .O(N__3772),
            .I(N__3766));
    LocalMux I__591 (
            .O(N__3769),
            .I(clk_divider_18));
    Odrv4 I__590 (
            .O(N__3766),
            .I(clk_divider_18));
    InMux I__589 (
            .O(N__3761),
            .I(N__3757));
    InMux I__588 (
            .O(N__3760),
            .I(N__3754));
    LocalMux I__587 (
            .O(N__3757),
            .I(clk_divider_13));
    LocalMux I__586 (
            .O(N__3754),
            .I(clk_divider_13));
    InMux I__585 (
            .O(N__3749),
            .I(N__3745));
    InMux I__584 (
            .O(N__3748),
            .I(N__3742));
    LocalMux I__583 (
            .O(N__3745),
            .I(N__3739));
    LocalMux I__582 (
            .O(N__3742),
            .I(clk_divider_29));
    Odrv4 I__581 (
            .O(N__3739),
            .I(clk_divider_29));
    CascadeMux I__580 (
            .O(N__3734),
            .I(N__3731));
    InMux I__579 (
            .O(N__3731),
            .I(N__3728));
    LocalMux I__578 (
            .O(N__3728),
            .I(N__3724));
    InMux I__577 (
            .O(N__3727),
            .I(N__3721));
    Span4Mux_h I__576 (
            .O(N__3724),
            .I(N__3718));
    LocalMux I__575 (
            .O(N__3721),
            .I(clk_divider_23));
    Odrv4 I__574 (
            .O(N__3718),
            .I(clk_divider_23));
    InMux I__573 (
            .O(N__3713),
            .I(N__3709));
    InMux I__572 (
            .O(N__3712),
            .I(N__3706));
    LocalMux I__571 (
            .O(N__3709),
            .I(N__3703));
    LocalMux I__570 (
            .O(N__3706),
            .I(clk_divider_16));
    Odrv4 I__569 (
            .O(N__3703),
            .I(clk_divider_16));
    InMux I__568 (
            .O(N__3698),
            .I(N__3695));
    LocalMux I__567 (
            .O(N__3695),
            .I(n43_adj_359));
    CascadeMux I__566 (
            .O(N__3692),
            .I(N__3688));
    InMux I__565 (
            .O(N__3691),
            .I(N__3683));
    InMux I__564 (
            .O(N__3688),
            .I(N__3683));
    LocalMux I__563 (
            .O(N__3683),
            .I(N__3679));
    InMux I__562 (
            .O(N__3682),
            .I(N__3676));
    Span4Mux_h I__561 (
            .O(N__3679),
            .I(N__3673));
    LocalMux I__560 (
            .O(N__3676),
            .I(clk_divider_31));
    Odrv4 I__559 (
            .O(N__3673),
            .I(clk_divider_31));
    CascadeMux I__558 (
            .O(N__3668),
            .I(N__3665));
    InMux I__557 (
            .O(N__3665),
            .I(N__3659));
    InMux I__556 (
            .O(N__3664),
            .I(N__3659));
    LocalMux I__555 (
            .O(N__3659),
            .I(n50));
    InMux I__554 (
            .O(N__3656),
            .I(N__3650));
    InMux I__553 (
            .O(N__3655),
            .I(N__3650));
    LocalMux I__552 (
            .O(N__3650),
            .I(N__3647));
    Odrv4 I__551 (
            .O(N__3647),
            .I(n10));
    InMux I__550 (
            .O(N__3644),
            .I(N__3640));
    InMux I__549 (
            .O(N__3643),
            .I(N__3637));
    LocalMux I__548 (
            .O(N__3640),
            .I(\uart.r_Clock_Count_20 ));
    LocalMux I__547 (
            .O(N__3637),
            .I(\uart.r_Clock_Count_20 ));
    InMux I__546 (
            .O(N__3632),
            .I(N__3628));
    InMux I__545 (
            .O(N__3631),
            .I(N__3625));
    LocalMux I__544 (
            .O(N__3628),
            .I(\uart.r_Clock_Count_15 ));
    LocalMux I__543 (
            .O(N__3625),
            .I(\uart.r_Clock_Count_15 ));
    CascadeMux I__542 (
            .O(N__3620),
            .I(N__3616));
    InMux I__541 (
            .O(N__3619),
            .I(N__3613));
    InMux I__540 (
            .O(N__3616),
            .I(N__3610));
    LocalMux I__539 (
            .O(N__3613),
            .I(\uart.r_Clock_Count_25 ));
    LocalMux I__538 (
            .O(N__3610),
            .I(\uart.r_Clock_Count_25 ));
    InMux I__537 (
            .O(N__3605),
            .I(N__3601));
    InMux I__536 (
            .O(N__3604),
            .I(N__3598));
    LocalMux I__535 (
            .O(N__3601),
            .I(\uart.r_Clock_Count_9 ));
    LocalMux I__534 (
            .O(N__3598),
            .I(\uart.r_Clock_Count_9 ));
    InMux I__533 (
            .O(N__3593),
            .I(N__3589));
    InMux I__532 (
            .O(N__3592),
            .I(N__3586));
    LocalMux I__531 (
            .O(N__3589),
            .I(N__3583));
    LocalMux I__530 (
            .O(N__3586),
            .I(\uart.r_Clock_Count_27 ));
    Odrv4 I__529 (
            .O(N__3583),
            .I(\uart.r_Clock_Count_27 ));
    InMux I__528 (
            .O(N__3578),
            .I(N__3574));
    InMux I__527 (
            .O(N__3577),
            .I(N__3571));
    LocalMux I__526 (
            .O(N__3574),
            .I(\uart.r_Clock_Count_19 ));
    LocalMux I__525 (
            .O(N__3571),
            .I(\uart.r_Clock_Count_19 ));
    CascadeMux I__524 (
            .O(N__3566),
            .I(N__3562));
    InMux I__523 (
            .O(N__3565),
            .I(N__3559));
    InMux I__522 (
            .O(N__3562),
            .I(N__3556));
    LocalMux I__521 (
            .O(N__3559),
            .I(\uart.r_Clock_Count_16 ));
    LocalMux I__520 (
            .O(N__3556),
            .I(\uart.r_Clock_Count_16 ));
    InMux I__519 (
            .O(N__3551),
            .I(N__3547));
    InMux I__518 (
            .O(N__3550),
            .I(N__3544));
    LocalMux I__517 (
            .O(N__3547),
            .I(\uart.r_Clock_Count_31 ));
    LocalMux I__516 (
            .O(N__3544),
            .I(\uart.r_Clock_Count_31 ));
    InMux I__515 (
            .O(N__3539),
            .I(N__3536));
    LocalMux I__514 (
            .O(N__3536),
            .I(\uart.n39 ));
    InMux I__513 (
            .O(N__3533),
            .I(N__3530));
    LocalMux I__512 (
            .O(N__3530),
            .I(\uart.n40 ));
    CascadeMux I__511 (
            .O(N__3527),
            .I(\uart.n37_cascade_ ));
    InMux I__510 (
            .O(N__3524),
            .I(N__3521));
    LocalMux I__509 (
            .O(N__3521),
            .I(\uart.n38 ));
    InMux I__508 (
            .O(N__3518),
            .I(N__3515));
    LocalMux I__507 (
            .O(N__3515),
            .I(N__3512));
    Odrv4 I__506 (
            .O(N__3512),
            .I(\uart.n46 ));
    InMux I__505 (
            .O(N__3509),
            .I(N__3506));
    LocalMux I__504 (
            .O(N__3506),
            .I(N__3502));
    InMux I__503 (
            .O(N__3505),
            .I(N__3499));
    Span4Mux_h I__502 (
            .O(N__3502),
            .I(N__3496));
    LocalMux I__501 (
            .O(N__3499),
            .I(clk_divider_26));
    Odrv4 I__500 (
            .O(N__3496),
            .I(clk_divider_26));
    InMux I__499 (
            .O(N__3491),
            .I(N__3487));
    InMux I__498 (
            .O(N__3490),
            .I(N__3484));
    LocalMux I__497 (
            .O(N__3487),
            .I(N__3481));
    LocalMux I__496 (
            .O(N__3484),
            .I(clk_divider_9));
    Odrv4 I__495 (
            .O(N__3481),
            .I(clk_divider_9));
    CascadeMux I__494 (
            .O(N__3476),
            .I(N__3473));
    InMux I__493 (
            .O(N__3473),
            .I(N__3469));
    InMux I__492 (
            .O(N__3472),
            .I(N__3466));
    LocalMux I__491 (
            .O(N__3469),
            .I(N__3463));
    LocalMux I__490 (
            .O(N__3466),
            .I(clk_divider_14));
    Odrv4 I__489 (
            .O(N__3463),
            .I(clk_divider_14));
    InMux I__488 (
            .O(N__3458),
            .I(N__3455));
    LocalMux I__487 (
            .O(N__3455),
            .I(N__3451));
    InMux I__486 (
            .O(N__3454),
            .I(N__3448));
    Span4Mux_h I__485 (
            .O(N__3451),
            .I(N__3445));
    LocalMux I__484 (
            .O(N__3448),
            .I(clk_divider_17));
    Odrv4 I__483 (
            .O(N__3445),
            .I(clk_divider_17));
    InMux I__482 (
            .O(N__3440),
            .I(N__3436));
    InMux I__481 (
            .O(N__3439),
            .I(N__3433));
    LocalMux I__480 (
            .O(N__3436),
            .I(N__3430));
    LocalMux I__479 (
            .O(N__3433),
            .I(clk_divider_21));
    Odrv4 I__478 (
            .O(N__3430),
            .I(clk_divider_21));
    InMux I__477 (
            .O(N__3425),
            .I(N__3422));
    LocalMux I__476 (
            .O(N__3422),
            .I(N__3418));
    InMux I__475 (
            .O(N__3421),
            .I(N__3415));
    Span4Mux_h I__474 (
            .O(N__3418),
            .I(N__3412));
    LocalMux I__473 (
            .O(N__3415),
            .I(clk_divider_22));
    Odrv4 I__472 (
            .O(N__3412),
            .I(clk_divider_22));
    CascadeMux I__471 (
            .O(N__3407),
            .I(N__3404));
    InMux I__470 (
            .O(N__3404),
            .I(N__3401));
    LocalMux I__469 (
            .O(N__3401),
            .I(N__3397));
    InMux I__468 (
            .O(N__3400),
            .I(N__3394));
    Span4Mux_h I__467 (
            .O(N__3397),
            .I(N__3391));
    LocalMux I__466 (
            .O(N__3394),
            .I(clk_divider_28));
    Odrv4 I__465 (
            .O(N__3391),
            .I(clk_divider_28));
    InMux I__464 (
            .O(N__3386),
            .I(N__3382));
    InMux I__463 (
            .O(N__3385),
            .I(N__3379));
    LocalMux I__462 (
            .O(N__3382),
            .I(clk_divider_6));
    LocalMux I__461 (
            .O(N__3379),
            .I(clk_divider_6));
    InMux I__460 (
            .O(N__3374),
            .I(N__3371));
    LocalMux I__459 (
            .O(N__3371),
            .I(N__3367));
    InMux I__458 (
            .O(N__3370),
            .I(N__3364));
    Span4Mux_v I__457 (
            .O(N__3367),
            .I(N__3361));
    LocalMux I__456 (
            .O(N__3364),
            .I(clk_divider_30));
    Odrv4 I__455 (
            .O(N__3361),
            .I(clk_divider_30));
    InMux I__454 (
            .O(N__3356),
            .I(N__3353));
    LocalMux I__453 (
            .O(N__3353),
            .I(N__3349));
    InMux I__452 (
            .O(N__3352),
            .I(N__3346));
    Span4Mux_h I__451 (
            .O(N__3349),
            .I(N__3343));
    LocalMux I__450 (
            .O(N__3346),
            .I(clk_divider_27));
    Odrv4 I__449 (
            .O(N__3343),
            .I(clk_divider_27));
    CascadeMux I__448 (
            .O(N__3338),
            .I(N__3335));
    InMux I__447 (
            .O(N__3335),
            .I(N__3331));
    InMux I__446 (
            .O(N__3334),
            .I(N__3328));
    LocalMux I__445 (
            .O(N__3331),
            .I(N__3325));
    LocalMux I__444 (
            .O(N__3328),
            .I(clk_divider_20));
    Odrv4 I__443 (
            .O(N__3325),
            .I(clk_divider_20));
    InMux I__442 (
            .O(N__3320),
            .I(N__3316));
    InMux I__441 (
            .O(N__3319),
            .I(N__3313));
    LocalMux I__440 (
            .O(N__3316),
            .I(N__3310));
    LocalMux I__439 (
            .O(N__3313),
            .I(clk_divider_19));
    Odrv4 I__438 (
            .O(N__3310),
            .I(clk_divider_19));
    InMux I__437 (
            .O(N__3305),
            .I(N__3302));
    LocalMux I__436 (
            .O(N__3302),
            .I(n44_adj_358));
    CascadeMux I__435 (
            .O(N__3299),
            .I(n42_adj_360_cascade_));
    InMux I__434 (
            .O(N__3296),
            .I(N__3293));
    LocalMux I__433 (
            .O(N__3293),
            .I(n41_adj_361));
    InMux I__432 (
            .O(N__3290),
            .I(N__3286));
    InMux I__431 (
            .O(N__3289),
            .I(N__3283));
    LocalMux I__430 (
            .O(N__3286),
            .I(\uart.r_Clock_Count_13 ));
    LocalMux I__429 (
            .O(N__3283),
            .I(\uart.r_Clock_Count_13 ));
    InMux I__428 (
            .O(N__3278),
            .I(N__3274));
    InMux I__427 (
            .O(N__3277),
            .I(N__3271));
    LocalMux I__426 (
            .O(N__3274),
            .I(\uart.r_Clock_Count_12 ));
    LocalMux I__425 (
            .O(N__3271),
            .I(\uart.r_Clock_Count_12 ));
    InMux I__424 (
            .O(N__3266),
            .I(N__3262));
    InMux I__423 (
            .O(N__3265),
            .I(N__3259));
    LocalMux I__422 (
            .O(N__3262),
            .I(N__3256));
    LocalMux I__421 (
            .O(N__3259),
            .I(\uart.r_Clock_Count_29 ));
    Odrv4 I__420 (
            .O(N__3256),
            .I(\uart.r_Clock_Count_29 ));
    CascadeMux I__419 (
            .O(N__3251),
            .I(\uart.n42_cascade_ ));
    InMux I__418 (
            .O(N__3248),
            .I(N__3244));
    InMux I__417 (
            .O(N__3247),
            .I(N__3241));
    LocalMux I__416 (
            .O(N__3244),
            .I(\uart.r_Clock_Count_7 ));
    LocalMux I__415 (
            .O(N__3241),
            .I(\uart.r_Clock_Count_7 ));
    CascadeMux I__414 (
            .O(N__3236),
            .I(\uart.n45_cascade_ ));
    InMux I__413 (
            .O(N__3233),
            .I(N__3230));
    LocalMux I__412 (
            .O(N__3230),
            .I(\uart.n2385 ));
    CascadeMux I__411 (
            .O(N__3227),
            .I(r_SM_Main_2_N_233_1_cascade_));
    SRMux I__410 (
            .O(N__3224),
            .I(N__3221));
    LocalMux I__409 (
            .O(N__3221),
            .I(N__3218));
    Span4Mux_s1_h I__408 (
            .O(N__3218),
            .I(N__3212));
    SRMux I__407 (
            .O(N__3217),
            .I(N__3209));
    SRMux I__406 (
            .O(N__3216),
            .I(N__3206));
    SRMux I__405 (
            .O(N__3215),
            .I(N__3203));
    Odrv4 I__404 (
            .O(N__3212),
            .I(\uart.n1796 ));
    LocalMux I__403 (
            .O(N__3209),
            .I(\uart.n1796 ));
    LocalMux I__402 (
            .O(N__3206),
            .I(\uart.n1796 ));
    LocalMux I__401 (
            .O(N__3203),
            .I(\uart.n1796 ));
    CascadeMux I__400 (
            .O(N__3194),
            .I(N__3190));
    InMux I__399 (
            .O(N__3193),
            .I(N__3187));
    InMux I__398 (
            .O(N__3190),
            .I(N__3184));
    LocalMux I__397 (
            .O(N__3187),
            .I(\uart.r_Clock_Count_8 ));
    LocalMux I__396 (
            .O(N__3184),
            .I(\uart.r_Clock_Count_8 ));
    InMux I__395 (
            .O(N__3179),
            .I(N__3175));
    InMux I__394 (
            .O(N__3178),
            .I(N__3172));
    LocalMux I__393 (
            .O(N__3175),
            .I(\uart.r_Clock_Count_14 ));
    LocalMux I__392 (
            .O(N__3172),
            .I(\uart.r_Clock_Count_14 ));
    InMux I__391 (
            .O(N__3167),
            .I(N__3164));
    LocalMux I__390 (
            .O(N__3164),
            .I(\uart.n34 ));
    InMux I__389 (
            .O(N__3161),
            .I(N__3157));
    InMux I__388 (
            .O(N__3160),
            .I(N__3154));
    LocalMux I__387 (
            .O(N__3157),
            .I(\uart.r_Clock_Count_30 ));
    LocalMux I__386 (
            .O(N__3154),
            .I(\uart.r_Clock_Count_30 ));
    InMux I__385 (
            .O(N__3149),
            .I(N__3145));
    InMux I__384 (
            .O(N__3148),
            .I(N__3142));
    LocalMux I__383 (
            .O(N__3145),
            .I(\uart.r_Clock_Count_28 ));
    LocalMux I__382 (
            .O(N__3142),
            .I(\uart.r_Clock_Count_28 ));
    CascadeMux I__381 (
            .O(N__3137),
            .I(N__3134));
    InMux I__380 (
            .O(N__3134),
            .I(N__3130));
    InMux I__379 (
            .O(N__3133),
            .I(N__3127));
    LocalMux I__378 (
            .O(N__3130),
            .I(N__3124));
    LocalMux I__377 (
            .O(N__3127),
            .I(\uart.r_Clock_Count_24 ));
    Odrv4 I__376 (
            .O(N__3124),
            .I(\uart.r_Clock_Count_24 ));
    InMux I__375 (
            .O(N__3119),
            .I(N__3115));
    InMux I__374 (
            .O(N__3118),
            .I(N__3112));
    LocalMux I__373 (
            .O(N__3115),
            .I(\uart.r_Clock_Count_23 ));
    LocalMux I__372 (
            .O(N__3112),
            .I(\uart.r_Clock_Count_23 ));
    CEMux I__371 (
            .O(N__3107),
            .I(N__3103));
    CEMux I__370 (
            .O(N__3106),
            .I(N__3100));
    LocalMux I__369 (
            .O(N__3103),
            .I(N__3097));
    LocalMux I__368 (
            .O(N__3100),
            .I(N__3091));
    Span4Mux_s2_v I__367 (
            .O(N__3097),
            .I(N__3088));
    CEMux I__366 (
            .O(N__3096),
            .I(N__3085));
    CEMux I__365 (
            .O(N__3095),
            .I(N__3082));
    CEMux I__364 (
            .O(N__3094),
            .I(N__3079));
    Sp12to4 I__363 (
            .O(N__3091),
            .I(N__3074));
    Sp12to4 I__362 (
            .O(N__3088),
            .I(N__3074));
    LocalMux I__361 (
            .O(N__3085),
            .I(\uart.n1 ));
    LocalMux I__360 (
            .O(N__3082),
            .I(\uart.n1 ));
    LocalMux I__359 (
            .O(N__3079),
            .I(\uart.n1 ));
    Odrv12 I__358 (
            .O(N__3074),
            .I(\uart.n1 ));
    InMux I__357 (
            .O(N__3065),
            .I(N__3061));
    InMux I__356 (
            .O(N__3064),
            .I(N__3058));
    LocalMux I__355 (
            .O(N__3061),
            .I(\uart.r_Clock_Count_11 ));
    LocalMux I__354 (
            .O(N__3058),
            .I(\uart.r_Clock_Count_11 ));
    InMux I__353 (
            .O(N__3053),
            .I(N__3049));
    InMux I__352 (
            .O(N__3052),
            .I(N__3046));
    LocalMux I__351 (
            .O(N__3049),
            .I(\uart.r_Clock_Count_21 ));
    LocalMux I__350 (
            .O(N__3046),
            .I(\uart.r_Clock_Count_21 ));
    CascadeMux I__349 (
            .O(N__3041),
            .I(N__3037));
    InMux I__348 (
            .O(N__3040),
            .I(N__3034));
    InMux I__347 (
            .O(N__3037),
            .I(N__3031));
    LocalMux I__346 (
            .O(N__3034),
            .I(\uart.r_Clock_Count_17 ));
    LocalMux I__345 (
            .O(N__3031),
            .I(\uart.r_Clock_Count_17 ));
    InMux I__344 (
            .O(N__3026),
            .I(N__3022));
    InMux I__343 (
            .O(N__3025),
            .I(N__3019));
    LocalMux I__342 (
            .O(N__3022),
            .I(\uart.r_Clock_Count_18 ));
    LocalMux I__341 (
            .O(N__3019),
            .I(\uart.r_Clock_Count_18 ));
    InMux I__340 (
            .O(N__3014),
            .I(n2252));
    InMux I__339 (
            .O(N__3011),
            .I(n2253));
    InMux I__338 (
            .O(N__3008),
            .I(n2254));
    InMux I__337 (
            .O(N__3005),
            .I(n2255));
    InMux I__336 (
            .O(N__3002),
            .I(n2256));
    InMux I__335 (
            .O(N__2999),
            .I(N__2995));
    InMux I__334 (
            .O(N__2998),
            .I(N__2992));
    LocalMux I__333 (
            .O(N__2995),
            .I(\uart.r_Clock_Count_2 ));
    LocalMux I__332 (
            .O(N__2992),
            .I(\uart.r_Clock_Count_2 ));
    InMux I__331 (
            .O(N__2987),
            .I(N__2983));
    InMux I__330 (
            .O(N__2986),
            .I(N__2980));
    LocalMux I__329 (
            .O(N__2983),
            .I(\uart.r_Clock_Count_0 ));
    LocalMux I__328 (
            .O(N__2980),
            .I(\uart.r_Clock_Count_0 ));
    CascadeMux I__327 (
            .O(N__2975),
            .I(N__2971));
    InMux I__326 (
            .O(N__2974),
            .I(N__2968));
    InMux I__325 (
            .O(N__2971),
            .I(N__2965));
    LocalMux I__324 (
            .O(N__2968),
            .I(\uart.r_Clock_Count_1 ));
    LocalMux I__323 (
            .O(N__2965),
            .I(\uart.r_Clock_Count_1 ));
    InMux I__322 (
            .O(N__2960),
            .I(N__2956));
    InMux I__321 (
            .O(N__2959),
            .I(N__2953));
    LocalMux I__320 (
            .O(N__2956),
            .I(\uart.r_Clock_Count_3 ));
    LocalMux I__319 (
            .O(N__2953),
            .I(\uart.r_Clock_Count_3 ));
    InMux I__318 (
            .O(N__2948),
            .I(N__2944));
    InMux I__317 (
            .O(N__2947),
            .I(N__2941));
    LocalMux I__316 (
            .O(N__2944),
            .I(\uart.r_Clock_Count_5 ));
    LocalMux I__315 (
            .O(N__2941),
            .I(\uart.r_Clock_Count_5 ));
    InMux I__314 (
            .O(N__2936),
            .I(N__2932));
    InMux I__313 (
            .O(N__2935),
            .I(N__2929));
    LocalMux I__312 (
            .O(N__2932),
            .I(\uart.r_Clock_Count_4 ));
    LocalMux I__311 (
            .O(N__2929),
            .I(\uart.r_Clock_Count_4 ));
    CascadeMux I__310 (
            .O(N__2924),
            .I(\uart.n2006_cascade_ ));
    InMux I__309 (
            .O(N__2921),
            .I(N__2917));
    InMux I__308 (
            .O(N__2920),
            .I(N__2914));
    LocalMux I__307 (
            .O(N__2917),
            .I(\uart.r_Clock_Count_6 ));
    LocalMux I__306 (
            .O(N__2914),
            .I(\uart.r_Clock_Count_6 ));
    InMux I__305 (
            .O(N__2909),
            .I(N__2905));
    InMux I__304 (
            .O(N__2908),
            .I(N__2902));
    LocalMux I__303 (
            .O(N__2905),
            .I(\uart.r_Clock_Count_10 ));
    LocalMux I__302 (
            .O(N__2902),
            .I(\uart.r_Clock_Count_10 ));
    InMux I__301 (
            .O(N__2897),
            .I(N__2893));
    InMux I__300 (
            .O(N__2896),
            .I(N__2890));
    LocalMux I__299 (
            .O(N__2893),
            .I(\uart.r_Clock_Count_22 ));
    LocalMux I__298 (
            .O(N__2890),
            .I(\uart.r_Clock_Count_22 ));
    CascadeMux I__297 (
            .O(N__2885),
            .I(N__2882));
    InMux I__296 (
            .O(N__2882),
            .I(N__2879));
    LocalMux I__295 (
            .O(N__2879),
            .I(N__2875));
    InMux I__294 (
            .O(N__2878),
            .I(N__2872));
    Span4Mux_v I__293 (
            .O(N__2875),
            .I(N__2869));
    LocalMux I__292 (
            .O(N__2872),
            .I(\uart.r_Clock_Count_26 ));
    Odrv4 I__291 (
            .O(N__2869),
            .I(\uart.r_Clock_Count_26 ));
    InMux I__290 (
            .O(N__2864),
            .I(n2243));
    InMux I__289 (
            .O(N__2861),
            .I(n2244));
    InMux I__288 (
            .O(N__2858),
            .I(n2245));
    InMux I__287 (
            .O(N__2855),
            .I(n2246));
    InMux I__286 (
            .O(N__2852),
            .I(n2247));
    InMux I__285 (
            .O(N__2849),
            .I(n2248));
    InMux I__284 (
            .O(N__2846),
            .I(bfn_1_25_0_));
    InMux I__283 (
            .O(N__2843),
            .I(n2250));
    InMux I__282 (
            .O(N__2840),
            .I(n2251));
    InMux I__281 (
            .O(N__2837),
            .I(n2234));
    InMux I__280 (
            .O(N__2834),
            .I(n2235));
    InMux I__279 (
            .O(N__2831),
            .I(n2236));
    InMux I__278 (
            .O(N__2828),
            .I(n2237));
    InMux I__277 (
            .O(N__2825),
            .I(n2238));
    InMux I__276 (
            .O(N__2822),
            .I(n2239));
    InMux I__275 (
            .O(N__2819),
            .I(n2240));
    InMux I__274 (
            .O(N__2816),
            .I(bfn_1_24_0_));
    InMux I__273 (
            .O(N__2813),
            .I(n2242));
    InMux I__272 (
            .O(N__2810),
            .I(bfn_1_22_0_));
    InMux I__271 (
            .O(N__2807),
            .I(n2226));
    InMux I__270 (
            .O(N__2804),
            .I(n2227));
    InMux I__269 (
            .O(N__2801),
            .I(n2228));
    InMux I__268 (
            .O(N__2798),
            .I(n2229));
    InMux I__267 (
            .O(N__2795),
            .I(n2230));
    InMux I__266 (
            .O(N__2792),
            .I(n2231));
    InMux I__265 (
            .O(N__2789),
            .I(n2232));
    InMux I__264 (
            .O(N__2786),
            .I(bfn_1_23_0_));
    InMux I__263 (
            .O(N__2783),
            .I(\uart.n2154 ));
    InMux I__262 (
            .O(N__2780),
            .I(bfn_1_21_0_));
    InMux I__261 (
            .O(N__2777),
            .I(\uart.n2156 ));
    InMux I__260 (
            .O(N__2774),
            .I(\uart.n2157 ));
    InMux I__259 (
            .O(N__2771),
            .I(\uart.n2158 ));
    InMux I__258 (
            .O(N__2768),
            .I(\uart.n2159 ));
    InMux I__257 (
            .O(N__2765),
            .I(\uart.n2160 ));
    InMux I__256 (
            .O(N__2762),
            .I(\uart.n2161 ));
    InMux I__255 (
            .O(N__2759),
            .I(\uart.n2162 ));
    InMux I__254 (
            .O(N__2756),
            .I(\uart.n2145 ));
    InMux I__253 (
            .O(N__2753),
            .I(\uart.n2146 ));
    InMux I__252 (
            .O(N__2750),
            .I(bfn_1_20_0_));
    InMux I__251 (
            .O(N__2747),
            .I(\uart.n2148 ));
    InMux I__250 (
            .O(N__2744),
            .I(\uart.n2149 ));
    InMux I__249 (
            .O(N__2741),
            .I(\uart.n2150 ));
    InMux I__248 (
            .O(N__2738),
            .I(\uart.n2151 ));
    InMux I__247 (
            .O(N__2735),
            .I(\uart.n2152 ));
    InMux I__246 (
            .O(N__2732),
            .I(\uart.n2153 ));
    InMux I__245 (
            .O(N__2729),
            .I(\uart.n2135 ));
    InMux I__244 (
            .O(N__2726),
            .I(\uart.n2136 ));
    InMux I__243 (
            .O(N__2723),
            .I(\uart.n2137 ));
    InMux I__242 (
            .O(N__2720),
            .I(\uart.n2138 ));
    InMux I__241 (
            .O(N__2717),
            .I(bfn_1_19_0_));
    InMux I__240 (
            .O(N__2714),
            .I(\uart.n2140 ));
    InMux I__239 (
            .O(N__2711),
            .I(\uart.n2141 ));
    InMux I__238 (
            .O(N__2708),
            .I(\uart.n2142 ));
    InMux I__237 (
            .O(N__2705),
            .I(\uart.n2143 ));
    InMux I__236 (
            .O(N__2702),
            .I(\uart.n2144 ));
    IoInMux I__235 (
            .O(N__2699),
            .I(N__2696));
    LocalMux I__234 (
            .O(N__2696),
            .I(N__2693));
    IoSpan4Mux I__233 (
            .O(N__2693),
            .I(N__2690));
    IoSpan4Mux I__232 (
            .O(N__2690),
            .I(N__2687));
    IoSpan4Mux I__231 (
            .O(N__2687),
            .I(N__2684));
    Odrv4 I__230 (
            .O(N__2684),
            .I(CLK_pad_gb_input));
    InMux I__229 (
            .O(N__2681),
            .I(bfn_1_18_0_));
    InMux I__228 (
            .O(N__2678),
            .I(\uart.n2132 ));
    InMux I__227 (
            .O(N__2675),
            .I(\uart.n2133 ));
    InMux I__226 (
            .O(N__2672),
            .I(\uart.n2134 ));
    defparam IN_MUX_bfv_1_18_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_18_0_ (
            .carryinitin(),
            .carryinitout(bfn_1_18_0_));
    defparam IN_MUX_bfv_1_19_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_19_0_ (
            .carryinitin(\uart.n2139 ),
            .carryinitout(bfn_1_19_0_));
    defparam IN_MUX_bfv_1_20_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_20_0_ (
            .carryinitin(\uart.n2147 ),
            .carryinitout(bfn_1_20_0_));
    defparam IN_MUX_bfv_1_21_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_21_0_ (
            .carryinitin(\uart.n2155 ),
            .carryinitout(bfn_1_21_0_));
    defparam IN_MUX_bfv_5_23_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_5_23_0_ (
            .carryinitin(),
            .carryinitout(bfn_5_23_0_));
    defparam IN_MUX_bfv_3_22_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_3_22_0_ (
            .carryinitin(),
            .carryinitout(bfn_3_22_0_));
    defparam IN_MUX_bfv_3_23_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_3_23_0_ (
            .carryinitin(n2202),
            .carryinitout(bfn_3_23_0_));
    defparam IN_MUX_bfv_3_24_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_3_24_0_ (
            .carryinitin(n2210),
            .carryinitout(bfn_3_24_0_));
    defparam IN_MUX_bfv_3_25_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_3_25_0_ (
            .carryinitin(n2218),
            .carryinitout(bfn_3_25_0_));
    defparam IN_MUX_bfv_1_22_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_22_0_ (
            .carryinitin(),
            .carryinitout(bfn_1_22_0_));
    defparam IN_MUX_bfv_1_23_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_23_0_ (
            .carryinitin(n2233),
            .carryinitout(bfn_1_23_0_));
    defparam IN_MUX_bfv_1_24_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_24_0_ (
            .carryinitin(n2241),
            .carryinitout(bfn_1_24_0_));
    defparam IN_MUX_bfv_1_25_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_25_0_ (
            .carryinitin(n2249),
            .carryinitout(bfn_1_25_0_));
    defparam IN_MUX_bfv_2_23_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_23_0_ (
            .carryinitin(),
            .carryinitout(bfn_2_23_0_));
    defparam IN_MUX_bfv_2_24_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_24_0_ (
            .carryinitin(n2170),
            .carryinitout(bfn_2_24_0_));
    defparam IN_MUX_bfv_2_25_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_25_0_ (
            .carryinitin(n2178),
            .carryinitout(bfn_2_25_0_));
    defparam IN_MUX_bfv_2_26_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_26_0_ (
            .carryinitin(n2186),
            .carryinitout(bfn_2_26_0_));
    ICE_GB CLK_pad_gb (
            .USERSIGNALTOGLOBALBUFFER(N__2699),
            .GLOBALBUFFEROUTPUT(CLK_c));
    VCC VCC (
            .Y(VCCG0));
    GND GND (
            .Y(GNDG0));
    GND GND_Inst (
            .Y(_gnd_net_));
    defparam \uart.r_Clock_Count_121__i0_LC_1_18_0 .C_ON=1'b1;
    defparam \uart.r_Clock_Count_121__i0_LC_1_18_0 .SEQ_MODE=4'b1000;
    defparam \uart.r_Clock_Count_121__i0_LC_1_18_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \uart.r_Clock_Count_121__i0_LC_1_18_0  (
            .in0(_gnd_net_),
            .in1(N__2986),
            .in2(_gnd_net_),
            .in3(N__2681),
            .lcout(\uart.r_Clock_Count_0 ),
            .ltout(),
            .carryin(bfn_1_18_0_),
            .carryout(\uart.n2132 ),
            .clk(N__5379),
            .ce(N__3106),
            .sr(N__3216));
    defparam \uart.r_Clock_Count_121__i1_LC_1_18_1 .C_ON=1'b1;
    defparam \uart.r_Clock_Count_121__i1_LC_1_18_1 .SEQ_MODE=4'b1000;
    defparam \uart.r_Clock_Count_121__i1_LC_1_18_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \uart.r_Clock_Count_121__i1_LC_1_18_1  (
            .in0(_gnd_net_),
            .in1(N__2974),
            .in2(_gnd_net_),
            .in3(N__2678),
            .lcout(\uart.r_Clock_Count_1 ),
            .ltout(),
            .carryin(\uart.n2132 ),
            .carryout(\uart.n2133 ),
            .clk(N__5379),
            .ce(N__3106),
            .sr(N__3216));
    defparam \uart.r_Clock_Count_121__i2_LC_1_18_2 .C_ON=1'b1;
    defparam \uart.r_Clock_Count_121__i2_LC_1_18_2 .SEQ_MODE=4'b1000;
    defparam \uart.r_Clock_Count_121__i2_LC_1_18_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \uart.r_Clock_Count_121__i2_LC_1_18_2  (
            .in0(_gnd_net_),
            .in1(N__2998),
            .in2(_gnd_net_),
            .in3(N__2675),
            .lcout(\uart.r_Clock_Count_2 ),
            .ltout(),
            .carryin(\uart.n2133 ),
            .carryout(\uart.n2134 ),
            .clk(N__5379),
            .ce(N__3106),
            .sr(N__3216));
    defparam \uart.r_Clock_Count_121__i3_LC_1_18_3 .C_ON=1'b1;
    defparam \uart.r_Clock_Count_121__i3_LC_1_18_3 .SEQ_MODE=4'b1000;
    defparam \uart.r_Clock_Count_121__i3_LC_1_18_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \uart.r_Clock_Count_121__i3_LC_1_18_3  (
            .in0(_gnd_net_),
            .in1(N__2960),
            .in2(_gnd_net_),
            .in3(N__2672),
            .lcout(\uart.r_Clock_Count_3 ),
            .ltout(),
            .carryin(\uart.n2134 ),
            .carryout(\uart.n2135 ),
            .clk(N__5379),
            .ce(N__3106),
            .sr(N__3216));
    defparam \uart.r_Clock_Count_121__i4_LC_1_18_4 .C_ON=1'b1;
    defparam \uart.r_Clock_Count_121__i4_LC_1_18_4 .SEQ_MODE=4'b1000;
    defparam \uart.r_Clock_Count_121__i4_LC_1_18_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \uart.r_Clock_Count_121__i4_LC_1_18_4  (
            .in0(_gnd_net_),
            .in1(N__2936),
            .in2(_gnd_net_),
            .in3(N__2729),
            .lcout(\uart.r_Clock_Count_4 ),
            .ltout(),
            .carryin(\uart.n2135 ),
            .carryout(\uart.n2136 ),
            .clk(N__5379),
            .ce(N__3106),
            .sr(N__3216));
    defparam \uart.r_Clock_Count_121__i5_LC_1_18_5 .C_ON=1'b1;
    defparam \uart.r_Clock_Count_121__i5_LC_1_18_5 .SEQ_MODE=4'b1000;
    defparam \uart.r_Clock_Count_121__i5_LC_1_18_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \uart.r_Clock_Count_121__i5_LC_1_18_5  (
            .in0(_gnd_net_),
            .in1(N__2948),
            .in2(_gnd_net_),
            .in3(N__2726),
            .lcout(\uart.r_Clock_Count_5 ),
            .ltout(),
            .carryin(\uart.n2136 ),
            .carryout(\uart.n2137 ),
            .clk(N__5379),
            .ce(N__3106),
            .sr(N__3216));
    defparam \uart.r_Clock_Count_121__i6_LC_1_18_6 .C_ON=1'b1;
    defparam \uart.r_Clock_Count_121__i6_LC_1_18_6 .SEQ_MODE=4'b1000;
    defparam \uart.r_Clock_Count_121__i6_LC_1_18_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \uart.r_Clock_Count_121__i6_LC_1_18_6  (
            .in0(_gnd_net_),
            .in1(N__2921),
            .in2(_gnd_net_),
            .in3(N__2723),
            .lcout(\uart.r_Clock_Count_6 ),
            .ltout(),
            .carryin(\uart.n2137 ),
            .carryout(\uart.n2138 ),
            .clk(N__5379),
            .ce(N__3106),
            .sr(N__3216));
    defparam \uart.r_Clock_Count_121__i7_LC_1_18_7 .C_ON=1'b1;
    defparam \uart.r_Clock_Count_121__i7_LC_1_18_7 .SEQ_MODE=4'b1000;
    defparam \uart.r_Clock_Count_121__i7_LC_1_18_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \uart.r_Clock_Count_121__i7_LC_1_18_7  (
            .in0(_gnd_net_),
            .in1(N__3248),
            .in2(_gnd_net_),
            .in3(N__2720),
            .lcout(\uart.r_Clock_Count_7 ),
            .ltout(),
            .carryin(\uart.n2138 ),
            .carryout(\uart.n2139 ),
            .clk(N__5379),
            .ce(N__3106),
            .sr(N__3216));
    defparam \uart.r_Clock_Count_121__i8_LC_1_19_0 .C_ON=1'b1;
    defparam \uart.r_Clock_Count_121__i8_LC_1_19_0 .SEQ_MODE=4'b1000;
    defparam \uart.r_Clock_Count_121__i8_LC_1_19_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \uart.r_Clock_Count_121__i8_LC_1_19_0  (
            .in0(_gnd_net_),
            .in1(N__3193),
            .in2(_gnd_net_),
            .in3(N__2717),
            .lcout(\uart.r_Clock_Count_8 ),
            .ltout(),
            .carryin(bfn_1_19_0_),
            .carryout(\uart.n2140 ),
            .clk(N__5380),
            .ce(N__3095),
            .sr(N__3215));
    defparam \uart.r_Clock_Count_121__i9_LC_1_19_1 .C_ON=1'b1;
    defparam \uart.r_Clock_Count_121__i9_LC_1_19_1 .SEQ_MODE=4'b1000;
    defparam \uart.r_Clock_Count_121__i9_LC_1_19_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \uart.r_Clock_Count_121__i9_LC_1_19_1  (
            .in0(_gnd_net_),
            .in1(N__3605),
            .in2(_gnd_net_),
            .in3(N__2714),
            .lcout(\uart.r_Clock_Count_9 ),
            .ltout(),
            .carryin(\uart.n2140 ),
            .carryout(\uart.n2141 ),
            .clk(N__5380),
            .ce(N__3095),
            .sr(N__3215));
    defparam \uart.r_Clock_Count_121__i10_LC_1_19_2 .C_ON=1'b1;
    defparam \uart.r_Clock_Count_121__i10_LC_1_19_2 .SEQ_MODE=4'b1000;
    defparam \uart.r_Clock_Count_121__i10_LC_1_19_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \uart.r_Clock_Count_121__i10_LC_1_19_2  (
            .in0(_gnd_net_),
            .in1(N__2909),
            .in2(_gnd_net_),
            .in3(N__2711),
            .lcout(\uart.r_Clock_Count_10 ),
            .ltout(),
            .carryin(\uart.n2141 ),
            .carryout(\uart.n2142 ),
            .clk(N__5380),
            .ce(N__3095),
            .sr(N__3215));
    defparam \uart.r_Clock_Count_121__i11_LC_1_19_3 .C_ON=1'b1;
    defparam \uart.r_Clock_Count_121__i11_LC_1_19_3 .SEQ_MODE=4'b1000;
    defparam \uart.r_Clock_Count_121__i11_LC_1_19_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \uart.r_Clock_Count_121__i11_LC_1_19_3  (
            .in0(_gnd_net_),
            .in1(N__3065),
            .in2(_gnd_net_),
            .in3(N__2708),
            .lcout(\uart.r_Clock_Count_11 ),
            .ltout(),
            .carryin(\uart.n2142 ),
            .carryout(\uart.n2143 ),
            .clk(N__5380),
            .ce(N__3095),
            .sr(N__3215));
    defparam \uart.r_Clock_Count_121__i12_LC_1_19_4 .C_ON=1'b1;
    defparam \uart.r_Clock_Count_121__i12_LC_1_19_4 .SEQ_MODE=4'b1000;
    defparam \uart.r_Clock_Count_121__i12_LC_1_19_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \uart.r_Clock_Count_121__i12_LC_1_19_4  (
            .in0(_gnd_net_),
            .in1(N__3278),
            .in2(_gnd_net_),
            .in3(N__2705),
            .lcout(\uart.r_Clock_Count_12 ),
            .ltout(),
            .carryin(\uart.n2143 ),
            .carryout(\uart.n2144 ),
            .clk(N__5380),
            .ce(N__3095),
            .sr(N__3215));
    defparam \uart.r_Clock_Count_121__i13_LC_1_19_5 .C_ON=1'b1;
    defparam \uart.r_Clock_Count_121__i13_LC_1_19_5 .SEQ_MODE=4'b1000;
    defparam \uart.r_Clock_Count_121__i13_LC_1_19_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \uart.r_Clock_Count_121__i13_LC_1_19_5  (
            .in0(_gnd_net_),
            .in1(N__3290),
            .in2(_gnd_net_),
            .in3(N__2702),
            .lcout(\uart.r_Clock_Count_13 ),
            .ltout(),
            .carryin(\uart.n2144 ),
            .carryout(\uart.n2145 ),
            .clk(N__5380),
            .ce(N__3095),
            .sr(N__3215));
    defparam \uart.r_Clock_Count_121__i14_LC_1_19_6 .C_ON=1'b1;
    defparam \uart.r_Clock_Count_121__i14_LC_1_19_6 .SEQ_MODE=4'b1000;
    defparam \uart.r_Clock_Count_121__i14_LC_1_19_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \uart.r_Clock_Count_121__i14_LC_1_19_6  (
            .in0(_gnd_net_),
            .in1(N__3179),
            .in2(_gnd_net_),
            .in3(N__2756),
            .lcout(\uart.r_Clock_Count_14 ),
            .ltout(),
            .carryin(\uart.n2145 ),
            .carryout(\uart.n2146 ),
            .clk(N__5380),
            .ce(N__3095),
            .sr(N__3215));
    defparam \uart.r_Clock_Count_121__i15_LC_1_19_7 .C_ON=1'b1;
    defparam \uart.r_Clock_Count_121__i15_LC_1_19_7 .SEQ_MODE=4'b1000;
    defparam \uart.r_Clock_Count_121__i15_LC_1_19_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \uart.r_Clock_Count_121__i15_LC_1_19_7  (
            .in0(_gnd_net_),
            .in1(N__3632),
            .in2(_gnd_net_),
            .in3(N__2753),
            .lcout(\uart.r_Clock_Count_15 ),
            .ltout(),
            .carryin(\uart.n2146 ),
            .carryout(\uart.n2147 ),
            .clk(N__5380),
            .ce(N__3095),
            .sr(N__3215));
    defparam \uart.r_Clock_Count_121__i16_LC_1_20_0 .C_ON=1'b1;
    defparam \uart.r_Clock_Count_121__i16_LC_1_20_0 .SEQ_MODE=4'b1000;
    defparam \uart.r_Clock_Count_121__i16_LC_1_20_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \uart.r_Clock_Count_121__i16_LC_1_20_0  (
            .in0(_gnd_net_),
            .in1(N__3565),
            .in2(_gnd_net_),
            .in3(N__2750),
            .lcout(\uart.r_Clock_Count_16 ),
            .ltout(),
            .carryin(bfn_1_20_0_),
            .carryout(\uart.n2148 ),
            .clk(N__5381),
            .ce(N__3094),
            .sr(N__3217));
    defparam \uart.r_Clock_Count_121__i17_LC_1_20_1 .C_ON=1'b1;
    defparam \uart.r_Clock_Count_121__i17_LC_1_20_1 .SEQ_MODE=4'b1000;
    defparam \uart.r_Clock_Count_121__i17_LC_1_20_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \uart.r_Clock_Count_121__i17_LC_1_20_1  (
            .in0(_gnd_net_),
            .in1(N__3040),
            .in2(_gnd_net_),
            .in3(N__2747),
            .lcout(\uart.r_Clock_Count_17 ),
            .ltout(),
            .carryin(\uart.n2148 ),
            .carryout(\uart.n2149 ),
            .clk(N__5381),
            .ce(N__3094),
            .sr(N__3217));
    defparam \uart.r_Clock_Count_121__i18_LC_1_20_2 .C_ON=1'b1;
    defparam \uart.r_Clock_Count_121__i18_LC_1_20_2 .SEQ_MODE=4'b1000;
    defparam \uart.r_Clock_Count_121__i18_LC_1_20_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \uart.r_Clock_Count_121__i18_LC_1_20_2  (
            .in0(_gnd_net_),
            .in1(N__3026),
            .in2(_gnd_net_),
            .in3(N__2744),
            .lcout(\uart.r_Clock_Count_18 ),
            .ltout(),
            .carryin(\uart.n2149 ),
            .carryout(\uart.n2150 ),
            .clk(N__5381),
            .ce(N__3094),
            .sr(N__3217));
    defparam \uart.r_Clock_Count_121__i19_LC_1_20_3 .C_ON=1'b1;
    defparam \uart.r_Clock_Count_121__i19_LC_1_20_3 .SEQ_MODE=4'b1000;
    defparam \uart.r_Clock_Count_121__i19_LC_1_20_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \uart.r_Clock_Count_121__i19_LC_1_20_3  (
            .in0(_gnd_net_),
            .in1(N__3578),
            .in2(_gnd_net_),
            .in3(N__2741),
            .lcout(\uart.r_Clock_Count_19 ),
            .ltout(),
            .carryin(\uart.n2150 ),
            .carryout(\uart.n2151 ),
            .clk(N__5381),
            .ce(N__3094),
            .sr(N__3217));
    defparam \uart.r_Clock_Count_121__i20_LC_1_20_4 .C_ON=1'b1;
    defparam \uart.r_Clock_Count_121__i20_LC_1_20_4 .SEQ_MODE=4'b1000;
    defparam \uart.r_Clock_Count_121__i20_LC_1_20_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \uart.r_Clock_Count_121__i20_LC_1_20_4  (
            .in0(_gnd_net_),
            .in1(N__3644),
            .in2(_gnd_net_),
            .in3(N__2738),
            .lcout(\uart.r_Clock_Count_20 ),
            .ltout(),
            .carryin(\uart.n2151 ),
            .carryout(\uart.n2152 ),
            .clk(N__5381),
            .ce(N__3094),
            .sr(N__3217));
    defparam \uart.r_Clock_Count_121__i21_LC_1_20_5 .C_ON=1'b1;
    defparam \uart.r_Clock_Count_121__i21_LC_1_20_5 .SEQ_MODE=4'b1000;
    defparam \uart.r_Clock_Count_121__i21_LC_1_20_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \uart.r_Clock_Count_121__i21_LC_1_20_5  (
            .in0(_gnd_net_),
            .in1(N__3053),
            .in2(_gnd_net_),
            .in3(N__2735),
            .lcout(\uart.r_Clock_Count_21 ),
            .ltout(),
            .carryin(\uart.n2152 ),
            .carryout(\uart.n2153 ),
            .clk(N__5381),
            .ce(N__3094),
            .sr(N__3217));
    defparam \uart.r_Clock_Count_121__i22_LC_1_20_6 .C_ON=1'b1;
    defparam \uart.r_Clock_Count_121__i22_LC_1_20_6 .SEQ_MODE=4'b1000;
    defparam \uart.r_Clock_Count_121__i22_LC_1_20_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \uart.r_Clock_Count_121__i22_LC_1_20_6  (
            .in0(_gnd_net_),
            .in1(N__2897),
            .in2(_gnd_net_),
            .in3(N__2732),
            .lcout(\uart.r_Clock_Count_22 ),
            .ltout(),
            .carryin(\uart.n2153 ),
            .carryout(\uart.n2154 ),
            .clk(N__5381),
            .ce(N__3094),
            .sr(N__3217));
    defparam \uart.r_Clock_Count_121__i23_LC_1_20_7 .C_ON=1'b1;
    defparam \uart.r_Clock_Count_121__i23_LC_1_20_7 .SEQ_MODE=4'b1000;
    defparam \uart.r_Clock_Count_121__i23_LC_1_20_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \uart.r_Clock_Count_121__i23_LC_1_20_7  (
            .in0(_gnd_net_),
            .in1(N__3119),
            .in2(_gnd_net_),
            .in3(N__2783),
            .lcout(\uart.r_Clock_Count_23 ),
            .ltout(),
            .carryin(\uart.n2154 ),
            .carryout(\uart.n2155 ),
            .clk(N__5381),
            .ce(N__3094),
            .sr(N__3217));
    defparam \uart.r_Clock_Count_121__i24_LC_1_21_0 .C_ON=1'b1;
    defparam \uart.r_Clock_Count_121__i24_LC_1_21_0 .SEQ_MODE=4'b1000;
    defparam \uart.r_Clock_Count_121__i24_LC_1_21_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \uart.r_Clock_Count_121__i24_LC_1_21_0  (
            .in0(_gnd_net_),
            .in1(N__3133),
            .in2(_gnd_net_),
            .in3(N__2780),
            .lcout(\uart.r_Clock_Count_24 ),
            .ltout(),
            .carryin(bfn_1_21_0_),
            .carryout(\uart.n2156 ),
            .clk(N__5383),
            .ce(N__3096),
            .sr(N__3224));
    defparam \uart.r_Clock_Count_121__i25_LC_1_21_1 .C_ON=1'b1;
    defparam \uart.r_Clock_Count_121__i25_LC_1_21_1 .SEQ_MODE=4'b1000;
    defparam \uart.r_Clock_Count_121__i25_LC_1_21_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \uart.r_Clock_Count_121__i25_LC_1_21_1  (
            .in0(_gnd_net_),
            .in1(N__3619),
            .in2(_gnd_net_),
            .in3(N__2777),
            .lcout(\uart.r_Clock_Count_25 ),
            .ltout(),
            .carryin(\uart.n2156 ),
            .carryout(\uart.n2157 ),
            .clk(N__5383),
            .ce(N__3096),
            .sr(N__3224));
    defparam \uart.r_Clock_Count_121__i26_LC_1_21_2 .C_ON=1'b1;
    defparam \uart.r_Clock_Count_121__i26_LC_1_21_2 .SEQ_MODE=4'b1000;
    defparam \uart.r_Clock_Count_121__i26_LC_1_21_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \uart.r_Clock_Count_121__i26_LC_1_21_2  (
            .in0(_gnd_net_),
            .in1(N__2878),
            .in2(_gnd_net_),
            .in3(N__2774),
            .lcout(\uart.r_Clock_Count_26 ),
            .ltout(),
            .carryin(\uart.n2157 ),
            .carryout(\uart.n2158 ),
            .clk(N__5383),
            .ce(N__3096),
            .sr(N__3224));
    defparam \uart.r_Clock_Count_121__i27_LC_1_21_3 .C_ON=1'b1;
    defparam \uart.r_Clock_Count_121__i27_LC_1_21_3 .SEQ_MODE=4'b1000;
    defparam \uart.r_Clock_Count_121__i27_LC_1_21_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \uart.r_Clock_Count_121__i27_LC_1_21_3  (
            .in0(_gnd_net_),
            .in1(N__3592),
            .in2(_gnd_net_),
            .in3(N__2771),
            .lcout(\uart.r_Clock_Count_27 ),
            .ltout(),
            .carryin(\uart.n2158 ),
            .carryout(\uart.n2159 ),
            .clk(N__5383),
            .ce(N__3096),
            .sr(N__3224));
    defparam \uart.r_Clock_Count_121__i28_LC_1_21_4 .C_ON=1'b1;
    defparam \uart.r_Clock_Count_121__i28_LC_1_21_4 .SEQ_MODE=4'b1000;
    defparam \uart.r_Clock_Count_121__i28_LC_1_21_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \uart.r_Clock_Count_121__i28_LC_1_21_4  (
            .in0(_gnd_net_),
            .in1(N__3149),
            .in2(_gnd_net_),
            .in3(N__2768),
            .lcout(\uart.r_Clock_Count_28 ),
            .ltout(),
            .carryin(\uart.n2159 ),
            .carryout(\uart.n2160 ),
            .clk(N__5383),
            .ce(N__3096),
            .sr(N__3224));
    defparam \uart.r_Clock_Count_121__i29_LC_1_21_5 .C_ON=1'b1;
    defparam \uart.r_Clock_Count_121__i29_LC_1_21_5 .SEQ_MODE=4'b1000;
    defparam \uart.r_Clock_Count_121__i29_LC_1_21_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \uart.r_Clock_Count_121__i29_LC_1_21_5  (
            .in0(_gnd_net_),
            .in1(N__3265),
            .in2(_gnd_net_),
            .in3(N__2765),
            .lcout(\uart.r_Clock_Count_29 ),
            .ltout(),
            .carryin(\uart.n2160 ),
            .carryout(\uart.n2161 ),
            .clk(N__5383),
            .ce(N__3096),
            .sr(N__3224));
    defparam \uart.r_Clock_Count_121__i30_LC_1_21_6 .C_ON=1'b1;
    defparam \uart.r_Clock_Count_121__i30_LC_1_21_6 .SEQ_MODE=4'b1000;
    defparam \uart.r_Clock_Count_121__i30_LC_1_21_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \uart.r_Clock_Count_121__i30_LC_1_21_6  (
            .in0(_gnd_net_),
            .in1(N__3161),
            .in2(_gnd_net_),
            .in3(N__2762),
            .lcout(\uart.r_Clock_Count_30 ),
            .ltout(),
            .carryin(\uart.n2161 ),
            .carryout(\uart.n2162 ),
            .clk(N__5383),
            .ce(N__3096),
            .sr(N__3224));
    defparam \uart.r_Clock_Count_121__i31_LC_1_21_7 .C_ON=1'b0;
    defparam \uart.r_Clock_Count_121__i31_LC_1_21_7 .SEQ_MODE=4'b1000;
    defparam \uart.r_Clock_Count_121__i31_LC_1_21_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \uart.r_Clock_Count_121__i31_LC_1_21_7  (
            .in0(_gnd_net_),
            .in1(N__3551),
            .in2(_gnd_net_),
            .in3(N__2759),
            .lcout(\uart.r_Clock_Count_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__5383),
            .ce(N__3096),
            .sr(N__3224));
    defparam clk_divider_116__i0_LC_1_22_0.C_ON=1'b1;
    defparam clk_divider_116__i0_LC_1_22_0.SEQ_MODE=4'b1000;
    defparam clk_divider_116__i0_LC_1_22_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 clk_divider_116__i0_LC_1_22_0 (
            .in0(_gnd_net_),
            .in1(N__3974),
            .in2(_gnd_net_),
            .in3(N__2810),
            .lcout(clk_divider_0),
            .ltout(),
            .carryin(bfn_1_22_0_),
            .carryout(n2226),
            .clk(N__5385),
            .ce(),
            .sr(N__3938));
    defparam clk_divider_116__i1_LC_1_22_1.C_ON=1'b1;
    defparam clk_divider_116__i1_LC_1_22_1.SEQ_MODE=4'b1000;
    defparam clk_divider_116__i1_LC_1_22_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 clk_divider_116__i1_LC_1_22_1 (
            .in0(_gnd_net_),
            .in1(N__3899),
            .in2(_gnd_net_),
            .in3(N__2807),
            .lcout(clk_divider_1),
            .ltout(),
            .carryin(n2226),
            .carryout(n2227),
            .clk(N__5385),
            .ce(),
            .sr(N__3938));
    defparam clk_divider_116__i2_LC_1_22_2.C_ON=1'b1;
    defparam clk_divider_116__i2_LC_1_22_2.SEQ_MODE=4'b1000;
    defparam clk_divider_116__i2_LC_1_22_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 clk_divider_116__i2_LC_1_22_2 (
            .in0(_gnd_net_),
            .in1(N__3887),
            .in2(_gnd_net_),
            .in3(N__2804),
            .lcout(clk_divider_2),
            .ltout(),
            .carryin(n2227),
            .carryout(n2228),
            .clk(N__5385),
            .ce(),
            .sr(N__3938));
    defparam clk_divider_116__i3_LC_1_22_3.C_ON=1'b1;
    defparam clk_divider_116__i3_LC_1_22_3.SEQ_MODE=4'b1000;
    defparam clk_divider_116__i3_LC_1_22_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 clk_divider_116__i3_LC_1_22_3 (
            .in0(_gnd_net_),
            .in1(N__3961),
            .in2(_gnd_net_),
            .in3(N__2801),
            .lcout(clk_divider_3),
            .ltout(),
            .carryin(n2228),
            .carryout(n2229),
            .clk(N__5385),
            .ce(),
            .sr(N__3938));
    defparam clk_divider_116__i4_LC_1_22_4.C_ON=1'b1;
    defparam clk_divider_116__i4_LC_1_22_4.SEQ_MODE=4'b1000;
    defparam clk_divider_116__i4_LC_1_22_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 clk_divider_116__i4_LC_1_22_4 (
            .in0(_gnd_net_),
            .in1(N__3988),
            .in2(_gnd_net_),
            .in3(N__2798),
            .lcout(clk_divider_4),
            .ltout(),
            .carryin(n2229),
            .carryout(n2230),
            .clk(N__5385),
            .ce(),
            .sr(N__3938));
    defparam clk_divider_116__i5_LC_1_22_5.C_ON=1'b1;
    defparam clk_divider_116__i5_LC_1_22_5.SEQ_MODE=4'b1000;
    defparam clk_divider_116__i5_LC_1_22_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 clk_divider_116__i5_LC_1_22_5 (
            .in0(_gnd_net_),
            .in1(N__3815),
            .in2(_gnd_net_),
            .in3(N__2795),
            .lcout(clk_divider_5),
            .ltout(),
            .carryin(n2230),
            .carryout(n2231),
            .clk(N__5385),
            .ce(),
            .sr(N__3938));
    defparam clk_divider_116__i6_LC_1_22_6.C_ON=1'b1;
    defparam clk_divider_116__i6_LC_1_22_6.SEQ_MODE=4'b1000;
    defparam clk_divider_116__i6_LC_1_22_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 clk_divider_116__i6_LC_1_22_6 (
            .in0(_gnd_net_),
            .in1(N__3386),
            .in2(_gnd_net_),
            .in3(N__2792),
            .lcout(clk_divider_6),
            .ltout(),
            .carryin(n2231),
            .carryout(n2232),
            .clk(N__5385),
            .ce(),
            .sr(N__3938));
    defparam clk_divider_116__i7_LC_1_22_7.C_ON=1'b1;
    defparam clk_divider_116__i7_LC_1_22_7.SEQ_MODE=4'b1000;
    defparam clk_divider_116__i7_LC_1_22_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 clk_divider_116__i7_LC_1_22_7 (
            .in0(_gnd_net_),
            .in1(N__4246),
            .in2(_gnd_net_),
            .in3(N__2789),
            .lcout(clk_divider_7),
            .ltout(),
            .carryin(n2232),
            .carryout(n2233),
            .clk(N__5385),
            .ce(),
            .sr(N__3938));
    defparam clk_divider_116__i8_LC_1_23_0.C_ON=1'b1;
    defparam clk_divider_116__i8_LC_1_23_0.SEQ_MODE=4'b1000;
    defparam clk_divider_116__i8_LC_1_23_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 clk_divider_116__i8_LC_1_23_0 (
            .in0(_gnd_net_),
            .in1(N__3869),
            .in2(_gnd_net_),
            .in3(N__2786),
            .lcout(clk_divider_8),
            .ltout(),
            .carryin(bfn_1_23_0_),
            .carryout(n2234),
            .clk(N__5388),
            .ce(),
            .sr(N__3942));
    defparam clk_divider_116__i9_LC_1_23_1.C_ON=1'b1;
    defparam clk_divider_116__i9_LC_1_23_1.SEQ_MODE=4'b1000;
    defparam clk_divider_116__i9_LC_1_23_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 clk_divider_116__i9_LC_1_23_1 (
            .in0(_gnd_net_),
            .in1(N__3490),
            .in2(_gnd_net_),
            .in3(N__2837),
            .lcout(clk_divider_9),
            .ltout(),
            .carryin(n2234),
            .carryout(n2235),
            .clk(N__5388),
            .ce(),
            .sr(N__3942));
    defparam clk_divider_116__i10_LC_1_23_2.C_ON=1'b1;
    defparam clk_divider_116__i10_LC_1_23_2.SEQ_MODE=4'b1000;
    defparam clk_divider_116__i10_LC_1_23_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 clk_divider_116__i10_LC_1_23_2 (
            .in0(_gnd_net_),
            .in1(N__3803),
            .in2(_gnd_net_),
            .in3(N__2834),
            .lcout(clk_divider_10),
            .ltout(),
            .carryin(n2235),
            .carryout(n2236),
            .clk(N__5388),
            .ce(),
            .sr(N__3942));
    defparam clk_divider_116__i11_LC_1_23_3.C_ON=1'b1;
    defparam clk_divider_116__i11_LC_1_23_3.SEQ_MODE=4'b1000;
    defparam clk_divider_116__i11_LC_1_23_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 clk_divider_116__i11_LC_1_23_3 (
            .in0(_gnd_net_),
            .in1(N__3827),
            .in2(_gnd_net_),
            .in3(N__2831),
            .lcout(clk_divider_11),
            .ltout(),
            .carryin(n2236),
            .carryout(n2237),
            .clk(N__5388),
            .ce(),
            .sr(N__3942));
    defparam clk_divider_116__i12_LC_1_23_4.C_ON=1'b1;
    defparam clk_divider_116__i12_LC_1_23_4.SEQ_MODE=4'b1000;
    defparam clk_divider_116__i12_LC_1_23_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 clk_divider_116__i12_LC_1_23_4 (
            .in0(_gnd_net_),
            .in1(N__3790),
            .in2(_gnd_net_),
            .in3(N__2828),
            .lcout(clk_divider_12),
            .ltout(),
            .carryin(n2237),
            .carryout(n2238),
            .clk(N__5388),
            .ce(),
            .sr(N__3942));
    defparam clk_divider_116__i13_LC_1_23_5.C_ON=1'b1;
    defparam clk_divider_116__i13_LC_1_23_5.SEQ_MODE=4'b1000;
    defparam clk_divider_116__i13_LC_1_23_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 clk_divider_116__i13_LC_1_23_5 (
            .in0(_gnd_net_),
            .in1(N__3761),
            .in2(_gnd_net_),
            .in3(N__2825),
            .lcout(clk_divider_13),
            .ltout(),
            .carryin(n2238),
            .carryout(n2239),
            .clk(N__5388),
            .ce(),
            .sr(N__3942));
    defparam clk_divider_116__i14_LC_1_23_6.C_ON=1'b1;
    defparam clk_divider_116__i14_LC_1_23_6.SEQ_MODE=4'b1000;
    defparam clk_divider_116__i14_LC_1_23_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 clk_divider_116__i14_LC_1_23_6 (
            .in0(_gnd_net_),
            .in1(N__3472),
            .in2(_gnd_net_),
            .in3(N__2822),
            .lcout(clk_divider_14),
            .ltout(),
            .carryin(n2239),
            .carryout(n2240),
            .clk(N__5388),
            .ce(),
            .sr(N__3942));
    defparam clk_divider_116__i15_LC_1_23_7.C_ON=1'b1;
    defparam clk_divider_116__i15_LC_1_23_7.SEQ_MODE=4'b1000;
    defparam clk_divider_116__i15_LC_1_23_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 clk_divider_116__i15_LC_1_23_7 (
            .in0(_gnd_net_),
            .in1(N__3857),
            .in2(_gnd_net_),
            .in3(N__2819),
            .lcout(clk_divider_15),
            .ltout(),
            .carryin(n2240),
            .carryout(n2241),
            .clk(N__5388),
            .ce(),
            .sr(N__3942));
    defparam clk_divider_116__i16_LC_1_24_0.C_ON=1'b1;
    defparam clk_divider_116__i16_LC_1_24_0.SEQ_MODE=4'b1000;
    defparam clk_divider_116__i16_LC_1_24_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 clk_divider_116__i16_LC_1_24_0 (
            .in0(_gnd_net_),
            .in1(N__3712),
            .in2(_gnd_net_),
            .in3(N__2816),
            .lcout(clk_divider_16),
            .ltout(),
            .carryin(bfn_1_24_0_),
            .carryout(n2242),
            .clk(N__5392),
            .ce(),
            .sr(N__3946));
    defparam clk_divider_116__i17_LC_1_24_1.C_ON=1'b1;
    defparam clk_divider_116__i17_LC_1_24_1.SEQ_MODE=4'b1000;
    defparam clk_divider_116__i17_LC_1_24_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 clk_divider_116__i17_LC_1_24_1 (
            .in0(_gnd_net_),
            .in1(N__3454),
            .in2(_gnd_net_),
            .in3(N__2813),
            .lcout(clk_divider_17),
            .ltout(),
            .carryin(n2242),
            .carryout(n2243),
            .clk(N__5392),
            .ce(),
            .sr(N__3946));
    defparam clk_divider_116__i18_LC_1_24_2.C_ON=1'b1;
    defparam clk_divider_116__i18_LC_1_24_2.SEQ_MODE=4'b1000;
    defparam clk_divider_116__i18_LC_1_24_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 clk_divider_116__i18_LC_1_24_2 (
            .in0(_gnd_net_),
            .in1(N__3775),
            .in2(_gnd_net_),
            .in3(N__2864),
            .lcout(clk_divider_18),
            .ltout(),
            .carryin(n2243),
            .carryout(n2244),
            .clk(N__5392),
            .ce(),
            .sr(N__3946));
    defparam clk_divider_116__i19_LC_1_24_3.C_ON=1'b1;
    defparam clk_divider_116__i19_LC_1_24_3.SEQ_MODE=4'b1000;
    defparam clk_divider_116__i19_LC_1_24_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 clk_divider_116__i19_LC_1_24_3 (
            .in0(_gnd_net_),
            .in1(N__3319),
            .in2(_gnd_net_),
            .in3(N__2861),
            .lcout(clk_divider_19),
            .ltout(),
            .carryin(n2244),
            .carryout(n2245),
            .clk(N__5392),
            .ce(),
            .sr(N__3946));
    defparam clk_divider_116__i20_LC_1_24_4.C_ON=1'b1;
    defparam clk_divider_116__i20_LC_1_24_4.SEQ_MODE=4'b1000;
    defparam clk_divider_116__i20_LC_1_24_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 clk_divider_116__i20_LC_1_24_4 (
            .in0(_gnd_net_),
            .in1(N__3334),
            .in2(_gnd_net_),
            .in3(N__2858),
            .lcout(clk_divider_20),
            .ltout(),
            .carryin(n2245),
            .carryout(n2246),
            .clk(N__5392),
            .ce(),
            .sr(N__3946));
    defparam clk_divider_116__i21_LC_1_24_5.C_ON=1'b1;
    defparam clk_divider_116__i21_LC_1_24_5.SEQ_MODE=4'b1000;
    defparam clk_divider_116__i21_LC_1_24_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 clk_divider_116__i21_LC_1_24_5 (
            .in0(_gnd_net_),
            .in1(N__3439),
            .in2(_gnd_net_),
            .in3(N__2855),
            .lcout(clk_divider_21),
            .ltout(),
            .carryin(n2246),
            .carryout(n2247),
            .clk(N__5392),
            .ce(),
            .sr(N__3946));
    defparam clk_divider_116__i22_LC_1_24_6.C_ON=1'b1;
    defparam clk_divider_116__i22_LC_1_24_6.SEQ_MODE=4'b1000;
    defparam clk_divider_116__i22_LC_1_24_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 clk_divider_116__i22_LC_1_24_6 (
            .in0(_gnd_net_),
            .in1(N__3421),
            .in2(_gnd_net_),
            .in3(N__2852),
            .lcout(clk_divider_22),
            .ltout(),
            .carryin(n2247),
            .carryout(n2248),
            .clk(N__5392),
            .ce(),
            .sr(N__3946));
    defparam clk_divider_116__i23_LC_1_24_7.C_ON=1'b1;
    defparam clk_divider_116__i23_LC_1_24_7.SEQ_MODE=4'b1000;
    defparam clk_divider_116__i23_LC_1_24_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 clk_divider_116__i23_LC_1_24_7 (
            .in0(_gnd_net_),
            .in1(N__3727),
            .in2(_gnd_net_),
            .in3(N__2849),
            .lcout(clk_divider_23),
            .ltout(),
            .carryin(n2248),
            .carryout(n2249),
            .clk(N__5392),
            .ce(),
            .sr(N__3946));
    defparam clk_divider_116__i24_LC_1_25_0.C_ON=1'b1;
    defparam clk_divider_116__i24_LC_1_25_0.SEQ_MODE=4'b1000;
    defparam clk_divider_116__i24_LC_1_25_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 clk_divider_116__i24_LC_1_25_0 (
            .in0(_gnd_net_),
            .in1(N__3841),
            .in2(_gnd_net_),
            .in3(N__2846),
            .lcout(clk_divider_24),
            .ltout(),
            .carryin(bfn_1_25_0_),
            .carryout(n2250),
            .clk(N__5395),
            .ce(),
            .sr(N__3947));
    defparam clk_divider_116__i25_LC_1_25_1.C_ON=1'b1;
    defparam clk_divider_116__i25_LC_1_25_1.SEQ_MODE=4'b1000;
    defparam clk_divider_116__i25_LC_1_25_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 clk_divider_116__i25_LC_1_25_1 (
            .in0(_gnd_net_),
            .in1(N__4219),
            .in2(_gnd_net_),
            .in3(N__2843),
            .lcout(clk_divider_25),
            .ltout(),
            .carryin(n2250),
            .carryout(n2251),
            .clk(N__5395),
            .ce(),
            .sr(N__3947));
    defparam clk_divider_116__i26_LC_1_25_2.C_ON=1'b1;
    defparam clk_divider_116__i26_LC_1_25_2.SEQ_MODE=4'b1000;
    defparam clk_divider_116__i26_LC_1_25_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 clk_divider_116__i26_LC_1_25_2 (
            .in0(_gnd_net_),
            .in1(N__3505),
            .in2(_gnd_net_),
            .in3(N__2840),
            .lcout(clk_divider_26),
            .ltout(),
            .carryin(n2251),
            .carryout(n2252),
            .clk(N__5395),
            .ce(),
            .sr(N__3947));
    defparam clk_divider_116__i27_LC_1_25_3.C_ON=1'b1;
    defparam clk_divider_116__i27_LC_1_25_3.SEQ_MODE=4'b1000;
    defparam clk_divider_116__i27_LC_1_25_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 clk_divider_116__i27_LC_1_25_3 (
            .in0(_gnd_net_),
            .in1(N__3352),
            .in2(_gnd_net_),
            .in3(N__3014),
            .lcout(clk_divider_27),
            .ltout(),
            .carryin(n2252),
            .carryout(n2253),
            .clk(N__5395),
            .ce(),
            .sr(N__3947));
    defparam clk_divider_116__i28_LC_1_25_4.C_ON=1'b1;
    defparam clk_divider_116__i28_LC_1_25_4.SEQ_MODE=4'b1000;
    defparam clk_divider_116__i28_LC_1_25_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 clk_divider_116__i28_LC_1_25_4 (
            .in0(_gnd_net_),
            .in1(N__3400),
            .in2(_gnd_net_),
            .in3(N__3011),
            .lcout(clk_divider_28),
            .ltout(),
            .carryin(n2253),
            .carryout(n2254),
            .clk(N__5395),
            .ce(),
            .sr(N__3947));
    defparam clk_divider_116__i29_LC_1_25_5.C_ON=1'b1;
    defparam clk_divider_116__i29_LC_1_25_5.SEQ_MODE=4'b1000;
    defparam clk_divider_116__i29_LC_1_25_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 clk_divider_116__i29_LC_1_25_5 (
            .in0(_gnd_net_),
            .in1(N__3748),
            .in2(_gnd_net_),
            .in3(N__3008),
            .lcout(clk_divider_29),
            .ltout(),
            .carryin(n2254),
            .carryout(n2255),
            .clk(N__5395),
            .ce(),
            .sr(N__3947));
    defparam clk_divider_116__i30_LC_1_25_6.C_ON=1'b1;
    defparam clk_divider_116__i30_LC_1_25_6.SEQ_MODE=4'b1000;
    defparam clk_divider_116__i30_LC_1_25_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 clk_divider_116__i30_LC_1_25_6 (
            .in0(_gnd_net_),
            .in1(N__3370),
            .in2(_gnd_net_),
            .in3(N__3005),
            .lcout(clk_divider_30),
            .ltout(),
            .carryin(n2255),
            .carryout(n2256),
            .clk(N__5395),
            .ce(),
            .sr(N__3947));
    defparam clk_divider_116__i31_LC_1_25_7.C_ON=1'b0;
    defparam clk_divider_116__i31_LC_1_25_7.SEQ_MODE=4'b1000;
    defparam clk_divider_116__i31_LC_1_25_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 clk_divider_116__i31_LC_1_25_7 (
            .in0(_gnd_net_),
            .in1(N__3682),
            .in2(_gnd_net_),
            .in3(N__3002),
            .lcout(clk_divider_31),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__5395),
            .ce(),
            .sr(N__3947));
    defparam \uart.i806_4_lut_LC_2_18_0 .C_ON=1'b0;
    defparam \uart.i806_4_lut_LC_2_18_0 .SEQ_MODE=4'b0000;
    defparam \uart.i806_4_lut_LC_2_18_0 .LUT_INIT=16'b1111111000000000;
    LogicCell40 \uart.i806_4_lut_LC_2_18_0  (
            .in0(N__2999),
            .in1(N__2987),
            .in2(N__2975),
            .in3(N__2959),
            .lcout(),
            .ltout(\uart.n2006_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart.i3_4_lut_LC_2_18_1 .C_ON=1'b0;
    defparam \uart.i3_4_lut_LC_2_18_1 .SEQ_MODE=4'b0000;
    defparam \uart.i3_4_lut_LC_2_18_1 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \uart.i3_4_lut_LC_2_18_1  (
            .in0(N__2947),
            .in1(N__2935),
            .in2(N__2924),
            .in3(N__2920),
            .lcout(\uart.n2385 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart.r_SM_Main_i2_LC_2_19_0 .C_ON=1'b0;
    defparam \uart.r_SM_Main_i2_LC_2_19_0 .SEQ_MODE=4'b1000;
    defparam \uart.r_SM_Main_i2_LC_2_19_0 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \uart.r_SM_Main_i2_LC_2_19_0  (
            .in0(N__4547),
            .in1(N__4678),
            .in2(N__4732),
            .in3(N__4630),
            .lcout(r_SM_Main_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__5382),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart.i18_4_lut_LC_2_19_1 .C_ON=1'b0;
    defparam \uart.i18_4_lut_LC_2_19_1 .SEQ_MODE=4'b0000;
    defparam \uart.i18_4_lut_LC_2_19_1 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \uart.i18_4_lut_LC_2_19_1  (
            .in0(N__2908),
            .in1(N__2896),
            .in2(N__2885),
            .in3(N__3289),
            .lcout(),
            .ltout(\uart.n42_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart.i21_4_lut_LC_2_19_2 .C_ON=1'b0;
    defparam \uart.i21_4_lut_LC_2_19_2 .SEQ_MODE=4'b0000;
    defparam \uart.i21_4_lut_LC_2_19_2 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \uart.i21_4_lut_LC_2_19_2  (
            .in0(N__3277),
            .in1(N__3266),
            .in2(N__3251),
            .in3(N__3167),
            .lcout(),
            .ltout(\uart.n45_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart.i1_4_lut_LC_2_19_3 .C_ON=1'b0;
    defparam \uart.i1_4_lut_LC_2_19_3 .SEQ_MODE=4'b0000;
    defparam \uart.i1_4_lut_LC_2_19_3 .LUT_INIT=16'b1111111011111010;
    LogicCell40 \uart.i1_4_lut_LC_2_19_3  (
            .in0(N__3518),
            .in1(N__3247),
            .in2(N__3236),
            .in3(N__3233),
            .lcout(r_SM_Main_2_N_233_1),
            .ltout(r_SM_Main_2_N_233_1_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart.i1088_4_lut_LC_2_19_4 .C_ON=1'b0;
    defparam \uart.i1088_4_lut_LC_2_19_4 .SEQ_MODE=4'b0000;
    defparam \uart.i1088_4_lut_LC_2_19_4 .LUT_INIT=16'b0000000011110001;
    LogicCell40 \uart.i1088_4_lut_LC_2_19_4  (
            .in0(N__4721),
            .in1(N__4677),
            .in2(N__3227),
            .in3(N__4629),
            .lcout(\uart.n1796 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart.i10_2_lut_LC_2_19_5 .C_ON=1'b0;
    defparam \uart.i10_2_lut_LC_2_19_5 .SEQ_MODE=4'b0000;
    defparam \uart.i10_2_lut_LC_2_19_5 .LUT_INIT=16'b1111111111110000;
    LogicCell40 \uart.i10_2_lut_LC_2_19_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__3194),
            .in3(N__3178),
            .lcout(\uart.n34 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart.i515_4_lut_LC_2_19_7 .C_ON=1'b0;
    defparam \uart.i515_4_lut_LC_2_19_7 .SEQ_MODE=4'b0000;
    defparam \uart.i515_4_lut_LC_2_19_7 .LUT_INIT=16'b1011100000110000;
    LogicCell40 \uart.i515_4_lut_LC_2_19_7  (
            .in0(N__4520),
            .in1(N__4720),
            .in2(N__5099),
            .in3(N__4546),
            .lcout(\uart.n1711 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart.i15_4_lut_LC_2_20_0 .C_ON=1'b0;
    defparam \uart.i15_4_lut_LC_2_20_0 .SEQ_MODE=4'b0000;
    defparam \uart.i15_4_lut_LC_2_20_0 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \uart.i15_4_lut_LC_2_20_0  (
            .in0(N__3160),
            .in1(N__3148),
            .in2(N__3137),
            .in3(N__3118),
            .lcout(\uart.n39 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart.i1_1_lut_LC_2_20_2 .C_ON=1'b0;
    defparam \uart.i1_1_lut_LC_2_20_2 .SEQ_MODE=4'b0000;
    defparam \uart.i1_1_lut_LC_2_20_2 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \uart.i1_1_lut_LC_2_20_2  (
            .in0(N__4631),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\uart.n1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart.i16_4_lut_LC_2_20_3 .C_ON=1'b0;
    defparam \uart.i16_4_lut_LC_2_20_3 .SEQ_MODE=4'b0000;
    defparam \uart.i16_4_lut_LC_2_20_3 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \uart.i16_4_lut_LC_2_20_3  (
            .in0(N__3064),
            .in1(N__3052),
            .in2(N__3041),
            .in3(N__3025),
            .lcout(\uart.n40 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart.i14_4_lut_LC_2_20_4 .C_ON=1'b0;
    defparam \uart.i14_4_lut_LC_2_20_4 .SEQ_MODE=4'b0000;
    defparam \uart.i14_4_lut_LC_2_20_4 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \uart.i14_4_lut_LC_2_20_4  (
            .in0(N__3643),
            .in1(N__3631),
            .in2(N__3620),
            .in3(N__3604),
            .lcout(\uart.n38 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart.i13_4_lut_LC_2_20_5 .C_ON=1'b0;
    defparam \uart.i13_4_lut_LC_2_20_5 .SEQ_MODE=4'b0000;
    defparam \uart.i13_4_lut_LC_2_20_5 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \uart.i13_4_lut_LC_2_20_5  (
            .in0(N__3593),
            .in1(N__3577),
            .in2(N__3566),
            .in3(N__3550),
            .lcout(),
            .ltout(\uart.n37_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart.i22_4_lut_LC_2_20_6 .C_ON=1'b0;
    defparam \uart.i22_4_lut_LC_2_20_6 .SEQ_MODE=4'b0000;
    defparam \uart.i22_4_lut_LC_2_20_6 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \uart.i22_4_lut_LC_2_20_6  (
            .in0(N__3539),
            .in1(N__3533),
            .in2(N__3527),
            .in3(N__3524),
            .lcout(\uart.n46 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i18_4_lut_LC_2_21_1.C_ON=1'b0;
    defparam i18_4_lut_LC_2_21_1.SEQ_MODE=4'b0000;
    defparam i18_4_lut_LC_2_21_1.LUT_INIT=16'b1111111111111110;
    LogicCell40 i18_4_lut_LC_2_21_1 (
            .in0(N__3509),
            .in1(N__3491),
            .in2(N__3476),
            .in3(N__3458),
            .lcout(n44_adj_358),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i15_4_lut_adj_1_LC_2_21_2.C_ON=1'b0;
    defparam i15_4_lut_adj_1_LC_2_21_2.SEQ_MODE=4'b0000;
    defparam i15_4_lut_adj_1_LC_2_21_2.LUT_INIT=16'b1111111111111110;
    LogicCell40 i15_4_lut_adj_1_LC_2_21_2 (
            .in0(N__3440),
            .in1(N__3425),
            .in2(N__3407),
            .in3(N__3385),
            .lcout(n41_adj_361),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i16_4_lut_adj_2_LC_2_21_3.C_ON=1'b0;
    defparam i16_4_lut_adj_2_LC_2_21_3.SEQ_MODE=4'b0000;
    defparam i16_4_lut_adj_2_LC_2_21_3.LUT_INIT=16'b1111111111111110;
    LogicCell40 i16_4_lut_adj_2_LC_2_21_3 (
            .in0(N__3374),
            .in1(N__3356),
            .in2(N__3338),
            .in3(N__3320),
            .lcout(),
            .ltout(n42_adj_360_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i24_4_lut_LC_2_21_4.C_ON=1'b0;
    defparam i24_4_lut_LC_2_21_4.SEQ_MODE=4'b0000;
    defparam i24_4_lut_LC_2_21_4.LUT_INIT=16'b1111111111111110;
    LogicCell40 i24_4_lut_LC_2_21_4 (
            .in0(N__3305),
            .in1(N__3698),
            .in2(N__3299),
            .in3(N__3296),
            .lcout(n50),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i291_4_lut_LC_2_21_5.C_ON=1'b0;
    defparam i291_4_lut_LC_2_21_5.SEQ_MODE=4'b0000;
    defparam i291_4_lut_LC_2_21_5.LUT_INIT=16'b1010101010101000;
    LogicCell40 i291_4_lut_LC_2_21_5 (
            .in0(N__3989),
            .in1(N__3973),
            .in2(N__3962),
            .in3(N__3875),
            .lcout(n10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i708_4_lut_LC_2_22_0.C_ON=1'b0;
    defparam i708_4_lut_LC_2_22_0.SEQ_MODE=4'b0000;
    defparam i708_4_lut_LC_2_22_0.LUT_INIT=16'b0000111100001110;
    LogicCell40 i708_4_lut_LC_2_22_0 (
            .in0(N__3655),
            .in1(N__3664),
            .in2(N__3692),
            .in3(N__4198),
            .lcout(clk_divider_31__N_139),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart.r_SM_Main_2__I_0_62_i3_3_lut_LC_2_22_1 .C_ON=1'b0;
    defparam \uart.r_SM_Main_2__I_0_62_i3_3_lut_LC_2_22_1 .SEQ_MODE=4'b0000;
    defparam \uart.r_SM_Main_2__I_0_62_i3_3_lut_LC_2_22_1 .LUT_INIT=16'b1010101011011101;
    LogicCell40 \uart.r_SM_Main_2__I_0_62_i3_3_lut_LC_2_22_1  (
            .in0(N__4736),
            .in1(N__4256),
            .in2(_gnd_net_),
            .in3(N__4679),
            .lcout(\uart.n3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i2_2_lut_LC_2_22_2.C_ON=1'b0;
    defparam i2_2_lut_LC_2_22_2.SEQ_MODE=4'b0000;
    defparam i2_2_lut_LC_2_22_2.LUT_INIT=16'b1111111111001100;
    LogicCell40 i2_2_lut_LC_2_22_2 (
            .in0(_gnd_net_),
            .in1(N__3898),
            .in2(_gnd_net_),
            .in3(N__3886),
            .lcout(n6_adj_324),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i14_4_lut_adj_4_LC_2_22_3.C_ON=1'b0;
    defparam i14_4_lut_adj_4_LC_2_22_3.SEQ_MODE=4'b0000;
    defparam i14_4_lut_adj_4_LC_2_22_3.LUT_INIT=16'b1111111111111110;
    LogicCell40 i14_4_lut_adj_4_LC_2_22_3 (
            .in0(N__3868),
            .in1(N__3856),
            .in2(N__3845),
            .in3(N__3826),
            .lcout(n40_adj_362),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i19_4_lut_LC_2_22_4.C_ON=1'b0;
    defparam i19_4_lut_LC_2_22_4.SEQ_MODE=4'b0000;
    defparam i19_4_lut_LC_2_22_4.LUT_INIT=16'b1111111111111110;
    LogicCell40 i19_4_lut_LC_2_22_4 (
            .in0(N__3814),
            .in1(N__3802),
            .in2(N__3791),
            .in3(N__3776),
            .lcout(n45_adj_357),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i17_4_lut_adj_3_LC_2_22_6.C_ON=1'b0;
    defparam i17_4_lut_adj_3_LC_2_22_6.SEQ_MODE=4'b0000;
    defparam i17_4_lut_adj_3_LC_2_22_6.LUT_INIT=16'b1111111111111110;
    LogicCell40 i17_4_lut_adj_3_LC_2_22_6 (
            .in0(N__3760),
            .in1(N__3749),
            .in2(N__3734),
            .in3(N__3713),
            .lcout(n43_adj_359),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam clk_slow_25_LC_2_22_7.C_ON=1'b0;
    defparam clk_slow_25_LC_2_22_7.SEQ_MODE=4'b1000;
    defparam clk_slow_25_LC_2_22_7.LUT_INIT=16'b0011001100110010;
    LogicCell40 clk_slow_25_LC_2_22_7 (
            .in0(N__4199),
            .in1(N__3691),
            .in2(N__3668),
            .in3(N__3656),
            .lcout(clk_slow),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__5389),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_119__i0_LC_2_23_0.C_ON=1'b1;
    defparam blink_counter_119__i0_LC_2_23_0.SEQ_MODE=4'b1000;
    defparam blink_counter_119__i0_LC_2_23_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_119__i0_LC_2_23_0 (
            .in0(_gnd_net_),
            .in1(N__4061),
            .in2(_gnd_net_),
            .in3(N__4055),
            .lcout(n26),
            .ltout(),
            .carryin(bfn_2_23_0_),
            .carryout(n2163),
            .clk(N__5393),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_119__i1_LC_2_23_1.C_ON=1'b1;
    defparam blink_counter_119__i1_LC_2_23_1.SEQ_MODE=4'b1000;
    defparam blink_counter_119__i1_LC_2_23_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_119__i1_LC_2_23_1 (
            .in0(_gnd_net_),
            .in1(N__4052),
            .in2(_gnd_net_),
            .in3(N__4046),
            .lcout(n25),
            .ltout(),
            .carryin(n2163),
            .carryout(n2164),
            .clk(N__5393),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_119__i2_LC_2_23_2.C_ON=1'b1;
    defparam blink_counter_119__i2_LC_2_23_2.SEQ_MODE=4'b1000;
    defparam blink_counter_119__i2_LC_2_23_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_119__i2_LC_2_23_2 (
            .in0(_gnd_net_),
            .in1(N__4043),
            .in2(_gnd_net_),
            .in3(N__4037),
            .lcout(n24),
            .ltout(),
            .carryin(n2164),
            .carryout(n2165),
            .clk(N__5393),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_119__i3_LC_2_23_3.C_ON=1'b1;
    defparam blink_counter_119__i3_LC_2_23_3.SEQ_MODE=4'b1000;
    defparam blink_counter_119__i3_LC_2_23_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_119__i3_LC_2_23_3 (
            .in0(_gnd_net_),
            .in1(N__4034),
            .in2(_gnd_net_),
            .in3(N__4028),
            .lcout(n23),
            .ltout(),
            .carryin(n2165),
            .carryout(n2166),
            .clk(N__5393),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_119__i4_LC_2_23_4.C_ON=1'b1;
    defparam blink_counter_119__i4_LC_2_23_4.SEQ_MODE=4'b1000;
    defparam blink_counter_119__i4_LC_2_23_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_119__i4_LC_2_23_4 (
            .in0(_gnd_net_),
            .in1(N__4025),
            .in2(_gnd_net_),
            .in3(N__4019),
            .lcout(n22),
            .ltout(),
            .carryin(n2166),
            .carryout(n2167),
            .clk(N__5393),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_119__i5_LC_2_23_5.C_ON=1'b1;
    defparam blink_counter_119__i5_LC_2_23_5.SEQ_MODE=4'b1000;
    defparam blink_counter_119__i5_LC_2_23_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_119__i5_LC_2_23_5 (
            .in0(_gnd_net_),
            .in1(N__4016),
            .in2(_gnd_net_),
            .in3(N__4010),
            .lcout(n21),
            .ltout(),
            .carryin(n2167),
            .carryout(n2168),
            .clk(N__5393),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_119__i6_LC_2_23_6.C_ON=1'b1;
    defparam blink_counter_119__i6_LC_2_23_6.SEQ_MODE=4'b1000;
    defparam blink_counter_119__i6_LC_2_23_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_119__i6_LC_2_23_6 (
            .in0(_gnd_net_),
            .in1(N__4007),
            .in2(_gnd_net_),
            .in3(N__4001),
            .lcout(n20),
            .ltout(),
            .carryin(n2168),
            .carryout(n2169),
            .clk(N__5393),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_119__i7_LC_2_23_7.C_ON=1'b1;
    defparam blink_counter_119__i7_LC_2_23_7.SEQ_MODE=4'b1000;
    defparam blink_counter_119__i7_LC_2_23_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_119__i7_LC_2_23_7 (
            .in0(_gnd_net_),
            .in1(N__3998),
            .in2(_gnd_net_),
            .in3(N__3992),
            .lcout(n19),
            .ltout(),
            .carryin(n2169),
            .carryout(n2170),
            .clk(N__5393),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_119__i8_LC_2_24_0.C_ON=1'b1;
    defparam blink_counter_119__i8_LC_2_24_0.SEQ_MODE=4'b1000;
    defparam blink_counter_119__i8_LC_2_24_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_119__i8_LC_2_24_0 (
            .in0(_gnd_net_),
            .in1(N__4142),
            .in2(_gnd_net_),
            .in3(N__4136),
            .lcout(n18),
            .ltout(),
            .carryin(bfn_2_24_0_),
            .carryout(n2171),
            .clk(N__5396),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_119__i9_LC_2_24_1.C_ON=1'b1;
    defparam blink_counter_119__i9_LC_2_24_1.SEQ_MODE=4'b1000;
    defparam blink_counter_119__i9_LC_2_24_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_119__i9_LC_2_24_1 (
            .in0(_gnd_net_),
            .in1(N__4133),
            .in2(_gnd_net_),
            .in3(N__4127),
            .lcout(n17),
            .ltout(),
            .carryin(n2171),
            .carryout(n2172),
            .clk(N__5396),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_119__i10_LC_2_24_2.C_ON=1'b1;
    defparam blink_counter_119__i10_LC_2_24_2.SEQ_MODE=4'b1000;
    defparam blink_counter_119__i10_LC_2_24_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_119__i10_LC_2_24_2 (
            .in0(_gnd_net_),
            .in1(N__4124),
            .in2(_gnd_net_),
            .in3(N__4118),
            .lcout(n16),
            .ltout(),
            .carryin(n2172),
            .carryout(n2173),
            .clk(N__5396),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_119__i11_LC_2_24_3.C_ON=1'b1;
    defparam blink_counter_119__i11_LC_2_24_3.SEQ_MODE=4'b1000;
    defparam blink_counter_119__i11_LC_2_24_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_119__i11_LC_2_24_3 (
            .in0(_gnd_net_),
            .in1(N__4115),
            .in2(_gnd_net_),
            .in3(N__4109),
            .lcout(n15),
            .ltout(),
            .carryin(n2173),
            .carryout(n2174),
            .clk(N__5396),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_119__i12_LC_2_24_4.C_ON=1'b1;
    defparam blink_counter_119__i12_LC_2_24_4.SEQ_MODE=4'b1000;
    defparam blink_counter_119__i12_LC_2_24_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_119__i12_LC_2_24_4 (
            .in0(_gnd_net_),
            .in1(N__4106),
            .in2(_gnd_net_),
            .in3(N__4100),
            .lcout(n14),
            .ltout(),
            .carryin(n2174),
            .carryout(n2175),
            .clk(N__5396),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_119__i13_LC_2_24_5.C_ON=1'b1;
    defparam blink_counter_119__i13_LC_2_24_5.SEQ_MODE=4'b1000;
    defparam blink_counter_119__i13_LC_2_24_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_119__i13_LC_2_24_5 (
            .in0(_gnd_net_),
            .in1(N__4097),
            .in2(_gnd_net_),
            .in3(N__4091),
            .lcout(n13),
            .ltout(),
            .carryin(n2175),
            .carryout(n2176),
            .clk(N__5396),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_119__i14_LC_2_24_6.C_ON=1'b1;
    defparam blink_counter_119__i14_LC_2_24_6.SEQ_MODE=4'b1000;
    defparam blink_counter_119__i14_LC_2_24_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_119__i14_LC_2_24_6 (
            .in0(_gnd_net_),
            .in1(N__4088),
            .in2(_gnd_net_),
            .in3(N__4082),
            .lcout(n12),
            .ltout(),
            .carryin(n2176),
            .carryout(n2177),
            .clk(N__5396),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_119__i15_LC_2_24_7.C_ON=1'b1;
    defparam blink_counter_119__i15_LC_2_24_7.SEQ_MODE=4'b1000;
    defparam blink_counter_119__i15_LC_2_24_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_119__i15_LC_2_24_7 (
            .in0(_gnd_net_),
            .in1(N__4079),
            .in2(_gnd_net_),
            .in3(N__4073),
            .lcout(n11),
            .ltout(),
            .carryin(n2177),
            .carryout(n2178),
            .clk(N__5396),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_119__i16_LC_2_25_0.C_ON=1'b1;
    defparam blink_counter_119__i16_LC_2_25_0.SEQ_MODE=4'b1000;
    defparam blink_counter_119__i16_LC_2_25_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_119__i16_LC_2_25_0 (
            .in0(_gnd_net_),
            .in1(N__4070),
            .in2(_gnd_net_),
            .in3(N__4064),
            .lcout(n10_adj_317),
            .ltout(),
            .carryin(bfn_2_25_0_),
            .carryout(n2179),
            .clk(N__5397),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_119__i17_LC_2_25_1.C_ON=1'b1;
    defparam blink_counter_119__i17_LC_2_25_1.SEQ_MODE=4'b1000;
    defparam blink_counter_119__i17_LC_2_25_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_119__i17_LC_2_25_1 (
            .in0(_gnd_net_),
            .in1(N__4190),
            .in2(_gnd_net_),
            .in3(N__4184),
            .lcout(n9),
            .ltout(),
            .carryin(n2179),
            .carryout(n2180),
            .clk(N__5397),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_119__i18_LC_2_25_2.C_ON=1'b1;
    defparam blink_counter_119__i18_LC_2_25_2.SEQ_MODE=4'b1000;
    defparam blink_counter_119__i18_LC_2_25_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_119__i18_LC_2_25_2 (
            .in0(_gnd_net_),
            .in1(N__4181),
            .in2(_gnd_net_),
            .in3(N__4175),
            .lcout(n8),
            .ltout(),
            .carryin(n2180),
            .carryout(n2181),
            .clk(N__5397),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_119__i19_LC_2_25_3.C_ON=1'b1;
    defparam blink_counter_119__i19_LC_2_25_3.SEQ_MODE=4'b1000;
    defparam blink_counter_119__i19_LC_2_25_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_119__i19_LC_2_25_3 (
            .in0(_gnd_net_),
            .in1(N__4172),
            .in2(_gnd_net_),
            .in3(N__4166),
            .lcout(n7),
            .ltout(),
            .carryin(n2181),
            .carryout(n2182),
            .clk(N__5397),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_119__i20_LC_2_25_4.C_ON=1'b1;
    defparam blink_counter_119__i20_LC_2_25_4.SEQ_MODE=4'b1000;
    defparam blink_counter_119__i20_LC_2_25_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_119__i20_LC_2_25_4 (
            .in0(_gnd_net_),
            .in1(N__4163),
            .in2(_gnd_net_),
            .in3(N__4157),
            .lcout(n6),
            .ltout(),
            .carryin(n2182),
            .carryout(n2183),
            .clk(N__5397),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_119__i21_LC_2_25_5.C_ON=1'b1;
    defparam blink_counter_119__i21_LC_2_25_5.SEQ_MODE=4'b1000;
    defparam blink_counter_119__i21_LC_2_25_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_119__i21_LC_2_25_5 (
            .in0(_gnd_net_),
            .in1(N__4336),
            .in2(_gnd_net_),
            .in3(N__4154),
            .lcout(blink_counter_21),
            .ltout(),
            .carryin(n2183),
            .carryout(n2184),
            .clk(N__5397),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_119__i22_LC_2_25_6.C_ON=1'b1;
    defparam blink_counter_119__i22_LC_2_25_6.SEQ_MODE=4'b1000;
    defparam blink_counter_119__i22_LC_2_25_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_119__i22_LC_2_25_6 (
            .in0(_gnd_net_),
            .in1(N__4279),
            .in2(_gnd_net_),
            .in3(N__4151),
            .lcout(blink_counter_22),
            .ltout(),
            .carryin(n2184),
            .carryout(n2185),
            .clk(N__5397),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_119__i23_LC_2_25_7.C_ON=1'b1;
    defparam blink_counter_119__i23_LC_2_25_7.SEQ_MODE=4'b1000;
    defparam blink_counter_119__i23_LC_2_25_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_119__i23_LC_2_25_7 (
            .in0(_gnd_net_),
            .in1(N__4297),
            .in2(_gnd_net_),
            .in3(N__4148),
            .lcout(blink_counter_23),
            .ltout(),
            .carryin(n2185),
            .carryout(n2186),
            .clk(N__5397),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_119__i24_LC_2_26_0.C_ON=1'b1;
    defparam blink_counter_119__i24_LC_2_26_0.SEQ_MODE=4'b1000;
    defparam blink_counter_119__i24_LC_2_26_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_119__i24_LC_2_26_0 (
            .in0(_gnd_net_),
            .in1(N__4323),
            .in2(_gnd_net_),
            .in3(N__4145),
            .lcout(blink_counter_24),
            .ltout(),
            .carryin(bfn_2_26_0_),
            .carryout(n2187),
            .clk(N__5398),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_119__i25_LC_2_26_1.C_ON=1'b0;
    defparam blink_counter_119__i25_LC_2_26_1.SEQ_MODE=4'b1000;
    defparam blink_counter_119__i25_LC_2_26_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_119__i25_LC_2_26_1 (
            .in0(_gnd_net_),
            .in1(N__4372),
            .in2(_gnd_net_),
            .in3(N__4376),
            .lcout(blink_counter_25),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__5398),
            .ce(),
            .sr(_gnd_net_));
    defparam i1070_4_lut_LC_2_27_0.C_ON=1'b0;
    defparam i1070_4_lut_LC_2_27_0.SEQ_MODE=4'b0000;
    defparam i1070_4_lut_LC_2_27_0.LUT_INIT=16'b1110101011111000;
    LogicCell40 i1070_4_lut_LC_2_27_0 (
            .in0(N__4343),
            .in1(N__4325),
            .in2(N__4310),
            .in3(N__4286),
            .lcout(),
            .ltout(n2395_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1071_3_lut_LC_2_27_1.C_ON=1'b0;
    defparam i1071_3_lut_LC_2_27_1.SEQ_MODE=4'b0000;
    defparam i1071_3_lut_LC_2_27_1.LUT_INIT=16'b0000101001011111;
    LogicCell40 i1071_3_lut_LC_2_27_1 (
            .in0(N__4373),
            .in1(_gnd_net_),
            .in2(N__4361),
            .in3(N__4268),
            .lcout(LED_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1069_4_lut_LC_2_27_6.C_ON=1'b0;
    defparam i1069_4_lut_LC_2_27_6.SEQ_MODE=4'b0000;
    defparam i1069_4_lut_LC_2_27_6.LUT_INIT=16'b1011101000100010;
    LogicCell40 i1069_4_lut_LC_2_27_6 (
            .in0(N__4342),
            .in1(N__4324),
            .in2(N__4309),
            .in3(N__4285),
            .lcout(n2394),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart.r_SM_Main_i0_LC_3_19_0 .C_ON=1'b0;
    defparam \uart.r_SM_Main_i0_LC_3_19_0 .SEQ_MODE=4'b1000;
    defparam \uart.r_SM_Main_i0_LC_3_19_0 .LUT_INIT=16'b0111011101000100;
    LogicCell40 \uart.r_SM_Main_i0_LC_3_19_0  (
            .in0(N__4549),
            .in1(N__4672),
            .in2(_gnd_net_),
            .in3(N__4262),
            .lcout(r_SM_Main_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__5384),
            .ce(),
            .sr(N__4636));
    defparam \uart.r_SM_Main_i1_LC_3_19_1 .C_ON=1'b0;
    defparam \uart.r_SM_Main_i1_LC_3_19_1 .SEQ_MODE=4'b1000;
    defparam \uart.r_SM_Main_i1_LC_3_19_1 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \uart.r_SM_Main_i1_LC_3_19_1  (
            .in0(N__4673),
            .in1(N__4729),
            .in2(_gnd_net_),
            .in3(N__4548),
            .lcout(r_SM_Main_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__5384),
            .ce(),
            .sr(N__4636));
    defparam \uart.r_Bit_Index_i2_LC_3_20_3 .C_ON=1'b0;
    defparam \uart.r_Bit_Index_i2_LC_3_20_3 .SEQ_MODE=4'b1000;
    defparam \uart.r_Bit_Index_i2_LC_3_20_3 .LUT_INIT=16'b0110011010101010;
    LogicCell40 \uart.r_Bit_Index_i2_LC_3_20_3  (
            .in0(N__4571),
            .in1(N__5447),
            .in2(_gnd_net_),
            .in3(N__5477),
            .lcout(\uart.r_Bit_Index_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__5386),
            .ce(N__5329),
            .sr(N__5302));
    defparam \uart.i8225_i1_3_lut_LC_3_21_0 .C_ON=1'b0;
    defparam \uart.i8225_i1_3_lut_LC_3_21_0 .SEQ_MODE=4'b0000;
    defparam \uart.i8225_i1_3_lut_LC_3_21_0 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \uart.i8225_i1_3_lut_LC_3_21_0  (
            .in0(N__4570),
            .in1(N__4751),
            .in2(_gnd_net_),
            .in3(N__4778),
            .lcout(\uart.o_Tx_Serial_N_312 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i23_4_lut_LC_3_21_5.C_ON=1'b0;
    defparam i23_4_lut_LC_3_21_5.SEQ_MODE=4'b0000;
    defparam i23_4_lut_LC_3_21_5.LUT_INIT=16'b1111111111111110;
    LogicCell40 i23_4_lut_LC_3_21_5 (
            .in0(N__4250),
            .in1(N__4232),
            .in2(N__4226),
            .in3(N__4205),
            .lcout(n49),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam counter_117__i0_LC_3_22_0.C_ON=1'b1;
    defparam counter_117__i0_LC_3_22_0.SEQ_MODE=4'b1000;
    defparam counter_117__i0_LC_3_22_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 counter_117__i0_LC_3_22_0 (
            .in0(_gnd_net_),
            .in1(N__4448),
            .in2(_gnd_net_),
            .in3(N__4442),
            .lcout(counter_0),
            .ltout(),
            .carryin(bfn_3_22_0_),
            .carryout(n2195),
            .clk(N__5754),
            .ce(),
            .sr(N__5709));
    defparam counter_117__i1_LC_3_22_1.C_ON=1'b1;
    defparam counter_117__i1_LC_3_22_1.SEQ_MODE=4'b1000;
    defparam counter_117__i1_LC_3_22_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 counter_117__i1_LC_3_22_1 (
            .in0(_gnd_net_),
            .in1(N__4439),
            .in2(_gnd_net_),
            .in3(N__4433),
            .lcout(counter_1),
            .ltout(),
            .carryin(n2195),
            .carryout(n2196),
            .clk(N__5754),
            .ce(),
            .sr(N__5709));
    defparam counter_117__i2_LC_3_22_2.C_ON=1'b1;
    defparam counter_117__i2_LC_3_22_2.SEQ_MODE=4'b1000;
    defparam counter_117__i2_LC_3_22_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 counter_117__i2_LC_3_22_2 (
            .in0(_gnd_net_),
            .in1(N__4430),
            .in2(_gnd_net_),
            .in3(N__4424),
            .lcout(counter_2),
            .ltout(),
            .carryin(n2196),
            .carryout(n2197),
            .clk(N__5754),
            .ce(),
            .sr(N__5709));
    defparam counter_117__i3_LC_3_22_3.C_ON=1'b1;
    defparam counter_117__i3_LC_3_22_3.SEQ_MODE=4'b1000;
    defparam counter_117__i3_LC_3_22_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 counter_117__i3_LC_3_22_3 (
            .in0(_gnd_net_),
            .in1(N__4421),
            .in2(_gnd_net_),
            .in3(N__4415),
            .lcout(counter_3),
            .ltout(),
            .carryin(n2197),
            .carryout(n2198),
            .clk(N__5754),
            .ce(),
            .sr(N__5709));
    defparam counter_117__i4_LC_3_22_4.C_ON=1'b1;
    defparam counter_117__i4_LC_3_22_4.SEQ_MODE=4'b1000;
    defparam counter_117__i4_LC_3_22_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 counter_117__i4_LC_3_22_4 (
            .in0(_gnd_net_),
            .in1(N__4412),
            .in2(_gnd_net_),
            .in3(N__4406),
            .lcout(counter_4),
            .ltout(),
            .carryin(n2198),
            .carryout(n2199),
            .clk(N__5754),
            .ce(),
            .sr(N__5709));
    defparam counter_117__i5_LC_3_22_5.C_ON=1'b1;
    defparam counter_117__i5_LC_3_22_5.SEQ_MODE=4'b1000;
    defparam counter_117__i5_LC_3_22_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 counter_117__i5_LC_3_22_5 (
            .in0(_gnd_net_),
            .in1(N__4403),
            .in2(_gnd_net_),
            .in3(N__4397),
            .lcout(counter_5),
            .ltout(),
            .carryin(n2199),
            .carryout(n2200),
            .clk(N__5754),
            .ce(),
            .sr(N__5709));
    defparam counter_117__i6_LC_3_22_6.C_ON=1'b1;
    defparam counter_117__i6_LC_3_22_6.SEQ_MODE=4'b1000;
    defparam counter_117__i6_LC_3_22_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 counter_117__i6_LC_3_22_6 (
            .in0(_gnd_net_),
            .in1(N__4394),
            .in2(_gnd_net_),
            .in3(N__4388),
            .lcout(counter_6),
            .ltout(),
            .carryin(n2200),
            .carryout(n2201),
            .clk(N__5754),
            .ce(),
            .sr(N__5709));
    defparam counter_117__i7_LC_3_22_7.C_ON=1'b1;
    defparam counter_117__i7_LC_3_22_7.SEQ_MODE=4'b1000;
    defparam counter_117__i7_LC_3_22_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 counter_117__i7_LC_3_22_7 (
            .in0(_gnd_net_),
            .in1(N__4385),
            .in2(_gnd_net_),
            .in3(N__4379),
            .lcout(counter_7),
            .ltout(),
            .carryin(n2201),
            .carryout(n2202),
            .clk(N__5754),
            .ce(),
            .sr(N__5709));
    defparam counter_117__i8_LC_3_23_0.C_ON=1'b1;
    defparam counter_117__i8_LC_3_23_0.SEQ_MODE=4'b1000;
    defparam counter_117__i8_LC_3_23_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 counter_117__i8_LC_3_23_0 (
            .in0(_gnd_net_),
            .in1(N__4988),
            .in2(_gnd_net_),
            .in3(N__4475),
            .lcout(counter_8),
            .ltout(),
            .carryin(bfn_3_23_0_),
            .carryout(n2203),
            .clk(N__5812),
            .ce(),
            .sr(N__5707));
    defparam counter_117__i9_LC_3_23_1.C_ON=1'b1;
    defparam counter_117__i9_LC_3_23_1.SEQ_MODE=4'b1000;
    defparam counter_117__i9_LC_3_23_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 counter_117__i9_LC_3_23_1 (
            .in0(_gnd_net_),
            .in1(N__5510),
            .in2(_gnd_net_),
            .in3(N__4472),
            .lcout(counter_9),
            .ltout(),
            .carryin(n2203),
            .carryout(n2204),
            .clk(N__5812),
            .ce(),
            .sr(N__5707));
    defparam counter_117__i10_LC_3_23_2.C_ON=1'b1;
    defparam counter_117__i10_LC_3_23_2.SEQ_MODE=4'b1000;
    defparam counter_117__i10_LC_3_23_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 counter_117__i10_LC_3_23_2 (
            .in0(_gnd_net_),
            .in1(N__5579),
            .in2(_gnd_net_),
            .in3(N__4469),
            .lcout(counter_10),
            .ltout(),
            .carryin(n2204),
            .carryout(n2205),
            .clk(N__5812),
            .ce(),
            .sr(N__5707));
    defparam counter_117__i11_LC_3_23_3.C_ON=1'b1;
    defparam counter_117__i11_LC_3_23_3.SEQ_MODE=4'b1000;
    defparam counter_117__i11_LC_3_23_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 counter_117__i11_LC_3_23_3 (
            .in0(_gnd_net_),
            .in1(N__5176),
            .in2(_gnd_net_),
            .in3(N__4466),
            .lcout(counter_11),
            .ltout(),
            .carryin(n2205),
            .carryout(n2206),
            .clk(N__5812),
            .ce(),
            .sr(N__5707));
    defparam counter_117__i12_LC_3_23_4.C_ON=1'b1;
    defparam counter_117__i12_LC_3_23_4.SEQ_MODE=4'b1000;
    defparam counter_117__i12_LC_3_23_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 counter_117__i12_LC_3_23_4 (
            .in0(_gnd_net_),
            .in1(N__5000),
            .in2(_gnd_net_),
            .in3(N__4463),
            .lcout(counter_12),
            .ltout(),
            .carryin(n2206),
            .carryout(n2207),
            .clk(N__5812),
            .ce(),
            .sr(N__5707));
    defparam counter_117__i13_LC_3_23_5.C_ON=1'b1;
    defparam counter_117__i13_LC_3_23_5.SEQ_MODE=4'b1000;
    defparam counter_117__i13_LC_3_23_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 counter_117__i13_LC_3_23_5 (
            .in0(_gnd_net_),
            .in1(N__5203),
            .in2(_gnd_net_),
            .in3(N__4460),
            .lcout(counter_13),
            .ltout(),
            .carryin(n2207),
            .carryout(n2208),
            .clk(N__5812),
            .ce(),
            .sr(N__5707));
    defparam counter_117__i14_LC_3_23_6.C_ON=1'b1;
    defparam counter_117__i14_LC_3_23_6.SEQ_MODE=4'b1000;
    defparam counter_117__i14_LC_3_23_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 counter_117__i14_LC_3_23_6 (
            .in0(_gnd_net_),
            .in1(N__5162),
            .in2(_gnd_net_),
            .in3(N__4457),
            .lcout(counter_14),
            .ltout(),
            .carryin(n2208),
            .carryout(n2209),
            .clk(N__5812),
            .ce(),
            .sr(N__5707));
    defparam counter_117__i15_LC_3_23_7.C_ON=1'b1;
    defparam counter_117__i15_LC_3_23_7.SEQ_MODE=4'b1000;
    defparam counter_117__i15_LC_3_23_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 counter_117__i15_LC_3_23_7 (
            .in0(_gnd_net_),
            .in1(N__4975),
            .in2(_gnd_net_),
            .in3(N__4454),
            .lcout(counter_15),
            .ltout(),
            .carryin(n2209),
            .carryout(n2210),
            .clk(N__5812),
            .ce(),
            .sr(N__5707));
    defparam counter_117__i16_LC_3_24_0.C_ON=1'b1;
    defparam counter_117__i16_LC_3_24_0.SEQ_MODE=4'b1000;
    defparam counter_117__i16_LC_3_24_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 counter_117__i16_LC_3_24_0 (
            .in0(_gnd_net_),
            .in1(N__5612),
            .in2(_gnd_net_),
            .in3(N__4451),
            .lcout(counter_16),
            .ltout(),
            .carryin(bfn_3_24_0_),
            .carryout(n2211),
            .clk(N__5814),
            .ce(),
            .sr(N__5710));
    defparam counter_117__i17_LC_3_24_1.C_ON=1'b1;
    defparam counter_117__i17_LC_3_24_1.SEQ_MODE=4'b1000;
    defparam counter_117__i17_LC_3_24_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 counter_117__i17_LC_3_24_1 (
            .in0(_gnd_net_),
            .in1(N__5651),
            .in2(_gnd_net_),
            .in3(N__4505),
            .lcout(counter_17),
            .ltout(),
            .carryin(n2211),
            .carryout(n2212),
            .clk(N__5814),
            .ce(),
            .sr(N__5710));
    defparam counter_117__i18_LC_3_24_2.C_ON=1'b1;
    defparam counter_117__i18_LC_3_24_2.SEQ_MODE=4'b1000;
    defparam counter_117__i18_LC_3_24_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 counter_117__i18_LC_3_24_2 (
            .in0(_gnd_net_),
            .in1(N__5534),
            .in2(_gnd_net_),
            .in3(N__4502),
            .lcout(counter_18),
            .ltout(),
            .carryin(n2212),
            .carryout(n2213),
            .clk(N__5814),
            .ce(),
            .sr(N__5710));
    defparam counter_117__i19_LC_3_24_3.C_ON=1'b1;
    defparam counter_117__i19_LC_3_24_3.SEQ_MODE=4'b1000;
    defparam counter_117__i19_LC_3_24_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 counter_117__i19_LC_3_24_3 (
            .in0(_gnd_net_),
            .in1(N__5032),
            .in2(_gnd_net_),
            .in3(N__4499),
            .lcout(counter_19),
            .ltout(),
            .carryin(n2213),
            .carryout(n2214),
            .clk(N__5814),
            .ce(),
            .sr(N__5710));
    defparam counter_117__i20_LC_3_24_4.C_ON=1'b1;
    defparam counter_117__i20_LC_3_24_4.SEQ_MODE=4'b1000;
    defparam counter_117__i20_LC_3_24_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 counter_117__i20_LC_3_24_4 (
            .in0(_gnd_net_),
            .in1(N__5591),
            .in2(_gnd_net_),
            .in3(N__4496),
            .lcout(counter_20),
            .ltout(),
            .carryin(n2214),
            .carryout(n2215),
            .clk(N__5814),
            .ce(),
            .sr(N__5710));
    defparam counter_117__i21_LC_3_24_5.C_ON=1'b1;
    defparam counter_117__i21_LC_3_24_5.SEQ_MODE=4'b1000;
    defparam counter_117__i21_LC_3_24_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 counter_117__i21_LC_3_24_5 (
            .in0(_gnd_net_),
            .in1(N__5626),
            .in2(_gnd_net_),
            .in3(N__4493),
            .lcout(counter_21),
            .ltout(),
            .carryin(n2215),
            .carryout(n2216),
            .clk(N__5814),
            .ce(),
            .sr(N__5710));
    defparam counter_117__i22_LC_3_24_6.C_ON=1'b1;
    defparam counter_117__i22_LC_3_24_6.SEQ_MODE=4'b1000;
    defparam counter_117__i22_LC_3_24_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 counter_117__i22_LC_3_24_6 (
            .in0(_gnd_net_),
            .in1(N__5057),
            .in2(_gnd_net_),
            .in3(N__4490),
            .lcout(counter_22),
            .ltout(),
            .carryin(n2216),
            .carryout(n2217),
            .clk(N__5814),
            .ce(),
            .sr(N__5710));
    defparam counter_117__i23_LC_3_24_7.C_ON=1'b1;
    defparam counter_117__i23_LC_3_24_7.SEQ_MODE=4'b1000;
    defparam counter_117__i23_LC_3_24_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 counter_117__i23_LC_3_24_7 (
            .in0(_gnd_net_),
            .in1(N__5189),
            .in2(_gnd_net_),
            .in3(N__4487),
            .lcout(counter_23),
            .ltout(),
            .carryin(n2217),
            .carryout(n2218),
            .clk(N__5814),
            .ce(),
            .sr(N__5710));
    defparam counter_117__i24_LC_3_25_0.C_ON=1'b1;
    defparam counter_117__i24_LC_3_25_0.SEQ_MODE=4'b1000;
    defparam counter_117__i24_LC_3_25_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 counter_117__i24_LC_3_25_0 (
            .in0(_gnd_net_),
            .in1(N__5639),
            .in2(_gnd_net_),
            .in3(N__4484),
            .lcout(counter_24),
            .ltout(),
            .carryin(bfn_3_25_0_),
            .carryout(n2219),
            .clk(N__5813),
            .ce(),
            .sr(N__5717));
    defparam counter_117__i25_LC_3_25_1.C_ON=1'b1;
    defparam counter_117__i25_LC_3_25_1.SEQ_MODE=4'b1000;
    defparam counter_117__i25_LC_3_25_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 counter_117__i25_LC_3_25_1 (
            .in0(_gnd_net_),
            .in1(N__4961),
            .in2(_gnd_net_),
            .in3(N__4481),
            .lcout(counter_25),
            .ltout(),
            .carryin(n2219),
            .carryout(n2220),
            .clk(N__5813),
            .ce(),
            .sr(N__5717));
    defparam counter_117__i26_LC_3_25_2.C_ON=1'b1;
    defparam counter_117__i26_LC_3_25_2.SEQ_MODE=4'b1000;
    defparam counter_117__i26_LC_3_25_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 counter_117__i26_LC_3_25_2 (
            .in0(_gnd_net_),
            .in1(N__5018),
            .in2(_gnd_net_),
            .in3(N__4478),
            .lcout(counter_26),
            .ltout(),
            .carryin(n2220),
            .carryout(n2221),
            .clk(N__5813),
            .ce(),
            .sr(N__5717));
    defparam counter_117__i27_LC_3_25_3.C_ON=1'b1;
    defparam counter_117__i27_LC_3_25_3.SEQ_MODE=4'b1000;
    defparam counter_117__i27_LC_3_25_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 counter_117__i27_LC_3_25_3 (
            .in0(_gnd_net_),
            .in1(N__5522),
            .in2(_gnd_net_),
            .in3(N__4586),
            .lcout(counter_27),
            .ltout(),
            .carryin(n2221),
            .carryout(n2222),
            .clk(N__5813),
            .ce(),
            .sr(N__5717));
    defparam counter_117__i28_LC_3_25_4.C_ON=1'b1;
    defparam counter_117__i28_LC_3_25_4.SEQ_MODE=4'b1000;
    defparam counter_117__i28_LC_3_25_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 counter_117__i28_LC_3_25_4 (
            .in0(_gnd_net_),
            .in1(N__5552),
            .in2(_gnd_net_),
            .in3(N__4583),
            .lcout(counter_28),
            .ltout(),
            .carryin(n2222),
            .carryout(n2223),
            .clk(N__5813),
            .ce(),
            .sr(N__5717));
    defparam counter_117__i29_LC_3_25_5.C_ON=1'b1;
    defparam counter_117__i29_LC_3_25_5.SEQ_MODE=4'b1000;
    defparam counter_117__i29_LC_3_25_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 counter_117__i29_LC_3_25_5 (
            .in0(_gnd_net_),
            .in1(N__5566),
            .in2(_gnd_net_),
            .in3(N__4580),
            .lcout(counter_29),
            .ltout(),
            .carryin(n2223),
            .carryout(n2224),
            .clk(N__5813),
            .ce(),
            .sr(N__5717));
    defparam counter_117__i30_LC_3_25_6.C_ON=1'b1;
    defparam counter_117__i30_LC_3_25_6.SEQ_MODE=4'b1000;
    defparam counter_117__i30_LC_3_25_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 counter_117__i30_LC_3_25_6 (
            .in0(_gnd_net_),
            .in1(N__5045),
            .in2(_gnd_net_),
            .in3(N__4577),
            .lcout(counter_30),
            .ltout(),
            .carryin(n2224),
            .carryout(n2225),
            .clk(N__5813),
            .ce(),
            .sr(N__5717));
    defparam counter_117__i31_LC_3_25_7.C_ON=1'b0;
    defparam counter_117__i31_LC_3_25_7.SEQ_MODE=4'b1000;
    defparam counter_117__i31_LC_3_25_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 counter_117__i31_LC_3_25_7 (
            .in0(_gnd_net_),
            .in1(N__5119),
            .in2(_gnd_net_),
            .in3(N__4574),
            .lcout(counter_31),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__5813),
            .ce(),
            .sr(N__5717));
    defparam \uart.i2_3_lut_LC_4_19_3 .C_ON=1'b0;
    defparam \uart.i2_3_lut_LC_4_19_3 .SEQ_MODE=4'b0000;
    defparam \uart.i2_3_lut_LC_4_19_3 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \uart.i2_3_lut_LC_4_19_3  (
            .in0(N__4569),
            .in1(N__5437),
            .in2(_gnd_net_),
            .in3(N__5474),
            .lcout(n2002),
            .ltout(n2002_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart.r_Bit_Index_i0_LC_4_19_4 .C_ON=1'b0;
    defparam \uart.r_Bit_Index_i0_LC_4_19_4 .SEQ_MODE=4'b1000;
    defparam \uart.r_Bit_Index_i0_LC_4_19_4 .LUT_INIT=16'b0000010010101010;
    LogicCell40 \uart.r_Bit_Index_i0_LC_4_19_4  (
            .in0(N__5475),
            .in1(N__4730),
            .in2(N__4553),
            .in3(N__5319),
            .lcout(r_Bit_Index_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__5387),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart.i1095_3_lut_4_lut_LC_4_19_6 .C_ON=1'b0;
    defparam \uart.i1095_3_lut_4_lut_LC_4_19_6 .SEQ_MODE=4'b0000;
    defparam \uart.i1095_3_lut_4_lut_LC_4_19_6 .LUT_INIT=16'b0001000100000001;
    LogicCell40 \uart.i1095_3_lut_4_lut_LC_4_19_6  (
            .in0(N__4662),
            .in1(N__4632),
            .in2(N__4731),
            .in3(N__4550),
            .lcout(n2308),
            .ltout(n2308_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart.i1091_2_lut_3_lut_LC_4_19_7 .C_ON=1'b0;
    defparam \uart.i1091_2_lut_3_lut_LC_4_19_7 .SEQ_MODE=4'b0000;
    defparam \uart.i1091_2_lut_3_lut_LC_4_19_7 .LUT_INIT=16'b1111000000110000;
    LogicCell40 \uart.i1091_2_lut_3_lut_LC_4_19_7  (
            .in0(_gnd_net_),
            .in1(N__4719),
            .in2(N__4523),
            .in3(N__4519),
            .lcout(\uart.n2310 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart.r_Tx_Data_i4_LC_4_20_0 .C_ON=1'b0;
    defparam \uart.r_Tx_Data_i4_LC_4_20_0 .SEQ_MODE=4'b1000;
    defparam \uart.r_Tx_Data_i4_LC_4_20_0 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \uart.r_Tx_Data_i4_LC_4_20_0  (
            .in0(N__5141),
            .in1(N__4888),
            .in2(_gnd_net_),
            .in3(N__4772),
            .lcout(r_Tx_Data_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__5390),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart.r_Bit_Index_0__bdd_4_lut_LC_4_20_1 .C_ON=1'b0;
    defparam \uart.r_Bit_Index_0__bdd_4_lut_LC_4_20_1 .SEQ_MODE=4'b0000;
    defparam \uart.r_Bit_Index_0__bdd_4_lut_LC_4_20_1 .LUT_INIT=16'b1010111111000000;
    LogicCell40 \uart.r_Bit_Index_0__bdd_4_lut_LC_4_20_1  (
            .in0(N__4930),
            .in1(N__4864),
            .in2(N__5442),
            .in3(N__5472),
            .lcout(),
            .ltout(\uart.n2428_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart.n2428_bdd_4_lut_LC_4_20_2 .C_ON=1'b0;
    defparam \uart.n2428_bdd_4_lut_LC_4_20_2 .SEQ_MODE=4'b0000;
    defparam \uart.n2428_bdd_4_lut_LC_4_20_2 .LUT_INIT=16'b1111001011000010;
    LogicCell40 \uart.n2428_bdd_4_lut_LC_4_20_2  (
            .in0(N__4906),
            .in1(N__5432),
            .in2(N__4781),
            .in3(N__4597),
            .lcout(\uart.n2431 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart.r_Tx_Data_i5_LC_4_20_3 .C_ON=1'b0;
    defparam \uart.r_Tx_Data_i5_LC_4_20_3 .SEQ_MODE=4'b1000;
    defparam \uart.r_Tx_Data_i5_LC_4_20_3 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \uart.r_Tx_Data_i5_LC_4_20_3  (
            .in0(N__4889),
            .in1(N__4853),
            .in2(_gnd_net_),
            .in3(N__4763),
            .lcout(r_Tx_Data_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__5390),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart.r_Bit_Index_0__bdd_4_lut_1104_LC_4_20_4 .C_ON=1'b0;
    defparam \uart.r_Bit_Index_0__bdd_4_lut_1104_LC_4_20_4 .SEQ_MODE=4'b0000;
    defparam \uart.r_Bit_Index_0__bdd_4_lut_1104_LC_4_20_4 .LUT_INIT=16'b1101101010001010;
    LogicCell40 \uart.r_Bit_Index_0__bdd_4_lut_1104_LC_4_20_4  (
            .in0(N__5473),
            .in1(N__4918),
            .in2(N__5443),
            .in3(N__4744),
            .lcout(),
            .ltout(\uart.n2422_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart.n2422_bdd_4_lut_LC_4_20_5 .C_ON=1'b0;
    defparam \uart.n2422_bdd_4_lut_LC_4_20_5 .SEQ_MODE=4'b0000;
    defparam \uart.n2422_bdd_4_lut_LC_4_20_5 .LUT_INIT=16'b1111000011001010;
    LogicCell40 \uart.n2422_bdd_4_lut_LC_4_20_5  (
            .in0(N__4771),
            .in1(N__4762),
            .in2(N__4754),
            .in3(N__5436),
            .lcout(\uart.n2425 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart.r_Tx_Data_i6_LC_4_20_6 .C_ON=1'b0;
    defparam \uart.r_Tx_Data_i6_LC_4_20_6 .SEQ_MODE=4'b1000;
    defparam \uart.r_Tx_Data_i6_LC_4_20_6 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \uart.r_Tx_Data_i6_LC_4_20_6  (
            .in0(N__5072),
            .in1(N__4890),
            .in2(_gnd_net_),
            .in3(N__4745),
            .lcout(r_Tx_Data_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__5390),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart.i2_3_lut_4_lut_LC_4_20_7 .C_ON=1'b0;
    defparam \uart.i2_3_lut_4_lut_LC_4_20_7 .SEQ_MODE=4'b0000;
    defparam \uart.i2_3_lut_4_lut_LC_4_20_7 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \uart.i2_3_lut_4_lut_LC_4_20_7  (
            .in0(N__4725),
            .in1(N__4663),
            .in2(N__5092),
            .in3(N__4637),
            .lcout(n1757),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart.r_Tx_Data_i1_LC_4_21_2 .C_ON=1'b0;
    defparam \uart.r_Tx_Data_i1_LC_4_21_2 .SEQ_MODE=4'b1000;
    defparam \uart.r_Tx_Data_i1_LC_4_21_2 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \uart.r_Tx_Data_i1_LC_4_21_2  (
            .in0(N__4811),
            .in1(N__4892),
            .in2(_gnd_net_),
            .in3(N__4598),
            .lcout(r_Tx_Data_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__5394),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart.r_Tx_Data_i3_LC_4_21_3 .C_ON=1'b0;
    defparam \uart.r_Tx_Data_i3_LC_4_21_3 .SEQ_MODE=4'b1000;
    defparam \uart.r_Tx_Data_i3_LC_4_21_3 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \uart.r_Tx_Data_i3_LC_4_21_3  (
            .in0(N__4894),
            .in1(N__4823),
            .in2(_gnd_net_),
            .in3(N__4931),
            .lcout(r_Tx_Data_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__5394),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart.r_Tx_Data_i7_LC_4_21_5 .C_ON=1'b0;
    defparam \uart.r_Tx_Data_i7_LC_4_21_5 .SEQ_MODE=4'b1000;
    defparam \uart.r_Tx_Data_i7_LC_4_21_5 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \uart.r_Tx_Data_i7_LC_4_21_5  (
            .in0(N__4895),
            .in1(N__5492),
            .in2(_gnd_net_),
            .in3(N__4919),
            .lcout(r_Tx_Data_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__5394),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart.r_Tx_Data_i0_LC_4_21_6 .C_ON=1'b0;
    defparam \uart.r_Tx_Data_i0_LC_4_21_6 .SEQ_MODE=4'b1000;
    defparam \uart.r_Tx_Data_i0_LC_4_21_6 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \uart.r_Tx_Data_i0_LC_4_21_6  (
            .in0(N__4838),
            .in1(N__4891),
            .in2(_gnd_net_),
            .in3(N__4907),
            .lcout(r_Tx_Data_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__5394),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart.r_Tx_Data_i2_LC_4_21_7 .C_ON=1'b0;
    defparam \uart.r_Tx_Data_i2_LC_4_21_7 .SEQ_MODE=4'b1000;
    defparam \uart.r_Tx_Data_i2_LC_4_21_7 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \uart.r_Tx_Data_i2_LC_4_21_7  (
            .in0(N__4893),
            .in1(N__4796),
            .in2(_gnd_net_),
            .in3(N__4865),
            .lcout(r_Tx_Data_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__5394),
            .ce(),
            .sr(_gnd_net_));
    defparam data_out_i0_i5_LC_4_22_0.C_ON=1'b0;
    defparam data_out_i0_i5_LC_4_22_0.SEQ_MODE=4'b1000;
    defparam data_out_i0_i5_LC_4_22_0.LUT_INIT=16'b1110111001000100;
    LogicCell40 data_out_i0_i5_LC_4_22_0 (
            .in0(N__5705),
            .in1(N__4849),
            .in2(_gnd_net_),
            .in3(N__5870),
            .lcout(data_out_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__5774),
            .ce(),
            .sr(_gnd_net_));
    defparam data_out_i0_i0_LC_4_22_5.C_ON=1'b0;
    defparam data_out_i0_i0_LC_4_22_5.SEQ_MODE=4'b1000;
    defparam data_out_i0_i0_LC_4_22_5.LUT_INIT=16'b1100110010101010;
    LogicCell40 data_out_i0_i0_LC_4_22_5 (
            .in0(N__4834),
            .in1(N__5231),
            .in2(_gnd_net_),
            .in3(N__5703),
            .lcout(data_out_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__5774),
            .ce(),
            .sr(_gnd_net_));
    defparam data_out_i0_i3_LC_4_22_6.C_ON=1'b0;
    defparam data_out_i0_i3_LC_4_22_6.SEQ_MODE=4'b1000;
    defparam data_out_i0_i3_LC_4_22_6.LUT_INIT=16'b1110111001000100;
    LogicCell40 data_out_i0_i3_LC_4_22_6 (
            .in0(N__5704),
            .in1(N__4822),
            .in2(_gnd_net_),
            .in3(N__5900),
            .lcout(data_out_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__5774),
            .ce(),
            .sr(_gnd_net_));
    defparam data_out_i0_i1_LC_4_23_0.C_ON=1'b0;
    defparam data_out_i0_i1_LC_4_23_0.SEQ_MODE=4'b1000;
    defparam data_out_i0_i1_LC_4_23_0.LUT_INIT=16'b1100110010101010;
    LogicCell40 data_out_i0_i1_LC_4_23_0 (
            .in0(N__4807),
            .in1(N__5219),
            .in2(_gnd_net_),
            .in3(N__5700),
            .lcout(data_out_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__5805),
            .ce(),
            .sr(_gnd_net_));
    defparam data_out_i0_i2_LC_4_23_1.C_ON=1'b0;
    defparam data_out_i0_i2_LC_4_23_1.SEQ_MODE=4'b1000;
    defparam data_out_i0_i2_LC_4_23_1.LUT_INIT=16'b1110111001000100;
    LogicCell40 data_out_i0_i2_LC_4_23_1 (
            .in0(N__5701),
            .in1(N__4792),
            .in2(_gnd_net_),
            .in3(N__5915),
            .lcout(data_out_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__5805),
            .ce(),
            .sr(_gnd_net_));
    defparam i15_4_lut_LC_4_23_2.C_ON=1'b0;
    defparam i15_4_lut_LC_4_23_2.SEQ_MODE=4'b0000;
    defparam i15_4_lut_LC_4_23_2.LUT_INIT=16'b1111111111111110;
    LogicCell40 i15_4_lut_LC_4_23_2 (
            .in0(N__5204),
            .in1(N__5188),
            .in2(N__5177),
            .in3(N__5161),
            .lcout(),
            .ltout(n38_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i21_4_lut_LC_4_23_3.C_ON=1'b0;
    defparam i21_4_lut_LC_4_23_3.SEQ_MODE=4'b0000;
    defparam i21_4_lut_LC_4_23_3.LUT_INIT=16'b1111111111111110;
    LogicCell40 i21_4_lut_LC_4_23_3 (
            .in0(N__5006),
            .in1(N__5540),
            .in2(N__5150),
            .in3(N__5498),
            .lcout(n44),
            .ltout(n44_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i710_4_lut_LC_4_23_4.C_ON=1'b0;
    defparam i710_4_lut_LC_4_23_4.SEQ_MODE=4'b0000;
    defparam i710_4_lut_LC_4_23_4.LUT_INIT=16'b0011001100110010;
    LogicCell40 i710_4_lut_LC_4_23_4 (
            .in0(N__5599),
            .in1(N__5125),
            .in2(N__5147),
            .in3(N__4945),
            .lcout(counter_31__N_172),
            .ltout(counter_31__N_172_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam data_out_i0_i4_LC_4_23_5.C_ON=1'b0;
    defparam data_out_i0_i4_LC_4_23_5.SEQ_MODE=4'b1000;
    defparam data_out_i0_i4_LC_4_23_5.LUT_INIT=16'b1111110000001100;
    LogicCell40 data_out_i0_i4_LC_4_23_5 (
            .in0(_gnd_net_),
            .in1(N__5137),
            .in2(N__5144),
            .in3(N__5885),
            .lcout(data_out_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__5805),
            .ce(),
            .sr(_gnd_net_));
    defparam send_29_LC_4_23_6.C_ON=1'b0;
    defparam send_29_LC_4_23_6.SEQ_MODE=4'b1000;
    defparam send_29_LC_4_23_6.LUT_INIT=16'b0011001100110010;
    LogicCell40 send_29_LC_4_23_6 (
            .in0(N__5600),
            .in1(N__5126),
            .in2(N__4949),
            .in3(N__5105),
            .lcout(r_SM_Main_2_N_236_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__5805),
            .ce(),
            .sr(_gnd_net_));
    defparam data_out_i0_i6_LC_4_23_7.C_ON=1'b0;
    defparam data_out_i0_i6_LC_4_23_7.SEQ_MODE=4'b1000;
    defparam data_out_i0_i6_LC_4_23_7.LUT_INIT=16'b1110111001000100;
    LogicCell40 data_out_i0_i6_LC_4_23_7 (
            .in0(N__5702),
            .in1(N__5068),
            .in2(_gnd_net_),
            .in3(N__5855),
            .lcout(data_out_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__5805),
            .ce(),
            .sr(_gnd_net_));
    defparam i13_4_lut_LC_4_24_0.C_ON=1'b0;
    defparam i13_4_lut_LC_4_24_0.SEQ_MODE=4'b0000;
    defparam i13_4_lut_LC_4_24_0.LUT_INIT=16'b1111111111111110;
    LogicCell40 i13_4_lut_LC_4_24_0 (
            .in0(N__5056),
            .in1(N__5044),
            .in2(N__5033),
            .in3(N__5017),
            .lcout(n36),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i17_4_lut_LC_4_24_3.C_ON=1'b0;
    defparam i17_4_lut_LC_4_24_3.SEQ_MODE=4'b0000;
    defparam i17_4_lut_LC_4_24_3.LUT_INIT=16'b1111111111111110;
    LogicCell40 i17_4_lut_LC_4_24_3 (
            .in0(N__4999),
            .in1(N__4987),
            .in2(N__4976),
            .in3(N__4960),
            .lcout(n40),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i16_4_lut_LC_4_24_4.C_ON=1'b0;
    defparam i16_4_lut_LC_4_24_4.SEQ_MODE=4'b0000;
    defparam i16_4_lut_LC_4_24_4.LUT_INIT=16'b1111111111111110;
    LogicCell40 i16_4_lut_LC_4_24_4 (
            .in0(N__5650),
            .in1(N__5638),
            .in2(N__5627),
            .in3(N__5611),
            .lcout(n39),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i14_4_lut_LC_4_24_5.C_ON=1'b0;
    defparam i14_4_lut_LC_4_24_5.SEQ_MODE=4'b0000;
    defparam i14_4_lut_LC_4_24_5.LUT_INIT=16'b1111111111111110;
    LogicCell40 i14_4_lut_LC_4_24_5 (
            .in0(N__5590),
            .in1(N__5578),
            .in2(N__5567),
            .in3(N__5551),
            .lcout(n37),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12_3_lut_LC_4_24_6.C_ON=1'b0;
    defparam i12_3_lut_LC_4_24_6.SEQ_MODE=4'b0000;
    defparam i12_3_lut_LC_4_24_6.LUT_INIT=16'b1111111111101110;
    LogicCell40 i12_3_lut_LC_4_24_6 (
            .in0(N__5533),
            .in1(N__5521),
            .in2(_gnd_net_),
            .in3(N__5509),
            .lcout(n35),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam data_out_i0_i7_LC_4_24_7.C_ON=1'b0;
    defparam data_out_i0_i7_LC_4_24_7.SEQ_MODE=4'b1000;
    defparam data_out_i0_i7_LC_4_24_7.LUT_INIT=16'b1010101011001100;
    LogicCell40 data_out_i0_i7_LC_4_24_7 (
            .in0(N__5836),
            .in1(N__5488),
            .in2(_gnd_net_),
            .in3(N__5706),
            .lcout(data_out_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__5804),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart.r_Bit_Index_i1_LC_5_19_1 .C_ON=1'b0;
    defparam \uart.r_Bit_Index_i1_LC_5_19_1 .SEQ_MODE=4'b1000;
    defparam \uart.r_Bit_Index_i1_LC_5_19_1 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \uart.r_Bit_Index_i1_LC_5_19_1  (
            .in0(_gnd_net_),
            .in1(N__5438),
            .in2(_gnd_net_),
            .in3(N__5476),
            .lcout(\uart.r_Bit_Index_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__5391),
            .ce(N__5330),
            .sr(N__5303));
    defparam integrator_118__i0_LC_5_23_0.C_ON=1'b1;
    defparam integrator_118__i0_LC_5_23_0.SEQ_MODE=4'b1000;
    defparam integrator_118__i0_LC_5_23_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 integrator_118__i0_LC_5_23_0 (
            .in0(_gnd_net_),
            .in1(N__5230),
            .in2(N__5275),
            .in3(_gnd_net_),
            .lcout(integrator_0),
            .ltout(),
            .carryin(bfn_5_23_0_),
            .carryout(n2188),
            .clk(N__5815),
            .ce(),
            .sr(N__5708));
    defparam integrator_118__i1_LC_5_23_1.C_ON=1'b1;
    defparam integrator_118__i1_LC_5_23_1.SEQ_MODE=4'b1000;
    defparam integrator_118__i1_LC_5_23_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 integrator_118__i1_LC_5_23_1 (
            .in0(_gnd_net_),
            .in1(N__5218),
            .in2(_gnd_net_),
            .in3(N__5207),
            .lcout(integrator_1),
            .ltout(),
            .carryin(n2188),
            .carryout(n2189),
            .clk(N__5815),
            .ce(),
            .sr(N__5708));
    defparam integrator_118__i2_LC_5_23_2.C_ON=1'b1;
    defparam integrator_118__i2_LC_5_23_2.SEQ_MODE=4'b1000;
    defparam integrator_118__i2_LC_5_23_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 integrator_118__i2_LC_5_23_2 (
            .in0(_gnd_net_),
            .in1(N__5914),
            .in2(_gnd_net_),
            .in3(N__5903),
            .lcout(integrator_2),
            .ltout(),
            .carryin(n2189),
            .carryout(n2190),
            .clk(N__5815),
            .ce(),
            .sr(N__5708));
    defparam integrator_118__i3_LC_5_23_3.C_ON=1'b1;
    defparam integrator_118__i3_LC_5_23_3.SEQ_MODE=4'b1000;
    defparam integrator_118__i3_LC_5_23_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 integrator_118__i3_LC_5_23_3 (
            .in0(_gnd_net_),
            .in1(N__5899),
            .in2(_gnd_net_),
            .in3(N__5888),
            .lcout(integrator_3),
            .ltout(),
            .carryin(n2190),
            .carryout(n2191),
            .clk(N__5815),
            .ce(),
            .sr(N__5708));
    defparam integrator_118__i4_LC_5_23_4.C_ON=1'b1;
    defparam integrator_118__i4_LC_5_23_4.SEQ_MODE=4'b1000;
    defparam integrator_118__i4_LC_5_23_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 integrator_118__i4_LC_5_23_4 (
            .in0(_gnd_net_),
            .in1(N__5884),
            .in2(_gnd_net_),
            .in3(N__5873),
            .lcout(integrator_4),
            .ltout(),
            .carryin(n2191),
            .carryout(n2192),
            .clk(N__5815),
            .ce(),
            .sr(N__5708));
    defparam integrator_118__i5_LC_5_23_5.C_ON=1'b1;
    defparam integrator_118__i5_LC_5_23_5.SEQ_MODE=4'b1000;
    defparam integrator_118__i5_LC_5_23_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 integrator_118__i5_LC_5_23_5 (
            .in0(_gnd_net_),
            .in1(N__5869),
            .in2(_gnd_net_),
            .in3(N__5858),
            .lcout(integrator_5),
            .ltout(),
            .carryin(n2192),
            .carryout(n2193),
            .clk(N__5815),
            .ce(),
            .sr(N__5708));
    defparam integrator_118__i6_LC_5_23_6.C_ON=1'b1;
    defparam integrator_118__i6_LC_5_23_6.SEQ_MODE=4'b1000;
    defparam integrator_118__i6_LC_5_23_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 integrator_118__i6_LC_5_23_6 (
            .in0(_gnd_net_),
            .in1(N__5854),
            .in2(_gnd_net_),
            .in3(N__5843),
            .lcout(integrator_6),
            .ltout(),
            .carryin(n2193),
            .carryout(n2194),
            .clk(N__5815),
            .ce(),
            .sr(N__5708));
    defparam integrator_118__i7_LC_5_23_7.C_ON=1'b0;
    defparam integrator_118__i7_LC_5_23_7.SEQ_MODE=4'b1000;
    defparam integrator_118__i7_LC_5_23_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 integrator_118__i7_LC_5_23_7 (
            .in0(_gnd_net_),
            .in1(N__5837),
            .in2(_gnd_net_),
            .in3(N__5840),
            .lcout(integrator_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__5815),
            .ce(),
            .sr(N__5708));
endmodule // TinyFPGA_B
