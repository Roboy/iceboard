-- ******************************************************************************

-- iCEcube Netlister

-- Version:            2017.08.27940

-- Build Date:         Sep 12 2017 08:26:01

-- File Generated:     Feb 24 2020 16:03:39

-- Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

-- Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

-- ******************************************************************************

-- VHDL file for cell "TinyFPGA_B" view "INTERFACE"

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library ice;
use ice.vcomponent_vital.all;

-- Entity of TinyFPGA_B
entity TinyFPGA_B is
port (
    USBPU : inout std_logic;
    TX : inout std_logic;
    SDA : inout std_logic;
    SCL : inout std_logic;
    RX : inout std_logic;
    NEOPXL : out std_logic;
    LED : out std_logic;
    INLC : inout std_logic;
    INLB : inout std_logic;
    INLA : inout std_logic;
    INHC : inout std_logic;
    INHB : inout std_logic;
    INHA : inout std_logic;
    HALL3 : inout std_logic;
    HALL2 : inout std_logic;
    HALL1 : inout std_logic;
    FAULT_N : inout std_logic;
    ENCODER1_B : inout std_logic;
    ENCODER1_A : inout std_logic;
    ENCODER0_B : inout std_logic;
    ENCODER0_A : inout std_logic;
    DE : inout std_logic;
    CS_MISO : inout std_logic;
    CS_CLK : inout std_logic;
    CS : inout std_logic;
    CLK : in std_logic);
end TinyFPGA_B;

-- Architecture of TinyFPGA_B
-- View name is \INTERFACE\
architecture \INTERFACE\ of TinyFPGA_B is

signal \N__47950\ : std_logic;
signal \N__47949\ : std_logic;
signal \N__47948\ : std_logic;
signal \N__47941\ : std_logic;
signal \N__47940\ : std_logic;
signal \N__47939\ : std_logic;
signal \N__47932\ : std_logic;
signal \N__47931\ : std_logic;
signal \N__47930\ : std_logic;
signal \N__47923\ : std_logic;
signal \N__47922\ : std_logic;
signal \N__47921\ : std_logic;
signal \N__47914\ : std_logic;
signal \N__47913\ : std_logic;
signal \N__47912\ : std_logic;
signal \N__47905\ : std_logic;
signal \N__47904\ : std_logic;
signal \N__47903\ : std_logic;
signal \N__47896\ : std_logic;
signal \N__47895\ : std_logic;
signal \N__47894\ : std_logic;
signal \N__47887\ : std_logic;
signal \N__47886\ : std_logic;
signal \N__47885\ : std_logic;
signal \N__47878\ : std_logic;
signal \N__47877\ : std_logic;
signal \N__47876\ : std_logic;
signal \N__47869\ : std_logic;
signal \N__47868\ : std_logic;
signal \N__47867\ : std_logic;
signal \N__47860\ : std_logic;
signal \N__47859\ : std_logic;
signal \N__47858\ : std_logic;
signal \N__47851\ : std_logic;
signal \N__47850\ : std_logic;
signal \N__47849\ : std_logic;
signal \N__47842\ : std_logic;
signal \N__47841\ : std_logic;
signal \N__47840\ : std_logic;
signal \N__47833\ : std_logic;
signal \N__47832\ : std_logic;
signal \N__47831\ : std_logic;
signal \N__47824\ : std_logic;
signal \N__47823\ : std_logic;
signal \N__47822\ : std_logic;
signal \N__47815\ : std_logic;
signal \N__47814\ : std_logic;
signal \N__47813\ : std_logic;
signal \N__47806\ : std_logic;
signal \N__47805\ : std_logic;
signal \N__47804\ : std_logic;
signal \N__47797\ : std_logic;
signal \N__47796\ : std_logic;
signal \N__47795\ : std_logic;
signal \N__47788\ : std_logic;
signal \N__47787\ : std_logic;
signal \N__47786\ : std_logic;
signal \N__47779\ : std_logic;
signal \N__47778\ : std_logic;
signal \N__47777\ : std_logic;
signal \N__47770\ : std_logic;
signal \N__47769\ : std_logic;
signal \N__47768\ : std_logic;
signal \N__47761\ : std_logic;
signal \N__47760\ : std_logic;
signal \N__47759\ : std_logic;
signal \N__47752\ : std_logic;
signal \N__47751\ : std_logic;
signal \N__47750\ : std_logic;
signal \N__47743\ : std_logic;
signal \N__47742\ : std_logic;
signal \N__47741\ : std_logic;
signal \N__47734\ : std_logic;
signal \N__47733\ : std_logic;
signal \N__47732\ : std_logic;
signal \N__47725\ : std_logic;
signal \N__47724\ : std_logic;
signal \N__47723\ : std_logic;
signal \N__47706\ : std_logic;
signal \N__47703\ : std_logic;
signal \N__47700\ : std_logic;
signal \N__47697\ : std_logic;
signal \N__47696\ : std_logic;
signal \N__47695\ : std_logic;
signal \N__47694\ : std_logic;
signal \N__47693\ : std_logic;
signal \N__47690\ : std_logic;
signal \N__47687\ : std_logic;
signal \N__47684\ : std_logic;
signal \N__47681\ : std_logic;
signal \N__47678\ : std_logic;
signal \N__47677\ : std_logic;
signal \N__47676\ : std_logic;
signal \N__47675\ : std_logic;
signal \N__47674\ : std_logic;
signal \N__47673\ : std_logic;
signal \N__47672\ : std_logic;
signal \N__47669\ : std_logic;
signal \N__47668\ : std_logic;
signal \N__47667\ : std_logic;
signal \N__47666\ : std_logic;
signal \N__47665\ : std_logic;
signal \N__47664\ : std_logic;
signal \N__47663\ : std_logic;
signal \N__47660\ : std_logic;
signal \N__47659\ : std_logic;
signal \N__47658\ : std_logic;
signal \N__47657\ : std_logic;
signal \N__47654\ : std_logic;
signal \N__47651\ : std_logic;
signal \N__47648\ : std_logic;
signal \N__47647\ : std_logic;
signal \N__47646\ : std_logic;
signal \N__47643\ : std_logic;
signal \N__47642\ : std_logic;
signal \N__47641\ : std_logic;
signal \N__47638\ : std_logic;
signal \N__47637\ : std_logic;
signal \N__47636\ : std_logic;
signal \N__47635\ : std_logic;
signal \N__47632\ : std_logic;
signal \N__47631\ : std_logic;
signal \N__47628\ : std_logic;
signal \N__47625\ : std_logic;
signal \N__47624\ : std_logic;
signal \N__47621\ : std_logic;
signal \N__47618\ : std_logic;
signal \N__47611\ : std_logic;
signal \N__47610\ : std_logic;
signal \N__47607\ : std_logic;
signal \N__47604\ : std_logic;
signal \N__47601\ : std_logic;
signal \N__47600\ : std_logic;
signal \N__47599\ : std_logic;
signal \N__47598\ : std_logic;
signal \N__47595\ : std_logic;
signal \N__47594\ : std_logic;
signal \N__47591\ : std_logic;
signal \N__47590\ : std_logic;
signal \N__47587\ : std_logic;
signal \N__47586\ : std_logic;
signal \N__47585\ : std_logic;
signal \N__47584\ : std_logic;
signal \N__47583\ : std_logic;
signal \N__47582\ : std_logic;
signal \N__47581\ : std_logic;
signal \N__47578\ : std_logic;
signal \N__47577\ : std_logic;
signal \N__47570\ : std_logic;
signal \N__47563\ : std_logic;
signal \N__47560\ : std_logic;
signal \N__47555\ : std_logic;
signal \N__47550\ : std_logic;
signal \N__47549\ : std_logic;
signal \N__47546\ : std_logic;
signal \N__47543\ : std_logic;
signal \N__47540\ : std_logic;
signal \N__47539\ : std_logic;
signal \N__47536\ : std_logic;
signal \N__47533\ : std_logic;
signal \N__47530\ : std_logic;
signal \N__47523\ : std_logic;
signal \N__47520\ : std_logic;
signal \N__47519\ : std_logic;
signal \N__47518\ : std_logic;
signal \N__47517\ : std_logic;
signal \N__47516\ : std_logic;
signal \N__47515\ : std_logic;
signal \N__47514\ : std_logic;
signal \N__47509\ : std_logic;
signal \N__47506\ : std_logic;
signal \N__47503\ : std_logic;
signal \N__47502\ : std_logic;
signal \N__47499\ : std_logic;
signal \N__47496\ : std_logic;
signal \N__47493\ : std_logic;
signal \N__47490\ : std_logic;
signal \N__47489\ : std_logic;
signal \N__47488\ : std_logic;
signal \N__47485\ : std_logic;
signal \N__47484\ : std_logic;
signal \N__47483\ : std_logic;
signal \N__47482\ : std_logic;
signal \N__47481\ : std_logic;
signal \N__47480\ : std_logic;
signal \N__47479\ : std_logic;
signal \N__47478\ : std_logic;
signal \N__47475\ : std_logic;
signal \N__47470\ : std_logic;
signal \N__47461\ : std_logic;
signal \N__47460\ : std_logic;
signal \N__47459\ : std_logic;
signal \N__47456\ : std_logic;
signal \N__47453\ : std_logic;
signal \N__47450\ : std_logic;
signal \N__47447\ : std_logic;
signal \N__47444\ : std_logic;
signal \N__47437\ : std_logic;
signal \N__47432\ : std_logic;
signal \N__47431\ : std_logic;
signal \N__47428\ : std_logic;
signal \N__47425\ : std_logic;
signal \N__47422\ : std_logic;
signal \N__47415\ : std_logic;
signal \N__47412\ : std_logic;
signal \N__47407\ : std_logic;
signal \N__47402\ : std_logic;
signal \N__47397\ : std_logic;
signal \N__47394\ : std_logic;
signal \N__47391\ : std_logic;
signal \N__47388\ : std_logic;
signal \N__47385\ : std_logic;
signal \N__47380\ : std_logic;
signal \N__47377\ : std_logic;
signal \N__47372\ : std_logic;
signal \N__47369\ : std_logic;
signal \N__47368\ : std_logic;
signal \N__47367\ : std_logic;
signal \N__47364\ : std_logic;
signal \N__47363\ : std_logic;
signal \N__47360\ : std_logic;
signal \N__47355\ : std_logic;
signal \N__47350\ : std_logic;
signal \N__47347\ : std_logic;
signal \N__47344\ : std_logic;
signal \N__47341\ : std_logic;
signal \N__47336\ : std_logic;
signal \N__47333\ : std_logic;
signal \N__47330\ : std_logic;
signal \N__47329\ : std_logic;
signal \N__47326\ : std_logic;
signal \N__47325\ : std_logic;
signal \N__47324\ : std_logic;
signal \N__47323\ : std_logic;
signal \N__47318\ : std_logic;
signal \N__47315\ : std_logic;
signal \N__47308\ : std_logic;
signal \N__47305\ : std_logic;
signal \N__47302\ : std_logic;
signal \N__47301\ : std_logic;
signal \N__47300\ : std_logic;
signal \N__47299\ : std_logic;
signal \N__47296\ : std_logic;
signal \N__47277\ : std_logic;
signal \N__47272\ : std_logic;
signal \N__47269\ : std_logic;
signal \N__47264\ : std_logic;
signal \N__47259\ : std_logic;
signal \N__47256\ : std_logic;
signal \N__47251\ : std_logic;
signal \N__47234\ : std_logic;
signal \N__47229\ : std_logic;
signal \N__47226\ : std_logic;
signal \N__47221\ : std_logic;
signal \N__47218\ : std_logic;
signal \N__47215\ : std_logic;
signal \N__47208\ : std_logic;
signal \N__47199\ : std_logic;
signal \N__47194\ : std_logic;
signal \N__47183\ : std_logic;
signal \N__47176\ : std_logic;
signal \N__47157\ : std_logic;
signal \N__47156\ : std_logic;
signal \N__47155\ : std_logic;
signal \N__47154\ : std_logic;
signal \N__47153\ : std_logic;
signal \N__47150\ : std_logic;
signal \N__47149\ : std_logic;
signal \N__47148\ : std_logic;
signal \N__47147\ : std_logic;
signal \N__47146\ : std_logic;
signal \N__47143\ : std_logic;
signal \N__47140\ : std_logic;
signal \N__47137\ : std_logic;
signal \N__47134\ : std_logic;
signal \N__47131\ : std_logic;
signal \N__47130\ : std_logic;
signal \N__47127\ : std_logic;
signal \N__47126\ : std_logic;
signal \N__47125\ : std_logic;
signal \N__47124\ : std_logic;
signal \N__47123\ : std_logic;
signal \N__47122\ : std_logic;
signal \N__47121\ : std_logic;
signal \N__47120\ : std_logic;
signal \N__47119\ : std_logic;
signal \N__47116\ : std_logic;
signal \N__47113\ : std_logic;
signal \N__47110\ : std_logic;
signal \N__47107\ : std_logic;
signal \N__47102\ : std_logic;
signal \N__47099\ : std_logic;
signal \N__47096\ : std_logic;
signal \N__47093\ : std_logic;
signal \N__47090\ : std_logic;
signal \N__47085\ : std_logic;
signal \N__47082\ : std_logic;
signal \N__47079\ : std_logic;
signal \N__47076\ : std_logic;
signal \N__47073\ : std_logic;
signal \N__47072\ : std_logic;
signal \N__47069\ : std_logic;
signal \N__47066\ : std_logic;
signal \N__47061\ : std_logic;
signal \N__47058\ : std_logic;
signal \N__47053\ : std_logic;
signal \N__47048\ : std_logic;
signal \N__47043\ : std_logic;
signal \N__47040\ : std_logic;
signal \N__47039\ : std_logic;
signal \N__47038\ : std_logic;
signal \N__47037\ : std_logic;
signal \N__47034\ : std_logic;
signal \N__47031\ : std_logic;
signal \N__47028\ : std_logic;
signal \N__47025\ : std_logic;
signal \N__47022\ : std_logic;
signal \N__47019\ : std_logic;
signal \N__47014\ : std_logic;
signal \N__47005\ : std_logic;
signal \N__47002\ : std_logic;
signal \N__46999\ : std_logic;
signal \N__46996\ : std_logic;
signal \N__46993\ : std_logic;
signal \N__46990\ : std_logic;
signal \N__46985\ : std_logic;
signal \N__46982\ : std_logic;
signal \N__46975\ : std_logic;
signal \N__46972\ : std_logic;
signal \N__46969\ : std_logic;
signal \N__46950\ : std_logic;
signal \N__46947\ : std_logic;
signal \N__46944\ : std_logic;
signal \N__46941\ : std_logic;
signal \N__46938\ : std_logic;
signal \N__46935\ : std_logic;
signal \N__46934\ : std_logic;
signal \N__46931\ : std_logic;
signal \N__46928\ : std_logic;
signal \N__46923\ : std_logic;
signal \N__46922\ : std_logic;
signal \N__46921\ : std_logic;
signal \N__46920\ : std_logic;
signal \N__46919\ : std_logic;
signal \N__46918\ : std_logic;
signal \N__46917\ : std_logic;
signal \N__46916\ : std_logic;
signal \N__46915\ : std_logic;
signal \N__46914\ : std_logic;
signal \N__46913\ : std_logic;
signal \N__46912\ : std_logic;
signal \N__46911\ : std_logic;
signal \N__46910\ : std_logic;
signal \N__46909\ : std_logic;
signal \N__46908\ : std_logic;
signal \N__46907\ : std_logic;
signal \N__46906\ : std_logic;
signal \N__46905\ : std_logic;
signal \N__46904\ : std_logic;
signal \N__46903\ : std_logic;
signal \N__46902\ : std_logic;
signal \N__46901\ : std_logic;
signal \N__46900\ : std_logic;
signal \N__46899\ : std_logic;
signal \N__46898\ : std_logic;
signal \N__46897\ : std_logic;
signal \N__46896\ : std_logic;
signal \N__46895\ : std_logic;
signal \N__46894\ : std_logic;
signal \N__46893\ : std_logic;
signal \N__46892\ : std_logic;
signal \N__46891\ : std_logic;
signal \N__46890\ : std_logic;
signal \N__46889\ : std_logic;
signal \N__46888\ : std_logic;
signal \N__46887\ : std_logic;
signal \N__46886\ : std_logic;
signal \N__46885\ : std_logic;
signal \N__46884\ : std_logic;
signal \N__46883\ : std_logic;
signal \N__46882\ : std_logic;
signal \N__46881\ : std_logic;
signal \N__46880\ : std_logic;
signal \N__46879\ : std_logic;
signal \N__46878\ : std_logic;
signal \N__46877\ : std_logic;
signal \N__46876\ : std_logic;
signal \N__46875\ : std_logic;
signal \N__46874\ : std_logic;
signal \N__46873\ : std_logic;
signal \N__46872\ : std_logic;
signal \N__46871\ : std_logic;
signal \N__46870\ : std_logic;
signal \N__46869\ : std_logic;
signal \N__46868\ : std_logic;
signal \N__46867\ : std_logic;
signal \N__46866\ : std_logic;
signal \N__46865\ : std_logic;
signal \N__46864\ : std_logic;
signal \N__46863\ : std_logic;
signal \N__46862\ : std_logic;
signal \N__46861\ : std_logic;
signal \N__46860\ : std_logic;
signal \N__46859\ : std_logic;
signal \N__46858\ : std_logic;
signal \N__46857\ : std_logic;
signal \N__46856\ : std_logic;
signal \N__46855\ : std_logic;
signal \N__46854\ : std_logic;
signal \N__46853\ : std_logic;
signal \N__46852\ : std_logic;
signal \N__46851\ : std_logic;
signal \N__46850\ : std_logic;
signal \N__46849\ : std_logic;
signal \N__46848\ : std_logic;
signal \N__46847\ : std_logic;
signal \N__46846\ : std_logic;
signal \N__46845\ : std_logic;
signal \N__46844\ : std_logic;
signal \N__46843\ : std_logic;
signal \N__46842\ : std_logic;
signal \N__46841\ : std_logic;
signal \N__46840\ : std_logic;
signal \N__46839\ : std_logic;
signal \N__46668\ : std_logic;
signal \N__46665\ : std_logic;
signal \N__46662\ : std_logic;
signal \N__46659\ : std_logic;
signal \N__46656\ : std_logic;
signal \N__46653\ : std_logic;
signal \N__46650\ : std_logic;
signal \N__46647\ : std_logic;
signal \N__46644\ : std_logic;
signal \N__46641\ : std_logic;
signal \N__46638\ : std_logic;
signal \N__46635\ : std_logic;
signal \N__46632\ : std_logic;
signal \N__46629\ : std_logic;
signal \N__46626\ : std_logic;
signal \N__46623\ : std_logic;
signal \N__46620\ : std_logic;
signal \N__46617\ : std_logic;
signal \N__46614\ : std_logic;
signal \N__46611\ : std_logic;
signal \N__46608\ : std_logic;
signal \N__46605\ : std_logic;
signal \N__46602\ : std_logic;
signal \N__46599\ : std_logic;
signal \N__46596\ : std_logic;
signal \N__46593\ : std_logic;
signal \N__46590\ : std_logic;
signal \N__46587\ : std_logic;
signal \N__46584\ : std_logic;
signal \N__46581\ : std_logic;
signal \N__46578\ : std_logic;
signal \N__46575\ : std_logic;
signal \N__46572\ : std_logic;
signal \N__46571\ : std_logic;
signal \N__46568\ : std_logic;
signal \N__46567\ : std_logic;
signal \N__46566\ : std_logic;
signal \N__46565\ : std_logic;
signal \N__46564\ : std_logic;
signal \N__46563\ : std_logic;
signal \N__46560\ : std_logic;
signal \N__46559\ : std_logic;
signal \N__46556\ : std_logic;
signal \N__46555\ : std_logic;
signal \N__46552\ : std_logic;
signal \N__46549\ : std_logic;
signal \N__46546\ : std_logic;
signal \N__46545\ : std_logic;
signal \N__46542\ : std_logic;
signal \N__46539\ : std_logic;
signal \N__46536\ : std_logic;
signal \N__46533\ : std_logic;
signal \N__46530\ : std_logic;
signal \N__46527\ : std_logic;
signal \N__46524\ : std_logic;
signal \N__46523\ : std_logic;
signal \N__46522\ : std_logic;
signal \N__46517\ : std_logic;
signal \N__46514\ : std_logic;
signal \N__46513\ : std_logic;
signal \N__46512\ : std_logic;
signal \N__46511\ : std_logic;
signal \N__46510\ : std_logic;
signal \N__46509\ : std_logic;
signal \N__46508\ : std_logic;
signal \N__46505\ : std_logic;
signal \N__46498\ : std_logic;
signal \N__46491\ : std_logic;
signal \N__46486\ : std_logic;
signal \N__46481\ : std_logic;
signal \N__46478\ : std_logic;
signal \N__46473\ : std_logic;
signal \N__46470\ : std_logic;
signal \N__46467\ : std_logic;
signal \N__46464\ : std_logic;
signal \N__46459\ : std_logic;
signal \N__46454\ : std_logic;
signal \N__46451\ : std_logic;
signal \N__46448\ : std_logic;
signal \N__46445\ : std_logic;
signal \N__46428\ : std_logic;
signal \N__46425\ : std_logic;
signal \N__46422\ : std_logic;
signal \N__46419\ : std_logic;
signal \N__46416\ : std_logic;
signal \N__46413\ : std_logic;
signal \N__46412\ : std_logic;
signal \N__46411\ : std_logic;
signal \N__46410\ : std_logic;
signal \N__46409\ : std_logic;
signal \N__46408\ : std_logic;
signal \N__46407\ : std_logic;
signal \N__46406\ : std_logic;
signal \N__46405\ : std_logic;
signal \N__46402\ : std_logic;
signal \N__46397\ : std_logic;
signal \N__46396\ : std_logic;
signal \N__46393\ : std_logic;
signal \N__46392\ : std_logic;
signal \N__46387\ : std_logic;
signal \N__46386\ : std_logic;
signal \N__46385\ : std_logic;
signal \N__46384\ : std_logic;
signal \N__46383\ : std_logic;
signal \N__46378\ : std_logic;
signal \N__46375\ : std_logic;
signal \N__46372\ : std_logic;
signal \N__46369\ : std_logic;
signal \N__46366\ : std_logic;
signal \N__46363\ : std_logic;
signal \N__46360\ : std_logic;
signal \N__46357\ : std_logic;
signal \N__46352\ : std_logic;
signal \N__46349\ : std_logic;
signal \N__46346\ : std_logic;
signal \N__46345\ : std_logic;
signal \N__46344\ : std_logic;
signal \N__46343\ : std_logic;
signal \N__46338\ : std_logic;
signal \N__46337\ : std_logic;
signal \N__46336\ : std_logic;
signal \N__46335\ : std_logic;
signal \N__46332\ : std_logic;
signal \N__46329\ : std_logic;
signal \N__46324\ : std_logic;
signal \N__46323\ : std_logic;
signal \N__46322\ : std_logic;
signal \N__46321\ : std_logic;
signal \N__46320\ : std_logic;
signal \N__46315\ : std_logic;
signal \N__46308\ : std_logic;
signal \N__46303\ : std_logic;
signal \N__46300\ : std_logic;
signal \N__46297\ : std_logic;
signal \N__46294\ : std_logic;
signal \N__46289\ : std_logic;
signal \N__46284\ : std_logic;
signal \N__46281\ : std_logic;
signal \N__46278\ : std_logic;
signal \N__46275\ : std_logic;
signal \N__46272\ : std_logic;
signal \N__46269\ : std_logic;
signal \N__46264\ : std_logic;
signal \N__46257\ : std_logic;
signal \N__46248\ : std_logic;
signal \N__46233\ : std_logic;
signal \N__46230\ : std_logic;
signal \N__46227\ : std_logic;
signal \N__46224\ : std_logic;
signal \N__46221\ : std_logic;
signal \N__46218\ : std_logic;
signal \N__46215\ : std_logic;
signal \N__46212\ : std_logic;
signal \N__46209\ : std_logic;
signal \N__46206\ : std_logic;
signal \N__46203\ : std_logic;
signal \N__46200\ : std_logic;
signal \N__46197\ : std_logic;
signal \N__46194\ : std_logic;
signal \N__46191\ : std_logic;
signal \N__46188\ : std_logic;
signal \N__46185\ : std_logic;
signal \N__46182\ : std_logic;
signal \N__46179\ : std_logic;
signal \N__46176\ : std_logic;
signal \N__46173\ : std_logic;
signal \N__46170\ : std_logic;
signal \N__46167\ : std_logic;
signal \N__46166\ : std_logic;
signal \N__46165\ : std_logic;
signal \N__46162\ : std_logic;
signal \N__46157\ : std_logic;
signal \N__46152\ : std_logic;
signal \N__46151\ : std_logic;
signal \N__46148\ : std_logic;
signal \N__46147\ : std_logic;
signal \N__46146\ : std_logic;
signal \N__46145\ : std_logic;
signal \N__46144\ : std_logic;
signal \N__46143\ : std_logic;
signal \N__46142\ : std_logic;
signal \N__46141\ : std_logic;
signal \N__46140\ : std_logic;
signal \N__46139\ : std_logic;
signal \N__46138\ : std_logic;
signal \N__46137\ : std_logic;
signal \N__46136\ : std_logic;
signal \N__46133\ : std_logic;
signal \N__46132\ : std_logic;
signal \N__46129\ : std_logic;
signal \N__46126\ : std_logic;
signal \N__46121\ : std_logic;
signal \N__46118\ : std_logic;
signal \N__46115\ : std_logic;
signal \N__46112\ : std_logic;
signal \N__46111\ : std_logic;
signal \N__46110\ : std_logic;
signal \N__46107\ : std_logic;
signal \N__46104\ : std_logic;
signal \N__46099\ : std_logic;
signal \N__46098\ : std_logic;
signal \N__46097\ : std_logic;
signal \N__46096\ : std_logic;
signal \N__46095\ : std_logic;
signal \N__46094\ : std_logic;
signal \N__46089\ : std_logic;
signal \N__46086\ : std_logic;
signal \N__46083\ : std_logic;
signal \N__46080\ : std_logic;
signal \N__46077\ : std_logic;
signal \N__46074\ : std_logic;
signal \N__46067\ : std_logic;
signal \N__46064\ : std_logic;
signal \N__46061\ : std_logic;
signal \N__46054\ : std_logic;
signal \N__46049\ : std_logic;
signal \N__46046\ : std_logic;
signal \N__46041\ : std_logic;
signal \N__46026\ : std_logic;
signal \N__46019\ : std_logic;
signal \N__46008\ : std_logic;
signal \N__46005\ : std_logic;
signal \N__46002\ : std_logic;
signal \N__45999\ : std_logic;
signal \N__45996\ : std_logic;
signal \N__45995\ : std_logic;
signal \N__45994\ : std_logic;
signal \N__45993\ : std_logic;
signal \N__45992\ : std_logic;
signal \N__45987\ : std_logic;
signal \N__45982\ : std_logic;
signal \N__45981\ : std_logic;
signal \N__45980\ : std_logic;
signal \N__45979\ : std_logic;
signal \N__45978\ : std_logic;
signal \N__45975\ : std_logic;
signal \N__45974\ : std_logic;
signal \N__45973\ : std_logic;
signal \N__45972\ : std_logic;
signal \N__45971\ : std_logic;
signal \N__45970\ : std_logic;
signal \N__45965\ : std_logic;
signal \N__45962\ : std_logic;
signal \N__45961\ : std_logic;
signal \N__45960\ : std_logic;
signal \N__45959\ : std_logic;
signal \N__45958\ : std_logic;
signal \N__45957\ : std_logic;
signal \N__45956\ : std_logic;
signal \N__45953\ : std_logic;
signal \N__45952\ : std_logic;
signal \N__45949\ : std_logic;
signal \N__45944\ : std_logic;
signal \N__45941\ : std_logic;
signal \N__45936\ : std_logic;
signal \N__45931\ : std_logic;
signal \N__45926\ : std_logic;
signal \N__45923\ : std_logic;
signal \N__45920\ : std_logic;
signal \N__45917\ : std_logic;
signal \N__45912\ : std_logic;
signal \N__45909\ : std_logic;
signal \N__45906\ : std_logic;
signal \N__45903\ : std_logic;
signal \N__45902\ : std_logic;
signal \N__45901\ : std_logic;
signal \N__45900\ : std_logic;
signal \N__45899\ : std_logic;
signal \N__45898\ : std_logic;
signal \N__45893\ : std_logic;
signal \N__45886\ : std_logic;
signal \N__45883\ : std_logic;
signal \N__45880\ : std_logic;
signal \N__45867\ : std_logic;
signal \N__45864\ : std_logic;
signal \N__45861\ : std_logic;
signal \N__45856\ : std_logic;
signal \N__45853\ : std_logic;
signal \N__45848\ : std_logic;
signal \N__45845\ : std_logic;
signal \N__45842\ : std_logic;
signal \N__45839\ : std_logic;
signal \N__45836\ : std_logic;
signal \N__45819\ : std_logic;
signal \N__45816\ : std_logic;
signal \N__45813\ : std_logic;
signal \N__45812\ : std_logic;
signal \N__45811\ : std_logic;
signal \N__45808\ : std_logic;
signal \N__45803\ : std_logic;
signal \N__45798\ : std_logic;
signal \N__45795\ : std_logic;
signal \N__45792\ : std_logic;
signal \N__45789\ : std_logic;
signal \N__45788\ : std_logic;
signal \N__45787\ : std_logic;
signal \N__45784\ : std_logic;
signal \N__45781\ : std_logic;
signal \N__45778\ : std_logic;
signal \N__45773\ : std_logic;
signal \N__45768\ : std_logic;
signal \N__45765\ : std_logic;
signal \N__45762\ : std_logic;
signal \N__45759\ : std_logic;
signal \N__45756\ : std_logic;
signal \N__45753\ : std_logic;
signal \N__45752\ : std_logic;
signal \N__45751\ : std_logic;
signal \N__45748\ : std_logic;
signal \N__45745\ : std_logic;
signal \N__45742\ : std_logic;
signal \N__45735\ : std_logic;
signal \N__45732\ : std_logic;
signal \N__45729\ : std_logic;
signal \N__45726\ : std_logic;
signal \N__45723\ : std_logic;
signal \N__45720\ : std_logic;
signal \N__45717\ : std_logic;
signal \N__45714\ : std_logic;
signal \N__45711\ : std_logic;
signal \N__45708\ : std_logic;
signal \N__45707\ : std_logic;
signal \N__45704\ : std_logic;
signal \N__45701\ : std_logic;
signal \N__45696\ : std_logic;
signal \N__45695\ : std_logic;
signal \N__45692\ : std_logic;
signal \N__45689\ : std_logic;
signal \N__45686\ : std_logic;
signal \N__45683\ : std_logic;
signal \N__45682\ : std_logic;
signal \N__45681\ : std_logic;
signal \N__45678\ : std_logic;
signal \N__45675\ : std_logic;
signal \N__45672\ : std_logic;
signal \N__45671\ : std_logic;
signal \N__45670\ : std_logic;
signal \N__45669\ : std_logic;
signal \N__45668\ : std_logic;
signal \N__45665\ : std_logic;
signal \N__45664\ : std_logic;
signal \N__45661\ : std_logic;
signal \N__45658\ : std_logic;
signal \N__45655\ : std_logic;
signal \N__45654\ : std_logic;
signal \N__45653\ : std_logic;
signal \N__45652\ : std_logic;
signal \N__45651\ : std_logic;
signal \N__45650\ : std_logic;
signal \N__45649\ : std_logic;
signal \N__45646\ : std_logic;
signal \N__45645\ : std_logic;
signal \N__45644\ : std_logic;
signal \N__45643\ : std_logic;
signal \N__45642\ : std_logic;
signal \N__45641\ : std_logic;
signal \N__45638\ : std_logic;
signal \N__45635\ : std_logic;
signal \N__45634\ : std_logic;
signal \N__45631\ : std_logic;
signal \N__45628\ : std_logic;
signal \N__45627\ : std_logic;
signal \N__45624\ : std_logic;
signal \N__45619\ : std_logic;
signal \N__45616\ : std_logic;
signal \N__45615\ : std_logic;
signal \N__45612\ : std_logic;
signal \N__45611\ : std_logic;
signal \N__45608\ : std_logic;
signal \N__45605\ : std_logic;
signal \N__45602\ : std_logic;
signal \N__45599\ : std_logic;
signal \N__45598\ : std_logic;
signal \N__45597\ : std_logic;
signal \N__45596\ : std_logic;
signal \N__45593\ : std_logic;
signal \N__45592\ : std_logic;
signal \N__45589\ : std_logic;
signal \N__45588\ : std_logic;
signal \N__45587\ : std_logic;
signal \N__45584\ : std_logic;
signal \N__45581\ : std_logic;
signal \N__45578\ : std_logic;
signal \N__45575\ : std_logic;
signal \N__45574\ : std_logic;
signal \N__45571\ : std_logic;
signal \N__45570\ : std_logic;
signal \N__45569\ : std_logic;
signal \N__45568\ : std_logic;
signal \N__45567\ : std_logic;
signal \N__45564\ : std_logic;
signal \N__45561\ : std_logic;
signal \N__45560\ : std_logic;
signal \N__45557\ : std_logic;
signal \N__45556\ : std_logic;
signal \N__45553\ : std_logic;
signal \N__45550\ : std_logic;
signal \N__45547\ : std_logic;
signal \N__45544\ : std_logic;
signal \N__45539\ : std_logic;
signal \N__45538\ : std_logic;
signal \N__45535\ : std_logic;
signal \N__45534\ : std_logic;
signal \N__45531\ : std_logic;
signal \N__45526\ : std_logic;
signal \N__45523\ : std_logic;
signal \N__45520\ : std_logic;
signal \N__45515\ : std_logic;
signal \N__45512\ : std_logic;
signal \N__45509\ : std_logic;
signal \N__45508\ : std_logic;
signal \N__45507\ : std_logic;
signal \N__45502\ : std_logic;
signal \N__45499\ : std_logic;
signal \N__45498\ : std_logic;
signal \N__45497\ : std_logic;
signal \N__45494\ : std_logic;
signal \N__45493\ : std_logic;
signal \N__45492\ : std_logic;
signal \N__45489\ : std_logic;
signal \N__45488\ : std_logic;
signal \N__45487\ : std_logic;
signal \N__45482\ : std_logic;
signal \N__45481\ : std_logic;
signal \N__45478\ : std_logic;
signal \N__45475\ : std_logic;
signal \N__45472\ : std_logic;
signal \N__45467\ : std_logic;
signal \N__45466\ : std_logic;
signal \N__45463\ : std_logic;
signal \N__45462\ : std_logic;
signal \N__45461\ : std_logic;
signal \N__45458\ : std_logic;
signal \N__45455\ : std_logic;
signal \N__45454\ : std_logic;
signal \N__45453\ : std_logic;
signal \N__45452\ : std_logic;
signal \N__45449\ : std_logic;
signal \N__45446\ : std_logic;
signal \N__45443\ : std_logic;
signal \N__45438\ : std_logic;
signal \N__45431\ : std_logic;
signal \N__45426\ : std_logic;
signal \N__45419\ : std_logic;
signal \N__45408\ : std_logic;
signal \N__45403\ : std_logic;
signal \N__45398\ : std_logic;
signal \N__45393\ : std_logic;
signal \N__45388\ : std_logic;
signal \N__45383\ : std_logic;
signal \N__45380\ : std_logic;
signal \N__45377\ : std_logic;
signal \N__45372\ : std_logic;
signal \N__45369\ : std_logic;
signal \N__45366\ : std_logic;
signal \N__45361\ : std_logic;
signal \N__45356\ : std_logic;
signal \N__45351\ : std_logic;
signal \N__45348\ : std_logic;
signal \N__45345\ : std_logic;
signal \N__45338\ : std_logic;
signal \N__45333\ : std_logic;
signal \N__45316\ : std_logic;
signal \N__45305\ : std_logic;
signal \N__45302\ : std_logic;
signal \N__45295\ : std_logic;
signal \N__45270\ : std_logic;
signal \N__45269\ : std_logic;
signal \N__45268\ : std_logic;
signal \N__45267\ : std_logic;
signal \N__45264\ : std_logic;
signal \N__45263\ : std_logic;
signal \N__45262\ : std_logic;
signal \N__45261\ : std_logic;
signal \N__45258\ : std_logic;
signal \N__45255\ : std_logic;
signal \N__45254\ : std_logic;
signal \N__45253\ : std_logic;
signal \N__45252\ : std_logic;
signal \N__45251\ : std_logic;
signal \N__45250\ : std_logic;
signal \N__45247\ : std_logic;
signal \N__45240\ : std_logic;
signal \N__45237\ : std_logic;
signal \N__45234\ : std_logic;
signal \N__45231\ : std_logic;
signal \N__45226\ : std_logic;
signal \N__45219\ : std_logic;
signal \N__45210\ : std_logic;
signal \N__45201\ : std_logic;
signal \N__45198\ : std_logic;
signal \N__45195\ : std_logic;
signal \N__45192\ : std_logic;
signal \N__45189\ : std_logic;
signal \N__45186\ : std_logic;
signal \N__45183\ : std_logic;
signal \N__45180\ : std_logic;
signal \N__45177\ : std_logic;
signal \N__45174\ : std_logic;
signal \N__45171\ : std_logic;
signal \N__45168\ : std_logic;
signal \N__45165\ : std_logic;
signal \N__45162\ : std_logic;
signal \N__45159\ : std_logic;
signal \N__45156\ : std_logic;
signal \N__45153\ : std_logic;
signal \N__45150\ : std_logic;
signal \N__45147\ : std_logic;
signal \N__45144\ : std_logic;
signal \N__45141\ : std_logic;
signal \N__45138\ : std_logic;
signal \N__45135\ : std_logic;
signal \N__45132\ : std_logic;
signal \N__45129\ : std_logic;
signal \N__45126\ : std_logic;
signal \N__45123\ : std_logic;
signal \N__45120\ : std_logic;
signal \N__45117\ : std_logic;
signal \N__45114\ : std_logic;
signal \N__45111\ : std_logic;
signal \N__45108\ : std_logic;
signal \N__45107\ : std_logic;
signal \N__45106\ : std_logic;
signal \N__45105\ : std_logic;
signal \N__45102\ : std_logic;
signal \N__45101\ : std_logic;
signal \N__45100\ : std_logic;
signal \N__45099\ : std_logic;
signal \N__45098\ : std_logic;
signal \N__45095\ : std_logic;
signal \N__45092\ : std_logic;
signal \N__45091\ : std_logic;
signal \N__45090\ : std_logic;
signal \N__45089\ : std_logic;
signal \N__45086\ : std_logic;
signal \N__45083\ : std_logic;
signal \N__45080\ : std_logic;
signal \N__45077\ : std_logic;
signal \N__45072\ : std_logic;
signal \N__45069\ : std_logic;
signal \N__45066\ : std_logic;
signal \N__45063\ : std_logic;
signal \N__45062\ : std_logic;
signal \N__45059\ : std_logic;
signal \N__45056\ : std_logic;
signal \N__45053\ : std_logic;
signal \N__45046\ : std_logic;
signal \N__45037\ : std_logic;
signal \N__45034\ : std_logic;
signal \N__45021\ : std_logic;
signal \N__45020\ : std_logic;
signal \N__45019\ : std_logic;
signal \N__45014\ : std_logic;
signal \N__45011\ : std_logic;
signal \N__45010\ : std_logic;
signal \N__45007\ : std_logic;
signal \N__45006\ : std_logic;
signal \N__45003\ : std_logic;
signal \N__45000\ : std_logic;
signal \N__44997\ : std_logic;
signal \N__44996\ : std_logic;
signal \N__44995\ : std_logic;
signal \N__44992\ : std_logic;
signal \N__44991\ : std_logic;
signal \N__44990\ : std_logic;
signal \N__44985\ : std_logic;
signal \N__44982\ : std_logic;
signal \N__44981\ : std_logic;
signal \N__44978\ : std_logic;
signal \N__44975\ : std_logic;
signal \N__44972\ : std_logic;
signal \N__44969\ : std_logic;
signal \N__44968\ : std_logic;
signal \N__44965\ : std_logic;
signal \N__44964\ : std_logic;
signal \N__44959\ : std_logic;
signal \N__44956\ : std_logic;
signal \N__44953\ : std_logic;
signal \N__44946\ : std_logic;
signal \N__44943\ : std_logic;
signal \N__44940\ : std_logic;
signal \N__44937\ : std_logic;
signal \N__44934\ : std_logic;
signal \N__44929\ : std_logic;
signal \N__44926\ : std_logic;
signal \N__44913\ : std_logic;
signal \N__44912\ : std_logic;
signal \N__44911\ : std_logic;
signal \N__44910\ : std_logic;
signal \N__44909\ : std_logic;
signal \N__44908\ : std_logic;
signal \N__44907\ : std_logic;
signal \N__44904\ : std_logic;
signal \N__44903\ : std_logic;
signal \N__44902\ : std_logic;
signal \N__44899\ : std_logic;
signal \N__44896\ : std_logic;
signal \N__44893\ : std_logic;
signal \N__44892\ : std_logic;
signal \N__44891\ : std_logic;
signal \N__44890\ : std_logic;
signal \N__44887\ : std_logic;
signal \N__44886\ : std_logic;
signal \N__44883\ : std_logic;
signal \N__44880\ : std_logic;
signal \N__44879\ : std_logic;
signal \N__44878\ : std_logic;
signal \N__44875\ : std_logic;
signal \N__44874\ : std_logic;
signal \N__44873\ : std_logic;
signal \N__44872\ : std_logic;
signal \N__44871\ : std_logic;
signal \N__44868\ : std_logic;
signal \N__44863\ : std_logic;
signal \N__44860\ : std_logic;
signal \N__44855\ : std_logic;
signal \N__44854\ : std_logic;
signal \N__44853\ : std_logic;
signal \N__44848\ : std_logic;
signal \N__44845\ : std_logic;
signal \N__44842\ : std_logic;
signal \N__44837\ : std_logic;
signal \N__44832\ : std_logic;
signal \N__44831\ : std_logic;
signal \N__44830\ : std_logic;
signal \N__44827\ : std_logic;
signal \N__44824\ : std_logic;
signal \N__44819\ : std_logic;
signal \N__44816\ : std_logic;
signal \N__44807\ : std_logic;
signal \N__44802\ : std_logic;
signal \N__44799\ : std_logic;
signal \N__44790\ : std_logic;
signal \N__44787\ : std_logic;
signal \N__44784\ : std_logic;
signal \N__44777\ : std_logic;
signal \N__44770\ : std_logic;
signal \N__44765\ : std_logic;
signal \N__44754\ : std_logic;
signal \N__44751\ : std_logic;
signal \N__44748\ : std_logic;
signal \N__44745\ : std_logic;
signal \N__44742\ : std_logic;
signal \N__44739\ : std_logic;
signal \N__44738\ : std_logic;
signal \N__44737\ : std_logic;
signal \N__44734\ : std_logic;
signal \N__44729\ : std_logic;
signal \N__44724\ : std_logic;
signal \N__44721\ : std_logic;
signal \N__44718\ : std_logic;
signal \N__44715\ : std_logic;
signal \N__44712\ : std_logic;
signal \N__44709\ : std_logic;
signal \N__44708\ : std_logic;
signal \N__44705\ : std_logic;
signal \N__44702\ : std_logic;
signal \N__44699\ : std_logic;
signal \N__44698\ : std_logic;
signal \N__44695\ : std_logic;
signal \N__44692\ : std_logic;
signal \N__44689\ : std_logic;
signal \N__44686\ : std_logic;
signal \N__44679\ : std_logic;
signal \N__44676\ : std_logic;
signal \N__44673\ : std_logic;
signal \N__44670\ : std_logic;
signal \N__44667\ : std_logic;
signal \N__44664\ : std_logic;
signal \N__44661\ : std_logic;
signal \N__44658\ : std_logic;
signal \N__44655\ : std_logic;
signal \N__44652\ : std_logic;
signal \N__44649\ : std_logic;
signal \N__44646\ : std_logic;
signal \N__44643\ : std_logic;
signal \N__44642\ : std_logic;
signal \N__44639\ : std_logic;
signal \N__44636\ : std_logic;
signal \N__44635\ : std_logic;
signal \N__44632\ : std_logic;
signal \N__44629\ : std_logic;
signal \N__44626\ : std_logic;
signal \N__44619\ : std_logic;
signal \N__44616\ : std_logic;
signal \N__44615\ : std_logic;
signal \N__44612\ : std_logic;
signal \N__44609\ : std_logic;
signal \N__44608\ : std_logic;
signal \N__44605\ : std_logic;
signal \N__44600\ : std_logic;
signal \N__44595\ : std_logic;
signal \N__44592\ : std_logic;
signal \N__44589\ : std_logic;
signal \N__44586\ : std_logic;
signal \N__44585\ : std_logic;
signal \N__44582\ : std_logic;
signal \N__44581\ : std_logic;
signal \N__44578\ : std_logic;
signal \N__44575\ : std_logic;
signal \N__44572\ : std_logic;
signal \N__44569\ : std_logic;
signal \N__44562\ : std_logic;
signal \N__44559\ : std_logic;
signal \N__44556\ : std_logic;
signal \N__44553\ : std_logic;
signal \N__44550\ : std_logic;
signal \N__44547\ : std_logic;
signal \N__44544\ : std_logic;
signal \N__44541\ : std_logic;
signal \N__44540\ : std_logic;
signal \N__44539\ : std_logic;
signal \N__44538\ : std_logic;
signal \N__44537\ : std_logic;
signal \N__44536\ : std_logic;
signal \N__44535\ : std_logic;
signal \N__44534\ : std_logic;
signal \N__44533\ : std_logic;
signal \N__44532\ : std_logic;
signal \N__44531\ : std_logic;
signal \N__44530\ : std_logic;
signal \N__44529\ : std_logic;
signal \N__44526\ : std_logic;
signal \N__44523\ : std_logic;
signal \N__44520\ : std_logic;
signal \N__44517\ : std_logic;
signal \N__44514\ : std_logic;
signal \N__44509\ : std_logic;
signal \N__44504\ : std_logic;
signal \N__44503\ : std_logic;
signal \N__44500\ : std_logic;
signal \N__44497\ : std_logic;
signal \N__44494\ : std_logic;
signal \N__44491\ : std_logic;
signal \N__44488\ : std_logic;
signal \N__44485\ : std_logic;
signal \N__44474\ : std_logic;
signal \N__44471\ : std_logic;
signal \N__44468\ : std_logic;
signal \N__44463\ : std_logic;
signal \N__44460\ : std_logic;
signal \N__44453\ : std_logic;
signal \N__44442\ : std_logic;
signal \N__44439\ : std_logic;
signal \N__44436\ : std_logic;
signal \N__44435\ : std_logic;
signal \N__44432\ : std_logic;
signal \N__44431\ : std_logic;
signal \N__44430\ : std_logic;
signal \N__44427\ : std_logic;
signal \N__44426\ : std_logic;
signal \N__44423\ : std_logic;
signal \N__44422\ : std_logic;
signal \N__44421\ : std_logic;
signal \N__44418\ : std_logic;
signal \N__44415\ : std_logic;
signal \N__44412\ : std_logic;
signal \N__44409\ : std_logic;
signal \N__44406\ : std_logic;
signal \N__44405\ : std_logic;
signal \N__44402\ : std_logic;
signal \N__44399\ : std_logic;
signal \N__44396\ : std_logic;
signal \N__44393\ : std_logic;
signal \N__44390\ : std_logic;
signal \N__44389\ : std_logic;
signal \N__44388\ : std_logic;
signal \N__44387\ : std_logic;
signal \N__44384\ : std_logic;
signal \N__44381\ : std_logic;
signal \N__44378\ : std_logic;
signal \N__44375\ : std_logic;
signal \N__44372\ : std_logic;
signal \N__44367\ : std_logic;
signal \N__44364\ : std_logic;
signal \N__44361\ : std_logic;
signal \N__44358\ : std_logic;
signal \N__44355\ : std_logic;
signal \N__44350\ : std_logic;
signal \N__44339\ : std_logic;
signal \N__44328\ : std_logic;
signal \N__44325\ : std_logic;
signal \N__44322\ : std_logic;
signal \N__44319\ : std_logic;
signal \N__44316\ : std_logic;
signal \N__44313\ : std_logic;
signal \N__44310\ : std_logic;
signal \N__44309\ : std_logic;
signal \N__44308\ : std_logic;
signal \N__44305\ : std_logic;
signal \N__44302\ : std_logic;
signal \N__44299\ : std_logic;
signal \N__44292\ : std_logic;
signal \N__44289\ : std_logic;
signal \N__44286\ : std_logic;
signal \N__44283\ : std_logic;
signal \N__44282\ : std_logic;
signal \N__44279\ : std_logic;
signal \N__44278\ : std_logic;
signal \N__44275\ : std_logic;
signal \N__44272\ : std_logic;
signal \N__44269\ : std_logic;
signal \N__44266\ : std_logic;
signal \N__44263\ : std_logic;
signal \N__44260\ : std_logic;
signal \N__44257\ : std_logic;
signal \N__44250\ : std_logic;
signal \N__44247\ : std_logic;
signal \N__44244\ : std_logic;
signal \N__44241\ : std_logic;
signal \N__44238\ : std_logic;
signal \N__44235\ : std_logic;
signal \N__44232\ : std_logic;
signal \N__44231\ : std_logic;
signal \N__44228\ : std_logic;
signal \N__44225\ : std_logic;
signal \N__44220\ : std_logic;
signal \N__44219\ : std_logic;
signal \N__44216\ : std_logic;
signal \N__44213\ : std_logic;
signal \N__44210\ : std_logic;
signal \N__44207\ : std_logic;
signal \N__44204\ : std_logic;
signal \N__44199\ : std_logic;
signal \N__44196\ : std_logic;
signal \N__44193\ : std_logic;
signal \N__44190\ : std_logic;
signal \N__44187\ : std_logic;
signal \N__44184\ : std_logic;
signal \N__44181\ : std_logic;
signal \N__44178\ : std_logic;
signal \N__44175\ : std_logic;
signal \N__44172\ : std_logic;
signal \N__44169\ : std_logic;
signal \N__44168\ : std_logic;
signal \N__44165\ : std_logic;
signal \N__44162\ : std_logic;
signal \N__44157\ : std_logic;
signal \N__44154\ : std_logic;
signal \N__44151\ : std_logic;
signal \N__44148\ : std_logic;
signal \N__44145\ : std_logic;
signal \N__44142\ : std_logic;
signal \N__44139\ : std_logic;
signal \N__44136\ : std_logic;
signal \N__44133\ : std_logic;
signal \N__44130\ : std_logic;
signal \N__44127\ : std_logic;
signal \N__44124\ : std_logic;
signal \N__44121\ : std_logic;
signal \N__44118\ : std_logic;
signal \N__44115\ : std_logic;
signal \N__44114\ : std_logic;
signal \N__44113\ : std_logic;
signal \N__44112\ : std_logic;
signal \N__44111\ : std_logic;
signal \N__44108\ : std_logic;
signal \N__44107\ : std_logic;
signal \N__44106\ : std_logic;
signal \N__44105\ : std_logic;
signal \N__44102\ : std_logic;
signal \N__44099\ : std_logic;
signal \N__44096\ : std_logic;
signal \N__44095\ : std_logic;
signal \N__44092\ : std_logic;
signal \N__44091\ : std_logic;
signal \N__44088\ : std_logic;
signal \N__44085\ : std_logic;
signal \N__44082\ : std_logic;
signal \N__44079\ : std_logic;
signal \N__44076\ : std_logic;
signal \N__44073\ : std_logic;
signal \N__44070\ : std_logic;
signal \N__44067\ : std_logic;
signal \N__44064\ : std_logic;
signal \N__44063\ : std_logic;
signal \N__44060\ : std_logic;
signal \N__44055\ : std_logic;
signal \N__44052\ : std_logic;
signal \N__44047\ : std_logic;
signal \N__44044\ : std_logic;
signal \N__44041\ : std_logic;
signal \N__44036\ : std_logic;
signal \N__44033\ : std_logic;
signal \N__44028\ : std_logic;
signal \N__44021\ : std_logic;
signal \N__44016\ : std_logic;
signal \N__44007\ : std_logic;
signal \N__44004\ : std_logic;
signal \N__44001\ : std_logic;
signal \N__43998\ : std_logic;
signal \N__43995\ : std_logic;
signal \N__43992\ : std_logic;
signal \N__43989\ : std_logic;
signal \N__43988\ : std_logic;
signal \N__43985\ : std_logic;
signal \N__43982\ : std_logic;
signal \N__43977\ : std_logic;
signal \N__43976\ : std_logic;
signal \N__43971\ : std_logic;
signal \N__43968\ : std_logic;
signal \N__43965\ : std_logic;
signal \N__43962\ : std_logic;
signal \N__43959\ : std_logic;
signal \N__43956\ : std_logic;
signal \N__43955\ : std_logic;
signal \N__43952\ : std_logic;
signal \N__43951\ : std_logic;
signal \N__43948\ : std_logic;
signal \N__43947\ : std_logic;
signal \N__43944\ : std_logic;
signal \N__43941\ : std_logic;
signal \N__43940\ : std_logic;
signal \N__43939\ : std_logic;
signal \N__43936\ : std_logic;
signal \N__43933\ : std_logic;
signal \N__43932\ : std_logic;
signal \N__43929\ : std_logic;
signal \N__43926\ : std_logic;
signal \N__43925\ : std_logic;
signal \N__43922\ : std_logic;
signal \N__43919\ : std_logic;
signal \N__43916\ : std_logic;
signal \N__43913\ : std_logic;
signal \N__43912\ : std_logic;
signal \N__43911\ : std_logic;
signal \N__43910\ : std_logic;
signal \N__43907\ : std_logic;
signal \N__43902\ : std_logic;
signal \N__43899\ : std_logic;
signal \N__43898\ : std_logic;
signal \N__43897\ : std_logic;
signal \N__43896\ : std_logic;
signal \N__43895\ : std_logic;
signal \N__43894\ : std_logic;
signal \N__43893\ : std_logic;
signal \N__43892\ : std_logic;
signal \N__43891\ : std_logic;
signal \N__43890\ : std_logic;
signal \N__43887\ : std_logic;
signal \N__43884\ : std_logic;
signal \N__43879\ : std_logic;
signal \N__43876\ : std_logic;
signal \N__43875\ : std_logic;
signal \N__43874\ : std_logic;
signal \N__43869\ : std_logic;
signal \N__43866\ : std_logic;
signal \N__43861\ : std_logic;
signal \N__43858\ : std_logic;
signal \N__43853\ : std_logic;
signal \N__43846\ : std_logic;
signal \N__43843\ : std_logic;
signal \N__43840\ : std_logic;
signal \N__43837\ : std_logic;
signal \N__43836\ : std_logic;
signal \N__43833\ : std_logic;
signal \N__43828\ : std_logic;
signal \N__43825\ : std_logic;
signal \N__43824\ : std_logic;
signal \N__43823\ : std_logic;
signal \N__43822\ : std_logic;
signal \N__43819\ : std_logic;
signal \N__43818\ : std_logic;
signal \N__43817\ : std_logic;
signal \N__43814\ : std_logic;
signal \N__43811\ : std_logic;
signal \N__43806\ : std_logic;
signal \N__43797\ : std_logic;
signal \N__43794\ : std_logic;
signal \N__43791\ : std_logic;
signal \N__43788\ : std_logic;
signal \N__43783\ : std_logic;
signal \N__43780\ : std_logic;
signal \N__43777\ : std_logic;
signal \N__43774\ : std_logic;
signal \N__43771\ : std_logic;
signal \N__43768\ : std_logic;
signal \N__43765\ : std_logic;
signal \N__43762\ : std_logic;
signal \N__43755\ : std_logic;
signal \N__43752\ : std_logic;
signal \N__43745\ : std_logic;
signal \N__43740\ : std_logic;
signal \N__43737\ : std_logic;
signal \N__43716\ : std_logic;
signal \N__43715\ : std_logic;
signal \N__43712\ : std_logic;
signal \N__43711\ : std_logic;
signal \N__43708\ : std_logic;
signal \N__43705\ : std_logic;
signal \N__43702\ : std_logic;
signal \N__43701\ : std_logic;
signal \N__43698\ : std_logic;
signal \N__43693\ : std_logic;
signal \N__43692\ : std_logic;
signal \N__43691\ : std_logic;
signal \N__43688\ : std_logic;
signal \N__43685\ : std_logic;
signal \N__43682\ : std_logic;
signal \N__43681\ : std_logic;
signal \N__43680\ : std_logic;
signal \N__43677\ : std_logic;
signal \N__43676\ : std_logic;
signal \N__43675\ : std_logic;
signal \N__43672\ : std_logic;
signal \N__43669\ : std_logic;
signal \N__43668\ : std_logic;
signal \N__43663\ : std_logic;
signal \N__43660\ : std_logic;
signal \N__43653\ : std_logic;
signal \N__43652\ : std_logic;
signal \N__43651\ : std_logic;
signal \N__43648\ : std_logic;
signal \N__43645\ : std_logic;
signal \N__43642\ : std_logic;
signal \N__43641\ : std_logic;
signal \N__43640\ : std_logic;
signal \N__43637\ : std_logic;
signal \N__43632\ : std_logic;
signal \N__43629\ : std_logic;
signal \N__43626\ : std_logic;
signal \N__43625\ : std_logic;
signal \N__43622\ : std_logic;
signal \N__43619\ : std_logic;
signal \N__43614\ : std_logic;
signal \N__43611\ : std_logic;
signal \N__43606\ : std_logic;
signal \N__43601\ : std_logic;
signal \N__43600\ : std_logic;
signal \N__43597\ : std_logic;
signal \N__43596\ : std_logic;
signal \N__43593\ : std_logic;
signal \N__43592\ : std_logic;
signal \N__43589\ : std_logic;
signal \N__43588\ : std_logic;
signal \N__43585\ : std_logic;
signal \N__43584\ : std_logic;
signal \N__43581\ : std_logic;
signal \N__43576\ : std_logic;
signal \N__43573\ : std_logic;
signal \N__43570\ : std_logic;
signal \N__43567\ : std_logic;
signal \N__43564\ : std_logic;
signal \N__43561\ : std_logic;
signal \N__43558\ : std_logic;
signal \N__43555\ : std_logic;
signal \N__43552\ : std_logic;
signal \N__43549\ : std_logic;
signal \N__43546\ : std_logic;
signal \N__43541\ : std_logic;
signal \N__43536\ : std_logic;
signal \N__43533\ : std_logic;
signal \N__43528\ : std_logic;
signal \N__43521\ : std_logic;
signal \N__43506\ : std_logic;
signal \N__43505\ : std_logic;
signal \N__43502\ : std_logic;
signal \N__43499\ : std_logic;
signal \N__43496\ : std_logic;
signal \N__43493\ : std_logic;
signal \N__43492\ : std_logic;
signal \N__43491\ : std_logic;
signal \N__43486\ : std_logic;
signal \N__43483\ : std_logic;
signal \N__43480\ : std_logic;
signal \N__43473\ : std_logic;
signal \N__43470\ : std_logic;
signal \N__43467\ : std_logic;
signal \N__43464\ : std_logic;
signal \N__43461\ : std_logic;
signal \N__43458\ : std_logic;
signal \N__43455\ : std_logic;
signal \N__43452\ : std_logic;
signal \N__43449\ : std_logic;
signal \N__43446\ : std_logic;
signal \N__43443\ : std_logic;
signal \N__43442\ : std_logic;
signal \N__43439\ : std_logic;
signal \N__43436\ : std_logic;
signal \N__43431\ : std_logic;
signal \N__43430\ : std_logic;
signal \N__43429\ : std_logic;
signal \N__43428\ : std_logic;
signal \N__43425\ : std_logic;
signal \N__43424\ : std_logic;
signal \N__43421\ : std_logic;
signal \N__43418\ : std_logic;
signal \N__43415\ : std_logic;
signal \N__43414\ : std_logic;
signal \N__43411\ : std_logic;
signal \N__43408\ : std_logic;
signal \N__43405\ : std_logic;
signal \N__43402\ : std_logic;
signal \N__43399\ : std_logic;
signal \N__43398\ : std_logic;
signal \N__43395\ : std_logic;
signal \N__43392\ : std_logic;
signal \N__43389\ : std_logic;
signal \N__43386\ : std_logic;
signal \N__43381\ : std_logic;
signal \N__43378\ : std_logic;
signal \N__43365\ : std_logic;
signal \N__43362\ : std_logic;
signal \N__43359\ : std_logic;
signal \N__43356\ : std_logic;
signal \N__43353\ : std_logic;
signal \N__43350\ : std_logic;
signal \N__43347\ : std_logic;
signal \N__43344\ : std_logic;
signal \N__43341\ : std_logic;
signal \N__43340\ : std_logic;
signal \N__43337\ : std_logic;
signal \N__43336\ : std_logic;
signal \N__43333\ : std_logic;
signal \N__43330\ : std_logic;
signal \N__43327\ : std_logic;
signal \N__43324\ : std_logic;
signal \N__43321\ : std_logic;
signal \N__43318\ : std_logic;
signal \N__43315\ : std_logic;
signal \N__43308\ : std_logic;
signal \N__43305\ : std_logic;
signal \N__43302\ : std_logic;
signal \N__43299\ : std_logic;
signal \N__43296\ : std_logic;
signal \N__43293\ : std_logic;
signal \N__43290\ : std_logic;
signal \N__43287\ : std_logic;
signal \N__43284\ : std_logic;
signal \N__43281\ : std_logic;
signal \N__43278\ : std_logic;
signal \N__43275\ : std_logic;
signal \N__43272\ : std_logic;
signal \N__43269\ : std_logic;
signal \N__43266\ : std_logic;
signal \N__43263\ : std_logic;
signal \N__43260\ : std_logic;
signal \N__43257\ : std_logic;
signal \N__43254\ : std_logic;
signal \N__43251\ : std_logic;
signal \N__43248\ : std_logic;
signal \N__43245\ : std_logic;
signal \N__43244\ : std_logic;
signal \N__43243\ : std_logic;
signal \N__43242\ : std_logic;
signal \N__43241\ : std_logic;
signal \N__43240\ : std_logic;
signal \N__43239\ : std_logic;
signal \N__43238\ : std_logic;
signal \N__43237\ : std_logic;
signal \N__43236\ : std_logic;
signal \N__43233\ : std_logic;
signal \N__43230\ : std_logic;
signal \N__43225\ : std_logic;
signal \N__43218\ : std_logic;
signal \N__43211\ : std_logic;
signal \N__43200\ : std_logic;
signal \N__43197\ : std_logic;
signal \N__43194\ : std_logic;
signal \N__43191\ : std_logic;
signal \N__43190\ : std_logic;
signal \N__43187\ : std_logic;
signal \N__43186\ : std_logic;
signal \N__43185\ : std_logic;
signal \N__43184\ : std_logic;
signal \N__43183\ : std_logic;
signal \N__43180\ : std_logic;
signal \N__43175\ : std_logic;
signal \N__43174\ : std_logic;
signal \N__43171\ : std_logic;
signal \N__43168\ : std_logic;
signal \N__43165\ : std_logic;
signal \N__43160\ : std_logic;
signal \N__43157\ : std_logic;
signal \N__43154\ : std_logic;
signal \N__43151\ : std_logic;
signal \N__43148\ : std_logic;
signal \N__43143\ : std_logic;
signal \N__43140\ : std_logic;
signal \N__43137\ : std_logic;
signal \N__43128\ : std_logic;
signal \N__43125\ : std_logic;
signal \N__43122\ : std_logic;
signal \N__43119\ : std_logic;
signal \N__43116\ : std_logic;
signal \N__43115\ : std_logic;
signal \N__43112\ : std_logic;
signal \N__43109\ : std_logic;
signal \N__43104\ : std_logic;
signal \N__43103\ : std_logic;
signal \N__43100\ : std_logic;
signal \N__43097\ : std_logic;
signal \N__43092\ : std_logic;
signal \N__43091\ : std_logic;
signal \N__43088\ : std_logic;
signal \N__43085\ : std_logic;
signal \N__43082\ : std_logic;
signal \N__43079\ : std_logic;
signal \N__43074\ : std_logic;
signal \N__43073\ : std_logic;
signal \N__43070\ : std_logic;
signal \N__43067\ : std_logic;
signal \N__43062\ : std_logic;
signal \N__43059\ : std_logic;
signal \N__43056\ : std_logic;
signal \N__43053\ : std_logic;
signal \N__43050\ : std_logic;
signal \N__43047\ : std_logic;
signal \N__43044\ : std_logic;
signal \N__43043\ : std_logic;
signal \N__43042\ : std_logic;
signal \N__43039\ : std_logic;
signal \N__43034\ : std_logic;
signal \N__43029\ : std_logic;
signal \N__43026\ : std_logic;
signal \N__43023\ : std_logic;
signal \N__43020\ : std_logic;
signal \N__43017\ : std_logic;
signal \N__43014\ : std_logic;
signal \N__43011\ : std_logic;
signal \N__43010\ : std_logic;
signal \N__43009\ : std_logic;
signal \N__43006\ : std_logic;
signal \N__43001\ : std_logic;
signal \N__42996\ : std_logic;
signal \N__42993\ : std_logic;
signal \N__42990\ : std_logic;
signal \N__42987\ : std_logic;
signal \N__42984\ : std_logic;
signal \N__42981\ : std_logic;
signal \N__42978\ : std_logic;
signal \N__42977\ : std_logic;
signal \N__42974\ : std_logic;
signal \N__42971\ : std_logic;
signal \N__42966\ : std_logic;
signal \N__42963\ : std_logic;
signal \N__42960\ : std_logic;
signal \N__42957\ : std_logic;
signal \N__42954\ : std_logic;
signal \N__42951\ : std_logic;
signal \N__42950\ : std_logic;
signal \N__42947\ : std_logic;
signal \N__42946\ : std_logic;
signal \N__42943\ : std_logic;
signal \N__42940\ : std_logic;
signal \N__42937\ : std_logic;
signal \N__42934\ : std_logic;
signal \N__42927\ : std_logic;
signal \N__42924\ : std_logic;
signal \N__42921\ : std_logic;
signal \N__42918\ : std_logic;
signal \N__42915\ : std_logic;
signal \N__42912\ : std_logic;
signal \N__42909\ : std_logic;
signal \N__42908\ : std_logic;
signal \N__42907\ : std_logic;
signal \N__42904\ : std_logic;
signal \N__42899\ : std_logic;
signal \N__42894\ : std_logic;
signal \N__42891\ : std_logic;
signal \N__42888\ : std_logic;
signal \N__42887\ : std_logic;
signal \N__42884\ : std_logic;
signal \N__42881\ : std_logic;
signal \N__42880\ : std_logic;
signal \N__42879\ : std_logic;
signal \N__42878\ : std_logic;
signal \N__42877\ : std_logic;
signal \N__42876\ : std_logic;
signal \N__42875\ : std_logic;
signal \N__42874\ : std_logic;
signal \N__42869\ : std_logic;
signal \N__42862\ : std_logic;
signal \N__42853\ : std_logic;
signal \N__42850\ : std_logic;
signal \N__42843\ : std_logic;
signal \N__42840\ : std_logic;
signal \N__42837\ : std_logic;
signal \N__42834\ : std_logic;
signal \N__42831\ : std_logic;
signal \N__42828\ : std_logic;
signal \N__42825\ : std_logic;
signal \N__42822\ : std_logic;
signal \N__42819\ : std_logic;
signal \N__42818\ : std_logic;
signal \N__42815\ : std_logic;
signal \N__42812\ : std_logic;
signal \N__42807\ : std_logic;
signal \N__42804\ : std_logic;
signal \N__42801\ : std_logic;
signal \N__42798\ : std_logic;
signal \N__42797\ : std_logic;
signal \N__42794\ : std_logic;
signal \N__42791\ : std_logic;
signal \N__42786\ : std_logic;
signal \N__42785\ : std_logic;
signal \N__42782\ : std_logic;
signal \N__42779\ : std_logic;
signal \N__42776\ : std_logic;
signal \N__42771\ : std_logic;
signal \N__42768\ : std_logic;
signal \N__42767\ : std_logic;
signal \N__42764\ : std_logic;
signal \N__42761\ : std_logic;
signal \N__42756\ : std_logic;
signal \N__42755\ : std_logic;
signal \N__42752\ : std_logic;
signal \N__42749\ : std_logic;
signal \N__42744\ : std_logic;
signal \N__42741\ : std_logic;
signal \N__42738\ : std_logic;
signal \N__42735\ : std_logic;
signal \N__42732\ : std_logic;
signal \N__42729\ : std_logic;
signal \N__42728\ : std_logic;
signal \N__42725\ : std_logic;
signal \N__42724\ : std_logic;
signal \N__42721\ : std_logic;
signal \N__42718\ : std_logic;
signal \N__42715\ : std_logic;
signal \N__42712\ : std_logic;
signal \N__42705\ : std_logic;
signal \N__42702\ : std_logic;
signal \N__42699\ : std_logic;
signal \N__42698\ : std_logic;
signal \N__42695\ : std_logic;
signal \N__42694\ : std_logic;
signal \N__42691\ : std_logic;
signal \N__42688\ : std_logic;
signal \N__42685\ : std_logic;
signal \N__42682\ : std_logic;
signal \N__42675\ : std_logic;
signal \N__42672\ : std_logic;
signal \N__42669\ : std_logic;
signal \N__42666\ : std_logic;
signal \N__42663\ : std_logic;
signal \N__42660\ : std_logic;
signal \N__42657\ : std_logic;
signal \N__42654\ : std_logic;
signal \N__42651\ : std_logic;
signal \N__42648\ : std_logic;
signal \N__42645\ : std_logic;
signal \N__42642\ : std_logic;
signal \N__42639\ : std_logic;
signal \N__42636\ : std_logic;
signal \N__42635\ : std_logic;
signal \N__42632\ : std_logic;
signal \N__42629\ : std_logic;
signal \N__42628\ : std_logic;
signal \N__42627\ : std_logic;
signal \N__42622\ : std_logic;
signal \N__42619\ : std_logic;
signal \N__42616\ : std_logic;
signal \N__42615\ : std_logic;
signal \N__42614\ : std_logic;
signal \N__42613\ : std_logic;
signal \N__42610\ : std_logic;
signal \N__42605\ : std_logic;
signal \N__42604\ : std_logic;
signal \N__42603\ : std_logic;
signal \N__42600\ : std_logic;
signal \N__42595\ : std_logic;
signal \N__42592\ : std_logic;
signal \N__42589\ : std_logic;
signal \N__42588\ : std_logic;
signal \N__42587\ : std_logic;
signal \N__42584\ : std_logic;
signal \N__42583\ : std_logic;
signal \N__42582\ : std_logic;
signal \N__42579\ : std_logic;
signal \N__42578\ : std_logic;
signal \N__42575\ : std_logic;
signal \N__42572\ : std_logic;
signal \N__42569\ : std_logic;
signal \N__42566\ : std_logic;
signal \N__42561\ : std_logic;
signal \N__42558\ : std_logic;
signal \N__42553\ : std_logic;
signal \N__42550\ : std_logic;
signal \N__42547\ : std_logic;
signal \N__42542\ : std_logic;
signal \N__42539\ : std_logic;
signal \N__42536\ : std_logic;
signal \N__42519\ : std_logic;
signal \N__42516\ : std_logic;
signal \N__42513\ : std_logic;
signal \N__42510\ : std_logic;
signal \N__42509\ : std_logic;
signal \N__42506\ : std_logic;
signal \N__42503\ : std_logic;
signal \N__42498\ : std_logic;
signal \N__42495\ : std_logic;
signal \N__42494\ : std_logic;
signal \N__42491\ : std_logic;
signal \N__42488\ : std_logic;
signal \N__42483\ : std_logic;
signal \N__42480\ : std_logic;
signal \N__42477\ : std_logic;
signal \N__42476\ : std_logic;
signal \N__42473\ : std_logic;
signal \N__42470\ : std_logic;
signal \N__42465\ : std_logic;
signal \N__42462\ : std_logic;
signal \N__42459\ : std_logic;
signal \N__42456\ : std_logic;
signal \N__42455\ : std_logic;
signal \N__42452\ : std_logic;
signal \N__42449\ : std_logic;
signal \N__42444\ : std_logic;
signal \N__42441\ : std_logic;
signal \N__42438\ : std_logic;
signal \N__42435\ : std_logic;
signal \N__42434\ : std_logic;
signal \N__42433\ : std_logic;
signal \N__42432\ : std_logic;
signal \N__42431\ : std_logic;
signal \N__42428\ : std_logic;
signal \N__42427\ : std_logic;
signal \N__42424\ : std_logic;
signal \N__42423\ : std_logic;
signal \N__42420\ : std_logic;
signal \N__42405\ : std_logic;
signal \N__42402\ : std_logic;
signal \N__42399\ : std_logic;
signal \N__42398\ : std_logic;
signal \N__42395\ : std_logic;
signal \N__42392\ : std_logic;
signal \N__42387\ : std_logic;
signal \N__42384\ : std_logic;
signal \N__42381\ : std_logic;
signal \N__42378\ : std_logic;
signal \N__42375\ : std_logic;
signal \N__42372\ : std_logic;
signal \N__42369\ : std_logic;
signal \N__42366\ : std_logic;
signal \N__42363\ : std_logic;
signal \N__42362\ : std_logic;
signal \N__42359\ : std_logic;
signal \N__42356\ : std_logic;
signal \N__42353\ : std_logic;
signal \N__42350\ : std_logic;
signal \N__42345\ : std_logic;
signal \N__42342\ : std_logic;
signal \N__42339\ : std_logic;
signal \N__42336\ : std_logic;
signal \N__42333\ : std_logic;
signal \N__42332\ : std_logic;
signal \N__42329\ : std_logic;
signal \N__42326\ : std_logic;
signal \N__42323\ : std_logic;
signal \N__42320\ : std_logic;
signal \N__42317\ : std_logic;
signal \N__42312\ : std_logic;
signal \N__42309\ : std_logic;
signal \N__42306\ : std_logic;
signal \N__42303\ : std_logic;
signal \N__42300\ : std_logic;
signal \N__42299\ : std_logic;
signal \N__42298\ : std_logic;
signal \N__42297\ : std_logic;
signal \N__42296\ : std_logic;
signal \N__42295\ : std_logic;
signal \N__42294\ : std_logic;
signal \N__42293\ : std_logic;
signal \N__42290\ : std_logic;
signal \N__42289\ : std_logic;
signal \N__42288\ : std_logic;
signal \N__42287\ : std_logic;
signal \N__42284\ : std_logic;
signal \N__42283\ : std_logic;
signal \N__42282\ : std_logic;
signal \N__42281\ : std_logic;
signal \N__42280\ : std_logic;
signal \N__42279\ : std_logic;
signal \N__42276\ : std_logic;
signal \N__42275\ : std_logic;
signal \N__42274\ : std_logic;
signal \N__42271\ : std_logic;
signal \N__42270\ : std_logic;
signal \N__42269\ : std_logic;
signal \N__42268\ : std_logic;
signal \N__42267\ : std_logic;
signal \N__42264\ : std_logic;
signal \N__42263\ : std_logic;
signal \N__42262\ : std_logic;
signal \N__42259\ : std_logic;
signal \N__42258\ : std_logic;
signal \N__42257\ : std_logic;
signal \N__42256\ : std_logic;
signal \N__42255\ : std_logic;
signal \N__42254\ : std_logic;
signal \N__42253\ : std_logic;
signal \N__42252\ : std_logic;
signal \N__42251\ : std_logic;
signal \N__42244\ : std_logic;
signal \N__42239\ : std_logic;
signal \N__42230\ : std_logic;
signal \N__42229\ : std_logic;
signal \N__42226\ : std_logic;
signal \N__42225\ : std_logic;
signal \N__42224\ : std_logic;
signal \N__42223\ : std_logic;
signal \N__42222\ : std_logic;
signal \N__42221\ : std_logic;
signal \N__42220\ : std_logic;
signal \N__42219\ : std_logic;
signal \N__42218\ : std_logic;
signal \N__42217\ : std_logic;
signal \N__42216\ : std_logic;
signal \N__42215\ : std_logic;
signal \N__42214\ : std_logic;
signal \N__42213\ : std_logic;
signal \N__42212\ : std_logic;
signal \N__42211\ : std_logic;
signal \N__42210\ : std_logic;
signal \N__42209\ : std_logic;
signal \N__42208\ : std_logic;
signal \N__42207\ : std_logic;
signal \N__42206\ : std_logic;
signal \N__42205\ : std_logic;
signal \N__42204\ : std_logic;
signal \N__42203\ : std_logic;
signal \N__42202\ : std_logic;
signal \N__42201\ : std_logic;
signal \N__42200\ : std_logic;
signal \N__42199\ : std_logic;
signal \N__42198\ : std_logic;
signal \N__42197\ : std_logic;
signal \N__42196\ : std_logic;
signal \N__42195\ : std_logic;
signal \N__42194\ : std_logic;
signal \N__42193\ : std_logic;
signal \N__42188\ : std_logic;
signal \N__42187\ : std_logic;
signal \N__42176\ : std_logic;
signal \N__42175\ : std_logic;
signal \N__42174\ : std_logic;
signal \N__42173\ : std_logic;
signal \N__42172\ : std_logic;
signal \N__42171\ : std_logic;
signal \N__42170\ : std_logic;
signal \N__42169\ : std_logic;
signal \N__42168\ : std_logic;
signal \N__42163\ : std_logic;
signal \N__42154\ : std_logic;
signal \N__42145\ : std_logic;
signal \N__42142\ : std_logic;
signal \N__42141\ : std_logic;
signal \N__42140\ : std_logic;
signal \N__42139\ : std_logic;
signal \N__42138\ : std_logic;
signal \N__42129\ : std_logic;
signal \N__42128\ : std_logic;
signal \N__42127\ : std_logic;
signal \N__42126\ : std_logic;
signal \N__42125\ : std_logic;
signal \N__42124\ : std_logic;
signal \N__42123\ : std_logic;
signal \N__42122\ : std_logic;
signal \N__42121\ : std_logic;
signal \N__42120\ : std_logic;
signal \N__42113\ : std_logic;
signal \N__42110\ : std_logic;
signal \N__42105\ : std_logic;
signal \N__42102\ : std_logic;
signal \N__42099\ : std_logic;
signal \N__42098\ : std_logic;
signal \N__42097\ : std_logic;
signal \N__42096\ : std_logic;
signal \N__42095\ : std_logic;
signal \N__42094\ : std_logic;
signal \N__42093\ : std_logic;
signal \N__42092\ : std_logic;
signal \N__42091\ : std_logic;
signal \N__42090\ : std_logic;
signal \N__42089\ : std_logic;
signal \N__42088\ : std_logic;
signal \N__42087\ : std_logic;
signal \N__42086\ : std_logic;
signal \N__42077\ : std_logic;
signal \N__42072\ : std_logic;
signal \N__42071\ : std_logic;
signal \N__42068\ : std_logic;
signal \N__42067\ : std_logic;
signal \N__42066\ : std_logic;
signal \N__42065\ : std_logic;
signal \N__42064\ : std_logic;
signal \N__42063\ : std_logic;
signal \N__42062\ : std_logic;
signal \N__42061\ : std_logic;
signal \N__42060\ : std_logic;
signal \N__42059\ : std_logic;
signal \N__42058\ : std_logic;
signal \N__42057\ : std_logic;
signal \N__42056\ : std_logic;
signal \N__42055\ : std_logic;
signal \N__42054\ : std_logic;
signal \N__42053\ : std_logic;
signal \N__42052\ : std_logic;
signal \N__42051\ : std_logic;
signal \N__42050\ : std_logic;
signal \N__42049\ : std_logic;
signal \N__42048\ : std_logic;
signal \N__42047\ : std_logic;
signal \N__42044\ : std_logic;
signal \N__42043\ : std_logic;
signal \N__42042\ : std_logic;
signal \N__42041\ : std_logic;
signal \N__42034\ : std_logic;
signal \N__42033\ : std_logic;
signal \N__42032\ : std_logic;
signal \N__42031\ : std_logic;
signal \N__42030\ : std_logic;
signal \N__42027\ : std_logic;
signal \N__42026\ : std_logic;
signal \N__42025\ : std_logic;
signal \N__42024\ : std_logic;
signal \N__42023\ : std_logic;
signal \N__42022\ : std_logic;
signal \N__42021\ : std_logic;
signal \N__42020\ : std_logic;
signal \N__42019\ : std_logic;
signal \N__42016\ : std_logic;
signal \N__42015\ : std_logic;
signal \N__42014\ : std_logic;
signal \N__42013\ : std_logic;
signal \N__42012\ : std_logic;
signal \N__42011\ : std_logic;
signal \N__42010\ : std_logic;
signal \N__42009\ : std_logic;
signal \N__42006\ : std_logic;
signal \N__42005\ : std_logic;
signal \N__42004\ : std_logic;
signal \N__42003\ : std_logic;
signal \N__42002\ : std_logic;
signal \N__42001\ : std_logic;
signal \N__42000\ : std_logic;
signal \N__41999\ : std_logic;
signal \N__41998\ : std_logic;
signal \N__41997\ : std_logic;
signal \N__41988\ : std_logic;
signal \N__41979\ : std_logic;
signal \N__41978\ : std_logic;
signal \N__41977\ : std_logic;
signal \N__41976\ : std_logic;
signal \N__41975\ : std_logic;
signal \N__41974\ : std_logic;
signal \N__41969\ : std_logic;
signal \N__41968\ : std_logic;
signal \N__41967\ : std_logic;
signal \N__41966\ : std_logic;
signal \N__41965\ : std_logic;
signal \N__41964\ : std_logic;
signal \N__41963\ : std_logic;
signal \N__41960\ : std_logic;
signal \N__41953\ : std_logic;
signal \N__41948\ : std_logic;
signal \N__41945\ : std_logic;
signal \N__41944\ : std_logic;
signal \N__41943\ : std_logic;
signal \N__41940\ : std_logic;
signal \N__41939\ : std_logic;
signal \N__41938\ : std_logic;
signal \N__41937\ : std_logic;
signal \N__41936\ : std_logic;
signal \N__41935\ : std_logic;
signal \N__41932\ : std_logic;
signal \N__41923\ : std_logic;
signal \N__41914\ : std_logic;
signal \N__41905\ : std_logic;
signal \N__41896\ : std_logic;
signal \N__41893\ : std_logic;
signal \N__41886\ : std_logic;
signal \N__41879\ : std_logic;
signal \N__41876\ : std_logic;
signal \N__41875\ : std_logic;
signal \N__41872\ : std_logic;
signal \N__41869\ : std_logic;
signal \N__41868\ : std_logic;
signal \N__41867\ : std_logic;
signal \N__41866\ : std_logic;
signal \N__41865\ : std_logic;
signal \N__41864\ : std_logic;
signal \N__41863\ : std_logic;
signal \N__41862\ : std_logic;
signal \N__41855\ : std_logic;
signal \N__41850\ : std_logic;
signal \N__41843\ : std_logic;
signal \N__41836\ : std_logic;
signal \N__41827\ : std_logic;
signal \N__41820\ : std_logic;
signal \N__41815\ : std_logic;
signal \N__41814\ : std_logic;
signal \N__41813\ : std_logic;
signal \N__41812\ : std_logic;
signal \N__41811\ : std_logic;
signal \N__41810\ : std_logic;
signal \N__41807\ : std_logic;
signal \N__41806\ : std_logic;
signal \N__41805\ : std_logic;
signal \N__41802\ : std_logic;
signal \N__41793\ : std_logic;
signal \N__41786\ : std_logic;
signal \N__41783\ : std_logic;
signal \N__41772\ : std_logic;
signal \N__41763\ : std_logic;
signal \N__41754\ : std_logic;
signal \N__41753\ : std_logic;
signal \N__41752\ : std_logic;
signal \N__41751\ : std_logic;
signal \N__41750\ : std_logic;
signal \N__41749\ : std_logic;
signal \N__41748\ : std_logic;
signal \N__41747\ : std_logic;
signal \N__41746\ : std_logic;
signal \N__41745\ : std_logic;
signal \N__41744\ : std_logic;
signal \N__41743\ : std_logic;
signal \N__41742\ : std_logic;
signal \N__41739\ : std_logic;
signal \N__41732\ : std_logic;
signal \N__41729\ : std_logic;
signal \N__41724\ : std_logic;
signal \N__41713\ : std_logic;
signal \N__41704\ : std_logic;
signal \N__41695\ : std_logic;
signal \N__41688\ : std_logic;
signal \N__41681\ : std_logic;
signal \N__41680\ : std_logic;
signal \N__41679\ : std_logic;
signal \N__41672\ : std_logic;
signal \N__41663\ : std_logic;
signal \N__41658\ : std_logic;
signal \N__41657\ : std_logic;
signal \N__41656\ : std_logic;
signal \N__41655\ : std_logic;
signal \N__41654\ : std_logic;
signal \N__41653\ : std_logic;
signal \N__41652\ : std_logic;
signal \N__41649\ : std_logic;
signal \N__41648\ : std_logic;
signal \N__41647\ : std_logic;
signal \N__41646\ : std_logic;
signal \N__41645\ : std_logic;
signal \N__41644\ : std_logic;
signal \N__41643\ : std_logic;
signal \N__41642\ : std_logic;
signal \N__41641\ : std_logic;
signal \N__41640\ : std_logic;
signal \N__41639\ : std_logic;
signal \N__41638\ : std_logic;
signal \N__41633\ : std_logic;
signal \N__41632\ : std_logic;
signal \N__41631\ : std_logic;
signal \N__41630\ : std_logic;
signal \N__41629\ : std_logic;
signal \N__41628\ : std_logic;
signal \N__41627\ : std_logic;
signal \N__41620\ : std_logic;
signal \N__41619\ : std_logic;
signal \N__41618\ : std_logic;
signal \N__41617\ : std_logic;
signal \N__41616\ : std_logic;
signal \N__41615\ : std_logic;
signal \N__41614\ : std_logic;
signal \N__41613\ : std_logic;
signal \N__41612\ : std_logic;
signal \N__41611\ : std_logic;
signal \N__41610\ : std_logic;
signal \N__41609\ : std_logic;
signal \N__41608\ : std_logic;
signal \N__41607\ : std_logic;
signal \N__41606\ : std_logic;
signal \N__41605\ : std_logic;
signal \N__41604\ : std_logic;
signal \N__41601\ : std_logic;
signal \N__41600\ : std_logic;
signal \N__41599\ : std_logic;
signal \N__41598\ : std_logic;
signal \N__41597\ : std_logic;
signal \N__41596\ : std_logic;
signal \N__41593\ : std_logic;
signal \N__41592\ : std_logic;
signal \N__41591\ : std_logic;
signal \N__41590\ : std_logic;
signal \N__41589\ : std_logic;
signal \N__41586\ : std_logic;
signal \N__41579\ : std_logic;
signal \N__41578\ : std_logic;
signal \N__41577\ : std_logic;
signal \N__41574\ : std_logic;
signal \N__41573\ : std_logic;
signal \N__41572\ : std_logic;
signal \N__41569\ : std_logic;
signal \N__41568\ : std_logic;
signal \N__41567\ : std_logic;
signal \N__41566\ : std_logic;
signal \N__41565\ : std_logic;
signal \N__41562\ : std_logic;
signal \N__41561\ : std_logic;
signal \N__41560\ : std_logic;
signal \N__41559\ : std_logic;
signal \N__41552\ : std_logic;
signal \N__41549\ : std_logic;
signal \N__41540\ : std_logic;
signal \N__41531\ : std_logic;
signal \N__41524\ : std_logic;
signal \N__41519\ : std_logic;
signal \N__41512\ : std_logic;
signal \N__41509\ : std_logic;
signal \N__41502\ : std_logic;
signal \N__41499\ : std_logic;
signal \N__41496\ : std_logic;
signal \N__41493\ : std_logic;
signal \N__41490\ : std_logic;
signal \N__41487\ : std_logic;
signal \N__41484\ : std_logic;
signal \N__41483\ : std_logic;
signal \N__41480\ : std_logic;
signal \N__41479\ : std_logic;
signal \N__41478\ : std_logic;
signal \N__41477\ : std_logic;
signal \N__41476\ : std_logic;
signal \N__41475\ : std_logic;
signal \N__41474\ : std_logic;
signal \N__41473\ : std_logic;
signal \N__41472\ : std_logic;
signal \N__41467\ : std_logic;
signal \N__41462\ : std_logic;
signal \N__41457\ : std_logic;
signal \N__41454\ : std_logic;
signal \N__41445\ : std_logic;
signal \N__41436\ : std_logic;
signal \N__41421\ : std_logic;
signal \N__41414\ : std_logic;
signal \N__41407\ : std_logic;
signal \N__41400\ : std_logic;
signal \N__41393\ : std_logic;
signal \N__41390\ : std_logic;
signal \N__41387\ : std_logic;
signal \N__41372\ : std_logic;
signal \N__41367\ : std_logic;
signal \N__41360\ : std_logic;
signal \N__41353\ : std_logic;
signal \N__41342\ : std_logic;
signal \N__41333\ : std_logic;
signal \N__41324\ : std_logic;
signal \N__41323\ : std_logic;
signal \N__41322\ : std_logic;
signal \N__41321\ : std_logic;
signal \N__41318\ : std_logic;
signal \N__41317\ : std_logic;
signal \N__41316\ : std_logic;
signal \N__41315\ : std_logic;
signal \N__41314\ : std_logic;
signal \N__41311\ : std_logic;
signal \N__41310\ : std_logic;
signal \N__41309\ : std_logic;
signal \N__41308\ : std_logic;
signal \N__41305\ : std_logic;
signal \N__41298\ : std_logic;
signal \N__41291\ : std_logic;
signal \N__41288\ : std_logic;
signal \N__41285\ : std_logic;
signal \N__41278\ : std_logic;
signal \N__41271\ : std_logic;
signal \N__41264\ : std_logic;
signal \N__41259\ : std_logic;
signal \N__41252\ : std_logic;
signal \N__41241\ : std_logic;
signal \N__41232\ : std_logic;
signal \N__41227\ : std_logic;
signal \N__41224\ : std_logic;
signal \N__41219\ : std_logic;
signal \N__41210\ : std_logic;
signal \N__41201\ : std_logic;
signal \N__41192\ : std_logic;
signal \N__41187\ : std_logic;
signal \N__41184\ : std_logic;
signal \N__41177\ : std_logic;
signal \N__41174\ : std_logic;
signal \N__41169\ : std_logic;
signal \N__41164\ : std_logic;
signal \N__41157\ : std_logic;
signal \N__41146\ : std_logic;
signal \N__41137\ : std_logic;
signal \N__41128\ : std_logic;
signal \N__41123\ : std_logic;
signal \N__41116\ : std_logic;
signal \N__41103\ : std_logic;
signal \N__41094\ : std_logic;
signal \N__41083\ : std_logic;
signal \N__41078\ : std_logic;
signal \N__41069\ : std_logic;
signal \N__41064\ : std_logic;
signal \N__41055\ : std_logic;
signal \N__41042\ : std_logic;
signal \N__41037\ : std_logic;
signal \N__41014\ : std_logic;
signal \N__41009\ : std_logic;
signal \N__40994\ : std_logic;
signal \N__40987\ : std_logic;
signal \N__40974\ : std_logic;
signal \N__40971\ : std_logic;
signal \N__40966\ : std_logic;
signal \N__40961\ : std_logic;
signal \N__40956\ : std_logic;
signal \N__40947\ : std_logic;
signal \N__40946\ : std_logic;
signal \N__40943\ : std_logic;
signal \N__40940\ : std_logic;
signal \N__40937\ : std_logic;
signal \N__40934\ : std_logic;
signal \N__40929\ : std_logic;
signal \N__40928\ : std_logic;
signal \N__40927\ : std_logic;
signal \N__40926\ : std_logic;
signal \N__40923\ : std_logic;
signal \N__40922\ : std_logic;
signal \N__40921\ : std_logic;
signal \N__40918\ : std_logic;
signal \N__40915\ : std_logic;
signal \N__40914\ : std_logic;
signal \N__40911\ : std_logic;
signal \N__40908\ : std_logic;
signal \N__40907\ : std_logic;
signal \N__40904\ : std_logic;
signal \N__40903\ : std_logic;
signal \N__40902\ : std_logic;
signal \N__40901\ : std_logic;
signal \N__40900\ : std_logic;
signal \N__40899\ : std_logic;
signal \N__40898\ : std_logic;
signal \N__40895\ : std_logic;
signal \N__40894\ : std_logic;
signal \N__40891\ : std_logic;
signal \N__40886\ : std_logic;
signal \N__40881\ : std_logic;
signal \N__40874\ : std_logic;
signal \N__40871\ : std_logic;
signal \N__40868\ : std_logic;
signal \N__40865\ : std_logic;
signal \N__40864\ : std_logic;
signal \N__40863\ : std_logic;
signal \N__40862\ : std_logic;
signal \N__40861\ : std_logic;
signal \N__40860\ : std_logic;
signal \N__40859\ : std_logic;
signal \N__40856\ : std_logic;
signal \N__40849\ : std_logic;
signal \N__40840\ : std_logic;
signal \N__40835\ : std_logic;
signal \N__40828\ : std_logic;
signal \N__40819\ : std_logic;
signal \N__40806\ : std_logic;
signal \N__40803\ : std_logic;
signal \N__40802\ : std_logic;
signal \N__40799\ : std_logic;
signal \N__40796\ : std_logic;
signal \N__40793\ : std_logic;
signal \N__40790\ : std_logic;
signal \N__40787\ : std_logic;
signal \N__40784\ : std_logic;
signal \N__40779\ : std_logic;
signal \N__40776\ : std_logic;
signal \N__40773\ : std_logic;
signal \N__40770\ : std_logic;
signal \N__40769\ : std_logic;
signal \N__40766\ : std_logic;
signal \N__40763\ : std_logic;
signal \N__40758\ : std_logic;
signal \N__40755\ : std_logic;
signal \N__40752\ : std_logic;
signal \N__40749\ : std_logic;
signal \N__40746\ : std_logic;
signal \N__40743\ : std_logic;
signal \N__40740\ : std_logic;
signal \N__40737\ : std_logic;
signal \N__40736\ : std_logic;
signal \N__40733\ : std_logic;
signal \N__40730\ : std_logic;
signal \N__40729\ : std_logic;
signal \N__40726\ : std_logic;
signal \N__40723\ : std_logic;
signal \N__40720\ : std_logic;
signal \N__40717\ : std_logic;
signal \N__40714\ : std_logic;
signal \N__40707\ : std_logic;
signal \N__40704\ : std_logic;
signal \N__40701\ : std_logic;
signal \N__40698\ : std_logic;
signal \N__40695\ : std_logic;
signal \N__40692\ : std_logic;
signal \N__40691\ : std_logic;
signal \N__40690\ : std_logic;
signal \N__40687\ : std_logic;
signal \N__40684\ : std_logic;
signal \N__40681\ : std_logic;
signal \N__40674\ : std_logic;
signal \N__40671\ : std_logic;
signal \N__40668\ : std_logic;
signal \N__40665\ : std_logic;
signal \N__40662\ : std_logic;
signal \N__40659\ : std_logic;
signal \N__40658\ : std_logic;
signal \N__40655\ : std_logic;
signal \N__40652\ : std_logic;
signal \N__40647\ : std_logic;
signal \N__40644\ : std_logic;
signal \N__40641\ : std_logic;
signal \N__40638\ : std_logic;
signal \N__40637\ : std_logic;
signal \N__40634\ : std_logic;
signal \N__40631\ : std_logic;
signal \N__40628\ : std_logic;
signal \N__40623\ : std_logic;
signal \N__40620\ : std_logic;
signal \N__40617\ : std_logic;
signal \N__40614\ : std_logic;
signal \N__40611\ : std_logic;
signal \N__40608\ : std_logic;
signal \N__40605\ : std_logic;
signal \N__40604\ : std_logic;
signal \N__40601\ : std_logic;
signal \N__40600\ : std_logic;
signal \N__40597\ : std_logic;
signal \N__40594\ : std_logic;
signal \N__40591\ : std_logic;
signal \N__40584\ : std_logic;
signal \N__40581\ : std_logic;
signal \N__40578\ : std_logic;
signal \N__40575\ : std_logic;
signal \N__40572\ : std_logic;
signal \N__40569\ : std_logic;
signal \N__40566\ : std_logic;
signal \N__40565\ : std_logic;
signal \N__40562\ : std_logic;
signal \N__40559\ : std_logic;
signal \N__40558\ : std_logic;
signal \N__40555\ : std_logic;
signal \N__40552\ : std_logic;
signal \N__40549\ : std_logic;
signal \N__40542\ : std_logic;
signal \N__40539\ : std_logic;
signal \N__40536\ : std_logic;
signal \N__40533\ : std_logic;
signal \N__40530\ : std_logic;
signal \N__40527\ : std_logic;
signal \N__40524\ : std_logic;
signal \N__40523\ : std_logic;
signal \N__40520\ : std_logic;
signal \N__40517\ : std_logic;
signal \N__40516\ : std_logic;
signal \N__40513\ : std_logic;
signal \N__40510\ : std_logic;
signal \N__40507\ : std_logic;
signal \N__40500\ : std_logic;
signal \N__40497\ : std_logic;
signal \N__40494\ : std_logic;
signal \N__40491\ : std_logic;
signal \N__40488\ : std_logic;
signal \N__40485\ : std_logic;
signal \N__40482\ : std_logic;
signal \N__40479\ : std_logic;
signal \N__40476\ : std_logic;
signal \N__40475\ : std_logic;
signal \N__40474\ : std_logic;
signal \N__40471\ : std_logic;
signal \N__40466\ : std_logic;
signal \N__40463\ : std_logic;
signal \N__40458\ : std_logic;
signal \N__40455\ : std_logic;
signal \N__40452\ : std_logic;
signal \N__40449\ : std_logic;
signal \N__40446\ : std_logic;
signal \N__40445\ : std_logic;
signal \N__40442\ : std_logic;
signal \N__40439\ : std_logic;
signal \N__40436\ : std_logic;
signal \N__40433\ : std_logic;
signal \N__40428\ : std_logic;
signal \N__40425\ : std_logic;
signal \N__40422\ : std_logic;
signal \N__40419\ : std_logic;
signal \N__40416\ : std_logic;
signal \N__40415\ : std_logic;
signal \N__40412\ : std_logic;
signal \N__40409\ : std_logic;
signal \N__40408\ : std_logic;
signal \N__40405\ : std_logic;
signal \N__40402\ : std_logic;
signal \N__40399\ : std_logic;
signal \N__40396\ : std_logic;
signal \N__40389\ : std_logic;
signal \N__40386\ : std_logic;
signal \N__40383\ : std_logic;
signal \N__40380\ : std_logic;
signal \N__40377\ : std_logic;
signal \N__40374\ : std_logic;
signal \N__40373\ : std_logic;
signal \N__40372\ : std_logic;
signal \N__40369\ : std_logic;
signal \N__40366\ : std_logic;
signal \N__40363\ : std_logic;
signal \N__40360\ : std_logic;
signal \N__40357\ : std_logic;
signal \N__40354\ : std_logic;
signal \N__40347\ : std_logic;
signal \N__40344\ : std_logic;
signal \N__40341\ : std_logic;
signal \N__40338\ : std_logic;
signal \N__40335\ : std_logic;
signal \N__40332\ : std_logic;
signal \N__40329\ : std_logic;
signal \N__40326\ : std_logic;
signal \N__40323\ : std_logic;
signal \N__40322\ : std_logic;
signal \N__40321\ : std_logic;
signal \N__40318\ : std_logic;
signal \N__40315\ : std_logic;
signal \N__40312\ : std_logic;
signal \N__40309\ : std_logic;
signal \N__40302\ : std_logic;
signal \N__40299\ : std_logic;
signal \N__40296\ : std_logic;
signal \N__40293\ : std_logic;
signal \N__40290\ : std_logic;
signal \N__40287\ : std_logic;
signal \N__40284\ : std_logic;
signal \N__40283\ : std_logic;
signal \N__40280\ : std_logic;
signal \N__40277\ : std_logic;
signal \N__40274\ : std_logic;
signal \N__40271\ : std_logic;
signal \N__40268\ : std_logic;
signal \N__40263\ : std_logic;
signal \N__40260\ : std_logic;
signal \N__40257\ : std_logic;
signal \N__40254\ : std_logic;
signal \N__40251\ : std_logic;
signal \N__40248\ : std_logic;
signal \N__40245\ : std_logic;
signal \N__40242\ : std_logic;
signal \N__40241\ : std_logic;
signal \N__40238\ : std_logic;
signal \N__40237\ : std_logic;
signal \N__40234\ : std_logic;
signal \N__40231\ : std_logic;
signal \N__40228\ : std_logic;
signal \N__40221\ : std_logic;
signal \N__40218\ : std_logic;
signal \N__40215\ : std_logic;
signal \N__40212\ : std_logic;
signal \N__40209\ : std_logic;
signal \N__40206\ : std_logic;
signal \N__40203\ : std_logic;
signal \N__40202\ : std_logic;
signal \N__40201\ : std_logic;
signal \N__40198\ : std_logic;
signal \N__40195\ : std_logic;
signal \N__40192\ : std_logic;
signal \N__40189\ : std_logic;
signal \N__40186\ : std_logic;
signal \N__40181\ : std_logic;
signal \N__40176\ : std_logic;
signal \N__40173\ : std_logic;
signal \N__40170\ : std_logic;
signal \N__40167\ : std_logic;
signal \N__40164\ : std_logic;
signal \N__40163\ : std_logic;
signal \N__40160\ : std_logic;
signal \N__40159\ : std_logic;
signal \N__40156\ : std_logic;
signal \N__40153\ : std_logic;
signal \N__40148\ : std_logic;
signal \N__40145\ : std_logic;
signal \N__40142\ : std_logic;
signal \N__40137\ : std_logic;
signal \N__40134\ : std_logic;
signal \N__40131\ : std_logic;
signal \N__40128\ : std_logic;
signal \N__40125\ : std_logic;
signal \N__40122\ : std_logic;
signal \N__40119\ : std_logic;
signal \N__40116\ : std_logic;
signal \N__40113\ : std_logic;
signal \N__40110\ : std_logic;
signal \N__40107\ : std_logic;
signal \N__40106\ : std_logic;
signal \N__40105\ : std_logic;
signal \N__40102\ : std_logic;
signal \N__40101\ : std_logic;
signal \N__40100\ : std_logic;
signal \N__40099\ : std_logic;
signal \N__40098\ : std_logic;
signal \N__40097\ : std_logic;
signal \N__40096\ : std_logic;
signal \N__40095\ : std_logic;
signal \N__40094\ : std_logic;
signal \N__40093\ : std_logic;
signal \N__40092\ : std_logic;
signal \N__40091\ : std_logic;
signal \N__40088\ : std_logic;
signal \N__40085\ : std_logic;
signal \N__40080\ : std_logic;
signal \N__40079\ : std_logic;
signal \N__40078\ : std_logic;
signal \N__40077\ : std_logic;
signal \N__40076\ : std_logic;
signal \N__40065\ : std_logic;
signal \N__40062\ : std_logic;
signal \N__40059\ : std_logic;
signal \N__40058\ : std_logic;
signal \N__40055\ : std_logic;
signal \N__40052\ : std_logic;
signal \N__40051\ : std_logic;
signal \N__40048\ : std_logic;
signal \N__40047\ : std_logic;
signal \N__40046\ : std_logic;
signal \N__40039\ : std_logic;
signal \N__40034\ : std_logic;
signal \N__40031\ : std_logic;
signal \N__40028\ : std_logic;
signal \N__40023\ : std_logic;
signal \N__40012\ : std_logic;
signal \N__40005\ : std_logic;
signal \N__40002\ : std_logic;
signal \N__39987\ : std_logic;
signal \N__39984\ : std_logic;
signal \N__39983\ : std_logic;
signal \N__39980\ : std_logic;
signal \N__39977\ : std_logic;
signal \N__39974\ : std_logic;
signal \N__39971\ : std_logic;
signal \N__39968\ : std_logic;
signal \N__39965\ : std_logic;
signal \N__39962\ : std_logic;
signal \N__39959\ : std_logic;
signal \N__39956\ : std_logic;
signal \N__39951\ : std_logic;
signal \N__39950\ : std_logic;
signal \N__39949\ : std_logic;
signal \N__39944\ : std_logic;
signal \N__39941\ : std_logic;
signal \N__39938\ : std_logic;
signal \N__39935\ : std_logic;
signal \N__39932\ : std_logic;
signal \N__39927\ : std_logic;
signal \N__39924\ : std_logic;
signal \N__39923\ : std_logic;
signal \N__39922\ : std_logic;
signal \N__39921\ : std_logic;
signal \N__39918\ : std_logic;
signal \N__39915\ : std_logic;
signal \N__39912\ : std_logic;
signal \N__39909\ : std_logic;
signal \N__39906\ : std_logic;
signal \N__39903\ : std_logic;
signal \N__39900\ : std_logic;
signal \N__39899\ : std_logic;
signal \N__39896\ : std_logic;
signal \N__39893\ : std_logic;
signal \N__39890\ : std_logic;
signal \N__39887\ : std_logic;
signal \N__39884\ : std_logic;
signal \N__39881\ : std_logic;
signal \N__39878\ : std_logic;
signal \N__39873\ : std_logic;
signal \N__39864\ : std_logic;
signal \N__39861\ : std_logic;
signal \N__39858\ : std_logic;
signal \N__39855\ : std_logic;
signal \N__39852\ : std_logic;
signal \N__39849\ : std_logic;
signal \N__39848\ : std_logic;
signal \N__39845\ : std_logic;
signal \N__39842\ : std_logic;
signal \N__39839\ : std_logic;
signal \N__39838\ : std_logic;
signal \N__39835\ : std_logic;
signal \N__39832\ : std_logic;
signal \N__39829\ : std_logic;
signal \N__39824\ : std_logic;
signal \N__39819\ : std_logic;
signal \N__39816\ : std_logic;
signal \N__39813\ : std_logic;
signal \N__39810\ : std_logic;
signal \N__39807\ : std_logic;
signal \N__39806\ : std_logic;
signal \N__39805\ : std_logic;
signal \N__39802\ : std_logic;
signal \N__39797\ : std_logic;
signal \N__39794\ : std_logic;
signal \N__39789\ : std_logic;
signal \N__39786\ : std_logic;
signal \N__39783\ : std_logic;
signal \N__39780\ : std_logic;
signal \N__39777\ : std_logic;
signal \N__39774\ : std_logic;
signal \N__39771\ : std_logic;
signal \N__39770\ : std_logic;
signal \N__39767\ : std_logic;
signal \N__39764\ : std_logic;
signal \N__39761\ : std_logic;
signal \N__39758\ : std_logic;
signal \N__39755\ : std_logic;
signal \N__39752\ : std_logic;
signal \N__39747\ : std_logic;
signal \N__39744\ : std_logic;
signal \N__39741\ : std_logic;
signal \N__39738\ : std_logic;
signal \N__39735\ : std_logic;
signal \N__39732\ : std_logic;
signal \N__39731\ : std_logic;
signal \N__39728\ : std_logic;
signal \N__39727\ : std_logic;
signal \N__39724\ : std_logic;
signal \N__39721\ : std_logic;
signal \N__39718\ : std_logic;
signal \N__39715\ : std_logic;
signal \N__39710\ : std_logic;
signal \N__39705\ : std_logic;
signal \N__39702\ : std_logic;
signal \N__39699\ : std_logic;
signal \N__39696\ : std_logic;
signal \N__39693\ : std_logic;
signal \N__39690\ : std_logic;
signal \N__39687\ : std_logic;
signal \N__39684\ : std_logic;
signal \N__39683\ : std_logic;
signal \N__39680\ : std_logic;
signal \N__39677\ : std_logic;
signal \N__39674\ : std_logic;
signal \N__39669\ : std_logic;
signal \N__39666\ : std_logic;
signal \N__39663\ : std_logic;
signal \N__39660\ : std_logic;
signal \N__39657\ : std_logic;
signal \N__39654\ : std_logic;
signal \N__39651\ : std_logic;
signal \N__39648\ : std_logic;
signal \N__39645\ : std_logic;
signal \N__39644\ : std_logic;
signal \N__39643\ : std_logic;
signal \N__39640\ : std_logic;
signal \N__39637\ : std_logic;
signal \N__39634\ : std_logic;
signal \N__39631\ : std_logic;
signal \N__39628\ : std_logic;
signal \N__39625\ : std_logic;
signal \N__39618\ : std_logic;
signal \N__39615\ : std_logic;
signal \N__39612\ : std_logic;
signal \N__39609\ : std_logic;
signal \N__39606\ : std_logic;
signal \N__39603\ : std_logic;
signal \N__39600\ : std_logic;
signal \N__39599\ : std_logic;
signal \N__39596\ : std_logic;
signal \N__39593\ : std_logic;
signal \N__39592\ : std_logic;
signal \N__39589\ : std_logic;
signal \N__39586\ : std_logic;
signal \N__39583\ : std_logic;
signal \N__39580\ : std_logic;
signal \N__39577\ : std_logic;
signal \N__39574\ : std_logic;
signal \N__39567\ : std_logic;
signal \N__39564\ : std_logic;
signal \N__39561\ : std_logic;
signal \N__39558\ : std_logic;
signal \N__39555\ : std_logic;
signal \N__39552\ : std_logic;
signal \N__39549\ : std_logic;
signal \N__39546\ : std_logic;
signal \N__39545\ : std_logic;
signal \N__39542\ : std_logic;
signal \N__39539\ : std_logic;
signal \N__39538\ : std_logic;
signal \N__39535\ : std_logic;
signal \N__39532\ : std_logic;
signal \N__39529\ : std_logic;
signal \N__39522\ : std_logic;
signal \N__39519\ : std_logic;
signal \N__39516\ : std_logic;
signal \N__39513\ : std_logic;
signal \N__39510\ : std_logic;
signal \N__39507\ : std_logic;
signal \N__39504\ : std_logic;
signal \N__39501\ : std_logic;
signal \N__39498\ : std_logic;
signal \N__39495\ : std_logic;
signal \N__39494\ : std_logic;
signal \N__39491\ : std_logic;
signal \N__39488\ : std_logic;
signal \N__39487\ : std_logic;
signal \N__39484\ : std_logic;
signal \N__39481\ : std_logic;
signal \N__39478\ : std_logic;
signal \N__39471\ : std_logic;
signal \N__39468\ : std_logic;
signal \N__39465\ : std_logic;
signal \N__39462\ : std_logic;
signal \N__39459\ : std_logic;
signal \N__39456\ : std_logic;
signal \N__39453\ : std_logic;
signal \N__39452\ : std_logic;
signal \N__39449\ : std_logic;
signal \N__39446\ : std_logic;
signal \N__39443\ : std_logic;
signal \N__39440\ : std_logic;
signal \N__39435\ : std_logic;
signal \N__39432\ : std_logic;
signal \N__39429\ : std_logic;
signal \N__39426\ : std_logic;
signal \N__39423\ : std_logic;
signal \N__39420\ : std_logic;
signal \N__39417\ : std_logic;
signal \N__39414\ : std_logic;
signal \N__39411\ : std_logic;
signal \N__39410\ : std_logic;
signal \N__39407\ : std_logic;
signal \N__39404\ : std_logic;
signal \N__39401\ : std_logic;
signal \N__39400\ : std_logic;
signal \N__39397\ : std_logic;
signal \N__39394\ : std_logic;
signal \N__39391\ : std_logic;
signal \N__39384\ : std_logic;
signal \N__39381\ : std_logic;
signal \N__39378\ : std_logic;
signal \N__39375\ : std_logic;
signal \N__39372\ : std_logic;
signal \N__39369\ : std_logic;
signal \N__39368\ : std_logic;
signal \N__39365\ : std_logic;
signal \N__39362\ : std_logic;
signal \N__39359\ : std_logic;
signal \N__39356\ : std_logic;
signal \N__39351\ : std_logic;
signal \N__39348\ : std_logic;
signal \N__39345\ : std_logic;
signal \N__39342\ : std_logic;
signal \N__39339\ : std_logic;
signal \N__39338\ : std_logic;
signal \N__39337\ : std_logic;
signal \N__39334\ : std_logic;
signal \N__39331\ : std_logic;
signal \N__39328\ : std_logic;
signal \N__39325\ : std_logic;
signal \N__39322\ : std_logic;
signal \N__39315\ : std_logic;
signal \N__39312\ : std_logic;
signal \N__39309\ : std_logic;
signal \N__39306\ : std_logic;
signal \N__39305\ : std_logic;
signal \N__39304\ : std_logic;
signal \N__39301\ : std_logic;
signal \N__39298\ : std_logic;
signal \N__39295\ : std_logic;
signal \N__39292\ : std_logic;
signal \N__39289\ : std_logic;
signal \N__39284\ : std_logic;
signal \N__39281\ : std_logic;
signal \N__39278\ : std_logic;
signal \N__39273\ : std_logic;
signal \N__39270\ : std_logic;
signal \N__39267\ : std_logic;
signal \N__39264\ : std_logic;
signal \N__39261\ : std_logic;
signal \N__39258\ : std_logic;
signal \N__39255\ : std_logic;
signal \N__39252\ : std_logic;
signal \N__39251\ : std_logic;
signal \N__39248\ : std_logic;
signal \N__39245\ : std_logic;
signal \N__39242\ : std_logic;
signal \N__39237\ : std_logic;
signal \N__39234\ : std_logic;
signal \N__39231\ : std_logic;
signal \N__39228\ : std_logic;
signal \N__39225\ : std_logic;
signal \N__39222\ : std_logic;
signal \N__39221\ : std_logic;
signal \N__39218\ : std_logic;
signal \N__39215\ : std_logic;
signal \N__39214\ : std_logic;
signal \N__39211\ : std_logic;
signal \N__39208\ : std_logic;
signal \N__39205\ : std_logic;
signal \N__39202\ : std_logic;
signal \N__39195\ : std_logic;
signal \N__39192\ : std_logic;
signal \N__39189\ : std_logic;
signal \N__39186\ : std_logic;
signal \N__39183\ : std_logic;
signal \N__39180\ : std_logic;
signal \N__39177\ : std_logic;
signal \N__39174\ : std_logic;
signal \N__39173\ : std_logic;
signal \N__39170\ : std_logic;
signal \N__39169\ : std_logic;
signal \N__39166\ : std_logic;
signal \N__39163\ : std_logic;
signal \N__39160\ : std_logic;
signal \N__39153\ : std_logic;
signal \N__39150\ : std_logic;
signal \N__39147\ : std_logic;
signal \N__39144\ : std_logic;
signal \N__39141\ : std_logic;
signal \N__39138\ : std_logic;
signal \N__39137\ : std_logic;
signal \N__39134\ : std_logic;
signal \N__39131\ : std_logic;
signal \N__39128\ : std_logic;
signal \N__39125\ : std_logic;
signal \N__39124\ : std_logic;
signal \N__39121\ : std_logic;
signal \N__39118\ : std_logic;
signal \N__39115\ : std_logic;
signal \N__39108\ : std_logic;
signal \N__39105\ : std_logic;
signal \N__39102\ : std_logic;
signal \N__39099\ : std_logic;
signal \N__39096\ : std_logic;
signal \N__39093\ : std_logic;
signal \N__39090\ : std_logic;
signal \N__39087\ : std_logic;
signal \N__39086\ : std_logic;
signal \N__39083\ : std_logic;
signal \N__39080\ : std_logic;
signal \N__39079\ : std_logic;
signal \N__39076\ : std_logic;
signal \N__39073\ : std_logic;
signal \N__39070\ : std_logic;
signal \N__39067\ : std_logic;
signal \N__39062\ : std_logic;
signal \N__39057\ : std_logic;
signal \N__39054\ : std_logic;
signal \N__39051\ : std_logic;
signal \N__39048\ : std_logic;
signal \N__39045\ : std_logic;
signal \N__39042\ : std_logic;
signal \N__39039\ : std_logic;
signal \N__39036\ : std_logic;
signal \N__39033\ : std_logic;
signal \N__39030\ : std_logic;
signal \N__39027\ : std_logic;
signal \N__39024\ : std_logic;
signal \N__39021\ : std_logic;
signal \N__39020\ : std_logic;
signal \N__39019\ : std_logic;
signal \N__39016\ : std_logic;
signal \N__39013\ : std_logic;
signal \N__39010\ : std_logic;
signal \N__39003\ : std_logic;
signal \N__39000\ : std_logic;
signal \N__38997\ : std_logic;
signal \N__38994\ : std_logic;
signal \N__38991\ : std_logic;
signal \N__38988\ : std_logic;
signal \N__38985\ : std_logic;
signal \N__38982\ : std_logic;
signal \N__38979\ : std_logic;
signal \N__38978\ : std_logic;
signal \N__38977\ : std_logic;
signal \N__38974\ : std_logic;
signal \N__38969\ : std_logic;
signal \N__38964\ : std_logic;
signal \N__38961\ : std_logic;
signal \N__38958\ : std_logic;
signal \N__38955\ : std_logic;
signal \N__38952\ : std_logic;
signal \N__38949\ : std_logic;
signal \N__38946\ : std_logic;
signal \N__38943\ : std_logic;
signal \N__38942\ : std_logic;
signal \N__38939\ : std_logic;
signal \N__38936\ : std_logic;
signal \N__38931\ : std_logic;
signal \N__38928\ : std_logic;
signal \N__38927\ : std_logic;
signal \N__38924\ : std_logic;
signal \N__38921\ : std_logic;
signal \N__38920\ : std_logic;
signal \N__38917\ : std_logic;
signal \N__38914\ : std_logic;
signal \N__38913\ : std_logic;
signal \N__38912\ : std_logic;
signal \N__38909\ : std_logic;
signal \N__38906\ : std_logic;
signal \N__38903\ : std_logic;
signal \N__38900\ : std_logic;
signal \N__38897\ : std_logic;
signal \N__38890\ : std_logic;
signal \N__38883\ : std_logic;
signal \N__38880\ : std_logic;
signal \N__38877\ : std_logic;
signal \N__38874\ : std_logic;
signal \N__38871\ : std_logic;
signal \N__38868\ : std_logic;
signal \N__38865\ : std_logic;
signal \N__38862\ : std_logic;
signal \N__38861\ : std_logic;
signal \N__38858\ : std_logic;
signal \N__38855\ : std_logic;
signal \N__38852\ : std_logic;
signal \N__38849\ : std_logic;
signal \N__38844\ : std_logic;
signal \N__38841\ : std_logic;
signal \N__38838\ : std_logic;
signal \N__38835\ : std_logic;
signal \N__38832\ : std_logic;
signal \N__38829\ : std_logic;
signal \N__38826\ : std_logic;
signal \N__38825\ : std_logic;
signal \N__38822\ : std_logic;
signal \N__38821\ : std_logic;
signal \N__38818\ : std_logic;
signal \N__38815\ : std_logic;
signal \N__38812\ : std_logic;
signal \N__38809\ : std_logic;
signal \N__38802\ : std_logic;
signal \N__38799\ : std_logic;
signal \N__38796\ : std_logic;
signal \N__38793\ : std_logic;
signal \N__38790\ : std_logic;
signal \N__38787\ : std_logic;
signal \N__38784\ : std_logic;
signal \N__38781\ : std_logic;
signal \N__38780\ : std_logic;
signal \N__38777\ : std_logic;
signal \N__38774\ : std_logic;
signal \N__38773\ : std_logic;
signal \N__38770\ : std_logic;
signal \N__38767\ : std_logic;
signal \N__38764\ : std_logic;
signal \N__38757\ : std_logic;
signal \N__38754\ : std_logic;
signal \N__38751\ : std_logic;
signal \N__38748\ : std_logic;
signal \N__38745\ : std_logic;
signal \N__38742\ : std_logic;
signal \N__38739\ : std_logic;
signal \N__38736\ : std_logic;
signal \N__38733\ : std_logic;
signal \N__38730\ : std_logic;
signal \N__38727\ : std_logic;
signal \N__38724\ : std_logic;
signal \N__38721\ : std_logic;
signal \N__38718\ : std_logic;
signal \N__38715\ : std_logic;
signal \N__38712\ : std_logic;
signal \N__38711\ : std_logic;
signal \N__38708\ : std_logic;
signal \N__38707\ : std_logic;
signal \N__38704\ : std_logic;
signal \N__38701\ : std_logic;
signal \N__38698\ : std_logic;
signal \N__38695\ : std_logic;
signal \N__38688\ : std_logic;
signal \N__38685\ : std_logic;
signal \N__38682\ : std_logic;
signal \N__38679\ : std_logic;
signal \N__38676\ : std_logic;
signal \N__38673\ : std_logic;
signal \N__38672\ : std_logic;
signal \N__38671\ : std_logic;
signal \N__38668\ : std_logic;
signal \N__38665\ : std_logic;
signal \N__38662\ : std_logic;
signal \N__38655\ : std_logic;
signal \N__38652\ : std_logic;
signal \N__38649\ : std_logic;
signal \N__38646\ : std_logic;
signal \N__38643\ : std_logic;
signal \N__38640\ : std_logic;
signal \N__38637\ : std_logic;
signal \N__38634\ : std_logic;
signal \N__38631\ : std_logic;
signal \N__38628\ : std_logic;
signal \N__38627\ : std_logic;
signal \N__38624\ : std_logic;
signal \N__38621\ : std_logic;
signal \N__38616\ : std_logic;
signal \N__38613\ : std_logic;
signal \N__38610\ : std_logic;
signal \N__38607\ : std_logic;
signal \N__38604\ : std_logic;
signal \N__38603\ : std_logic;
signal \N__38600\ : std_logic;
signal \N__38597\ : std_logic;
signal \N__38592\ : std_logic;
signal \N__38591\ : std_logic;
signal \N__38588\ : std_logic;
signal \N__38585\ : std_logic;
signal \N__38582\ : std_logic;
signal \N__38579\ : std_logic;
signal \N__38574\ : std_logic;
signal \N__38573\ : std_logic;
signal \N__38570\ : std_logic;
signal \N__38567\ : std_logic;
signal \N__38562\ : std_logic;
signal \N__38559\ : std_logic;
signal \N__38556\ : std_logic;
signal \N__38553\ : std_logic;
signal \N__38550\ : std_logic;
signal \N__38547\ : std_logic;
signal \N__38544\ : std_logic;
signal \N__38541\ : std_logic;
signal \N__38538\ : std_logic;
signal \N__38535\ : std_logic;
signal \N__38532\ : std_logic;
signal \N__38531\ : std_logic;
signal \N__38528\ : std_logic;
signal \N__38525\ : std_logic;
signal \N__38522\ : std_logic;
signal \N__38519\ : std_logic;
signal \N__38518\ : std_logic;
signal \N__38513\ : std_logic;
signal \N__38510\ : std_logic;
signal \N__38505\ : std_logic;
signal \N__38504\ : std_logic;
signal \N__38503\ : std_logic;
signal \N__38502\ : std_logic;
signal \N__38501\ : std_logic;
signal \N__38500\ : std_logic;
signal \N__38499\ : std_logic;
signal \N__38498\ : std_logic;
signal \N__38497\ : std_logic;
signal \N__38496\ : std_logic;
signal \N__38493\ : std_logic;
signal \N__38492\ : std_logic;
signal \N__38489\ : std_logic;
signal \N__38488\ : std_logic;
signal \N__38487\ : std_logic;
signal \N__38482\ : std_logic;
signal \N__38479\ : std_logic;
signal \N__38478\ : std_logic;
signal \N__38475\ : std_logic;
signal \N__38474\ : std_logic;
signal \N__38471\ : std_logic;
signal \N__38470\ : std_logic;
signal \N__38469\ : std_logic;
signal \N__38466\ : std_logic;
signal \N__38465\ : std_logic;
signal \N__38462\ : std_logic;
signal \N__38461\ : std_logic;
signal \N__38460\ : std_logic;
signal \N__38457\ : std_logic;
signal \N__38456\ : std_logic;
signal \N__38445\ : std_logic;
signal \N__38440\ : std_logic;
signal \N__38437\ : std_logic;
signal \N__38434\ : std_logic;
signal \N__38431\ : std_logic;
signal \N__38424\ : std_logic;
signal \N__38419\ : std_logic;
signal \N__38408\ : std_logic;
signal \N__38391\ : std_logic;
signal \N__38390\ : std_logic;
signal \N__38387\ : std_logic;
signal \N__38384\ : std_logic;
signal \N__38379\ : std_logic;
signal \N__38376\ : std_logic;
signal \N__38373\ : std_logic;
signal \N__38370\ : std_logic;
signal \N__38367\ : std_logic;
signal \N__38364\ : std_logic;
signal \N__38361\ : std_logic;
signal \N__38358\ : std_logic;
signal \N__38355\ : std_logic;
signal \N__38352\ : std_logic;
signal \N__38349\ : std_logic;
signal \N__38346\ : std_logic;
signal \N__38345\ : std_logic;
signal \N__38342\ : std_logic;
signal \N__38339\ : std_logic;
signal \N__38334\ : std_logic;
signal \N__38331\ : std_logic;
signal \N__38328\ : std_logic;
signal \N__38325\ : std_logic;
signal \N__38322\ : std_logic;
signal \N__38321\ : std_logic;
signal \N__38318\ : std_logic;
signal \N__38317\ : std_logic;
signal \N__38314\ : std_logic;
signal \N__38311\ : std_logic;
signal \N__38308\ : std_logic;
signal \N__38305\ : std_logic;
signal \N__38298\ : std_logic;
signal \N__38297\ : std_logic;
signal \N__38294\ : std_logic;
signal \N__38291\ : std_logic;
signal \N__38290\ : std_logic;
signal \N__38287\ : std_logic;
signal \N__38284\ : std_logic;
signal \N__38281\ : std_logic;
signal \N__38278\ : std_logic;
signal \N__38273\ : std_logic;
signal \N__38268\ : std_logic;
signal \N__38265\ : std_logic;
signal \N__38262\ : std_logic;
signal \N__38259\ : std_logic;
signal \N__38258\ : std_logic;
signal \N__38255\ : std_logic;
signal \N__38254\ : std_logic;
signal \N__38251\ : std_logic;
signal \N__38248\ : std_logic;
signal \N__38245\ : std_logic;
signal \N__38242\ : std_logic;
signal \N__38239\ : std_logic;
signal \N__38236\ : std_logic;
signal \N__38229\ : std_logic;
signal \N__38226\ : std_logic;
signal \N__38223\ : std_logic;
signal \N__38220\ : std_logic;
signal \N__38217\ : std_logic;
signal \N__38214\ : std_logic;
signal \N__38211\ : std_logic;
signal \N__38208\ : std_logic;
signal \N__38205\ : std_logic;
signal \N__38204\ : std_logic;
signal \N__38201\ : std_logic;
signal \N__38198\ : std_logic;
signal \N__38195\ : std_logic;
signal \N__38192\ : std_logic;
signal \N__38187\ : std_logic;
signal \N__38184\ : std_logic;
signal \N__38181\ : std_logic;
signal \N__38180\ : std_logic;
signal \N__38177\ : std_logic;
signal \N__38174\ : std_logic;
signal \N__38173\ : std_logic;
signal \N__38170\ : std_logic;
signal \N__38167\ : std_logic;
signal \N__38164\ : std_logic;
signal \N__38157\ : std_logic;
signal \N__38154\ : std_logic;
signal \N__38151\ : std_logic;
signal \N__38148\ : std_logic;
signal \N__38147\ : std_logic;
signal \N__38144\ : std_logic;
signal \N__38143\ : std_logic;
signal \N__38140\ : std_logic;
signal \N__38137\ : std_logic;
signal \N__38134\ : std_logic;
signal \N__38131\ : std_logic;
signal \N__38128\ : std_logic;
signal \N__38125\ : std_logic;
signal \N__38118\ : std_logic;
signal \N__38115\ : std_logic;
signal \N__38112\ : std_logic;
signal \N__38109\ : std_logic;
signal \N__38106\ : std_logic;
signal \N__38105\ : std_logic;
signal \N__38104\ : std_logic;
signal \N__38101\ : std_logic;
signal \N__38098\ : std_logic;
signal \N__38095\ : std_logic;
signal \N__38092\ : std_logic;
signal \N__38089\ : std_logic;
signal \N__38086\ : std_logic;
signal \N__38079\ : std_logic;
signal \N__38076\ : std_logic;
signal \N__38073\ : std_logic;
signal \N__38070\ : std_logic;
signal \N__38067\ : std_logic;
signal \N__38064\ : std_logic;
signal \N__38061\ : std_logic;
signal \N__38058\ : std_logic;
signal \N__38055\ : std_logic;
signal \N__38054\ : std_logic;
signal \N__38051\ : std_logic;
signal \N__38048\ : std_logic;
signal \N__38043\ : std_logic;
signal \N__38040\ : std_logic;
signal \N__38037\ : std_logic;
signal \N__38034\ : std_logic;
signal \N__38031\ : std_logic;
signal \N__38028\ : std_logic;
signal \N__38025\ : std_logic;
signal \N__38022\ : std_logic;
signal \N__38021\ : std_logic;
signal \N__38018\ : std_logic;
signal \N__38017\ : std_logic;
signal \N__38016\ : std_logic;
signal \N__38015\ : std_logic;
signal \N__38014\ : std_logic;
signal \N__38013\ : std_logic;
signal \N__38012\ : std_logic;
signal \N__38011\ : std_logic;
signal \N__38010\ : std_logic;
signal \N__38009\ : std_logic;
signal \N__38008\ : std_logic;
signal \N__38005\ : std_logic;
signal \N__38004\ : std_logic;
signal \N__38001\ : std_logic;
signal \N__38000\ : std_logic;
signal \N__37999\ : std_logic;
signal \N__37996\ : std_logic;
signal \N__37995\ : std_logic;
signal \N__37992\ : std_logic;
signal \N__37989\ : std_logic;
signal \N__37988\ : std_logic;
signal \N__37987\ : std_logic;
signal \N__37978\ : std_logic;
signal \N__37975\ : std_logic;
signal \N__37972\ : std_logic;
signal \N__37969\ : std_logic;
signal \N__37968\ : std_logic;
signal \N__37967\ : std_logic;
signal \N__37964\ : std_logic;
signal \N__37961\ : std_logic;
signal \N__37958\ : std_logic;
signal \N__37949\ : std_logic;
signal \N__37944\ : std_logic;
signal \N__37939\ : std_logic;
signal \N__37936\ : std_logic;
signal \N__37925\ : std_logic;
signal \N__37920\ : std_logic;
signal \N__37905\ : std_logic;
signal \N__37902\ : std_logic;
signal \N__37899\ : std_logic;
signal \N__37898\ : std_logic;
signal \N__37897\ : std_logic;
signal \N__37896\ : std_logic;
signal \N__37893\ : std_logic;
signal \N__37890\ : std_logic;
signal \N__37887\ : std_logic;
signal \N__37884\ : std_logic;
signal \N__37879\ : std_logic;
signal \N__37876\ : std_logic;
signal \N__37869\ : std_logic;
signal \N__37866\ : std_logic;
signal \N__37863\ : std_logic;
signal \N__37860\ : std_logic;
signal \N__37857\ : std_logic;
signal \N__37856\ : std_logic;
signal \N__37853\ : std_logic;
signal \N__37850\ : std_logic;
signal \N__37847\ : std_logic;
signal \N__37846\ : std_logic;
signal \N__37843\ : std_logic;
signal \N__37840\ : std_logic;
signal \N__37837\ : std_logic;
signal \N__37832\ : std_logic;
signal \N__37829\ : std_logic;
signal \N__37826\ : std_logic;
signal \N__37821\ : std_logic;
signal \N__37818\ : std_logic;
signal \N__37817\ : std_logic;
signal \N__37814\ : std_logic;
signal \N__37811\ : std_logic;
signal \N__37808\ : std_logic;
signal \N__37805\ : std_logic;
signal \N__37804\ : std_logic;
signal \N__37801\ : std_logic;
signal \N__37798\ : std_logic;
signal \N__37795\ : std_logic;
signal \N__37792\ : std_logic;
signal \N__37785\ : std_logic;
signal \N__37782\ : std_logic;
signal \N__37779\ : std_logic;
signal \N__37776\ : std_logic;
signal \N__37773\ : std_logic;
signal \N__37770\ : std_logic;
signal \N__37767\ : std_logic;
signal \N__37766\ : std_logic;
signal \N__37763\ : std_logic;
signal \N__37762\ : std_logic;
signal \N__37759\ : std_logic;
signal \N__37756\ : std_logic;
signal \N__37753\ : std_logic;
signal \N__37750\ : std_logic;
signal \N__37743\ : std_logic;
signal \N__37740\ : std_logic;
signal \N__37737\ : std_logic;
signal \N__37734\ : std_logic;
signal \N__37731\ : std_logic;
signal \N__37728\ : std_logic;
signal \N__37725\ : std_logic;
signal \N__37722\ : std_logic;
signal \N__37719\ : std_logic;
signal \N__37718\ : std_logic;
signal \N__37715\ : std_logic;
signal \N__37714\ : std_logic;
signal \N__37711\ : std_logic;
signal \N__37708\ : std_logic;
signal \N__37705\ : std_logic;
signal \N__37702\ : std_logic;
signal \N__37695\ : std_logic;
signal \N__37692\ : std_logic;
signal \N__37689\ : std_logic;
signal \N__37686\ : std_logic;
signal \N__37685\ : std_logic;
signal \N__37682\ : std_logic;
signal \N__37679\ : std_logic;
signal \N__37674\ : std_logic;
signal \N__37673\ : std_logic;
signal \N__37670\ : std_logic;
signal \N__37667\ : std_logic;
signal \N__37662\ : std_logic;
signal \N__37659\ : std_logic;
signal \N__37658\ : std_logic;
signal \N__37655\ : std_logic;
signal \N__37654\ : std_logic;
signal \N__37651\ : std_logic;
signal \N__37648\ : std_logic;
signal \N__37645\ : std_logic;
signal \N__37642\ : std_logic;
signal \N__37639\ : std_logic;
signal \N__37636\ : std_logic;
signal \N__37633\ : std_logic;
signal \N__37626\ : std_logic;
signal \N__37623\ : std_logic;
signal \N__37620\ : std_logic;
signal \N__37617\ : std_logic;
signal \N__37614\ : std_logic;
signal \N__37611\ : std_logic;
signal \N__37608\ : std_logic;
signal \N__37607\ : std_logic;
signal \N__37606\ : std_logic;
signal \N__37605\ : std_logic;
signal \N__37604\ : std_logic;
signal \N__37603\ : std_logic;
signal \N__37602\ : std_logic;
signal \N__37599\ : std_logic;
signal \N__37598\ : std_logic;
signal \N__37597\ : std_logic;
signal \N__37596\ : std_logic;
signal \N__37595\ : std_logic;
signal \N__37592\ : std_logic;
signal \N__37589\ : std_logic;
signal \N__37588\ : std_logic;
signal \N__37581\ : std_logic;
signal \N__37580\ : std_logic;
signal \N__37579\ : std_logic;
signal \N__37576\ : std_logic;
signal \N__37575\ : std_logic;
signal \N__37570\ : std_logic;
signal \N__37567\ : std_logic;
signal \N__37566\ : std_logic;
signal \N__37565\ : std_logic;
signal \N__37564\ : std_logic;
signal \N__37561\ : std_logic;
signal \N__37560\ : std_logic;
signal \N__37557\ : std_logic;
signal \N__37556\ : std_logic;
signal \N__37555\ : std_logic;
signal \N__37552\ : std_logic;
signal \N__37547\ : std_logic;
signal \N__37544\ : std_logic;
signal \N__37539\ : std_logic;
signal \N__37534\ : std_logic;
signal \N__37531\ : std_logic;
signal \N__37528\ : std_logic;
signal \N__37525\ : std_logic;
signal \N__37522\ : std_logic;
signal \N__37521\ : std_logic;
signal \N__37518\ : std_logic;
signal \N__37517\ : std_logic;
signal \N__37514\ : std_logic;
signal \N__37513\ : std_logic;
signal \N__37506\ : std_logic;
signal \N__37503\ : std_logic;
signal \N__37500\ : std_logic;
signal \N__37493\ : std_logic;
signal \N__37486\ : std_logic;
signal \N__37479\ : std_logic;
signal \N__37474\ : std_logic;
signal \N__37471\ : std_logic;
signal \N__37468\ : std_logic;
signal \N__37449\ : std_logic;
signal \N__37448\ : std_logic;
signal \N__37445\ : std_logic;
signal \N__37442\ : std_logic;
signal \N__37437\ : std_logic;
signal \N__37436\ : std_logic;
signal \N__37433\ : std_logic;
signal \N__37430\ : std_logic;
signal \N__37427\ : std_logic;
signal \N__37422\ : std_logic;
signal \N__37419\ : std_logic;
signal \N__37418\ : std_logic;
signal \N__37417\ : std_logic;
signal \N__37414\ : std_logic;
signal \N__37411\ : std_logic;
signal \N__37408\ : std_logic;
signal \N__37405\ : std_logic;
signal \N__37402\ : std_logic;
signal \N__37395\ : std_logic;
signal \N__37392\ : std_logic;
signal \N__37389\ : std_logic;
signal \N__37386\ : std_logic;
signal \N__37383\ : std_logic;
signal \N__37382\ : std_logic;
signal \N__37381\ : std_logic;
signal \N__37378\ : std_logic;
signal \N__37375\ : std_logic;
signal \N__37372\ : std_logic;
signal \N__37367\ : std_logic;
signal \N__37364\ : std_logic;
signal \N__37359\ : std_logic;
signal \N__37356\ : std_logic;
signal \N__37353\ : std_logic;
signal \N__37350\ : std_logic;
signal \N__37349\ : std_logic;
signal \N__37346\ : std_logic;
signal \N__37343\ : std_logic;
signal \N__37340\ : std_logic;
signal \N__37339\ : std_logic;
signal \N__37336\ : std_logic;
signal \N__37333\ : std_logic;
signal \N__37330\ : std_logic;
signal \N__37323\ : std_logic;
signal \N__37322\ : std_logic;
signal \N__37321\ : std_logic;
signal \N__37320\ : std_logic;
signal \N__37319\ : std_logic;
signal \N__37318\ : std_logic;
signal \N__37317\ : std_logic;
signal \N__37314\ : std_logic;
signal \N__37313\ : std_logic;
signal \N__37312\ : std_logic;
signal \N__37311\ : std_logic;
signal \N__37308\ : std_logic;
signal \N__37307\ : std_logic;
signal \N__37306\ : std_logic;
signal \N__37305\ : std_logic;
signal \N__37304\ : std_logic;
signal \N__37303\ : std_logic;
signal \N__37300\ : std_logic;
signal \N__37299\ : std_logic;
signal \N__37298\ : std_logic;
signal \N__37295\ : std_logic;
signal \N__37294\ : std_logic;
signal \N__37293\ : std_logic;
signal \N__37288\ : std_logic;
signal \N__37285\ : std_logic;
signal \N__37280\ : std_logic;
signal \N__37277\ : std_logic;
signal \N__37276\ : std_logic;
signal \N__37269\ : std_logic;
signal \N__37264\ : std_logic;
signal \N__37263\ : std_logic;
signal \N__37262\ : std_logic;
signal \N__37259\ : std_logic;
signal \N__37256\ : std_logic;
signal \N__37255\ : std_logic;
signal \N__37252\ : std_logic;
signal \N__37241\ : std_logic;
signal \N__37232\ : std_logic;
signal \N__37231\ : std_logic;
signal \N__37228\ : std_logic;
signal \N__37227\ : std_logic;
signal \N__37224\ : std_logic;
signal \N__37221\ : std_logic;
signal \N__37218\ : std_logic;
signal \N__37215\ : std_logic;
signal \N__37208\ : std_logic;
signal \N__37201\ : std_logic;
signal \N__37194\ : std_logic;
signal \N__37189\ : std_logic;
signal \N__37186\ : std_logic;
signal \N__37173\ : std_logic;
signal \N__37170\ : std_logic;
signal \N__37167\ : std_logic;
signal \N__37166\ : std_logic;
signal \N__37163\ : std_logic;
signal \N__37160\ : std_logic;
signal \N__37159\ : std_logic;
signal \N__37154\ : std_logic;
signal \N__37151\ : std_logic;
signal \N__37146\ : std_logic;
signal \N__37143\ : std_logic;
signal \N__37140\ : std_logic;
signal \N__37137\ : std_logic;
signal \N__37134\ : std_logic;
signal \N__37131\ : std_logic;
signal \N__37128\ : std_logic;
signal \N__37125\ : std_logic;
signal \N__37122\ : std_logic;
signal \N__37119\ : std_logic;
signal \N__37116\ : std_logic;
signal \N__37113\ : std_logic;
signal \N__37110\ : std_logic;
signal \N__37107\ : std_logic;
signal \N__37104\ : std_logic;
signal \N__37103\ : std_logic;
signal \N__37102\ : std_logic;
signal \N__37099\ : std_logic;
signal \N__37096\ : std_logic;
signal \N__37093\ : std_logic;
signal \N__37090\ : std_logic;
signal \N__37087\ : std_logic;
signal \N__37084\ : std_logic;
signal \N__37081\ : std_logic;
signal \N__37076\ : std_logic;
signal \N__37073\ : std_logic;
signal \N__37070\ : std_logic;
signal \N__37065\ : std_logic;
signal \N__37062\ : std_logic;
signal \N__37059\ : std_logic;
signal \N__37056\ : std_logic;
signal \N__37053\ : std_logic;
signal \N__37050\ : std_logic;
signal \N__37047\ : std_logic;
signal \N__37044\ : std_logic;
signal \N__37041\ : std_logic;
signal \N__37038\ : std_logic;
signal \N__37035\ : std_logic;
signal \N__37032\ : std_logic;
signal \N__37029\ : std_logic;
signal \N__37026\ : std_logic;
signal \N__37023\ : std_logic;
signal \N__37020\ : std_logic;
signal \N__37017\ : std_logic;
signal \N__37014\ : std_logic;
signal \N__37011\ : std_logic;
signal \N__37008\ : std_logic;
signal \N__37007\ : std_logic;
signal \N__37004\ : std_logic;
signal \N__37001\ : std_logic;
signal \N__36998\ : std_logic;
signal \N__36993\ : std_logic;
signal \N__36990\ : std_logic;
signal \N__36987\ : std_logic;
signal \N__36984\ : std_logic;
signal \N__36981\ : std_logic;
signal \N__36978\ : std_logic;
signal \N__36977\ : std_logic;
signal \N__36974\ : std_logic;
signal \N__36971\ : std_logic;
signal \N__36966\ : std_logic;
signal \N__36963\ : std_logic;
signal \N__36960\ : std_logic;
signal \N__36959\ : std_logic;
signal \N__36956\ : std_logic;
signal \N__36953\ : std_logic;
signal \N__36948\ : std_logic;
signal \N__36947\ : std_logic;
signal \N__36944\ : std_logic;
signal \N__36941\ : std_logic;
signal \N__36936\ : std_logic;
signal \N__36933\ : std_logic;
signal \N__36930\ : std_logic;
signal \N__36927\ : std_logic;
signal \N__36924\ : std_logic;
signal \N__36921\ : std_logic;
signal \N__36918\ : std_logic;
signal \N__36915\ : std_logic;
signal \N__36912\ : std_logic;
signal \N__36911\ : std_logic;
signal \N__36908\ : std_logic;
signal \N__36905\ : std_logic;
signal \N__36904\ : std_logic;
signal \N__36901\ : std_logic;
signal \N__36898\ : std_logic;
signal \N__36895\ : std_logic;
signal \N__36892\ : std_logic;
signal \N__36889\ : std_logic;
signal \N__36886\ : std_logic;
signal \N__36883\ : std_logic;
signal \N__36878\ : std_logic;
signal \N__36873\ : std_logic;
signal \N__36872\ : std_logic;
signal \N__36871\ : std_logic;
signal \N__36868\ : std_logic;
signal \N__36865\ : std_logic;
signal \N__36862\ : std_logic;
signal \N__36857\ : std_logic;
signal \N__36854\ : std_logic;
signal \N__36849\ : std_logic;
signal \N__36846\ : std_logic;
signal \N__36845\ : std_logic;
signal \N__36842\ : std_logic;
signal \N__36841\ : std_logic;
signal \N__36838\ : std_logic;
signal \N__36835\ : std_logic;
signal \N__36832\ : std_logic;
signal \N__36829\ : std_logic;
signal \N__36822\ : std_logic;
signal \N__36819\ : std_logic;
signal \N__36816\ : std_logic;
signal \N__36813\ : std_logic;
signal \N__36810\ : std_logic;
signal \N__36807\ : std_logic;
signal \N__36804\ : std_logic;
signal \N__36803\ : std_logic;
signal \N__36802\ : std_logic;
signal \N__36799\ : std_logic;
signal \N__36796\ : std_logic;
signal \N__36793\ : std_logic;
signal \N__36790\ : std_logic;
signal \N__36787\ : std_logic;
signal \N__36784\ : std_logic;
signal \N__36777\ : std_logic;
signal \N__36774\ : std_logic;
signal \N__36771\ : std_logic;
signal \N__36768\ : std_logic;
signal \N__36767\ : std_logic;
signal \N__36764\ : std_logic;
signal \N__36761\ : std_logic;
signal \N__36756\ : std_logic;
signal \N__36753\ : std_logic;
signal \N__36750\ : std_logic;
signal \N__36747\ : std_logic;
signal \N__36746\ : std_logic;
signal \N__36743\ : std_logic;
signal \N__36740\ : std_logic;
signal \N__36735\ : std_logic;
signal \N__36732\ : std_logic;
signal \N__36729\ : std_logic;
signal \N__36726\ : std_logic;
signal \N__36723\ : std_logic;
signal \N__36720\ : std_logic;
signal \N__36717\ : std_logic;
signal \N__36714\ : std_logic;
signal \N__36713\ : std_logic;
signal \N__36710\ : std_logic;
signal \N__36707\ : std_logic;
signal \N__36702\ : std_logic;
signal \N__36699\ : std_logic;
signal \N__36696\ : std_logic;
signal \N__36693\ : std_logic;
signal \N__36690\ : std_logic;
signal \N__36689\ : std_logic;
signal \N__36688\ : std_logic;
signal \N__36685\ : std_logic;
signal \N__36682\ : std_logic;
signal \N__36679\ : std_logic;
signal \N__36672\ : std_logic;
signal \N__36671\ : std_logic;
signal \N__36668\ : std_logic;
signal \N__36665\ : std_logic;
signal \N__36664\ : std_logic;
signal \N__36661\ : std_logic;
signal \N__36658\ : std_logic;
signal \N__36655\ : std_logic;
signal \N__36648\ : std_logic;
signal \N__36645\ : std_logic;
signal \N__36642\ : std_logic;
signal \N__36639\ : std_logic;
signal \N__36638\ : std_logic;
signal \N__36635\ : std_logic;
signal \N__36632\ : std_logic;
signal \N__36631\ : std_logic;
signal \N__36628\ : std_logic;
signal \N__36625\ : std_logic;
signal \N__36622\ : std_logic;
signal \N__36615\ : std_logic;
signal \N__36612\ : std_logic;
signal \N__36609\ : std_logic;
signal \N__36606\ : std_logic;
signal \N__36603\ : std_logic;
signal \N__36600\ : std_logic;
signal \N__36597\ : std_logic;
signal \N__36594\ : std_logic;
signal \N__36593\ : std_logic;
signal \N__36590\ : std_logic;
signal \N__36587\ : std_logic;
signal \N__36584\ : std_logic;
signal \N__36581\ : std_logic;
signal \N__36580\ : std_logic;
signal \N__36577\ : std_logic;
signal \N__36574\ : std_logic;
signal \N__36571\ : std_logic;
signal \N__36564\ : std_logic;
signal \N__36563\ : std_logic;
signal \N__36562\ : std_logic;
signal \N__36561\ : std_logic;
signal \N__36560\ : std_logic;
signal \N__36559\ : std_logic;
signal \N__36558\ : std_logic;
signal \N__36557\ : std_logic;
signal \N__36554\ : std_logic;
signal \N__36553\ : std_logic;
signal \N__36552\ : std_logic;
signal \N__36549\ : std_logic;
signal \N__36548\ : std_logic;
signal \N__36545\ : std_logic;
signal \N__36542\ : std_logic;
signal \N__36539\ : std_logic;
signal \N__36538\ : std_logic;
signal \N__36535\ : std_logic;
signal \N__36534\ : std_logic;
signal \N__36533\ : std_logic;
signal \N__36532\ : std_logic;
signal \N__36529\ : std_logic;
signal \N__36526\ : std_logic;
signal \N__36525\ : std_logic;
signal \N__36524\ : std_logic;
signal \N__36519\ : std_logic;
signal \N__36512\ : std_logic;
signal \N__36509\ : std_logic;
signal \N__36506\ : std_logic;
signal \N__36501\ : std_logic;
signal \N__36496\ : std_logic;
signal \N__36491\ : std_logic;
signal \N__36482\ : std_logic;
signal \N__36475\ : std_logic;
signal \N__36472\ : std_logic;
signal \N__36459\ : std_logic;
signal \N__36456\ : std_logic;
signal \N__36455\ : std_logic;
signal \N__36454\ : std_logic;
signal \N__36451\ : std_logic;
signal \N__36448\ : std_logic;
signal \N__36445\ : std_logic;
signal \N__36442\ : std_logic;
signal \N__36439\ : std_logic;
signal \N__36436\ : std_logic;
signal \N__36433\ : std_logic;
signal \N__36430\ : std_logic;
signal \N__36423\ : std_logic;
signal \N__36422\ : std_logic;
signal \N__36419\ : std_logic;
signal \N__36416\ : std_logic;
signal \N__36415\ : std_logic;
signal \N__36412\ : std_logic;
signal \N__36409\ : std_logic;
signal \N__36406\ : std_logic;
signal \N__36401\ : std_logic;
signal \N__36396\ : std_logic;
signal \N__36393\ : std_logic;
signal \N__36390\ : std_logic;
signal \N__36387\ : std_logic;
signal \N__36384\ : std_logic;
signal \N__36381\ : std_logic;
signal \N__36378\ : std_logic;
signal \N__36375\ : std_logic;
signal \N__36372\ : std_logic;
signal \N__36369\ : std_logic;
signal \N__36366\ : std_logic;
signal \N__36363\ : std_logic;
signal \N__36360\ : std_logic;
signal \N__36359\ : std_logic;
signal \N__36356\ : std_logic;
signal \N__36353\ : std_logic;
signal \N__36350\ : std_logic;
signal \N__36347\ : std_logic;
signal \N__36342\ : std_logic;
signal \N__36339\ : std_logic;
signal \N__36336\ : std_logic;
signal \N__36333\ : std_logic;
signal \N__36330\ : std_logic;
signal \N__36329\ : std_logic;
signal \N__36326\ : std_logic;
signal \N__36323\ : std_logic;
signal \N__36318\ : std_logic;
signal \N__36317\ : std_logic;
signal \N__36314\ : std_logic;
signal \N__36311\ : std_logic;
signal \N__36308\ : std_logic;
signal \N__36307\ : std_logic;
signal \N__36302\ : std_logic;
signal \N__36299\ : std_logic;
signal \N__36294\ : std_logic;
signal \N__36291\ : std_logic;
signal \N__36288\ : std_logic;
signal \N__36285\ : std_logic;
signal \N__36282\ : std_logic;
signal \N__36281\ : std_logic;
signal \N__36278\ : std_logic;
signal \N__36275\ : std_logic;
signal \N__36274\ : std_logic;
signal \N__36271\ : std_logic;
signal \N__36268\ : std_logic;
signal \N__36265\ : std_logic;
signal \N__36258\ : std_logic;
signal \N__36255\ : std_logic;
signal \N__36252\ : std_logic;
signal \N__36249\ : std_logic;
signal \N__36246\ : std_logic;
signal \N__36245\ : std_logic;
signal \N__36242\ : std_logic;
signal \N__36239\ : std_logic;
signal \N__36238\ : std_logic;
signal \N__36235\ : std_logic;
signal \N__36232\ : std_logic;
signal \N__36229\ : std_logic;
signal \N__36222\ : std_logic;
signal \N__36219\ : std_logic;
signal \N__36216\ : std_logic;
signal \N__36213\ : std_logic;
signal \N__36212\ : std_logic;
signal \N__36209\ : std_logic;
signal \N__36206\ : std_logic;
signal \N__36203\ : std_logic;
signal \N__36202\ : std_logic;
signal \N__36199\ : std_logic;
signal \N__36196\ : std_logic;
signal \N__36193\ : std_logic;
signal \N__36186\ : std_logic;
signal \N__36183\ : std_logic;
signal \N__36180\ : std_logic;
signal \N__36177\ : std_logic;
signal \N__36174\ : std_logic;
signal \N__36171\ : std_logic;
signal \N__36170\ : std_logic;
signal \N__36167\ : std_logic;
signal \N__36164\ : std_logic;
signal \N__36161\ : std_logic;
signal \N__36158\ : std_logic;
signal \N__36155\ : std_logic;
signal \N__36152\ : std_logic;
signal \N__36147\ : std_logic;
signal \N__36144\ : std_logic;
signal \N__36141\ : std_logic;
signal \N__36138\ : std_logic;
signal \N__36135\ : std_logic;
signal \N__36132\ : std_logic;
signal \N__36131\ : std_logic;
signal \N__36128\ : std_logic;
signal \N__36127\ : std_logic;
signal \N__36124\ : std_logic;
signal \N__36121\ : std_logic;
signal \N__36118\ : std_logic;
signal \N__36115\ : std_logic;
signal \N__36112\ : std_logic;
signal \N__36109\ : std_logic;
signal \N__36106\ : std_logic;
signal \N__36099\ : std_logic;
signal \N__36096\ : std_logic;
signal \N__36093\ : std_logic;
signal \N__36090\ : std_logic;
signal \N__36087\ : std_logic;
signal \N__36084\ : std_logic;
signal \N__36081\ : std_logic;
signal \N__36078\ : std_logic;
signal \N__36075\ : std_logic;
signal \N__36072\ : std_logic;
signal \N__36071\ : std_logic;
signal \N__36068\ : std_logic;
signal \N__36065\ : std_logic;
signal \N__36060\ : std_logic;
signal \N__36059\ : std_logic;
signal \N__36058\ : std_logic;
signal \N__36057\ : std_logic;
signal \N__36054\ : std_logic;
signal \N__36049\ : std_logic;
signal \N__36046\ : std_logic;
signal \N__36045\ : std_logic;
signal \N__36042\ : std_logic;
signal \N__36039\ : std_logic;
signal \N__36036\ : std_logic;
signal \N__36033\ : std_logic;
signal \N__36030\ : std_logic;
signal \N__36027\ : std_logic;
signal \N__36024\ : std_logic;
signal \N__36015\ : std_logic;
signal \N__36012\ : std_logic;
signal \N__36009\ : std_logic;
signal \N__36006\ : std_logic;
signal \N__36003\ : std_logic;
signal \N__36002\ : std_logic;
signal \N__35999\ : std_logic;
signal \N__35996\ : std_logic;
signal \N__35995\ : std_logic;
signal \N__35992\ : std_logic;
signal \N__35989\ : std_logic;
signal \N__35986\ : std_logic;
signal \N__35979\ : std_logic;
signal \N__35976\ : std_logic;
signal \N__35973\ : std_logic;
signal \N__35970\ : std_logic;
signal \N__35969\ : std_logic;
signal \N__35968\ : std_logic;
signal \N__35965\ : std_logic;
signal \N__35962\ : std_logic;
signal \N__35957\ : std_logic;
signal \N__35954\ : std_logic;
signal \N__35949\ : std_logic;
signal \N__35946\ : std_logic;
signal \N__35943\ : std_logic;
signal \N__35940\ : std_logic;
signal \N__35937\ : std_logic;
signal \N__35936\ : std_logic;
signal \N__35933\ : std_logic;
signal \N__35930\ : std_logic;
signal \N__35925\ : std_logic;
signal \N__35922\ : std_logic;
signal \N__35919\ : std_logic;
signal \N__35916\ : std_logic;
signal \N__35913\ : std_logic;
signal \N__35912\ : std_logic;
signal \N__35909\ : std_logic;
signal \N__35906\ : std_logic;
signal \N__35905\ : std_logic;
signal \N__35902\ : std_logic;
signal \N__35899\ : std_logic;
signal \N__35896\ : std_logic;
signal \N__35889\ : std_logic;
signal \N__35886\ : std_logic;
signal \N__35883\ : std_logic;
signal \N__35880\ : std_logic;
signal \N__35877\ : std_logic;
signal \N__35874\ : std_logic;
signal \N__35871\ : std_logic;
signal \N__35868\ : std_logic;
signal \N__35865\ : std_logic;
signal \N__35862\ : std_logic;
signal \N__35861\ : std_logic;
signal \N__35858\ : std_logic;
signal \N__35855\ : std_logic;
signal \N__35850\ : std_logic;
signal \N__35847\ : std_logic;
signal \N__35844\ : std_logic;
signal \N__35843\ : std_logic;
signal \N__35840\ : std_logic;
signal \N__35837\ : std_logic;
signal \N__35836\ : std_logic;
signal \N__35831\ : std_logic;
signal \N__35828\ : std_logic;
signal \N__35823\ : std_logic;
signal \N__35820\ : std_logic;
signal \N__35817\ : std_logic;
signal \N__35814\ : std_logic;
signal \N__35811\ : std_logic;
signal \N__35808\ : std_logic;
signal \N__35805\ : std_logic;
signal \N__35804\ : std_logic;
signal \N__35803\ : std_logic;
signal \N__35800\ : std_logic;
signal \N__35797\ : std_logic;
signal \N__35794\ : std_logic;
signal \N__35791\ : std_logic;
signal \N__35788\ : std_logic;
signal \N__35785\ : std_logic;
signal \N__35778\ : std_logic;
signal \N__35775\ : std_logic;
signal \N__35772\ : std_logic;
signal \N__35771\ : std_logic;
signal \N__35768\ : std_logic;
signal \N__35765\ : std_logic;
signal \N__35764\ : std_logic;
signal \N__35761\ : std_logic;
signal \N__35758\ : std_logic;
signal \N__35755\ : std_logic;
signal \N__35752\ : std_logic;
signal \N__35745\ : std_logic;
signal \N__35742\ : std_logic;
signal \N__35739\ : std_logic;
signal \N__35736\ : std_logic;
signal \N__35733\ : std_logic;
signal \N__35730\ : std_logic;
signal \N__35727\ : std_logic;
signal \N__35724\ : std_logic;
signal \N__35721\ : std_logic;
signal \N__35718\ : std_logic;
signal \N__35715\ : std_logic;
signal \N__35712\ : std_logic;
signal \N__35709\ : std_logic;
signal \N__35706\ : std_logic;
signal \N__35703\ : std_logic;
signal \N__35700\ : std_logic;
signal \N__35697\ : std_logic;
signal \N__35694\ : std_logic;
signal \N__35691\ : std_logic;
signal \N__35688\ : std_logic;
signal \N__35685\ : std_logic;
signal \N__35682\ : std_logic;
signal \N__35679\ : std_logic;
signal \N__35676\ : std_logic;
signal \N__35673\ : std_logic;
signal \N__35670\ : std_logic;
signal \N__35667\ : std_logic;
signal \N__35664\ : std_logic;
signal \N__35661\ : std_logic;
signal \N__35658\ : std_logic;
signal \N__35657\ : std_logic;
signal \N__35654\ : std_logic;
signal \N__35651\ : std_logic;
signal \N__35648\ : std_logic;
signal \N__35643\ : std_logic;
signal \N__35640\ : std_logic;
signal \N__35637\ : std_logic;
signal \N__35634\ : std_logic;
signal \N__35631\ : std_logic;
signal \N__35628\ : std_logic;
signal \N__35625\ : std_logic;
signal \N__35622\ : std_logic;
signal \N__35619\ : std_logic;
signal \N__35616\ : std_logic;
signal \N__35613\ : std_logic;
signal \N__35612\ : std_logic;
signal \N__35611\ : std_logic;
signal \N__35608\ : std_logic;
signal \N__35605\ : std_logic;
signal \N__35602\ : std_logic;
signal \N__35599\ : std_logic;
signal \N__35596\ : std_logic;
signal \N__35589\ : std_logic;
signal \N__35586\ : std_logic;
signal \N__35583\ : std_logic;
signal \N__35580\ : std_logic;
signal \N__35577\ : std_logic;
signal \N__35574\ : std_logic;
signal \N__35571\ : std_logic;
signal \N__35570\ : std_logic;
signal \N__35567\ : std_logic;
signal \N__35564\ : std_logic;
signal \N__35561\ : std_logic;
signal \N__35560\ : std_logic;
signal \N__35555\ : std_logic;
signal \N__35552\ : std_logic;
signal \N__35547\ : std_logic;
signal \N__35544\ : std_logic;
signal \N__35541\ : std_logic;
signal \N__35538\ : std_logic;
signal \N__35535\ : std_logic;
signal \N__35532\ : std_logic;
signal \N__35529\ : std_logic;
signal \N__35528\ : std_logic;
signal \N__35525\ : std_logic;
signal \N__35522\ : std_logic;
signal \N__35517\ : std_logic;
signal \N__35516\ : std_logic;
signal \N__35515\ : std_logic;
signal \N__35512\ : std_logic;
signal \N__35509\ : std_logic;
signal \N__35506\ : std_logic;
signal \N__35503\ : std_logic;
signal \N__35500\ : std_logic;
signal \N__35497\ : std_logic;
signal \N__35494\ : std_logic;
signal \N__35491\ : std_logic;
signal \N__35486\ : std_logic;
signal \N__35481\ : std_logic;
signal \N__35478\ : std_logic;
signal \N__35475\ : std_logic;
signal \N__35472\ : std_logic;
signal \N__35469\ : std_logic;
signal \N__35466\ : std_logic;
signal \N__35463\ : std_logic;
signal \N__35462\ : std_logic;
signal \N__35459\ : std_logic;
signal \N__35456\ : std_logic;
signal \N__35453\ : std_logic;
signal \N__35450\ : std_logic;
signal \N__35449\ : std_logic;
signal \N__35446\ : std_logic;
signal \N__35443\ : std_logic;
signal \N__35440\ : std_logic;
signal \N__35437\ : std_logic;
signal \N__35430\ : std_logic;
signal \N__35427\ : std_logic;
signal \N__35424\ : std_logic;
signal \N__35421\ : std_logic;
signal \N__35418\ : std_logic;
signal \N__35415\ : std_logic;
signal \N__35412\ : std_logic;
signal \N__35411\ : std_logic;
signal \N__35408\ : std_logic;
signal \N__35405\ : std_logic;
signal \N__35402\ : std_logic;
signal \N__35401\ : std_logic;
signal \N__35398\ : std_logic;
signal \N__35395\ : std_logic;
signal \N__35392\ : std_logic;
signal \N__35389\ : std_logic;
signal \N__35382\ : std_logic;
signal \N__35379\ : std_logic;
signal \N__35376\ : std_logic;
signal \N__35373\ : std_logic;
signal \N__35370\ : std_logic;
signal \N__35369\ : std_logic;
signal \N__35366\ : std_logic;
signal \N__35363\ : std_logic;
signal \N__35360\ : std_logic;
signal \N__35357\ : std_logic;
signal \N__35356\ : std_logic;
signal \N__35353\ : std_logic;
signal \N__35350\ : std_logic;
signal \N__35347\ : std_logic;
signal \N__35344\ : std_logic;
signal \N__35341\ : std_logic;
signal \N__35334\ : std_logic;
signal \N__35331\ : std_logic;
signal \N__35328\ : std_logic;
signal \N__35325\ : std_logic;
signal \N__35322\ : std_logic;
signal \N__35319\ : std_logic;
signal \N__35316\ : std_logic;
signal \N__35313\ : std_logic;
signal \N__35310\ : std_logic;
signal \N__35307\ : std_logic;
signal \N__35304\ : std_logic;
signal \N__35301\ : std_logic;
signal \N__35298\ : std_logic;
signal \N__35295\ : std_logic;
signal \N__35292\ : std_logic;
signal \N__35289\ : std_logic;
signal \N__35286\ : std_logic;
signal \N__35283\ : std_logic;
signal \N__35282\ : std_logic;
signal \N__35279\ : std_logic;
signal \N__35276\ : std_logic;
signal \N__35271\ : std_logic;
signal \N__35268\ : std_logic;
signal \N__35265\ : std_logic;
signal \N__35262\ : std_logic;
signal \N__35259\ : std_logic;
signal \N__35258\ : std_logic;
signal \N__35257\ : std_logic;
signal \N__35254\ : std_logic;
signal \N__35251\ : std_logic;
signal \N__35248\ : std_logic;
signal \N__35245\ : std_logic;
signal \N__35242\ : std_logic;
signal \N__35239\ : std_logic;
signal \N__35234\ : std_logic;
signal \N__35233\ : std_logic;
signal \N__35232\ : std_logic;
signal \N__35229\ : std_logic;
signal \N__35226\ : std_logic;
signal \N__35223\ : std_logic;
signal \N__35220\ : std_logic;
signal \N__35217\ : std_logic;
signal \N__35214\ : std_logic;
signal \N__35205\ : std_logic;
signal \N__35202\ : std_logic;
signal \N__35199\ : std_logic;
signal \N__35196\ : std_logic;
signal \N__35193\ : std_logic;
signal \N__35190\ : std_logic;
signal \N__35187\ : std_logic;
signal \N__35186\ : std_logic;
signal \N__35185\ : std_logic;
signal \N__35182\ : std_logic;
signal \N__35179\ : std_logic;
signal \N__35176\ : std_logic;
signal \N__35173\ : std_logic;
signal \N__35166\ : std_logic;
signal \N__35163\ : std_logic;
signal \N__35160\ : std_logic;
signal \N__35157\ : std_logic;
signal \N__35154\ : std_logic;
signal \N__35151\ : std_logic;
signal \N__35150\ : std_logic;
signal \N__35147\ : std_logic;
signal \N__35146\ : std_logic;
signal \N__35143\ : std_logic;
signal \N__35140\ : std_logic;
signal \N__35137\ : std_logic;
signal \N__35134\ : std_logic;
signal \N__35131\ : std_logic;
signal \N__35128\ : std_logic;
signal \N__35121\ : std_logic;
signal \N__35118\ : std_logic;
signal \N__35115\ : std_logic;
signal \N__35112\ : std_logic;
signal \N__35109\ : std_logic;
signal \N__35106\ : std_logic;
signal \N__35105\ : std_logic;
signal \N__35100\ : std_logic;
signal \N__35099\ : std_logic;
signal \N__35096\ : std_logic;
signal \N__35093\ : std_logic;
signal \N__35090\ : std_logic;
signal \N__35087\ : std_logic;
signal \N__35082\ : std_logic;
signal \N__35079\ : std_logic;
signal \N__35076\ : std_logic;
signal \N__35073\ : std_logic;
signal \N__35070\ : std_logic;
signal \N__35069\ : std_logic;
signal \N__35066\ : std_logic;
signal \N__35065\ : std_logic;
signal \N__35062\ : std_logic;
signal \N__35059\ : std_logic;
signal \N__35056\ : std_logic;
signal \N__35051\ : std_logic;
signal \N__35048\ : std_logic;
signal \N__35045\ : std_logic;
signal \N__35040\ : std_logic;
signal \N__35037\ : std_logic;
signal \N__35034\ : std_logic;
signal \N__35031\ : std_logic;
signal \N__35028\ : std_logic;
signal \N__35027\ : std_logic;
signal \N__35026\ : std_logic;
signal \N__35021\ : std_logic;
signal \N__35018\ : std_logic;
signal \N__35013\ : std_logic;
signal \N__35010\ : std_logic;
signal \N__35007\ : std_logic;
signal \N__35004\ : std_logic;
signal \N__35001\ : std_logic;
signal \N__34998\ : std_logic;
signal \N__34995\ : std_logic;
signal \N__34992\ : std_logic;
signal \N__34989\ : std_logic;
signal \N__34986\ : std_logic;
signal \N__34983\ : std_logic;
signal \N__34980\ : std_logic;
signal \N__34977\ : std_logic;
signal \N__34974\ : std_logic;
signal \N__34973\ : std_logic;
signal \N__34970\ : std_logic;
signal \N__34967\ : std_logic;
signal \N__34962\ : std_logic;
signal \N__34959\ : std_logic;
signal \N__34958\ : std_logic;
signal \N__34955\ : std_logic;
signal \N__34952\ : std_logic;
signal \N__34947\ : std_logic;
signal \N__34944\ : std_logic;
signal \N__34943\ : std_logic;
signal \N__34940\ : std_logic;
signal \N__34937\ : std_logic;
signal \N__34936\ : std_logic;
signal \N__34931\ : std_logic;
signal \N__34928\ : std_logic;
signal \N__34923\ : std_logic;
signal \N__34920\ : std_logic;
signal \N__34917\ : std_logic;
signal \N__34914\ : std_logic;
signal \N__34911\ : std_logic;
signal \N__34908\ : std_logic;
signal \N__34907\ : std_logic;
signal \N__34904\ : std_logic;
signal \N__34901\ : std_logic;
signal \N__34896\ : std_logic;
signal \N__34895\ : std_logic;
signal \N__34892\ : std_logic;
signal \N__34889\ : std_logic;
signal \N__34884\ : std_logic;
signal \N__34883\ : std_logic;
signal \N__34882\ : std_logic;
signal \N__34879\ : std_logic;
signal \N__34876\ : std_logic;
signal \N__34873\ : std_logic;
signal \N__34870\ : std_logic;
signal \N__34867\ : std_logic;
signal \N__34864\ : std_logic;
signal \N__34859\ : std_logic;
signal \N__34856\ : std_logic;
signal \N__34851\ : std_logic;
signal \N__34848\ : std_logic;
signal \N__34845\ : std_logic;
signal \N__34842\ : std_logic;
signal \N__34839\ : std_logic;
signal \N__34836\ : std_logic;
signal \N__34833\ : std_logic;
signal \N__34830\ : std_logic;
signal \N__34827\ : std_logic;
signal \N__34824\ : std_logic;
signal \N__34821\ : std_logic;
signal \N__34818\ : std_logic;
signal \N__34817\ : std_logic;
signal \N__34814\ : std_logic;
signal \N__34811\ : std_logic;
signal \N__34808\ : std_logic;
signal \N__34805\ : std_logic;
signal \N__34804\ : std_logic;
signal \N__34801\ : std_logic;
signal \N__34798\ : std_logic;
signal \N__34795\ : std_logic;
signal \N__34790\ : std_logic;
signal \N__34785\ : std_logic;
signal \N__34782\ : std_logic;
signal \N__34779\ : std_logic;
signal \N__34776\ : std_logic;
signal \N__34773\ : std_logic;
signal \N__34770\ : std_logic;
signal \N__34767\ : std_logic;
signal \N__34764\ : std_logic;
signal \N__34761\ : std_logic;
signal \N__34760\ : std_logic;
signal \N__34757\ : std_logic;
signal \N__34754\ : std_logic;
signal \N__34749\ : std_logic;
signal \N__34746\ : std_logic;
signal \N__34743\ : std_logic;
signal \N__34740\ : std_logic;
signal \N__34737\ : std_logic;
signal \N__34734\ : std_logic;
signal \N__34731\ : std_logic;
signal \N__34730\ : std_logic;
signal \N__34727\ : std_logic;
signal \N__34724\ : std_logic;
signal \N__34721\ : std_logic;
signal \N__34718\ : std_logic;
signal \N__34717\ : std_logic;
signal \N__34714\ : std_logic;
signal \N__34711\ : std_logic;
signal \N__34708\ : std_logic;
signal \N__34701\ : std_logic;
signal \N__34698\ : std_logic;
signal \N__34695\ : std_logic;
signal \N__34692\ : std_logic;
signal \N__34689\ : std_logic;
signal \N__34686\ : std_logic;
signal \N__34683\ : std_logic;
signal \N__34680\ : std_logic;
signal \N__34679\ : std_logic;
signal \N__34678\ : std_logic;
signal \N__34675\ : std_logic;
signal \N__34672\ : std_logic;
signal \N__34667\ : std_logic;
signal \N__34664\ : std_logic;
signal \N__34661\ : std_logic;
signal \N__34656\ : std_logic;
signal \N__34653\ : std_logic;
signal \N__34650\ : std_logic;
signal \N__34647\ : std_logic;
signal \N__34644\ : std_logic;
signal \N__34643\ : std_logic;
signal \N__34642\ : std_logic;
signal \N__34639\ : std_logic;
signal \N__34636\ : std_logic;
signal \N__34633\ : std_logic;
signal \N__34630\ : std_logic;
signal \N__34627\ : std_logic;
signal \N__34620\ : std_logic;
signal \N__34617\ : std_logic;
signal \N__34614\ : std_logic;
signal \N__34611\ : std_logic;
signal \N__34608\ : std_logic;
signal \N__34605\ : std_logic;
signal \N__34602\ : std_logic;
signal \N__34601\ : std_logic;
signal \N__34600\ : std_logic;
signal \N__34597\ : std_logic;
signal \N__34592\ : std_logic;
signal \N__34587\ : std_logic;
signal \N__34584\ : std_logic;
signal \N__34581\ : std_logic;
signal \N__34578\ : std_logic;
signal \N__34575\ : std_logic;
signal \N__34572\ : std_logic;
signal \N__34571\ : std_logic;
signal \N__34570\ : std_logic;
signal \N__34567\ : std_logic;
signal \N__34564\ : std_logic;
signal \N__34561\ : std_logic;
signal \N__34558\ : std_logic;
signal \N__34555\ : std_logic;
signal \N__34548\ : std_logic;
signal \N__34545\ : std_logic;
signal \N__34542\ : std_logic;
signal \N__34539\ : std_logic;
signal \N__34536\ : std_logic;
signal \N__34535\ : std_logic;
signal \N__34532\ : std_logic;
signal \N__34529\ : std_logic;
signal \N__34528\ : std_logic;
signal \N__34525\ : std_logic;
signal \N__34522\ : std_logic;
signal \N__34519\ : std_logic;
signal \N__34516\ : std_logic;
signal \N__34509\ : std_logic;
signal \N__34506\ : std_logic;
signal \N__34503\ : std_logic;
signal \N__34500\ : std_logic;
signal \N__34499\ : std_logic;
signal \N__34498\ : std_logic;
signal \N__34495\ : std_logic;
signal \N__34492\ : std_logic;
signal \N__34489\ : std_logic;
signal \N__34486\ : std_logic;
signal \N__34479\ : std_logic;
signal \N__34476\ : std_logic;
signal \N__34473\ : std_logic;
signal \N__34470\ : std_logic;
signal \N__34469\ : std_logic;
signal \N__34466\ : std_logic;
signal \N__34463\ : std_logic;
signal \N__34460\ : std_logic;
signal \N__34455\ : std_logic;
signal \N__34452\ : std_logic;
signal \N__34449\ : std_logic;
signal \N__34446\ : std_logic;
signal \N__34443\ : std_logic;
signal \N__34442\ : std_logic;
signal \N__34439\ : std_logic;
signal \N__34436\ : std_logic;
signal \N__34433\ : std_logic;
signal \N__34428\ : std_logic;
signal \N__34425\ : std_logic;
signal \N__34422\ : std_logic;
signal \N__34419\ : std_logic;
signal \N__34416\ : std_logic;
signal \N__34413\ : std_logic;
signal \N__34412\ : std_logic;
signal \N__34409\ : std_logic;
signal \N__34406\ : std_logic;
signal \N__34405\ : std_logic;
signal \N__34402\ : std_logic;
signal \N__34399\ : std_logic;
signal \N__34396\ : std_logic;
signal \N__34389\ : std_logic;
signal \N__34386\ : std_logic;
signal \N__34383\ : std_logic;
signal \N__34380\ : std_logic;
signal \N__34377\ : std_logic;
signal \N__34374\ : std_logic;
signal \N__34371\ : std_logic;
signal \N__34368\ : std_logic;
signal \N__34365\ : std_logic;
signal \N__34362\ : std_logic;
signal \N__34359\ : std_logic;
signal \N__34356\ : std_logic;
signal \N__34353\ : std_logic;
signal \N__34350\ : std_logic;
signal \N__34347\ : std_logic;
signal \N__34344\ : std_logic;
signal \N__34341\ : std_logic;
signal \N__34340\ : std_logic;
signal \N__34337\ : std_logic;
signal \N__34334\ : std_logic;
signal \N__34333\ : std_logic;
signal \N__34330\ : std_logic;
signal \N__34329\ : std_logic;
signal \N__34328\ : std_logic;
signal \N__34325\ : std_logic;
signal \N__34322\ : std_logic;
signal \N__34319\ : std_logic;
signal \N__34316\ : std_logic;
signal \N__34313\ : std_logic;
signal \N__34310\ : std_logic;
signal \N__34303\ : std_logic;
signal \N__34296\ : std_logic;
signal \N__34293\ : std_logic;
signal \N__34290\ : std_logic;
signal \N__34287\ : std_logic;
signal \N__34284\ : std_logic;
signal \N__34281\ : std_logic;
signal \N__34280\ : std_logic;
signal \N__34277\ : std_logic;
signal \N__34274\ : std_logic;
signal \N__34271\ : std_logic;
signal \N__34266\ : std_logic;
signal \N__34263\ : std_logic;
signal \N__34260\ : std_logic;
signal \N__34257\ : std_logic;
signal \N__34254\ : std_logic;
signal \N__34251\ : std_logic;
signal \N__34250\ : std_logic;
signal \N__34249\ : std_logic;
signal \N__34246\ : std_logic;
signal \N__34243\ : std_logic;
signal \N__34240\ : std_logic;
signal \N__34237\ : std_logic;
signal \N__34230\ : std_logic;
signal \N__34227\ : std_logic;
signal \N__34224\ : std_logic;
signal \N__34221\ : std_logic;
signal \N__34218\ : std_logic;
signal \N__34215\ : std_logic;
signal \N__34212\ : std_logic;
signal \N__34209\ : std_logic;
signal \N__34208\ : std_logic;
signal \N__34205\ : std_logic;
signal \N__34202\ : std_logic;
signal \N__34201\ : std_logic;
signal \N__34198\ : std_logic;
signal \N__34195\ : std_logic;
signal \N__34192\ : std_logic;
signal \N__34187\ : std_logic;
signal \N__34184\ : std_logic;
signal \N__34181\ : std_logic;
signal \N__34176\ : std_logic;
signal \N__34173\ : std_logic;
signal \N__34172\ : std_logic;
signal \N__34169\ : std_logic;
signal \N__34168\ : std_logic;
signal \N__34165\ : std_logic;
signal \N__34162\ : std_logic;
signal \N__34159\ : std_logic;
signal \N__34156\ : std_logic;
signal \N__34149\ : std_logic;
signal \N__34146\ : std_logic;
signal \N__34143\ : std_logic;
signal \N__34140\ : std_logic;
signal \N__34137\ : std_logic;
signal \N__34134\ : std_logic;
signal \N__34131\ : std_logic;
signal \N__34128\ : std_logic;
signal \N__34127\ : std_logic;
signal \N__34126\ : std_logic;
signal \N__34123\ : std_logic;
signal \N__34120\ : std_logic;
signal \N__34117\ : std_logic;
signal \N__34112\ : std_logic;
signal \N__34109\ : std_logic;
signal \N__34106\ : std_logic;
signal \N__34103\ : std_logic;
signal \N__34098\ : std_logic;
signal \N__34095\ : std_logic;
signal \N__34092\ : std_logic;
signal \N__34089\ : std_logic;
signal \N__34086\ : std_logic;
signal \N__34083\ : std_logic;
signal \N__34080\ : std_logic;
signal \N__34079\ : std_logic;
signal \N__34078\ : std_logic;
signal \N__34075\ : std_logic;
signal \N__34072\ : std_logic;
signal \N__34069\ : std_logic;
signal \N__34066\ : std_logic;
signal \N__34063\ : std_logic;
signal \N__34060\ : std_logic;
signal \N__34055\ : std_logic;
signal \N__34052\ : std_logic;
signal \N__34047\ : std_logic;
signal \N__34044\ : std_logic;
signal \N__34041\ : std_logic;
signal \N__34038\ : std_logic;
signal \N__34035\ : std_logic;
signal \N__34032\ : std_logic;
signal \N__34029\ : std_logic;
signal \N__34028\ : std_logic;
signal \N__34027\ : std_logic;
signal \N__34026\ : std_logic;
signal \N__34025\ : std_logic;
signal \N__34024\ : std_logic;
signal \N__34017\ : std_logic;
signal \N__34014\ : std_logic;
signal \N__34011\ : std_logic;
signal \N__34008\ : std_logic;
signal \N__34007\ : std_logic;
signal \N__34006\ : std_logic;
signal \N__34005\ : std_logic;
signal \N__34004\ : std_logic;
signal \N__34003\ : std_logic;
signal \N__34002\ : std_logic;
signal \N__34001\ : std_logic;
signal \N__33998\ : std_logic;
signal \N__33995\ : std_logic;
signal \N__33990\ : std_logic;
signal \N__33989\ : std_logic;
signal \N__33988\ : std_logic;
signal \N__33987\ : std_logic;
signal \N__33986\ : std_logic;
signal \N__33985\ : std_logic;
signal \N__33984\ : std_logic;
signal \N__33981\ : std_logic;
signal \N__33978\ : std_logic;
signal \N__33977\ : std_logic;
signal \N__33974\ : std_logic;
signal \N__33973\ : std_logic;
signal \N__33972\ : std_logic;
signal \N__33969\ : std_logic;
signal \N__33968\ : std_logic;
signal \N__33967\ : std_logic;
signal \N__33966\ : std_logic;
signal \N__33963\ : std_logic;
signal \N__33962\ : std_logic;
signal \N__33959\ : std_logic;
signal \N__33956\ : std_logic;
signal \N__33955\ : std_logic;
signal \N__33948\ : std_logic;
signal \N__33943\ : std_logic;
signal \N__33930\ : std_logic;
signal \N__33915\ : std_logic;
signal \N__33902\ : std_logic;
signal \N__33891\ : std_logic;
signal \N__33888\ : std_logic;
signal \N__33887\ : std_logic;
signal \N__33884\ : std_logic;
signal \N__33881\ : std_logic;
signal \N__33878\ : std_logic;
signal \N__33875\ : std_logic;
signal \N__33872\ : std_logic;
signal \N__33869\ : std_logic;
signal \N__33864\ : std_logic;
signal \N__33861\ : std_logic;
signal \N__33858\ : std_logic;
signal \N__33855\ : std_logic;
signal \N__33852\ : std_logic;
signal \N__33849\ : std_logic;
signal \N__33846\ : std_logic;
signal \N__33845\ : std_logic;
signal \N__33844\ : std_logic;
signal \N__33841\ : std_logic;
signal \N__33838\ : std_logic;
signal \N__33835\ : std_logic;
signal \N__33832\ : std_logic;
signal \N__33829\ : std_logic;
signal \N__33826\ : std_logic;
signal \N__33819\ : std_logic;
signal \N__33816\ : std_logic;
signal \N__33813\ : std_logic;
signal \N__33810\ : std_logic;
signal \N__33807\ : std_logic;
signal \N__33804\ : std_logic;
signal \N__33803\ : std_logic;
signal \N__33800\ : std_logic;
signal \N__33797\ : std_logic;
signal \N__33796\ : std_logic;
signal \N__33793\ : std_logic;
signal \N__33790\ : std_logic;
signal \N__33787\ : std_logic;
signal \N__33784\ : std_logic;
signal \N__33779\ : std_logic;
signal \N__33776\ : std_logic;
signal \N__33771\ : std_logic;
signal \N__33768\ : std_logic;
signal \N__33765\ : std_logic;
signal \N__33762\ : std_logic;
signal \N__33759\ : std_logic;
signal \N__33756\ : std_logic;
signal \N__33753\ : std_logic;
signal \N__33752\ : std_logic;
signal \N__33749\ : std_logic;
signal \N__33746\ : std_logic;
signal \N__33745\ : std_logic;
signal \N__33740\ : std_logic;
signal \N__33737\ : std_logic;
signal \N__33732\ : std_logic;
signal \N__33731\ : std_logic;
signal \N__33728\ : std_logic;
signal \N__33725\ : std_logic;
signal \N__33720\ : std_logic;
signal \N__33719\ : std_logic;
signal \N__33716\ : std_logic;
signal \N__33713\ : std_logic;
signal \N__33708\ : std_logic;
signal \N__33705\ : std_logic;
signal \N__33702\ : std_logic;
signal \N__33699\ : std_logic;
signal \N__33696\ : std_logic;
signal \N__33693\ : std_logic;
signal \N__33692\ : std_logic;
signal \N__33689\ : std_logic;
signal \N__33686\ : std_logic;
signal \N__33685\ : std_logic;
signal \N__33682\ : std_logic;
signal \N__33679\ : std_logic;
signal \N__33676\ : std_logic;
signal \N__33673\ : std_logic;
signal \N__33668\ : std_logic;
signal \N__33663\ : std_logic;
signal \N__33660\ : std_logic;
signal \N__33657\ : std_logic;
signal \N__33654\ : std_logic;
signal \N__33651\ : std_logic;
signal \N__33648\ : std_logic;
signal \N__33647\ : std_logic;
signal \N__33644\ : std_logic;
signal \N__33641\ : std_logic;
signal \N__33640\ : std_logic;
signal \N__33637\ : std_logic;
signal \N__33634\ : std_logic;
signal \N__33631\ : std_logic;
signal \N__33626\ : std_logic;
signal \N__33623\ : std_logic;
signal \N__33618\ : std_logic;
signal \N__33615\ : std_logic;
signal \N__33612\ : std_logic;
signal \N__33609\ : std_logic;
signal \N__33606\ : std_logic;
signal \N__33603\ : std_logic;
signal \N__33602\ : std_logic;
signal \N__33599\ : std_logic;
signal \N__33596\ : std_logic;
signal \N__33595\ : std_logic;
signal \N__33592\ : std_logic;
signal \N__33589\ : std_logic;
signal \N__33586\ : std_logic;
signal \N__33581\ : std_logic;
signal \N__33578\ : std_logic;
signal \N__33573\ : std_logic;
signal \N__33570\ : std_logic;
signal \N__33567\ : std_logic;
signal \N__33564\ : std_logic;
signal \N__33561\ : std_logic;
signal \N__33558\ : std_logic;
signal \N__33555\ : std_logic;
signal \N__33554\ : std_logic;
signal \N__33553\ : std_logic;
signal \N__33550\ : std_logic;
signal \N__33547\ : std_logic;
signal \N__33544\ : std_logic;
signal \N__33541\ : std_logic;
signal \N__33536\ : std_logic;
signal \N__33531\ : std_logic;
signal \N__33528\ : std_logic;
signal \N__33525\ : std_logic;
signal \N__33522\ : std_logic;
signal \N__33519\ : std_logic;
signal \N__33516\ : std_logic;
signal \N__33515\ : std_logic;
signal \N__33512\ : std_logic;
signal \N__33509\ : std_logic;
signal \N__33508\ : std_logic;
signal \N__33505\ : std_logic;
signal \N__33502\ : std_logic;
signal \N__33499\ : std_logic;
signal \N__33496\ : std_logic;
signal \N__33493\ : std_logic;
signal \N__33490\ : std_logic;
signal \N__33483\ : std_logic;
signal \N__33480\ : std_logic;
signal \N__33477\ : std_logic;
signal \N__33474\ : std_logic;
signal \N__33471\ : std_logic;
signal \N__33468\ : std_logic;
signal \N__33467\ : std_logic;
signal \N__33466\ : std_logic;
signal \N__33463\ : std_logic;
signal \N__33460\ : std_logic;
signal \N__33457\ : std_logic;
signal \N__33454\ : std_logic;
signal \N__33451\ : std_logic;
signal \N__33448\ : std_logic;
signal \N__33445\ : std_logic;
signal \N__33442\ : std_logic;
signal \N__33439\ : std_logic;
signal \N__33432\ : std_logic;
signal \N__33429\ : std_logic;
signal \N__33426\ : std_logic;
signal \N__33423\ : std_logic;
signal \N__33420\ : std_logic;
signal \N__33417\ : std_logic;
signal \N__33414\ : std_logic;
signal \N__33413\ : std_logic;
signal \N__33412\ : std_logic;
signal \N__33409\ : std_logic;
signal \N__33406\ : std_logic;
signal \N__33403\ : std_logic;
signal \N__33400\ : std_logic;
signal \N__33397\ : std_logic;
signal \N__33394\ : std_logic;
signal \N__33387\ : std_logic;
signal \N__33384\ : std_logic;
signal \N__33381\ : std_logic;
signal \N__33378\ : std_logic;
signal \N__33375\ : std_logic;
signal \N__33372\ : std_logic;
signal \N__33369\ : std_logic;
signal \N__33366\ : std_logic;
signal \N__33365\ : std_logic;
signal \N__33362\ : std_logic;
signal \N__33361\ : std_logic;
signal \N__33358\ : std_logic;
signal \N__33355\ : std_logic;
signal \N__33352\ : std_logic;
signal \N__33345\ : std_logic;
signal \N__33342\ : std_logic;
signal \N__33339\ : std_logic;
signal \N__33336\ : std_logic;
signal \N__33333\ : std_logic;
signal \N__33330\ : std_logic;
signal \N__33329\ : std_logic;
signal \N__33328\ : std_logic;
signal \N__33325\ : std_logic;
signal \N__33322\ : std_logic;
signal \N__33319\ : std_logic;
signal \N__33316\ : std_logic;
signal \N__33311\ : std_logic;
signal \N__33306\ : std_logic;
signal \N__33303\ : std_logic;
signal \N__33300\ : std_logic;
signal \N__33297\ : std_logic;
signal \N__33294\ : std_logic;
signal \N__33293\ : std_logic;
signal \N__33290\ : std_logic;
signal \N__33287\ : std_logic;
signal \N__33286\ : std_logic;
signal \N__33283\ : std_logic;
signal \N__33280\ : std_logic;
signal \N__33277\ : std_logic;
signal \N__33274\ : std_logic;
signal \N__33271\ : std_logic;
signal \N__33264\ : std_logic;
signal \N__33261\ : std_logic;
signal \N__33258\ : std_logic;
signal \N__33255\ : std_logic;
signal \N__33252\ : std_logic;
signal \N__33249\ : std_logic;
signal \N__33248\ : std_logic;
signal \N__33245\ : std_logic;
signal \N__33242\ : std_logic;
signal \N__33239\ : std_logic;
signal \N__33238\ : std_logic;
signal \N__33235\ : std_logic;
signal \N__33232\ : std_logic;
signal \N__33229\ : std_logic;
signal \N__33222\ : std_logic;
signal \N__33219\ : std_logic;
signal \N__33216\ : std_logic;
signal \N__33213\ : std_logic;
signal \N__33210\ : std_logic;
signal \N__33209\ : std_logic;
signal \N__33206\ : std_logic;
signal \N__33205\ : std_logic;
signal \N__33202\ : std_logic;
signal \N__33199\ : std_logic;
signal \N__33196\ : std_logic;
signal \N__33193\ : std_logic;
signal \N__33190\ : std_logic;
signal \N__33187\ : std_logic;
signal \N__33180\ : std_logic;
signal \N__33177\ : std_logic;
signal \N__33174\ : std_logic;
signal \N__33171\ : std_logic;
signal \N__33168\ : std_logic;
signal \N__33165\ : std_logic;
signal \N__33164\ : std_logic;
signal \N__33163\ : std_logic;
signal \N__33160\ : std_logic;
signal \N__33157\ : std_logic;
signal \N__33154\ : std_logic;
signal \N__33151\ : std_logic;
signal \N__33148\ : std_logic;
signal \N__33141\ : std_logic;
signal \N__33138\ : std_logic;
signal \N__33135\ : std_logic;
signal \N__33132\ : std_logic;
signal \N__33131\ : std_logic;
signal \N__33128\ : std_logic;
signal \N__33125\ : std_logic;
signal \N__33124\ : std_logic;
signal \N__33121\ : std_logic;
signal \N__33118\ : std_logic;
signal \N__33115\ : std_logic;
signal \N__33110\ : std_logic;
signal \N__33105\ : std_logic;
signal \N__33102\ : std_logic;
signal \N__33099\ : std_logic;
signal \N__33096\ : std_logic;
signal \N__33093\ : std_logic;
signal \N__33092\ : std_logic;
signal \N__33089\ : std_logic;
signal \N__33086\ : std_logic;
signal \N__33085\ : std_logic;
signal \N__33082\ : std_logic;
signal \N__33079\ : std_logic;
signal \N__33076\ : std_logic;
signal \N__33073\ : std_logic;
signal \N__33070\ : std_logic;
signal \N__33067\ : std_logic;
signal \N__33064\ : std_logic;
signal \N__33061\ : std_logic;
signal \N__33054\ : std_logic;
signal \N__33051\ : std_logic;
signal \N__33050\ : std_logic;
signal \N__33047\ : std_logic;
signal \N__33044\ : std_logic;
signal \N__33043\ : std_logic;
signal \N__33040\ : std_logic;
signal \N__33035\ : std_logic;
signal \N__33032\ : std_logic;
signal \N__33027\ : std_logic;
signal \N__33024\ : std_logic;
signal \N__33021\ : std_logic;
signal \N__33018\ : std_logic;
signal \N__33015\ : std_logic;
signal \N__33012\ : std_logic;
signal \N__33009\ : std_logic;
signal \N__33006\ : std_logic;
signal \N__33005\ : std_logic;
signal \N__33004\ : std_logic;
signal \N__33001\ : std_logic;
signal \N__32998\ : std_logic;
signal \N__32995\ : std_logic;
signal \N__32992\ : std_logic;
signal \N__32985\ : std_logic;
signal \N__32982\ : std_logic;
signal \N__32979\ : std_logic;
signal \N__32976\ : std_logic;
signal \N__32975\ : std_logic;
signal \N__32972\ : std_logic;
signal \N__32969\ : std_logic;
signal \N__32966\ : std_logic;
signal \N__32963\ : std_logic;
signal \N__32962\ : std_logic;
signal \N__32959\ : std_logic;
signal \N__32956\ : std_logic;
signal \N__32953\ : std_logic;
signal \N__32948\ : std_logic;
signal \N__32943\ : std_logic;
signal \N__32940\ : std_logic;
signal \N__32937\ : std_logic;
signal \N__32934\ : std_logic;
signal \N__32931\ : std_logic;
signal \N__32928\ : std_logic;
signal \N__32925\ : std_logic;
signal \N__32924\ : std_logic;
signal \N__32923\ : std_logic;
signal \N__32920\ : std_logic;
signal \N__32917\ : std_logic;
signal \N__32914\ : std_logic;
signal \N__32911\ : std_logic;
signal \N__32904\ : std_logic;
signal \N__32901\ : std_logic;
signal \N__32898\ : std_logic;
signal \N__32895\ : std_logic;
signal \N__32892\ : std_logic;
signal \N__32891\ : std_logic;
signal \N__32888\ : std_logic;
signal \N__32885\ : std_logic;
signal \N__32884\ : std_logic;
signal \N__32881\ : std_logic;
signal \N__32878\ : std_logic;
signal \N__32875\ : std_logic;
signal \N__32872\ : std_logic;
signal \N__32869\ : std_logic;
signal \N__32866\ : std_logic;
signal \N__32861\ : std_logic;
signal \N__32856\ : std_logic;
signal \N__32853\ : std_logic;
signal \N__32850\ : std_logic;
signal \N__32847\ : std_logic;
signal \N__32844\ : std_logic;
signal \N__32843\ : std_logic;
signal \N__32840\ : std_logic;
signal \N__32837\ : std_logic;
signal \N__32834\ : std_logic;
signal \N__32833\ : std_logic;
signal \N__32830\ : std_logic;
signal \N__32827\ : std_logic;
signal \N__32824\ : std_logic;
signal \N__32821\ : std_logic;
signal \N__32818\ : std_logic;
signal \N__32811\ : std_logic;
signal \N__32808\ : std_logic;
signal \N__32805\ : std_logic;
signal \N__32802\ : std_logic;
signal \N__32799\ : std_logic;
signal \N__32798\ : std_logic;
signal \N__32795\ : std_logic;
signal \N__32794\ : std_logic;
signal \N__32791\ : std_logic;
signal \N__32788\ : std_logic;
signal \N__32785\ : std_logic;
signal \N__32778\ : std_logic;
signal \N__32775\ : std_logic;
signal \N__32772\ : std_logic;
signal \N__32769\ : std_logic;
signal \N__32768\ : std_logic;
signal \N__32767\ : std_logic;
signal \N__32764\ : std_logic;
signal \N__32761\ : std_logic;
signal \N__32758\ : std_logic;
signal \N__32755\ : std_logic;
signal \N__32752\ : std_logic;
signal \N__32749\ : std_logic;
signal \N__32746\ : std_logic;
signal \N__32743\ : std_logic;
signal \N__32740\ : std_logic;
signal \N__32737\ : std_logic;
signal \N__32732\ : std_logic;
signal \N__32727\ : std_logic;
signal \N__32724\ : std_logic;
signal \N__32721\ : std_logic;
signal \N__32718\ : std_logic;
signal \N__32715\ : std_logic;
signal \N__32712\ : std_logic;
signal \N__32709\ : std_logic;
signal \N__32708\ : std_logic;
signal \N__32707\ : std_logic;
signal \N__32704\ : std_logic;
signal \N__32701\ : std_logic;
signal \N__32698\ : std_logic;
signal \N__32695\ : std_logic;
signal \N__32692\ : std_logic;
signal \N__32689\ : std_logic;
signal \N__32684\ : std_logic;
signal \N__32681\ : std_logic;
signal \N__32678\ : std_logic;
signal \N__32673\ : std_logic;
signal \N__32670\ : std_logic;
signal \N__32669\ : std_logic;
signal \N__32666\ : std_logic;
signal \N__32665\ : std_logic;
signal \N__32662\ : std_logic;
signal \N__32659\ : std_logic;
signal \N__32656\ : std_logic;
signal \N__32649\ : std_logic;
signal \N__32646\ : std_logic;
signal \N__32643\ : std_logic;
signal \N__32642\ : std_logic;
signal \N__32639\ : std_logic;
signal \N__32638\ : std_logic;
signal \N__32635\ : std_logic;
signal \N__32632\ : std_logic;
signal \N__32629\ : std_logic;
signal \N__32622\ : std_logic;
signal \N__32619\ : std_logic;
signal \N__32616\ : std_logic;
signal \N__32613\ : std_logic;
signal \N__32610\ : std_logic;
signal \N__32609\ : std_logic;
signal \N__32606\ : std_logic;
signal \N__32603\ : std_logic;
signal \N__32600\ : std_logic;
signal \N__32597\ : std_logic;
signal \N__32596\ : std_logic;
signal \N__32593\ : std_logic;
signal \N__32590\ : std_logic;
signal \N__32587\ : std_logic;
signal \N__32580\ : std_logic;
signal \N__32579\ : std_logic;
signal \N__32578\ : std_logic;
signal \N__32577\ : std_logic;
signal \N__32576\ : std_logic;
signal \N__32573\ : std_logic;
signal \N__32572\ : std_logic;
signal \N__32571\ : std_logic;
signal \N__32570\ : std_logic;
signal \N__32569\ : std_logic;
signal \N__32566\ : std_logic;
signal \N__32563\ : std_logic;
signal \N__32562\ : std_logic;
signal \N__32561\ : std_logic;
signal \N__32560\ : std_logic;
signal \N__32559\ : std_logic;
signal \N__32558\ : std_logic;
signal \N__32555\ : std_logic;
signal \N__32554\ : std_logic;
signal \N__32553\ : std_logic;
signal \N__32552\ : std_logic;
signal \N__32549\ : std_logic;
signal \N__32542\ : std_logic;
signal \N__32539\ : std_logic;
signal \N__32538\ : std_logic;
signal \N__32535\ : std_logic;
signal \N__32532\ : std_logic;
signal \N__32525\ : std_logic;
signal \N__32518\ : std_logic;
signal \N__32511\ : std_logic;
signal \N__32506\ : std_logic;
signal \N__32503\ : std_logic;
signal \N__32496\ : std_logic;
signal \N__32493\ : std_logic;
signal \N__32490\ : std_logic;
signal \N__32475\ : std_logic;
signal \N__32472\ : std_logic;
signal \N__32469\ : std_logic;
signal \N__32466\ : std_logic;
signal \N__32463\ : std_logic;
signal \N__32462\ : std_logic;
signal \N__32459\ : std_logic;
signal \N__32456\ : std_logic;
signal \N__32451\ : std_logic;
signal \N__32448\ : std_logic;
signal \N__32445\ : std_logic;
signal \N__32442\ : std_logic;
signal \N__32439\ : std_logic;
signal \N__32436\ : std_logic;
signal \N__32435\ : std_logic;
signal \N__32432\ : std_logic;
signal \N__32429\ : std_logic;
signal \N__32424\ : std_logic;
signal \N__32421\ : std_logic;
signal \N__32418\ : std_logic;
signal \N__32415\ : std_logic;
signal \N__32412\ : std_logic;
signal \N__32411\ : std_logic;
signal \N__32408\ : std_logic;
signal \N__32405\ : std_logic;
signal \N__32400\ : std_logic;
signal \N__32399\ : std_logic;
signal \N__32396\ : std_logic;
signal \N__32393\ : std_logic;
signal \N__32392\ : std_logic;
signal \N__32391\ : std_logic;
signal \N__32386\ : std_logic;
signal \N__32383\ : std_logic;
signal \N__32380\ : std_logic;
signal \N__32377\ : std_logic;
signal \N__32370\ : std_logic;
signal \N__32367\ : std_logic;
signal \N__32364\ : std_logic;
signal \N__32361\ : std_logic;
signal \N__32358\ : std_logic;
signal \N__32355\ : std_logic;
signal \N__32354\ : std_logic;
signal \N__32353\ : std_logic;
signal \N__32350\ : std_logic;
signal \N__32347\ : std_logic;
signal \N__32344\ : std_logic;
signal \N__32341\ : std_logic;
signal \N__32338\ : std_logic;
signal \N__32335\ : std_logic;
signal \N__32332\ : std_logic;
signal \N__32325\ : std_logic;
signal \N__32322\ : std_logic;
signal \N__32319\ : std_logic;
signal \N__32316\ : std_logic;
signal \N__32313\ : std_logic;
signal \N__32310\ : std_logic;
signal \N__32307\ : std_logic;
signal \N__32304\ : std_logic;
signal \N__32301\ : std_logic;
signal \N__32298\ : std_logic;
signal \N__32297\ : std_logic;
signal \N__32294\ : std_logic;
signal \N__32291\ : std_logic;
signal \N__32290\ : std_logic;
signal \N__32287\ : std_logic;
signal \N__32284\ : std_logic;
signal \N__32281\ : std_logic;
signal \N__32274\ : std_logic;
signal \N__32271\ : std_logic;
signal \N__32270\ : std_logic;
signal \N__32267\ : std_logic;
signal \N__32264\ : std_logic;
signal \N__32259\ : std_logic;
signal \N__32256\ : std_logic;
signal \N__32253\ : std_logic;
signal \N__32250\ : std_logic;
signal \N__32247\ : std_logic;
signal \N__32244\ : std_logic;
signal \N__32241\ : std_logic;
signal \N__32238\ : std_logic;
signal \N__32235\ : std_logic;
signal \N__32232\ : std_logic;
signal \N__32229\ : std_logic;
signal \N__32226\ : std_logic;
signal \N__32223\ : std_logic;
signal \N__32222\ : std_logic;
signal \N__32221\ : std_logic;
signal \N__32220\ : std_logic;
signal \N__32215\ : std_logic;
signal \N__32212\ : std_logic;
signal \N__32209\ : std_logic;
signal \N__32204\ : std_logic;
signal \N__32203\ : std_logic;
signal \N__32200\ : std_logic;
signal \N__32197\ : std_logic;
signal \N__32194\ : std_logic;
signal \N__32191\ : std_logic;
signal \N__32188\ : std_logic;
signal \N__32181\ : std_logic;
signal \N__32178\ : std_logic;
signal \N__32175\ : std_logic;
signal \N__32172\ : std_logic;
signal \N__32169\ : std_logic;
signal \N__32166\ : std_logic;
signal \N__32163\ : std_logic;
signal \N__32162\ : std_logic;
signal \N__32159\ : std_logic;
signal \N__32156\ : std_logic;
signal \N__32153\ : std_logic;
signal \N__32150\ : std_logic;
signal \N__32147\ : std_logic;
signal \N__32142\ : std_logic;
signal \N__32139\ : std_logic;
signal \N__32136\ : std_logic;
signal \N__32133\ : std_logic;
signal \N__32132\ : std_logic;
signal \N__32129\ : std_logic;
signal \N__32128\ : std_logic;
signal \N__32125\ : std_logic;
signal \N__32122\ : std_logic;
signal \N__32119\ : std_logic;
signal \N__32112\ : std_logic;
signal \N__32109\ : std_logic;
signal \N__32106\ : std_logic;
signal \N__32105\ : std_logic;
signal \N__32102\ : std_logic;
signal \N__32099\ : std_logic;
signal \N__32096\ : std_logic;
signal \N__32093\ : std_logic;
signal \N__32092\ : std_logic;
signal \N__32089\ : std_logic;
signal \N__32086\ : std_logic;
signal \N__32083\ : std_logic;
signal \N__32080\ : std_logic;
signal \N__32073\ : std_logic;
signal \N__32072\ : std_logic;
signal \N__32069\ : std_logic;
signal \N__32066\ : std_logic;
signal \N__32063\ : std_logic;
signal \N__32062\ : std_logic;
signal \N__32059\ : std_logic;
signal \N__32056\ : std_logic;
signal \N__32053\ : std_logic;
signal \N__32050\ : std_logic;
signal \N__32043\ : std_logic;
signal \N__32040\ : std_logic;
signal \N__32037\ : std_logic;
signal \N__32034\ : std_logic;
signal \N__32031\ : std_logic;
signal \N__32028\ : std_logic;
signal \N__32025\ : std_logic;
signal \N__32024\ : std_logic;
signal \N__32021\ : std_logic;
signal \N__32018\ : std_logic;
signal \N__32015\ : std_logic;
signal \N__32012\ : std_logic;
signal \N__32011\ : std_logic;
signal \N__32008\ : std_logic;
signal \N__32005\ : std_logic;
signal \N__32002\ : std_logic;
signal \N__31999\ : std_logic;
signal \N__31992\ : std_logic;
signal \N__31989\ : std_logic;
signal \N__31986\ : std_logic;
signal \N__31983\ : std_logic;
signal \N__31980\ : std_logic;
signal \N__31979\ : std_logic;
signal \N__31976\ : std_logic;
signal \N__31973\ : std_logic;
signal \N__31970\ : std_logic;
signal \N__31967\ : std_logic;
signal \N__31962\ : std_logic;
signal \N__31959\ : std_logic;
signal \N__31956\ : std_logic;
signal \N__31955\ : std_logic;
signal \N__31952\ : std_logic;
signal \N__31951\ : std_logic;
signal \N__31948\ : std_logic;
signal \N__31945\ : std_logic;
signal \N__31942\ : std_logic;
signal \N__31939\ : std_logic;
signal \N__31936\ : std_logic;
signal \N__31933\ : std_logic;
signal \N__31930\ : std_logic;
signal \N__31923\ : std_logic;
signal \N__31920\ : std_logic;
signal \N__31917\ : std_logic;
signal \N__31914\ : std_logic;
signal \N__31911\ : std_logic;
signal \N__31908\ : std_logic;
signal \N__31905\ : std_logic;
signal \N__31904\ : std_logic;
signal \N__31901\ : std_logic;
signal \N__31898\ : std_logic;
signal \N__31895\ : std_logic;
signal \N__31892\ : std_logic;
signal \N__31887\ : std_logic;
signal \N__31884\ : std_logic;
signal \N__31883\ : std_logic;
signal \N__31880\ : std_logic;
signal \N__31877\ : std_logic;
signal \N__31874\ : std_logic;
signal \N__31873\ : std_logic;
signal \N__31870\ : std_logic;
signal \N__31867\ : std_logic;
signal \N__31864\ : std_logic;
signal \N__31861\ : std_logic;
signal \N__31854\ : std_logic;
signal \N__31851\ : std_logic;
signal \N__31848\ : std_logic;
signal \N__31845\ : std_logic;
signal \N__31842\ : std_logic;
signal \N__31839\ : std_logic;
signal \N__31836\ : std_logic;
signal \N__31833\ : std_logic;
signal \N__31830\ : std_logic;
signal \N__31827\ : std_logic;
signal \N__31824\ : std_logic;
signal \N__31821\ : std_logic;
signal \N__31818\ : std_logic;
signal \N__31815\ : std_logic;
signal \N__31814\ : std_logic;
signal \N__31813\ : std_logic;
signal \N__31810\ : std_logic;
signal \N__31807\ : std_logic;
signal \N__31804\ : std_logic;
signal \N__31801\ : std_logic;
signal \N__31794\ : std_logic;
signal \N__31791\ : std_logic;
signal \N__31790\ : std_logic;
signal \N__31789\ : std_logic;
signal \N__31786\ : std_logic;
signal \N__31783\ : std_logic;
signal \N__31780\ : std_logic;
signal \N__31779\ : std_logic;
signal \N__31778\ : std_logic;
signal \N__31775\ : std_logic;
signal \N__31772\ : std_logic;
signal \N__31769\ : std_logic;
signal \N__31766\ : std_logic;
signal \N__31763\ : std_logic;
signal \N__31760\ : std_logic;
signal \N__31755\ : std_logic;
signal \N__31746\ : std_logic;
signal \N__31743\ : std_logic;
signal \N__31740\ : std_logic;
signal \N__31737\ : std_logic;
signal \N__31734\ : std_logic;
signal \N__31731\ : std_logic;
signal \N__31728\ : std_logic;
signal \N__31725\ : std_logic;
signal \N__31724\ : std_logic;
signal \N__31723\ : std_logic;
signal \N__31720\ : std_logic;
signal \N__31717\ : std_logic;
signal \N__31714\ : std_logic;
signal \N__31709\ : std_logic;
signal \N__31704\ : std_logic;
signal \N__31703\ : std_logic;
signal \N__31700\ : std_logic;
signal \N__31697\ : std_logic;
signal \N__31696\ : std_logic;
signal \N__31693\ : std_logic;
signal \N__31690\ : std_logic;
signal \N__31687\ : std_logic;
signal \N__31682\ : std_logic;
signal \N__31677\ : std_logic;
signal \N__31674\ : std_logic;
signal \N__31671\ : std_logic;
signal \N__31668\ : std_logic;
signal \N__31667\ : std_logic;
signal \N__31664\ : std_logic;
signal \N__31661\ : std_logic;
signal \N__31658\ : std_logic;
signal \N__31657\ : std_logic;
signal \N__31654\ : std_logic;
signal \N__31651\ : std_logic;
signal \N__31648\ : std_logic;
signal \N__31641\ : std_logic;
signal \N__31638\ : std_logic;
signal \N__31637\ : std_logic;
signal \N__31634\ : std_logic;
signal \N__31631\ : std_logic;
signal \N__31628\ : std_logic;
signal \N__31625\ : std_logic;
signal \N__31622\ : std_logic;
signal \N__31619\ : std_logic;
signal \N__31616\ : std_logic;
signal \N__31611\ : std_logic;
signal \N__31608\ : std_logic;
signal \N__31607\ : std_logic;
signal \N__31604\ : std_logic;
signal \N__31601\ : std_logic;
signal \N__31598\ : std_logic;
signal \N__31595\ : std_logic;
signal \N__31594\ : std_logic;
signal \N__31591\ : std_logic;
signal \N__31588\ : std_logic;
signal \N__31585\ : std_logic;
signal \N__31578\ : std_logic;
signal \N__31575\ : std_logic;
signal \N__31574\ : std_logic;
signal \N__31571\ : std_logic;
signal \N__31568\ : std_logic;
signal \N__31565\ : std_logic;
signal \N__31562\ : std_logic;
signal \N__31559\ : std_logic;
signal \N__31558\ : std_logic;
signal \N__31555\ : std_logic;
signal \N__31552\ : std_logic;
signal \N__31549\ : std_logic;
signal \N__31542\ : std_logic;
signal \N__31539\ : std_logic;
signal \N__31536\ : std_logic;
signal \N__31533\ : std_logic;
signal \N__31530\ : std_logic;
signal \N__31529\ : std_logic;
signal \N__31528\ : std_logic;
signal \N__31525\ : std_logic;
signal \N__31522\ : std_logic;
signal \N__31519\ : std_logic;
signal \N__31516\ : std_logic;
signal \N__31509\ : std_logic;
signal \N__31506\ : std_logic;
signal \N__31505\ : std_logic;
signal \N__31502\ : std_logic;
signal \N__31499\ : std_logic;
signal \N__31496\ : std_logic;
signal \N__31495\ : std_logic;
signal \N__31492\ : std_logic;
signal \N__31489\ : std_logic;
signal \N__31486\ : std_logic;
signal \N__31479\ : std_logic;
signal \N__31478\ : std_logic;
signal \N__31475\ : std_logic;
signal \N__31472\ : std_logic;
signal \N__31469\ : std_logic;
signal \N__31466\ : std_logic;
signal \N__31463\ : std_logic;
signal \N__31460\ : std_logic;
signal \N__31459\ : std_logic;
signal \N__31456\ : std_logic;
signal \N__31453\ : std_logic;
signal \N__31450\ : std_logic;
signal \N__31443\ : std_logic;
signal \N__31440\ : std_logic;
signal \N__31439\ : std_logic;
signal \N__31436\ : std_logic;
signal \N__31433\ : std_logic;
signal \N__31432\ : std_logic;
signal \N__31429\ : std_logic;
signal \N__31426\ : std_logic;
signal \N__31423\ : std_logic;
signal \N__31420\ : std_logic;
signal \N__31413\ : std_logic;
signal \N__31410\ : std_logic;
signal \N__31407\ : std_logic;
signal \N__31404\ : std_logic;
signal \N__31401\ : std_logic;
signal \N__31398\ : std_logic;
signal \N__31397\ : std_logic;
signal \N__31394\ : std_logic;
signal \N__31391\ : std_logic;
signal \N__31386\ : std_logic;
signal \N__31383\ : std_logic;
signal \N__31380\ : std_logic;
signal \N__31377\ : std_logic;
signal \N__31374\ : std_logic;
signal \N__31371\ : std_logic;
signal \N__31370\ : std_logic;
signal \N__31369\ : std_logic;
signal \N__31366\ : std_logic;
signal \N__31363\ : std_logic;
signal \N__31360\ : std_logic;
signal \N__31353\ : std_logic;
signal \N__31350\ : std_logic;
signal \N__31347\ : std_logic;
signal \N__31344\ : std_logic;
signal \N__31341\ : std_logic;
signal \N__31338\ : std_logic;
signal \N__31335\ : std_logic;
signal \N__31332\ : std_logic;
signal \N__31331\ : std_logic;
signal \N__31328\ : std_logic;
signal \N__31325\ : std_logic;
signal \N__31320\ : std_logic;
signal \N__31317\ : std_logic;
signal \N__31314\ : std_logic;
signal \N__31311\ : std_logic;
signal \N__31308\ : std_logic;
signal \N__31305\ : std_logic;
signal \N__31302\ : std_logic;
signal \N__31301\ : std_logic;
signal \N__31298\ : std_logic;
signal \N__31295\ : std_logic;
signal \N__31294\ : std_logic;
signal \N__31291\ : std_logic;
signal \N__31288\ : std_logic;
signal \N__31285\ : std_logic;
signal \N__31278\ : std_logic;
signal \N__31277\ : std_logic;
signal \N__31276\ : std_logic;
signal \N__31275\ : std_logic;
signal \N__31274\ : std_logic;
signal \N__31271\ : std_logic;
signal \N__31270\ : std_logic;
signal \N__31269\ : std_logic;
signal \N__31268\ : std_logic;
signal \N__31265\ : std_logic;
signal \N__31262\ : std_logic;
signal \N__31261\ : std_logic;
signal \N__31260\ : std_logic;
signal \N__31259\ : std_logic;
signal \N__31256\ : std_logic;
signal \N__31255\ : std_logic;
signal \N__31254\ : std_logic;
signal \N__31253\ : std_logic;
signal \N__31252\ : std_logic;
signal \N__31249\ : std_logic;
signal \N__31244\ : std_logic;
signal \N__31231\ : std_logic;
signal \N__31230\ : std_logic;
signal \N__31227\ : std_logic;
signal \N__31226\ : std_logic;
signal \N__31223\ : std_logic;
signal \N__31222\ : std_logic;
signal \N__31221\ : std_logic;
signal \N__31220\ : std_logic;
signal \N__31217\ : std_logic;
signal \N__31216\ : std_logic;
signal \N__31213\ : std_logic;
signal \N__31212\ : std_logic;
signal \N__31209\ : std_logic;
signal \N__31206\ : std_logic;
signal \N__31205\ : std_logic;
signal \N__31202\ : std_logic;
signal \N__31199\ : std_logic;
signal \N__31196\ : std_logic;
signal \N__31189\ : std_logic;
signal \N__31186\ : std_logic;
signal \N__31181\ : std_logic;
signal \N__31172\ : std_logic;
signal \N__31163\ : std_logic;
signal \N__31154\ : std_logic;
signal \N__31143\ : std_logic;
signal \N__31140\ : std_logic;
signal \N__31139\ : std_logic;
signal \N__31138\ : std_logic;
signal \N__31135\ : std_logic;
signal \N__31132\ : std_logic;
signal \N__31129\ : std_logic;
signal \N__31126\ : std_logic;
signal \N__31123\ : std_logic;
signal \N__31118\ : std_logic;
signal \N__31113\ : std_logic;
signal \N__31112\ : std_logic;
signal \N__31111\ : std_logic;
signal \N__31108\ : std_logic;
signal \N__31105\ : std_logic;
signal \N__31102\ : std_logic;
signal \N__31099\ : std_logic;
signal \N__31092\ : std_logic;
signal \N__31091\ : std_logic;
signal \N__31088\ : std_logic;
signal \N__31085\ : std_logic;
signal \N__31080\ : std_logic;
signal \N__31077\ : std_logic;
signal \N__31074\ : std_logic;
signal \N__31071\ : std_logic;
signal \N__31068\ : std_logic;
signal \N__31067\ : std_logic;
signal \N__31066\ : std_logic;
signal \N__31063\ : std_logic;
signal \N__31060\ : std_logic;
signal \N__31057\ : std_logic;
signal \N__31050\ : std_logic;
signal \N__31049\ : std_logic;
signal \N__31048\ : std_logic;
signal \N__31045\ : std_logic;
signal \N__31042\ : std_logic;
signal \N__31039\ : std_logic;
signal \N__31032\ : std_logic;
signal \N__31029\ : std_logic;
signal \N__31026\ : std_logic;
signal \N__31023\ : std_logic;
signal \N__31020\ : std_logic;
signal \N__31017\ : std_logic;
signal \N__31014\ : std_logic;
signal \N__31013\ : std_logic;
signal \N__31012\ : std_logic;
signal \N__31009\ : std_logic;
signal \N__31006\ : std_logic;
signal \N__31003\ : std_logic;
signal \N__31000\ : std_logic;
signal \N__30993\ : std_logic;
signal \N__30990\ : std_logic;
signal \N__30987\ : std_logic;
signal \N__30984\ : std_logic;
signal \N__30981\ : std_logic;
signal \N__30978\ : std_logic;
signal \N__30975\ : std_logic;
signal \N__30972\ : std_logic;
signal \N__30969\ : std_logic;
signal \N__30966\ : std_logic;
signal \N__30963\ : std_logic;
signal \N__30960\ : std_logic;
signal \N__30957\ : std_logic;
signal \N__30954\ : std_logic;
signal \N__30951\ : std_logic;
signal \N__30948\ : std_logic;
signal \N__30945\ : std_logic;
signal \N__30942\ : std_logic;
signal \N__30939\ : std_logic;
signal \N__30936\ : std_logic;
signal \N__30933\ : std_logic;
signal \N__30930\ : std_logic;
signal \N__30927\ : std_logic;
signal \N__30924\ : std_logic;
signal \N__30921\ : std_logic;
signal \N__30920\ : std_logic;
signal \N__30919\ : std_logic;
signal \N__30916\ : std_logic;
signal \N__30913\ : std_logic;
signal \N__30910\ : std_logic;
signal \N__30907\ : std_logic;
signal \N__30904\ : std_logic;
signal \N__30901\ : std_logic;
signal \N__30894\ : std_logic;
signal \N__30891\ : std_logic;
signal \N__30888\ : std_logic;
signal \N__30887\ : std_logic;
signal \N__30884\ : std_logic;
signal \N__30881\ : std_logic;
signal \N__30878\ : std_logic;
signal \N__30873\ : std_logic;
signal \N__30870\ : std_logic;
signal \N__30867\ : std_logic;
signal \N__30864\ : std_logic;
signal \N__30861\ : std_logic;
signal \N__30858\ : std_logic;
signal \N__30855\ : std_logic;
signal \N__30854\ : std_logic;
signal \N__30851\ : std_logic;
signal \N__30848\ : std_logic;
signal \N__30843\ : std_logic;
signal \N__30840\ : std_logic;
signal \N__30837\ : std_logic;
signal \N__30834\ : std_logic;
signal \N__30833\ : std_logic;
signal \N__30830\ : std_logic;
signal \N__30827\ : std_logic;
signal \N__30822\ : std_logic;
signal \N__30819\ : std_logic;
signal \N__30816\ : std_logic;
signal \N__30815\ : std_logic;
signal \N__30812\ : std_logic;
signal \N__30811\ : std_logic;
signal \N__30808\ : std_logic;
signal \N__30805\ : std_logic;
signal \N__30802\ : std_logic;
signal \N__30799\ : std_logic;
signal \N__30796\ : std_logic;
signal \N__30793\ : std_logic;
signal \N__30792\ : std_logic;
signal \N__30791\ : std_logic;
signal \N__30788\ : std_logic;
signal \N__30785\ : std_logic;
signal \N__30782\ : std_logic;
signal \N__30779\ : std_logic;
signal \N__30776\ : std_logic;
signal \N__30771\ : std_logic;
signal \N__30762\ : std_logic;
signal \N__30759\ : std_logic;
signal \N__30756\ : std_logic;
signal \N__30753\ : std_logic;
signal \N__30750\ : std_logic;
signal \N__30747\ : std_logic;
signal \N__30744\ : std_logic;
signal \N__30743\ : std_logic;
signal \N__30740\ : std_logic;
signal \N__30737\ : std_logic;
signal \N__30732\ : std_logic;
signal \N__30729\ : std_logic;
signal \N__30726\ : std_logic;
signal \N__30723\ : std_logic;
signal \N__30722\ : std_logic;
signal \N__30719\ : std_logic;
signal \N__30716\ : std_logic;
signal \N__30713\ : std_logic;
signal \N__30712\ : std_logic;
signal \N__30709\ : std_logic;
signal \N__30706\ : std_logic;
signal \N__30703\ : std_logic;
signal \N__30696\ : std_logic;
signal \N__30693\ : std_logic;
signal \N__30690\ : std_logic;
signal \N__30687\ : std_logic;
signal \N__30684\ : std_logic;
signal \N__30681\ : std_logic;
signal \N__30678\ : std_logic;
signal \N__30675\ : std_logic;
signal \N__30672\ : std_logic;
signal \N__30671\ : std_logic;
signal \N__30670\ : std_logic;
signal \N__30667\ : std_logic;
signal \N__30664\ : std_logic;
signal \N__30661\ : std_logic;
signal \N__30658\ : std_logic;
signal \N__30655\ : std_logic;
signal \N__30648\ : std_logic;
signal \N__30645\ : std_logic;
signal \N__30642\ : std_logic;
signal \N__30639\ : std_logic;
signal \N__30636\ : std_logic;
signal \N__30635\ : std_logic;
signal \N__30632\ : std_logic;
signal \N__30629\ : std_logic;
signal \N__30628\ : std_logic;
signal \N__30625\ : std_logic;
signal \N__30622\ : std_logic;
signal \N__30619\ : std_logic;
signal \N__30612\ : std_logic;
signal \N__30609\ : std_logic;
signal \N__30606\ : std_logic;
signal \N__30603\ : std_logic;
signal \N__30600\ : std_logic;
signal \N__30597\ : std_logic;
signal \N__30596\ : std_logic;
signal \N__30593\ : std_logic;
signal \N__30590\ : std_logic;
signal \N__30587\ : std_logic;
signal \N__30582\ : std_logic;
signal \N__30579\ : std_logic;
signal \N__30576\ : std_logic;
signal \N__30573\ : std_logic;
signal \N__30570\ : std_logic;
signal \N__30569\ : std_logic;
signal \N__30566\ : std_logic;
signal \N__30563\ : std_logic;
signal \N__30562\ : std_logic;
signal \N__30559\ : std_logic;
signal \N__30556\ : std_logic;
signal \N__30553\ : std_logic;
signal \N__30546\ : std_logic;
signal \N__30543\ : std_logic;
signal \N__30540\ : std_logic;
signal \N__30537\ : std_logic;
signal \N__30534\ : std_logic;
signal \N__30533\ : std_logic;
signal \N__30532\ : std_logic;
signal \N__30529\ : std_logic;
signal \N__30528\ : std_logic;
signal \N__30525\ : std_logic;
signal \N__30522\ : std_logic;
signal \N__30519\ : std_logic;
signal \N__30516\ : std_logic;
signal \N__30511\ : std_logic;
signal \N__30510\ : std_logic;
signal \N__30507\ : std_logic;
signal \N__30502\ : std_logic;
signal \N__30499\ : std_logic;
signal \N__30496\ : std_logic;
signal \N__30493\ : std_logic;
signal \N__30486\ : std_logic;
signal \N__30483\ : std_logic;
signal \N__30480\ : std_logic;
signal \N__30477\ : std_logic;
signal \N__30474\ : std_logic;
signal \N__30471\ : std_logic;
signal \N__30470\ : std_logic;
signal \N__30467\ : std_logic;
signal \N__30464\ : std_logic;
signal \N__30461\ : std_logic;
signal \N__30456\ : std_logic;
signal \N__30453\ : std_logic;
signal \N__30450\ : std_logic;
signal \N__30447\ : std_logic;
signal \N__30446\ : std_logic;
signal \N__30443\ : std_logic;
signal \N__30440\ : std_logic;
signal \N__30437\ : std_logic;
signal \N__30432\ : std_logic;
signal \N__30429\ : std_logic;
signal \N__30426\ : std_logic;
signal \N__30423\ : std_logic;
signal \N__30422\ : std_logic;
signal \N__30419\ : std_logic;
signal \N__30416\ : std_logic;
signal \N__30413\ : std_logic;
signal \N__30408\ : std_logic;
signal \N__30405\ : std_logic;
signal \N__30402\ : std_logic;
signal \N__30399\ : std_logic;
signal \N__30398\ : std_logic;
signal \N__30397\ : std_logic;
signal \N__30392\ : std_logic;
signal \N__30389\ : std_logic;
signal \N__30384\ : std_logic;
signal \N__30381\ : std_logic;
signal \N__30378\ : std_logic;
signal \N__30375\ : std_logic;
signal \N__30372\ : std_logic;
signal \N__30369\ : std_logic;
signal \N__30366\ : std_logic;
signal \N__30365\ : std_logic;
signal \N__30362\ : std_logic;
signal \N__30359\ : std_logic;
signal \N__30354\ : std_logic;
signal \N__30351\ : std_logic;
signal \N__30348\ : std_logic;
signal \N__30345\ : std_logic;
signal \N__30342\ : std_logic;
signal \N__30339\ : std_logic;
signal \N__30338\ : std_logic;
signal \N__30337\ : std_logic;
signal \N__30334\ : std_logic;
signal \N__30331\ : std_logic;
signal \N__30328\ : std_logic;
signal \N__30325\ : std_logic;
signal \N__30318\ : std_logic;
signal \N__30315\ : std_logic;
signal \N__30312\ : std_logic;
signal \N__30309\ : std_logic;
signal \N__30306\ : std_logic;
signal \N__30305\ : std_logic;
signal \N__30302\ : std_logic;
signal \N__30299\ : std_logic;
signal \N__30296\ : std_logic;
signal \N__30291\ : std_logic;
signal \N__30288\ : std_logic;
signal \N__30285\ : std_logic;
signal \N__30282\ : std_logic;
signal \N__30281\ : std_logic;
signal \N__30278\ : std_logic;
signal \N__30275\ : std_logic;
signal \N__30270\ : std_logic;
signal \N__30267\ : std_logic;
signal \N__30264\ : std_logic;
signal \N__30261\ : std_logic;
signal \N__30258\ : std_logic;
signal \N__30255\ : std_logic;
signal \N__30252\ : std_logic;
signal \N__30249\ : std_logic;
signal \N__30246\ : std_logic;
signal \N__30243\ : std_logic;
signal \N__30240\ : std_logic;
signal \N__30237\ : std_logic;
signal \N__30234\ : std_logic;
signal \N__30231\ : std_logic;
signal \N__30228\ : std_logic;
signal \N__30225\ : std_logic;
signal \N__30222\ : std_logic;
signal \N__30219\ : std_logic;
signal \N__30216\ : std_logic;
signal \N__30213\ : std_logic;
signal \N__30210\ : std_logic;
signal \N__30207\ : std_logic;
signal \N__30204\ : std_logic;
signal \N__30201\ : std_logic;
signal \N__30198\ : std_logic;
signal \N__30195\ : std_logic;
signal \N__30192\ : std_logic;
signal \N__30189\ : std_logic;
signal \N__30186\ : std_logic;
signal \N__30183\ : std_logic;
signal \N__30180\ : std_logic;
signal \N__30177\ : std_logic;
signal \N__30174\ : std_logic;
signal \N__30171\ : std_logic;
signal \N__30168\ : std_logic;
signal \N__30165\ : std_logic;
signal \N__30162\ : std_logic;
signal \N__30159\ : std_logic;
signal \N__30156\ : std_logic;
signal \N__30153\ : std_logic;
signal \N__30150\ : std_logic;
signal \N__30147\ : std_logic;
signal \N__30146\ : std_logic;
signal \N__30143\ : std_logic;
signal \N__30142\ : std_logic;
signal \N__30139\ : std_logic;
signal \N__30136\ : std_logic;
signal \N__30133\ : std_logic;
signal \N__30132\ : std_logic;
signal \N__30129\ : std_logic;
signal \N__30124\ : std_logic;
signal \N__30123\ : std_logic;
signal \N__30120\ : std_logic;
signal \N__30115\ : std_logic;
signal \N__30112\ : std_logic;
signal \N__30109\ : std_logic;
signal \N__30106\ : std_logic;
signal \N__30101\ : std_logic;
signal \N__30096\ : std_logic;
signal \N__30093\ : std_logic;
signal \N__30090\ : std_logic;
signal \N__30087\ : std_logic;
signal \N__30084\ : std_logic;
signal \N__30083\ : std_logic;
signal \N__30080\ : std_logic;
signal \N__30077\ : std_logic;
signal \N__30074\ : std_logic;
signal \N__30071\ : std_logic;
signal \N__30066\ : std_logic;
signal \N__30063\ : std_logic;
signal \N__30062\ : std_logic;
signal \N__30059\ : std_logic;
signal \N__30056\ : std_logic;
signal \N__30055\ : std_logic;
signal \N__30052\ : std_logic;
signal \N__30049\ : std_logic;
signal \N__30046\ : std_logic;
signal \N__30039\ : std_logic;
signal \N__30036\ : std_logic;
signal \N__30035\ : std_logic;
signal \N__30032\ : std_logic;
signal \N__30031\ : std_logic;
signal \N__30028\ : std_logic;
signal \N__30025\ : std_logic;
signal \N__30022\ : std_logic;
signal \N__30015\ : std_logic;
signal \N__30012\ : std_logic;
signal \N__30009\ : std_logic;
signal \N__30006\ : std_logic;
signal \N__30003\ : std_logic;
signal \N__30000\ : std_logic;
signal \N__29999\ : std_logic;
signal \N__29996\ : std_logic;
signal \N__29995\ : std_logic;
signal \N__29992\ : std_logic;
signal \N__29989\ : std_logic;
signal \N__29986\ : std_logic;
signal \N__29983\ : std_logic;
signal \N__29976\ : std_logic;
signal \N__29973\ : std_logic;
signal \N__29970\ : std_logic;
signal \N__29967\ : std_logic;
signal \N__29964\ : std_logic;
signal \N__29961\ : std_logic;
signal \N__29958\ : std_logic;
signal \N__29955\ : std_logic;
signal \N__29952\ : std_logic;
signal \N__29949\ : std_logic;
signal \N__29946\ : std_logic;
signal \N__29943\ : std_logic;
signal \N__29942\ : std_logic;
signal \N__29939\ : std_logic;
signal \N__29938\ : std_logic;
signal \N__29935\ : std_logic;
signal \N__29932\ : std_logic;
signal \N__29929\ : std_logic;
signal \N__29922\ : std_logic;
signal \N__29921\ : std_logic;
signal \N__29918\ : std_logic;
signal \N__29915\ : std_logic;
signal \N__29912\ : std_logic;
signal \N__29907\ : std_logic;
signal \N__29904\ : std_logic;
signal \N__29901\ : std_logic;
signal \N__29898\ : std_logic;
signal \N__29895\ : std_logic;
signal \N__29894\ : std_logic;
signal \N__29891\ : std_logic;
signal \N__29888\ : std_logic;
signal \N__29885\ : std_logic;
signal \N__29882\ : std_logic;
signal \N__29877\ : std_logic;
signal \N__29874\ : std_logic;
signal \N__29871\ : std_logic;
signal \N__29868\ : std_logic;
signal \N__29865\ : std_logic;
signal \N__29862\ : std_logic;
signal \N__29859\ : std_logic;
signal \N__29858\ : std_logic;
signal \N__29855\ : std_logic;
signal \N__29852\ : std_logic;
signal \N__29849\ : std_logic;
signal \N__29846\ : std_logic;
signal \N__29841\ : std_logic;
signal \N__29838\ : std_logic;
signal \N__29835\ : std_logic;
signal \N__29832\ : std_logic;
signal \N__29829\ : std_logic;
signal \N__29826\ : std_logic;
signal \N__29823\ : std_logic;
signal \N__29820\ : std_logic;
signal \N__29817\ : std_logic;
signal \N__29814\ : std_logic;
signal \N__29811\ : std_logic;
signal \N__29808\ : std_logic;
signal \N__29805\ : std_logic;
signal \N__29802\ : std_logic;
signal \N__29799\ : std_logic;
signal \N__29798\ : std_logic;
signal \N__29797\ : std_logic;
signal \N__29794\ : std_logic;
signal \N__29789\ : std_logic;
signal \N__29784\ : std_logic;
signal \N__29781\ : std_logic;
signal \N__29778\ : std_logic;
signal \N__29775\ : std_logic;
signal \N__29774\ : std_logic;
signal \N__29773\ : std_logic;
signal \N__29770\ : std_logic;
signal \N__29767\ : std_logic;
signal \N__29764\ : std_logic;
signal \N__29761\ : std_logic;
signal \N__29758\ : std_logic;
signal \N__29751\ : std_logic;
signal \N__29748\ : std_logic;
signal \N__29745\ : std_logic;
signal \N__29742\ : std_logic;
signal \N__29741\ : std_logic;
signal \N__29738\ : std_logic;
signal \N__29735\ : std_logic;
signal \N__29732\ : std_logic;
signal \N__29727\ : std_logic;
signal \N__29724\ : std_logic;
signal \N__29723\ : std_logic;
signal \N__29720\ : std_logic;
signal \N__29717\ : std_logic;
signal \N__29712\ : std_logic;
signal \N__29709\ : std_logic;
signal \N__29706\ : std_logic;
signal \N__29703\ : std_logic;
signal \N__29702\ : std_logic;
signal \N__29701\ : std_logic;
signal \N__29698\ : std_logic;
signal \N__29695\ : std_logic;
signal \N__29692\ : std_logic;
signal \N__29691\ : std_logic;
signal \N__29690\ : std_logic;
signal \N__29689\ : std_logic;
signal \N__29688\ : std_logic;
signal \N__29687\ : std_logic;
signal \N__29686\ : std_logic;
signal \N__29685\ : std_logic;
signal \N__29684\ : std_logic;
signal \N__29683\ : std_logic;
signal \N__29682\ : std_logic;
signal \N__29681\ : std_logic;
signal \N__29680\ : std_logic;
signal \N__29679\ : std_logic;
signal \N__29678\ : std_logic;
signal \N__29677\ : std_logic;
signal \N__29676\ : std_logic;
signal \N__29675\ : std_logic;
signal \N__29674\ : std_logic;
signal \N__29673\ : std_logic;
signal \N__29672\ : std_logic;
signal \N__29671\ : std_logic;
signal \N__29670\ : std_logic;
signal \N__29669\ : std_logic;
signal \N__29666\ : std_logic;
signal \N__29661\ : std_logic;
signal \N__29658\ : std_logic;
signal \N__29655\ : std_logic;
signal \N__29652\ : std_logic;
signal \N__29649\ : std_logic;
signal \N__29646\ : std_logic;
signal \N__29643\ : std_logic;
signal \N__29640\ : std_logic;
signal \N__29637\ : std_logic;
signal \N__29634\ : std_logic;
signal \N__29631\ : std_logic;
signal \N__29628\ : std_logic;
signal \N__29625\ : std_logic;
signal \N__29622\ : std_logic;
signal \N__29619\ : std_logic;
signal \N__29616\ : std_logic;
signal \N__29613\ : std_logic;
signal \N__29610\ : std_logic;
signal \N__29607\ : std_logic;
signal \N__29604\ : std_logic;
signal \N__29601\ : std_logic;
signal \N__29598\ : std_logic;
signal \N__29595\ : std_logic;
signal \N__29592\ : std_logic;
signal \N__29587\ : std_logic;
signal \N__29578\ : std_logic;
signal \N__29569\ : std_logic;
signal \N__29560\ : std_logic;
signal \N__29551\ : std_logic;
signal \N__29544\ : std_logic;
signal \N__29537\ : std_logic;
signal \N__29534\ : std_logic;
signal \N__29517\ : std_logic;
signal \N__29514\ : std_logic;
signal \N__29511\ : std_logic;
signal \N__29508\ : std_logic;
signal \N__29505\ : std_logic;
signal \N__29504\ : std_logic;
signal \N__29501\ : std_logic;
signal \N__29498\ : std_logic;
signal \N__29497\ : std_logic;
signal \N__29492\ : std_logic;
signal \N__29489\ : std_logic;
signal \N__29484\ : std_logic;
signal \N__29481\ : std_logic;
signal \N__29478\ : std_logic;
signal \N__29477\ : std_logic;
signal \N__29476\ : std_logic;
signal \N__29473\ : std_logic;
signal \N__29470\ : std_logic;
signal \N__29467\ : std_logic;
signal \N__29462\ : std_logic;
signal \N__29459\ : std_logic;
signal \N__29454\ : std_logic;
signal \N__29451\ : std_logic;
signal \N__29448\ : std_logic;
signal \N__29445\ : std_logic;
signal \N__29442\ : std_logic;
signal \N__29439\ : std_logic;
signal \N__29436\ : std_logic;
signal \N__29433\ : std_logic;
signal \N__29430\ : std_logic;
signal \N__29427\ : std_logic;
signal \N__29424\ : std_logic;
signal \N__29421\ : std_logic;
signal \N__29418\ : std_logic;
signal \N__29415\ : std_logic;
signal \N__29412\ : std_logic;
signal \N__29409\ : std_logic;
signal \N__29406\ : std_logic;
signal \N__29403\ : std_logic;
signal \N__29400\ : std_logic;
signal \N__29397\ : std_logic;
signal \N__29394\ : std_logic;
signal \N__29391\ : std_logic;
signal \N__29388\ : std_logic;
signal \N__29385\ : std_logic;
signal \N__29382\ : std_logic;
signal \N__29379\ : std_logic;
signal \N__29376\ : std_logic;
signal \N__29373\ : std_logic;
signal \N__29370\ : std_logic;
signal \N__29367\ : std_logic;
signal \N__29364\ : std_logic;
signal \N__29361\ : std_logic;
signal \N__29358\ : std_logic;
signal \N__29355\ : std_logic;
signal \N__29352\ : std_logic;
signal \N__29349\ : std_logic;
signal \N__29346\ : std_logic;
signal \N__29345\ : std_logic;
signal \N__29342\ : std_logic;
signal \N__29339\ : std_logic;
signal \N__29338\ : std_logic;
signal \N__29333\ : std_logic;
signal \N__29330\ : std_logic;
signal \N__29329\ : std_logic;
signal \N__29328\ : std_logic;
signal \N__29325\ : std_logic;
signal \N__29322\ : std_logic;
signal \N__29319\ : std_logic;
signal \N__29316\ : std_logic;
signal \N__29313\ : std_logic;
signal \N__29310\ : std_logic;
signal \N__29301\ : std_logic;
signal \N__29298\ : std_logic;
signal \N__29297\ : std_logic;
signal \N__29294\ : std_logic;
signal \N__29291\ : std_logic;
signal \N__29286\ : std_logic;
signal \N__29283\ : std_logic;
signal \N__29280\ : std_logic;
signal \N__29277\ : std_logic;
signal \N__29276\ : std_logic;
signal \N__29273\ : std_logic;
signal \N__29270\ : std_logic;
signal \N__29267\ : std_logic;
signal \N__29264\ : std_logic;
signal \N__29259\ : std_logic;
signal \N__29256\ : std_logic;
signal \N__29253\ : std_logic;
signal \N__29250\ : std_logic;
signal \N__29249\ : std_logic;
signal \N__29248\ : std_logic;
signal \N__29245\ : std_logic;
signal \N__29242\ : std_logic;
signal \N__29239\ : std_logic;
signal \N__29232\ : std_logic;
signal \N__29229\ : std_logic;
signal \N__29228\ : std_logic;
signal \N__29227\ : std_logic;
signal \N__29224\ : std_logic;
signal \N__29221\ : std_logic;
signal \N__29218\ : std_logic;
signal \N__29211\ : std_logic;
signal \N__29208\ : std_logic;
signal \N__29205\ : std_logic;
signal \N__29204\ : std_logic;
signal \N__29201\ : std_logic;
signal \N__29200\ : std_logic;
signal \N__29197\ : std_logic;
signal \N__29194\ : std_logic;
signal \N__29191\ : std_logic;
signal \N__29188\ : std_logic;
signal \N__29181\ : std_logic;
signal \N__29178\ : std_logic;
signal \N__29175\ : std_logic;
signal \N__29172\ : std_logic;
signal \N__29169\ : std_logic;
signal \N__29166\ : std_logic;
signal \N__29163\ : std_logic;
signal \N__29160\ : std_logic;
signal \N__29157\ : std_logic;
signal \N__29154\ : std_logic;
signal \N__29153\ : std_logic;
signal \N__29150\ : std_logic;
signal \N__29147\ : std_logic;
signal \N__29144\ : std_logic;
signal \N__29143\ : std_logic;
signal \N__29140\ : std_logic;
signal \N__29137\ : std_logic;
signal \N__29134\ : std_logic;
signal \N__29127\ : std_logic;
signal \N__29126\ : std_logic;
signal \N__29125\ : std_logic;
signal \N__29124\ : std_logic;
signal \N__29123\ : std_logic;
signal \N__29122\ : std_logic;
signal \N__29121\ : std_logic;
signal \N__29120\ : std_logic;
signal \N__29117\ : std_logic;
signal \N__29116\ : std_logic;
signal \N__29113\ : std_logic;
signal \N__29112\ : std_logic;
signal \N__29111\ : std_logic;
signal \N__29108\ : std_logic;
signal \N__29107\ : std_logic;
signal \N__29106\ : std_logic;
signal \N__29105\ : std_logic;
signal \N__29102\ : std_logic;
signal \N__29099\ : std_logic;
signal \N__29096\ : std_logic;
signal \N__29095\ : std_logic;
signal \N__29094\ : std_logic;
signal \N__29089\ : std_logic;
signal \N__29084\ : std_logic;
signal \N__29075\ : std_logic;
signal \N__29068\ : std_logic;
signal \N__29057\ : std_logic;
signal \N__29048\ : std_logic;
signal \N__29043\ : std_logic;
signal \N__29040\ : std_logic;
signal \N__29037\ : std_logic;
signal \N__29034\ : std_logic;
signal \N__29031\ : std_logic;
signal \N__29028\ : std_logic;
signal \N__29025\ : std_logic;
signal \N__29022\ : std_logic;
signal \N__29021\ : std_logic;
signal \N__29020\ : std_logic;
signal \N__29017\ : std_logic;
signal \N__29014\ : std_logic;
signal \N__29011\ : std_logic;
signal \N__29008\ : std_logic;
signal \N__29005\ : std_logic;
signal \N__29002\ : std_logic;
signal \N__28995\ : std_logic;
signal \N__28992\ : std_logic;
signal \N__28989\ : std_logic;
signal \N__28986\ : std_logic;
signal \N__28983\ : std_logic;
signal \N__28982\ : std_logic;
signal \N__28979\ : std_logic;
signal \N__28976\ : std_logic;
signal \N__28973\ : std_logic;
signal \N__28970\ : std_logic;
signal \N__28965\ : std_logic;
signal \N__28964\ : std_logic;
signal \N__28961\ : std_logic;
signal \N__28958\ : std_logic;
signal \N__28953\ : std_logic;
signal \N__28950\ : std_logic;
signal \N__28947\ : std_logic;
signal \N__28944\ : std_logic;
signal \N__28941\ : std_logic;
signal \N__28938\ : std_logic;
signal \N__28937\ : std_logic;
signal \N__28936\ : std_logic;
signal \N__28933\ : std_logic;
signal \N__28930\ : std_logic;
signal \N__28929\ : std_logic;
signal \N__28926\ : std_logic;
signal \N__28921\ : std_logic;
signal \N__28918\ : std_logic;
signal \N__28917\ : std_logic;
signal \N__28914\ : std_logic;
signal \N__28909\ : std_logic;
signal \N__28906\ : std_logic;
signal \N__28903\ : std_logic;
signal \N__28900\ : std_logic;
signal \N__28893\ : std_logic;
signal \N__28890\ : std_logic;
signal \N__28887\ : std_logic;
signal \N__28884\ : std_logic;
signal \N__28881\ : std_logic;
signal \N__28878\ : std_logic;
signal \N__28875\ : std_logic;
signal \N__28872\ : std_logic;
signal \N__28869\ : std_logic;
signal \N__28868\ : std_logic;
signal \N__28867\ : std_logic;
signal \N__28864\ : std_logic;
signal \N__28859\ : std_logic;
signal \N__28856\ : std_logic;
signal \N__28851\ : std_logic;
signal \N__28848\ : std_logic;
signal \N__28847\ : std_logic;
signal \N__28844\ : std_logic;
signal \N__28843\ : std_logic;
signal \N__28840\ : std_logic;
signal \N__28837\ : std_logic;
signal \N__28832\ : std_logic;
signal \N__28827\ : std_logic;
signal \N__28824\ : std_logic;
signal \N__28821\ : std_logic;
signal \N__28820\ : std_logic;
signal \N__28819\ : std_logic;
signal \N__28816\ : std_logic;
signal \N__28813\ : std_logic;
signal \N__28810\ : std_logic;
signal \N__28807\ : std_logic;
signal \N__28804\ : std_logic;
signal \N__28797\ : std_logic;
signal \N__28794\ : std_logic;
signal \N__28791\ : std_logic;
signal \N__28790\ : std_logic;
signal \N__28789\ : std_logic;
signal \N__28786\ : std_logic;
signal \N__28783\ : std_logic;
signal \N__28780\ : std_logic;
signal \N__28777\ : std_logic;
signal \N__28774\ : std_logic;
signal \N__28771\ : std_logic;
signal \N__28764\ : std_logic;
signal \N__28761\ : std_logic;
signal \N__28758\ : std_logic;
signal \N__28755\ : std_logic;
signal \N__28754\ : std_logic;
signal \N__28751\ : std_logic;
signal \N__28748\ : std_logic;
signal \N__28745\ : std_logic;
signal \N__28744\ : std_logic;
signal \N__28741\ : std_logic;
signal \N__28738\ : std_logic;
signal \N__28735\ : std_logic;
signal \N__28728\ : std_logic;
signal \N__28725\ : std_logic;
signal \N__28722\ : std_logic;
signal \N__28719\ : std_logic;
signal \N__28716\ : std_logic;
signal \N__28713\ : std_logic;
signal \N__28712\ : std_logic;
signal \N__28711\ : std_logic;
signal \N__28708\ : std_logic;
signal \N__28705\ : std_logic;
signal \N__28702\ : std_logic;
signal \N__28699\ : std_logic;
signal \N__28696\ : std_logic;
signal \N__28693\ : std_logic;
signal \N__28686\ : std_logic;
signal \N__28683\ : std_logic;
signal \N__28680\ : std_logic;
signal \N__28679\ : std_logic;
signal \N__28676\ : std_logic;
signal \N__28673\ : std_logic;
signal \N__28672\ : std_logic;
signal \N__28669\ : std_logic;
signal \N__28666\ : std_logic;
signal \N__28663\ : std_logic;
signal \N__28656\ : std_logic;
signal \N__28653\ : std_logic;
signal \N__28650\ : std_logic;
signal \N__28647\ : std_logic;
signal \N__28644\ : std_logic;
signal \N__28643\ : std_logic;
signal \N__28640\ : std_logic;
signal \N__28637\ : std_logic;
signal \N__28636\ : std_logic;
signal \N__28633\ : std_logic;
signal \N__28630\ : std_logic;
signal \N__28627\ : std_logic;
signal \N__28624\ : std_logic;
signal \N__28617\ : std_logic;
signal \N__28614\ : std_logic;
signal \N__28611\ : std_logic;
signal \N__28608\ : std_logic;
signal \N__28607\ : std_logic;
signal \N__28604\ : std_logic;
signal \N__28601\ : std_logic;
signal \N__28598\ : std_logic;
signal \N__28595\ : std_logic;
signal \N__28590\ : std_logic;
signal \N__28587\ : std_logic;
signal \N__28584\ : std_logic;
signal \N__28581\ : std_logic;
signal \N__28578\ : std_logic;
signal \N__28575\ : std_logic;
signal \N__28572\ : std_logic;
signal \N__28569\ : std_logic;
signal \N__28566\ : std_logic;
signal \N__28563\ : std_logic;
signal \N__28560\ : std_logic;
signal \N__28557\ : std_logic;
signal \N__28554\ : std_logic;
signal \N__28553\ : std_logic;
signal \N__28550\ : std_logic;
signal \N__28547\ : std_logic;
signal \N__28544\ : std_logic;
signal \N__28541\ : std_logic;
signal \N__28536\ : std_logic;
signal \N__28533\ : std_logic;
signal \N__28530\ : std_logic;
signal \N__28527\ : std_logic;
signal \N__28524\ : std_logic;
signal \N__28523\ : std_logic;
signal \N__28522\ : std_logic;
signal \N__28519\ : std_logic;
signal \N__28514\ : std_logic;
signal \N__28509\ : std_logic;
signal \N__28506\ : std_logic;
signal \N__28503\ : std_logic;
signal \N__28500\ : std_logic;
signal \N__28497\ : std_logic;
signal \N__28494\ : std_logic;
signal \N__28491\ : std_logic;
signal \N__28488\ : std_logic;
signal \N__28485\ : std_logic;
signal \N__28482\ : std_logic;
signal \N__28479\ : std_logic;
signal \N__28476\ : std_logic;
signal \N__28473\ : std_logic;
signal \N__28470\ : std_logic;
signal \N__28467\ : std_logic;
signal \N__28464\ : std_logic;
signal \N__28461\ : std_logic;
signal \N__28458\ : std_logic;
signal \N__28455\ : std_logic;
signal \N__28452\ : std_logic;
signal \N__28449\ : std_logic;
signal \N__28446\ : std_logic;
signal \N__28443\ : std_logic;
signal \N__28440\ : std_logic;
signal \N__28437\ : std_logic;
signal \N__28434\ : std_logic;
signal \N__28431\ : std_logic;
signal \N__28428\ : std_logic;
signal \N__28425\ : std_logic;
signal \N__28422\ : std_logic;
signal \N__28419\ : std_logic;
signal \N__28416\ : std_logic;
signal \N__28413\ : std_logic;
signal \N__28410\ : std_logic;
signal \N__28407\ : std_logic;
signal \N__28404\ : std_logic;
signal \N__28401\ : std_logic;
signal \N__28398\ : std_logic;
signal \N__28395\ : std_logic;
signal \N__28392\ : std_logic;
signal \N__28389\ : std_logic;
signal \N__28386\ : std_logic;
signal \N__28383\ : std_logic;
signal \N__28380\ : std_logic;
signal \N__28377\ : std_logic;
signal \N__28374\ : std_logic;
signal \N__28371\ : std_logic;
signal \N__28368\ : std_logic;
signal \N__28365\ : std_logic;
signal \N__28362\ : std_logic;
signal \N__28359\ : std_logic;
signal \N__28356\ : std_logic;
signal \N__28353\ : std_logic;
signal \N__28350\ : std_logic;
signal \N__28347\ : std_logic;
signal \N__28344\ : std_logic;
signal \N__28341\ : std_logic;
signal \N__28340\ : std_logic;
signal \N__28337\ : std_logic;
signal \N__28336\ : std_logic;
signal \N__28333\ : std_logic;
signal \N__28330\ : std_logic;
signal \N__28327\ : std_logic;
signal \N__28324\ : std_logic;
signal \N__28319\ : std_logic;
signal \N__28314\ : std_logic;
signal \N__28311\ : std_logic;
signal \N__28308\ : std_logic;
signal \N__28305\ : std_logic;
signal \N__28302\ : std_logic;
signal \N__28299\ : std_logic;
signal \N__28296\ : std_logic;
signal \N__28293\ : std_logic;
signal \N__28290\ : std_logic;
signal \N__28287\ : std_logic;
signal \N__28284\ : std_logic;
signal \N__28281\ : std_logic;
signal \N__28278\ : std_logic;
signal \N__28275\ : std_logic;
signal \N__28272\ : std_logic;
signal \N__28269\ : std_logic;
signal \N__28266\ : std_logic;
signal \N__28263\ : std_logic;
signal \N__28260\ : std_logic;
signal \N__28257\ : std_logic;
signal \N__28254\ : std_logic;
signal \N__28251\ : std_logic;
signal \N__28248\ : std_logic;
signal \N__28245\ : std_logic;
signal \N__28242\ : std_logic;
signal \N__28239\ : std_logic;
signal \N__28236\ : std_logic;
signal \N__28233\ : std_logic;
signal \N__28230\ : std_logic;
signal \N__28229\ : std_logic;
signal \N__28226\ : std_logic;
signal \N__28223\ : std_logic;
signal \N__28218\ : std_logic;
signal \N__28215\ : std_logic;
signal \N__28214\ : std_logic;
signal \N__28213\ : std_logic;
signal \N__28210\ : std_logic;
signal \N__28207\ : std_logic;
signal \N__28206\ : std_logic;
signal \N__28205\ : std_logic;
signal \N__28202\ : std_logic;
signal \N__28199\ : std_logic;
signal \N__28196\ : std_logic;
signal \N__28193\ : std_logic;
signal \N__28190\ : std_logic;
signal \N__28187\ : std_logic;
signal \N__28180\ : std_logic;
signal \N__28175\ : std_logic;
signal \N__28172\ : std_logic;
signal \N__28167\ : std_logic;
signal \N__28164\ : std_logic;
signal \N__28161\ : std_logic;
signal \N__28160\ : std_logic;
signal \N__28157\ : std_logic;
signal \N__28154\ : std_logic;
signal \N__28151\ : std_logic;
signal \N__28146\ : std_logic;
signal \N__28143\ : std_logic;
signal \N__28140\ : std_logic;
signal \N__28137\ : std_logic;
signal \N__28136\ : std_logic;
signal \N__28133\ : std_logic;
signal \N__28130\ : std_logic;
signal \N__28129\ : std_logic;
signal \N__28126\ : std_logic;
signal \N__28123\ : std_logic;
signal \N__28120\ : std_logic;
signal \N__28113\ : std_logic;
signal \N__28110\ : std_logic;
signal \N__28109\ : std_logic;
signal \N__28108\ : std_logic;
signal \N__28103\ : std_logic;
signal \N__28100\ : std_logic;
signal \N__28097\ : std_logic;
signal \N__28094\ : std_logic;
signal \N__28091\ : std_logic;
signal \N__28088\ : std_logic;
signal \N__28083\ : std_logic;
signal \N__28082\ : std_logic;
signal \N__28081\ : std_logic;
signal \N__28078\ : std_logic;
signal \N__28075\ : std_logic;
signal \N__28072\ : std_logic;
signal \N__28069\ : std_logic;
signal \N__28062\ : std_logic;
signal \N__28059\ : std_logic;
signal \N__28056\ : std_logic;
signal \N__28053\ : std_logic;
signal \N__28050\ : std_logic;
signal \N__28047\ : std_logic;
signal \N__28044\ : std_logic;
signal \N__28041\ : std_logic;
signal \N__28038\ : std_logic;
signal \N__28035\ : std_logic;
signal \N__28032\ : std_logic;
signal \N__28031\ : std_logic;
signal \N__28028\ : std_logic;
signal \N__28027\ : std_logic;
signal \N__28024\ : std_logic;
signal \N__28019\ : std_logic;
signal \N__28016\ : std_logic;
signal \N__28011\ : std_logic;
signal \N__28008\ : std_logic;
signal \N__28005\ : std_logic;
signal \N__28002\ : std_logic;
signal \N__27999\ : std_logic;
signal \N__27996\ : std_logic;
signal \N__27993\ : std_logic;
signal \N__27990\ : std_logic;
signal \N__27987\ : std_logic;
signal \N__27984\ : std_logic;
signal \N__27981\ : std_logic;
signal \N__27978\ : std_logic;
signal \N__27975\ : std_logic;
signal \N__27974\ : std_logic;
signal \N__27971\ : std_logic;
signal \N__27970\ : std_logic;
signal \N__27967\ : std_logic;
signal \N__27964\ : std_logic;
signal \N__27961\ : std_logic;
signal \N__27958\ : std_logic;
signal \N__27955\ : std_logic;
signal \N__27952\ : std_logic;
signal \N__27949\ : std_logic;
signal \N__27942\ : std_logic;
signal \N__27939\ : std_logic;
signal \N__27936\ : std_logic;
signal \N__27933\ : std_logic;
signal \N__27930\ : std_logic;
signal \N__27927\ : std_logic;
signal \N__27924\ : std_logic;
signal \N__27921\ : std_logic;
signal \N__27918\ : std_logic;
signal \N__27915\ : std_logic;
signal \N__27912\ : std_logic;
signal \N__27909\ : std_logic;
signal \N__27906\ : std_logic;
signal \N__27903\ : std_logic;
signal \N__27900\ : std_logic;
signal \N__27897\ : std_logic;
signal \N__27894\ : std_logic;
signal \N__27891\ : std_logic;
signal \N__27888\ : std_logic;
signal \N__27885\ : std_logic;
signal \N__27884\ : std_logic;
signal \N__27879\ : std_logic;
signal \N__27878\ : std_logic;
signal \N__27875\ : std_logic;
signal \N__27872\ : std_logic;
signal \N__27867\ : std_logic;
signal \N__27864\ : std_logic;
signal \N__27863\ : std_logic;
signal \N__27858\ : std_logic;
signal \N__27857\ : std_logic;
signal \N__27854\ : std_logic;
signal \N__27851\ : std_logic;
signal \N__27846\ : std_logic;
signal \N__27843\ : std_logic;
signal \N__27842\ : std_logic;
signal \N__27839\ : std_logic;
signal \N__27834\ : std_logic;
signal \N__27833\ : std_logic;
signal \N__27830\ : std_logic;
signal \N__27827\ : std_logic;
signal \N__27822\ : std_logic;
signal \N__27819\ : std_logic;
signal \N__27816\ : std_logic;
signal \N__27815\ : std_logic;
signal \N__27810\ : std_logic;
signal \N__27807\ : std_logic;
signal \N__27806\ : std_logic;
signal \N__27803\ : std_logic;
signal \N__27800\ : std_logic;
signal \N__27795\ : std_logic;
signal \N__27792\ : std_logic;
signal \N__27789\ : std_logic;
signal \N__27786\ : std_logic;
signal \N__27783\ : std_logic;
signal \N__27782\ : std_logic;
signal \N__27779\ : std_logic;
signal \N__27776\ : std_logic;
signal \N__27771\ : std_logic;
signal \N__27768\ : std_logic;
signal \N__27765\ : std_logic;
signal \N__27762\ : std_logic;
signal \N__27759\ : std_logic;
signal \N__27756\ : std_logic;
signal \N__27753\ : std_logic;
signal \N__27750\ : std_logic;
signal \N__27747\ : std_logic;
signal \N__27744\ : std_logic;
signal \N__27741\ : std_logic;
signal \N__27738\ : std_logic;
signal \N__27735\ : std_logic;
signal \N__27732\ : std_logic;
signal \N__27729\ : std_logic;
signal \N__27726\ : std_logic;
signal \N__27723\ : std_logic;
signal \N__27720\ : std_logic;
signal \N__27717\ : std_logic;
signal \N__27714\ : std_logic;
signal \N__27711\ : std_logic;
signal \N__27708\ : std_logic;
signal \N__27705\ : std_logic;
signal \N__27702\ : std_logic;
signal \N__27699\ : std_logic;
signal \N__27696\ : std_logic;
signal \N__27693\ : std_logic;
signal \N__27690\ : std_logic;
signal \N__27687\ : std_logic;
signal \N__27684\ : std_logic;
signal \N__27681\ : std_logic;
signal \N__27678\ : std_logic;
signal \N__27675\ : std_logic;
signal \N__27672\ : std_logic;
signal \N__27669\ : std_logic;
signal \N__27666\ : std_logic;
signal \N__27663\ : std_logic;
signal \N__27660\ : std_logic;
signal \N__27657\ : std_logic;
signal \N__27654\ : std_logic;
signal \N__27651\ : std_logic;
signal \N__27648\ : std_logic;
signal \N__27645\ : std_logic;
signal \N__27642\ : std_logic;
signal \N__27639\ : std_logic;
signal \N__27636\ : std_logic;
signal \N__27633\ : std_logic;
signal \N__27630\ : std_logic;
signal \N__27627\ : std_logic;
signal \N__27624\ : std_logic;
signal \N__27621\ : std_logic;
signal \N__27618\ : std_logic;
signal \N__27615\ : std_logic;
signal \N__27612\ : std_logic;
signal \N__27609\ : std_logic;
signal \N__27606\ : std_logic;
signal \N__27605\ : std_logic;
signal \N__27602\ : std_logic;
signal \N__27601\ : std_logic;
signal \N__27598\ : std_logic;
signal \N__27595\ : std_logic;
signal \N__27592\ : std_logic;
signal \N__27589\ : std_logic;
signal \N__27582\ : std_logic;
signal \N__27581\ : std_logic;
signal \N__27580\ : std_logic;
signal \N__27577\ : std_logic;
signal \N__27576\ : std_logic;
signal \N__27573\ : std_logic;
signal \N__27572\ : std_logic;
signal \N__27569\ : std_logic;
signal \N__27568\ : std_logic;
signal \N__27567\ : std_logic;
signal \N__27558\ : std_logic;
signal \N__27553\ : std_logic;
signal \N__27552\ : std_logic;
signal \N__27551\ : std_logic;
signal \N__27550\ : std_logic;
signal \N__27547\ : std_logic;
signal \N__27546\ : std_logic;
signal \N__27545\ : std_logic;
signal \N__27544\ : std_logic;
signal \N__27543\ : std_logic;
signal \N__27540\ : std_logic;
signal \N__27537\ : std_logic;
signal \N__27534\ : std_logic;
signal \N__27525\ : std_logic;
signal \N__27522\ : std_logic;
signal \N__27519\ : std_logic;
signal \N__27518\ : std_logic;
signal \N__27515\ : std_logic;
signal \N__27510\ : std_logic;
signal \N__27505\ : std_logic;
signal \N__27498\ : std_logic;
signal \N__27489\ : std_logic;
signal \N__27486\ : std_logic;
signal \N__27483\ : std_logic;
signal \N__27480\ : std_logic;
signal \N__27477\ : std_logic;
signal \N__27474\ : std_logic;
signal \N__27471\ : std_logic;
signal \N__27468\ : std_logic;
signal \N__27465\ : std_logic;
signal \N__27462\ : std_logic;
signal \N__27459\ : std_logic;
signal \N__27456\ : std_logic;
signal \N__27453\ : std_logic;
signal \N__27450\ : std_logic;
signal \N__27447\ : std_logic;
signal \N__27444\ : std_logic;
signal \N__27441\ : std_logic;
signal \N__27438\ : std_logic;
signal \N__27435\ : std_logic;
signal \N__27432\ : std_logic;
signal \N__27429\ : std_logic;
signal \N__27426\ : std_logic;
signal \N__27423\ : std_logic;
signal \N__27420\ : std_logic;
signal \N__27417\ : std_logic;
signal \N__27414\ : std_logic;
signal \N__27411\ : std_logic;
signal \N__27408\ : std_logic;
signal \N__27407\ : std_logic;
signal \N__27404\ : std_logic;
signal \N__27401\ : std_logic;
signal \N__27396\ : std_logic;
signal \N__27393\ : std_logic;
signal \N__27392\ : std_logic;
signal \N__27389\ : std_logic;
signal \N__27386\ : std_logic;
signal \N__27383\ : std_logic;
signal \N__27380\ : std_logic;
signal \N__27375\ : std_logic;
signal \N__27372\ : std_logic;
signal \N__27369\ : std_logic;
signal \N__27366\ : std_logic;
signal \N__27363\ : std_logic;
signal \N__27360\ : std_logic;
signal \N__27357\ : std_logic;
signal \N__27356\ : std_logic;
signal \N__27355\ : std_logic;
signal \N__27352\ : std_logic;
signal \N__27349\ : std_logic;
signal \N__27346\ : std_logic;
signal \N__27343\ : std_logic;
signal \N__27340\ : std_logic;
signal \N__27337\ : std_logic;
signal \N__27330\ : std_logic;
signal \N__27327\ : std_logic;
signal \N__27324\ : std_logic;
signal \N__27321\ : std_logic;
signal \N__27318\ : std_logic;
signal \N__27315\ : std_logic;
signal \N__27312\ : std_logic;
signal \N__27309\ : std_logic;
signal \N__27306\ : std_logic;
signal \N__27303\ : std_logic;
signal \N__27300\ : std_logic;
signal \N__27297\ : std_logic;
signal \N__27294\ : std_logic;
signal \N__27293\ : std_logic;
signal \N__27290\ : std_logic;
signal \N__27289\ : std_logic;
signal \N__27286\ : std_logic;
signal \N__27283\ : std_logic;
signal \N__27280\ : std_logic;
signal \N__27275\ : std_logic;
signal \N__27272\ : std_logic;
signal \N__27271\ : std_logic;
signal \N__27270\ : std_logic;
signal \N__27267\ : std_logic;
signal \N__27264\ : std_logic;
signal \N__27261\ : std_logic;
signal \N__27258\ : std_logic;
signal \N__27255\ : std_logic;
signal \N__27252\ : std_logic;
signal \N__27243\ : std_logic;
signal \N__27240\ : std_logic;
signal \N__27237\ : std_logic;
signal \N__27234\ : std_logic;
signal \N__27231\ : std_logic;
signal \N__27228\ : std_logic;
signal \N__27225\ : std_logic;
signal \N__27222\ : std_logic;
signal \N__27219\ : std_logic;
signal \N__27216\ : std_logic;
signal \N__27213\ : std_logic;
signal \N__27212\ : std_logic;
signal \N__27209\ : std_logic;
signal \N__27206\ : std_logic;
signal \N__27205\ : std_logic;
signal \N__27202\ : std_logic;
signal \N__27199\ : std_logic;
signal \N__27196\ : std_logic;
signal \N__27189\ : std_logic;
signal \N__27186\ : std_logic;
signal \N__27183\ : std_logic;
signal \N__27180\ : std_logic;
signal \N__27177\ : std_logic;
signal \N__27174\ : std_logic;
signal \N__27171\ : std_logic;
signal \N__27170\ : std_logic;
signal \N__27167\ : std_logic;
signal \N__27164\ : std_logic;
signal \N__27163\ : std_logic;
signal \N__27160\ : std_logic;
signal \N__27157\ : std_logic;
signal \N__27154\ : std_logic;
signal \N__27147\ : std_logic;
signal \N__27144\ : std_logic;
signal \N__27141\ : std_logic;
signal \N__27138\ : std_logic;
signal \N__27135\ : std_logic;
signal \N__27132\ : std_logic;
signal \N__27131\ : std_logic;
signal \N__27128\ : std_logic;
signal \N__27127\ : std_logic;
signal \N__27124\ : std_logic;
signal \N__27121\ : std_logic;
signal \N__27118\ : std_logic;
signal \N__27115\ : std_logic;
signal \N__27108\ : std_logic;
signal \N__27105\ : std_logic;
signal \N__27102\ : std_logic;
signal \N__27099\ : std_logic;
signal \N__27096\ : std_logic;
signal \N__27093\ : std_logic;
signal \N__27090\ : std_logic;
signal \N__27089\ : std_logic;
signal \N__27088\ : std_logic;
signal \N__27085\ : std_logic;
signal \N__27082\ : std_logic;
signal \N__27079\ : std_logic;
signal \N__27076\ : std_logic;
signal \N__27073\ : std_logic;
signal \N__27070\ : std_logic;
signal \N__27063\ : std_logic;
signal \N__27060\ : std_logic;
signal \N__27057\ : std_logic;
signal \N__27054\ : std_logic;
signal \N__27051\ : std_logic;
signal \N__27048\ : std_logic;
signal \N__27047\ : std_logic;
signal \N__27046\ : std_logic;
signal \N__27043\ : std_logic;
signal \N__27038\ : std_logic;
signal \N__27035\ : std_logic;
signal \N__27032\ : std_logic;
signal \N__27027\ : std_logic;
signal \N__27024\ : std_logic;
signal \N__27021\ : std_logic;
signal \N__27018\ : std_logic;
signal \N__27015\ : std_logic;
signal \N__27012\ : std_logic;
signal \N__27009\ : std_logic;
signal \N__27006\ : std_logic;
signal \N__27003\ : std_logic;
signal \N__27000\ : std_logic;
signal \N__26997\ : std_logic;
signal \N__26994\ : std_logic;
signal \N__26991\ : std_logic;
signal \N__26988\ : std_logic;
signal \N__26985\ : std_logic;
signal \N__26982\ : std_logic;
signal \N__26981\ : std_logic;
signal \N__26978\ : std_logic;
signal \N__26975\ : std_logic;
signal \N__26970\ : std_logic;
signal \N__26967\ : std_logic;
signal \N__26964\ : std_logic;
signal \N__26961\ : std_logic;
signal \N__26958\ : std_logic;
signal \N__26955\ : std_logic;
signal \N__26952\ : std_logic;
signal \N__26949\ : std_logic;
signal \N__26946\ : std_logic;
signal \N__26943\ : std_logic;
signal \N__26940\ : std_logic;
signal \N__26937\ : std_logic;
signal \N__26934\ : std_logic;
signal \N__26931\ : std_logic;
signal \N__26928\ : std_logic;
signal \N__26925\ : std_logic;
signal \N__26922\ : std_logic;
signal \N__26919\ : std_logic;
signal \N__26916\ : std_logic;
signal \N__26913\ : std_logic;
signal \N__26910\ : std_logic;
signal \N__26907\ : std_logic;
signal \N__26904\ : std_logic;
signal \N__26901\ : std_logic;
signal \N__26898\ : std_logic;
signal \N__26895\ : std_logic;
signal \N__26892\ : std_logic;
signal \N__26889\ : std_logic;
signal \N__26886\ : std_logic;
signal \N__26883\ : std_logic;
signal \N__26880\ : std_logic;
signal \N__26877\ : std_logic;
signal \N__26874\ : std_logic;
signal \N__26871\ : std_logic;
signal \N__26870\ : std_logic;
signal \N__26867\ : std_logic;
signal \N__26864\ : std_logic;
signal \N__26859\ : std_logic;
signal \N__26856\ : std_logic;
signal \N__26855\ : std_logic;
signal \N__26854\ : std_logic;
signal \N__26853\ : std_logic;
signal \N__26850\ : std_logic;
signal \N__26847\ : std_logic;
signal \N__26844\ : std_logic;
signal \N__26841\ : std_logic;
signal \N__26838\ : std_logic;
signal \N__26831\ : std_logic;
signal \N__26826\ : std_logic;
signal \N__26823\ : std_logic;
signal \N__26820\ : std_logic;
signal \N__26817\ : std_logic;
signal \N__26814\ : std_logic;
signal \N__26811\ : std_logic;
signal \N__26808\ : std_logic;
signal \N__26805\ : std_logic;
signal \N__26804\ : std_logic;
signal \N__26803\ : std_logic;
signal \N__26802\ : std_logic;
signal \N__26801\ : std_logic;
signal \N__26800\ : std_logic;
signal \N__26799\ : std_logic;
signal \N__26798\ : std_logic;
signal \N__26797\ : std_logic;
signal \N__26796\ : std_logic;
signal \N__26795\ : std_logic;
signal \N__26794\ : std_logic;
signal \N__26791\ : std_logic;
signal \N__26788\ : std_logic;
signal \N__26781\ : std_logic;
signal \N__26778\ : std_logic;
signal \N__26777\ : std_logic;
signal \N__26772\ : std_logic;
signal \N__26769\ : std_logic;
signal \N__26760\ : std_logic;
signal \N__26757\ : std_logic;
signal \N__26754\ : std_logic;
signal \N__26751\ : std_logic;
signal \N__26748\ : std_logic;
signal \N__26745\ : std_logic;
signal \N__26742\ : std_logic;
signal \N__26737\ : std_logic;
signal \N__26732\ : std_logic;
signal \N__26725\ : std_logic;
signal \N__26720\ : std_logic;
signal \N__26715\ : std_logic;
signal \N__26712\ : std_logic;
signal \N__26709\ : std_logic;
signal \N__26708\ : std_logic;
signal \N__26705\ : std_logic;
signal \N__26702\ : std_logic;
signal \N__26697\ : std_logic;
signal \N__26694\ : std_logic;
signal \N__26691\ : std_logic;
signal \N__26688\ : std_logic;
signal \N__26685\ : std_logic;
signal \N__26682\ : std_logic;
signal \N__26679\ : std_logic;
signal \N__26676\ : std_logic;
signal \N__26673\ : std_logic;
signal \N__26670\ : std_logic;
signal \N__26667\ : std_logic;
signal \N__26664\ : std_logic;
signal \N__26661\ : std_logic;
signal \N__26658\ : std_logic;
signal \N__26655\ : std_logic;
signal \N__26654\ : std_logic;
signal \N__26653\ : std_logic;
signal \N__26650\ : std_logic;
signal \N__26647\ : std_logic;
signal \N__26644\ : std_logic;
signal \N__26641\ : std_logic;
signal \N__26638\ : std_logic;
signal \N__26635\ : std_logic;
signal \N__26628\ : std_logic;
signal \N__26625\ : std_logic;
signal \N__26622\ : std_logic;
signal \N__26619\ : std_logic;
signal \N__26616\ : std_logic;
signal \N__26613\ : std_logic;
signal \N__26610\ : std_logic;
signal \N__26607\ : std_logic;
signal \N__26606\ : std_logic;
signal \N__26605\ : std_logic;
signal \N__26600\ : std_logic;
signal \N__26597\ : std_logic;
signal \N__26596\ : std_logic;
signal \N__26593\ : std_logic;
signal \N__26590\ : std_logic;
signal \N__26587\ : std_logic;
signal \N__26584\ : std_logic;
signal \N__26581\ : std_logic;
signal \N__26574\ : std_logic;
signal \N__26571\ : std_logic;
signal \N__26568\ : std_logic;
signal \N__26565\ : std_logic;
signal \N__26564\ : std_logic;
signal \N__26561\ : std_logic;
signal \N__26558\ : std_logic;
signal \N__26555\ : std_logic;
signal \N__26550\ : std_logic;
signal \N__26547\ : std_logic;
signal \N__26544\ : std_logic;
signal \N__26543\ : std_logic;
signal \N__26540\ : std_logic;
signal \N__26537\ : std_logic;
signal \N__26534\ : std_logic;
signal \N__26531\ : std_logic;
signal \N__26526\ : std_logic;
signal \N__26523\ : std_logic;
signal \N__26520\ : std_logic;
signal \N__26517\ : std_logic;
signal \N__26514\ : std_logic;
signal \N__26511\ : std_logic;
signal \N__26508\ : std_logic;
signal \N__26505\ : std_logic;
signal \N__26504\ : std_logic;
signal \N__26501\ : std_logic;
signal \N__26500\ : std_logic;
signal \N__26497\ : std_logic;
signal \N__26494\ : std_logic;
signal \N__26491\ : std_logic;
signal \N__26488\ : std_logic;
signal \N__26485\ : std_logic;
signal \N__26478\ : std_logic;
signal \N__26475\ : std_logic;
signal \N__26472\ : std_logic;
signal \N__26469\ : std_logic;
signal \N__26468\ : std_logic;
signal \N__26467\ : std_logic;
signal \N__26464\ : std_logic;
signal \N__26461\ : std_logic;
signal \N__26458\ : std_logic;
signal \N__26455\ : std_logic;
signal \N__26452\ : std_logic;
signal \N__26449\ : std_logic;
signal \N__26442\ : std_logic;
signal \N__26439\ : std_logic;
signal \N__26436\ : std_logic;
signal \N__26433\ : std_logic;
signal \N__26432\ : std_logic;
signal \N__26431\ : std_logic;
signal \N__26428\ : std_logic;
signal \N__26423\ : std_logic;
signal \N__26418\ : std_logic;
signal \N__26417\ : std_logic;
signal \N__26416\ : std_logic;
signal \N__26413\ : std_logic;
signal \N__26408\ : std_logic;
signal \N__26405\ : std_logic;
signal \N__26400\ : std_logic;
signal \N__26397\ : std_logic;
signal \N__26394\ : std_logic;
signal \N__26391\ : std_logic;
signal \N__26388\ : std_logic;
signal \N__26385\ : std_logic;
signal \N__26382\ : std_logic;
signal \N__26379\ : std_logic;
signal \N__26376\ : std_logic;
signal \N__26373\ : std_logic;
signal \N__26370\ : std_logic;
signal \N__26367\ : std_logic;
signal \N__26364\ : std_logic;
signal \N__26361\ : std_logic;
signal \N__26358\ : std_logic;
signal \N__26355\ : std_logic;
signal \N__26354\ : std_logic;
signal \N__26353\ : std_logic;
signal \N__26350\ : std_logic;
signal \N__26349\ : std_logic;
signal \N__26348\ : std_logic;
signal \N__26345\ : std_logic;
signal \N__26342\ : std_logic;
signal \N__26339\ : std_logic;
signal \N__26334\ : std_logic;
signal \N__26325\ : std_logic;
signal \N__26322\ : std_logic;
signal \N__26319\ : std_logic;
signal \N__26316\ : std_logic;
signal \N__26313\ : std_logic;
signal \N__26310\ : std_logic;
signal \N__26309\ : std_logic;
signal \N__26308\ : std_logic;
signal \N__26305\ : std_logic;
signal \N__26302\ : std_logic;
signal \N__26299\ : std_logic;
signal \N__26296\ : std_logic;
signal \N__26293\ : std_logic;
signal \N__26286\ : std_logic;
signal \N__26283\ : std_logic;
signal \N__26280\ : std_logic;
signal \N__26277\ : std_logic;
signal \N__26276\ : std_logic;
signal \N__26275\ : std_logic;
signal \N__26272\ : std_logic;
signal \N__26267\ : std_logic;
signal \N__26264\ : std_logic;
signal \N__26259\ : std_logic;
signal \N__26256\ : std_logic;
signal \N__26253\ : std_logic;
signal \N__26250\ : std_logic;
signal \N__26249\ : std_logic;
signal \N__26248\ : std_logic;
signal \N__26245\ : std_logic;
signal \N__26240\ : std_logic;
signal \N__26237\ : std_logic;
signal \N__26232\ : std_logic;
signal \N__26229\ : std_logic;
signal \N__26226\ : std_logic;
signal \N__26223\ : std_logic;
signal \N__26220\ : std_logic;
signal \N__26219\ : std_logic;
signal \N__26216\ : std_logic;
signal \N__26213\ : std_logic;
signal \N__26210\ : std_logic;
signal \N__26209\ : std_logic;
signal \N__26208\ : std_logic;
signal \N__26207\ : std_logic;
signal \N__26204\ : std_logic;
signal \N__26201\ : std_logic;
signal \N__26198\ : std_logic;
signal \N__26195\ : std_logic;
signal \N__26192\ : std_logic;
signal \N__26187\ : std_logic;
signal \N__26182\ : std_logic;
signal \N__26175\ : std_logic;
signal \N__26174\ : std_logic;
signal \N__26171\ : std_logic;
signal \N__26170\ : std_logic;
signal \N__26167\ : std_logic;
signal \N__26162\ : std_logic;
signal \N__26161\ : std_logic;
signal \N__26156\ : std_logic;
signal \N__26155\ : std_logic;
signal \N__26152\ : std_logic;
signal \N__26149\ : std_logic;
signal \N__26146\ : std_logic;
signal \N__26139\ : std_logic;
signal \N__26136\ : std_logic;
signal \N__26133\ : std_logic;
signal \N__26130\ : std_logic;
signal \N__26129\ : std_logic;
signal \N__26128\ : std_logic;
signal \N__26127\ : std_logic;
signal \N__26126\ : std_logic;
signal \N__26123\ : std_logic;
signal \N__26114\ : std_logic;
signal \N__26109\ : std_logic;
signal \N__26106\ : std_logic;
signal \N__26103\ : std_logic;
signal \N__26100\ : std_logic;
signal \N__26097\ : std_logic;
signal \N__26094\ : std_logic;
signal \N__26091\ : std_logic;
signal \N__26088\ : std_logic;
signal \N__26085\ : std_logic;
signal \N__26082\ : std_logic;
signal \N__26081\ : std_logic;
signal \N__26078\ : std_logic;
signal \N__26075\ : std_logic;
signal \N__26074\ : std_logic;
signal \N__26073\ : std_logic;
signal \N__26070\ : std_logic;
signal \N__26069\ : std_logic;
signal \N__26068\ : std_logic;
signal \N__26065\ : std_logic;
signal \N__26060\ : std_logic;
signal \N__26057\ : std_logic;
signal \N__26054\ : std_logic;
signal \N__26051\ : std_logic;
signal \N__26046\ : std_logic;
signal \N__26041\ : std_logic;
signal \N__26034\ : std_logic;
signal \N__26033\ : std_logic;
signal \N__26030\ : std_logic;
signal \N__26029\ : std_logic;
signal \N__26026\ : std_logic;
signal \N__26025\ : std_logic;
signal \N__26022\ : std_logic;
signal \N__26017\ : std_logic;
signal \N__26016\ : std_logic;
signal \N__26013\ : std_logic;
signal \N__26010\ : std_logic;
signal \N__26007\ : std_logic;
signal \N__26004\ : std_logic;
signal \N__26001\ : std_logic;
signal \N__25996\ : std_logic;
signal \N__25989\ : std_logic;
signal \N__25986\ : std_logic;
signal \N__25985\ : std_logic;
signal \N__25984\ : std_logic;
signal \N__25979\ : std_logic;
signal \N__25978\ : std_logic;
signal \N__25975\ : std_logic;
signal \N__25974\ : std_logic;
signal \N__25971\ : std_logic;
signal \N__25968\ : std_logic;
signal \N__25965\ : std_logic;
signal \N__25962\ : std_logic;
signal \N__25959\ : std_logic;
signal \N__25954\ : std_logic;
signal \N__25947\ : std_logic;
signal \N__25944\ : std_logic;
signal \N__25941\ : std_logic;
signal \N__25940\ : std_logic;
signal \N__25939\ : std_logic;
signal \N__25938\ : std_logic;
signal \N__25935\ : std_logic;
signal \N__25928\ : std_logic;
signal \N__25927\ : std_logic;
signal \N__25926\ : std_logic;
signal \N__25925\ : std_logic;
signal \N__25922\ : std_logic;
signal \N__25919\ : std_logic;
signal \N__25914\ : std_logic;
signal \N__25911\ : std_logic;
signal \N__25904\ : std_logic;
signal \N__25899\ : std_logic;
signal \N__25898\ : std_logic;
signal \N__25897\ : std_logic;
signal \N__25896\ : std_logic;
signal \N__25895\ : std_logic;
signal \N__25894\ : std_logic;
signal \N__25893\ : std_logic;
signal \N__25890\ : std_logic;
signal \N__25885\ : std_logic;
signal \N__25878\ : std_logic;
signal \N__25875\ : std_logic;
signal \N__25872\ : std_logic;
signal \N__25869\ : std_logic;
signal \N__25866\ : std_logic;
signal \N__25857\ : std_logic;
signal \N__25856\ : std_logic;
signal \N__25855\ : std_logic;
signal \N__25852\ : std_logic;
signal \N__25849\ : std_logic;
signal \N__25846\ : std_logic;
signal \N__25843\ : std_logic;
signal \N__25840\ : std_logic;
signal \N__25837\ : std_logic;
signal \N__25830\ : std_logic;
signal \N__25829\ : std_logic;
signal \N__25828\ : std_logic;
signal \N__25827\ : std_logic;
signal \N__25824\ : std_logic;
signal \N__25819\ : std_logic;
signal \N__25816\ : std_logic;
signal \N__25809\ : std_logic;
signal \N__25808\ : std_logic;
signal \N__25807\ : std_logic;
signal \N__25804\ : std_logic;
signal \N__25801\ : std_logic;
signal \N__25796\ : std_logic;
signal \N__25791\ : std_logic;
signal \N__25788\ : std_logic;
signal \N__25785\ : std_logic;
signal \N__25782\ : std_logic;
signal \N__25779\ : std_logic;
signal \N__25776\ : std_logic;
signal \N__25773\ : std_logic;
signal \N__25770\ : std_logic;
signal \N__25769\ : std_logic;
signal \N__25766\ : std_logic;
signal \N__25761\ : std_logic;
signal \N__25758\ : std_logic;
signal \N__25757\ : std_logic;
signal \N__25756\ : std_logic;
signal \N__25753\ : std_logic;
signal \N__25750\ : std_logic;
signal \N__25747\ : std_logic;
signal \N__25744\ : std_logic;
signal \N__25737\ : std_logic;
signal \N__25734\ : std_logic;
signal \N__25731\ : std_logic;
signal \N__25730\ : std_logic;
signal \N__25727\ : std_logic;
signal \N__25724\ : std_logic;
signal \N__25721\ : std_logic;
signal \N__25718\ : std_logic;
signal \N__25713\ : std_logic;
signal \N__25710\ : std_logic;
signal \N__25707\ : std_logic;
signal \N__25704\ : std_logic;
signal \N__25701\ : std_logic;
signal \N__25698\ : std_logic;
signal \N__25695\ : std_logic;
signal \N__25694\ : std_logic;
signal \N__25691\ : std_logic;
signal \N__25688\ : std_logic;
signal \N__25685\ : std_logic;
signal \N__25680\ : std_logic;
signal \N__25677\ : std_logic;
signal \N__25676\ : std_logic;
signal \N__25671\ : std_logic;
signal \N__25668\ : std_logic;
signal \N__25665\ : std_logic;
signal \N__25664\ : std_logic;
signal \N__25661\ : std_logic;
signal \N__25658\ : std_logic;
signal \N__25657\ : std_logic;
signal \N__25654\ : std_logic;
signal \N__25651\ : std_logic;
signal \N__25648\ : std_logic;
signal \N__25641\ : std_logic;
signal \N__25638\ : std_logic;
signal \N__25635\ : std_logic;
signal \N__25632\ : std_logic;
signal \N__25629\ : std_logic;
signal \N__25626\ : std_logic;
signal \N__25623\ : std_logic;
signal \N__25620\ : std_logic;
signal \N__25617\ : std_logic;
signal \N__25614\ : std_logic;
signal \N__25611\ : std_logic;
signal \N__25610\ : std_logic;
signal \N__25607\ : std_logic;
signal \N__25604\ : std_logic;
signal \N__25599\ : std_logic;
signal \N__25596\ : std_logic;
signal \N__25595\ : std_logic;
signal \N__25594\ : std_logic;
signal \N__25589\ : std_logic;
signal \N__25586\ : std_logic;
signal \N__25581\ : std_logic;
signal \N__25580\ : std_logic;
signal \N__25579\ : std_logic;
signal \N__25576\ : std_logic;
signal \N__25571\ : std_logic;
signal \N__25568\ : std_logic;
signal \N__25563\ : std_logic;
signal \N__25562\ : std_logic;
signal \N__25561\ : std_logic;
signal \N__25560\ : std_logic;
signal \N__25559\ : std_logic;
signal \N__25554\ : std_logic;
signal \N__25551\ : std_logic;
signal \N__25546\ : std_logic;
signal \N__25539\ : std_logic;
signal \N__25536\ : std_logic;
signal \N__25535\ : std_logic;
signal \N__25532\ : std_logic;
signal \N__25529\ : std_logic;
signal \N__25524\ : std_logic;
signal \N__25523\ : std_logic;
signal \N__25522\ : std_logic;
signal \N__25519\ : std_logic;
signal \N__25516\ : std_logic;
signal \N__25515\ : std_logic;
signal \N__25514\ : std_logic;
signal \N__25511\ : std_logic;
signal \N__25506\ : std_logic;
signal \N__25503\ : std_logic;
signal \N__25500\ : std_logic;
signal \N__25497\ : std_logic;
signal \N__25494\ : std_logic;
signal \N__25491\ : std_logic;
signal \N__25482\ : std_logic;
signal \N__25481\ : std_logic;
signal \N__25478\ : std_logic;
signal \N__25477\ : std_logic;
signal \N__25476\ : std_logic;
signal \N__25473\ : std_logic;
signal \N__25470\ : std_logic;
signal \N__25467\ : std_logic;
signal \N__25464\ : std_logic;
signal \N__25463\ : std_logic;
signal \N__25460\ : std_logic;
signal \N__25455\ : std_logic;
signal \N__25452\ : std_logic;
signal \N__25449\ : std_logic;
signal \N__25446\ : std_logic;
signal \N__25441\ : std_logic;
signal \N__25434\ : std_logic;
signal \N__25431\ : std_logic;
signal \N__25428\ : std_logic;
signal \N__25425\ : std_logic;
signal \N__25422\ : std_logic;
signal \N__25419\ : std_logic;
signal \N__25416\ : std_logic;
signal \N__25415\ : std_logic;
signal \N__25412\ : std_logic;
signal \N__25411\ : std_logic;
signal \N__25408\ : std_logic;
signal \N__25403\ : std_logic;
signal \N__25400\ : std_logic;
signal \N__25395\ : std_logic;
signal \N__25394\ : std_logic;
signal \N__25391\ : std_logic;
signal \N__25388\ : std_logic;
signal \N__25385\ : std_logic;
signal \N__25380\ : std_logic;
signal \N__25377\ : std_logic;
signal \N__25374\ : std_logic;
signal \N__25371\ : std_logic;
signal \N__25368\ : std_logic;
signal \N__25367\ : std_logic;
signal \N__25366\ : std_logic;
signal \N__25365\ : std_logic;
signal \N__25362\ : std_logic;
signal \N__25359\ : std_logic;
signal \N__25358\ : std_logic;
signal \N__25357\ : std_logic;
signal \N__25352\ : std_logic;
signal \N__25345\ : std_logic;
signal \N__25342\ : std_logic;
signal \N__25335\ : std_logic;
signal \N__25332\ : std_logic;
signal \N__25329\ : std_logic;
signal \N__25328\ : std_logic;
signal \N__25327\ : std_logic;
signal \N__25326\ : std_logic;
signal \N__25323\ : std_logic;
signal \N__25320\ : std_logic;
signal \N__25317\ : std_logic;
signal \N__25314\ : std_logic;
signal \N__25313\ : std_logic;
signal \N__25310\ : std_logic;
signal \N__25307\ : std_logic;
signal \N__25302\ : std_logic;
signal \N__25299\ : std_logic;
signal \N__25296\ : std_logic;
signal \N__25291\ : std_logic;
signal \N__25284\ : std_logic;
signal \N__25281\ : std_logic;
signal \N__25278\ : std_logic;
signal \N__25275\ : std_logic;
signal \N__25272\ : std_logic;
signal \N__25269\ : std_logic;
signal \N__25268\ : std_logic;
signal \N__25265\ : std_logic;
signal \N__25262\ : std_logic;
signal \N__25259\ : std_logic;
signal \N__25258\ : std_logic;
signal \N__25255\ : std_logic;
signal \N__25252\ : std_logic;
signal \N__25249\ : std_logic;
signal \N__25246\ : std_logic;
signal \N__25239\ : std_logic;
signal \N__25238\ : std_logic;
signal \N__25237\ : std_logic;
signal \N__25236\ : std_logic;
signal \N__25235\ : std_logic;
signal \N__25234\ : std_logic;
signal \N__25233\ : std_logic;
signal \N__25232\ : std_logic;
signal \N__25231\ : std_logic;
signal \N__25230\ : std_logic;
signal \N__25229\ : std_logic;
signal \N__25228\ : std_logic;
signal \N__25227\ : std_logic;
signal \N__25226\ : std_logic;
signal \N__25225\ : std_logic;
signal \N__25224\ : std_logic;
signal \N__25221\ : std_logic;
signal \N__25220\ : std_logic;
signal \N__25219\ : std_logic;
signal \N__25218\ : std_logic;
signal \N__25217\ : std_logic;
signal \N__25216\ : std_logic;
signal \N__25213\ : std_logic;
signal \N__25208\ : std_logic;
signal \N__25201\ : std_logic;
signal \N__25194\ : std_logic;
signal \N__25185\ : std_logic;
signal \N__25180\ : std_logic;
signal \N__25179\ : std_logic;
signal \N__25178\ : std_logic;
signal \N__25177\ : std_logic;
signal \N__25176\ : std_logic;
signal \N__25173\ : std_logic;
signal \N__25170\ : std_logic;
signal \N__25167\ : std_logic;
signal \N__25166\ : std_logic;
signal \N__25165\ : std_logic;
signal \N__25158\ : std_logic;
signal \N__25157\ : std_logic;
signal \N__25156\ : std_logic;
signal \N__25155\ : std_logic;
signal \N__25152\ : std_logic;
signal \N__25143\ : std_logic;
signal \N__25140\ : std_logic;
signal \N__25131\ : std_logic;
signal \N__25126\ : std_logic;
signal \N__25123\ : std_logic;
signal \N__25118\ : std_logic;
signal \N__25117\ : std_logic;
signal \N__25116\ : std_logic;
signal \N__25113\ : std_logic;
signal \N__25110\ : std_logic;
signal \N__25107\ : std_logic;
signal \N__25104\ : std_logic;
signal \N__25095\ : std_logic;
signal \N__25088\ : std_logic;
signal \N__25083\ : std_logic;
signal \N__25068\ : std_logic;
signal \N__25067\ : std_logic;
signal \N__25064\ : std_logic;
signal \N__25061\ : std_logic;
signal \N__25058\ : std_logic;
signal \N__25053\ : std_logic;
signal \N__25050\ : std_logic;
signal \N__25047\ : std_logic;
signal \N__25044\ : std_logic;
signal \N__25041\ : std_logic;
signal \N__25038\ : std_logic;
signal \N__25035\ : std_logic;
signal \N__25032\ : std_logic;
signal \N__25029\ : std_logic;
signal \N__25026\ : std_logic;
signal \N__25025\ : std_logic;
signal \N__25024\ : std_logic;
signal \N__25023\ : std_logic;
signal \N__25020\ : std_logic;
signal \N__25017\ : std_logic;
signal \N__25010\ : std_logic;
signal \N__25007\ : std_logic;
signal \N__25002\ : std_logic;
signal \N__24999\ : std_logic;
signal \N__24996\ : std_logic;
signal \N__24993\ : std_logic;
signal \N__24990\ : std_logic;
signal \N__24987\ : std_logic;
signal \N__24984\ : std_logic;
signal \N__24983\ : std_logic;
signal \N__24980\ : std_logic;
signal \N__24979\ : std_logic;
signal \N__24978\ : std_logic;
signal \N__24975\ : std_logic;
signal \N__24972\ : std_logic;
signal \N__24965\ : std_logic;
signal \N__24962\ : std_logic;
signal \N__24957\ : std_logic;
signal \N__24956\ : std_logic;
signal \N__24955\ : std_logic;
signal \N__24952\ : std_logic;
signal \N__24949\ : std_logic;
signal \N__24946\ : std_logic;
signal \N__24945\ : std_logic;
signal \N__24944\ : std_logic;
signal \N__24943\ : std_logic;
signal \N__24942\ : std_logic;
signal \N__24941\ : std_logic;
signal \N__24940\ : std_logic;
signal \N__24937\ : std_logic;
signal \N__24934\ : std_logic;
signal \N__24933\ : std_logic;
signal \N__24930\ : std_logic;
signal \N__24927\ : std_logic;
signal \N__24920\ : std_logic;
signal \N__24915\ : std_logic;
signal \N__24912\ : std_logic;
signal \N__24909\ : std_logic;
signal \N__24908\ : std_logic;
signal \N__24907\ : std_logic;
signal \N__24904\ : std_logic;
signal \N__24895\ : std_logic;
signal \N__24892\ : std_logic;
signal \N__24889\ : std_logic;
signal \N__24884\ : std_logic;
signal \N__24873\ : std_logic;
signal \N__24870\ : std_logic;
signal \N__24867\ : std_logic;
signal \N__24864\ : std_logic;
signal \N__24861\ : std_logic;
signal \N__24858\ : std_logic;
signal \N__24855\ : std_logic;
signal \N__24852\ : std_logic;
signal \N__24849\ : std_logic;
signal \N__24846\ : std_logic;
signal \N__24843\ : std_logic;
signal \N__24842\ : std_logic;
signal \N__24839\ : std_logic;
signal \N__24836\ : std_logic;
signal \N__24833\ : std_logic;
signal \N__24828\ : std_logic;
signal \N__24825\ : std_logic;
signal \N__24822\ : std_logic;
signal \N__24819\ : std_logic;
signal \N__24816\ : std_logic;
signal \N__24813\ : std_logic;
signal \N__24810\ : std_logic;
signal \N__24807\ : std_logic;
signal \N__24804\ : std_logic;
signal \N__24801\ : std_logic;
signal \N__24798\ : std_logic;
signal \N__24795\ : std_logic;
signal \N__24792\ : std_logic;
signal \N__24789\ : std_logic;
signal \N__24786\ : std_logic;
signal \N__24783\ : std_logic;
signal \N__24782\ : std_logic;
signal \N__24779\ : std_logic;
signal \N__24776\ : std_logic;
signal \N__24771\ : std_logic;
signal \N__24768\ : std_logic;
signal \N__24765\ : std_logic;
signal \N__24764\ : std_logic;
signal \N__24763\ : std_logic;
signal \N__24760\ : std_logic;
signal \N__24757\ : std_logic;
signal \N__24754\ : std_logic;
signal \N__24753\ : std_logic;
signal \N__24750\ : std_logic;
signal \N__24747\ : std_logic;
signal \N__24744\ : std_logic;
signal \N__24743\ : std_logic;
signal \N__24740\ : std_logic;
signal \N__24737\ : std_logic;
signal \N__24734\ : std_logic;
signal \N__24731\ : std_logic;
signal \N__24728\ : std_logic;
signal \N__24717\ : std_logic;
signal \N__24714\ : std_logic;
signal \N__24711\ : std_logic;
signal \N__24708\ : std_logic;
signal \N__24705\ : std_logic;
signal \N__24702\ : std_logic;
signal \N__24699\ : std_logic;
signal \N__24696\ : std_logic;
signal \N__24695\ : std_logic;
signal \N__24694\ : std_logic;
signal \N__24691\ : std_logic;
signal \N__24688\ : std_logic;
signal \N__24685\ : std_logic;
signal \N__24678\ : std_logic;
signal \N__24675\ : std_logic;
signal \N__24674\ : std_logic;
signal \N__24673\ : std_logic;
signal \N__24670\ : std_logic;
signal \N__24667\ : std_logic;
signal \N__24664\ : std_logic;
signal \N__24661\ : std_logic;
signal \N__24654\ : std_logic;
signal \N__24651\ : std_logic;
signal \N__24648\ : std_logic;
signal \N__24647\ : std_logic;
signal \N__24644\ : std_logic;
signal \N__24641\ : std_logic;
signal \N__24640\ : std_logic;
signal \N__24635\ : std_logic;
signal \N__24632\ : std_logic;
signal \N__24627\ : std_logic;
signal \N__24626\ : std_logic;
signal \N__24625\ : std_logic;
signal \N__24622\ : std_logic;
signal \N__24619\ : std_logic;
signal \N__24616\ : std_logic;
signal \N__24613\ : std_logic;
signal \N__24606\ : std_logic;
signal \N__24603\ : std_logic;
signal \N__24602\ : std_logic;
signal \N__24601\ : std_logic;
signal \N__24598\ : std_logic;
signal \N__24595\ : std_logic;
signal \N__24592\ : std_logic;
signal \N__24589\ : std_logic;
signal \N__24582\ : std_logic;
signal \N__24581\ : std_logic;
signal \N__24580\ : std_logic;
signal \N__24577\ : std_logic;
signal \N__24574\ : std_logic;
signal \N__24571\ : std_logic;
signal \N__24568\ : std_logic;
signal \N__24561\ : std_logic;
signal \N__24560\ : std_logic;
signal \N__24559\ : std_logic;
signal \N__24556\ : std_logic;
signal \N__24553\ : std_logic;
signal \N__24550\ : std_logic;
signal \N__24543\ : std_logic;
signal \N__24540\ : std_logic;
signal \N__24539\ : std_logic;
signal \N__24538\ : std_logic;
signal \N__24535\ : std_logic;
signal \N__24532\ : std_logic;
signal \N__24529\ : std_logic;
signal \N__24522\ : std_logic;
signal \N__24519\ : std_logic;
signal \N__24516\ : std_logic;
signal \N__24515\ : std_logic;
signal \N__24514\ : std_logic;
signal \N__24513\ : std_logic;
signal \N__24512\ : std_logic;
signal \N__24511\ : std_logic;
signal \N__24510\ : std_logic;
signal \N__24509\ : std_logic;
signal \N__24508\ : std_logic;
signal \N__24507\ : std_logic;
signal \N__24506\ : std_logic;
signal \N__24505\ : std_logic;
signal \N__24504\ : std_logic;
signal \N__24501\ : std_logic;
signal \N__24498\ : std_logic;
signal \N__24495\ : std_logic;
signal \N__24492\ : std_logic;
signal \N__24489\ : std_logic;
signal \N__24486\ : std_logic;
signal \N__24483\ : std_logic;
signal \N__24480\ : std_logic;
signal \N__24477\ : std_logic;
signal \N__24474\ : std_logic;
signal \N__24471\ : std_logic;
signal \N__24468\ : std_logic;
signal \N__24465\ : std_logic;
signal \N__24458\ : std_logic;
signal \N__24451\ : std_logic;
signal \N__24450\ : std_logic;
signal \N__24443\ : std_logic;
signal \N__24434\ : std_logic;
signal \N__24429\ : std_logic;
signal \N__24426\ : std_logic;
signal \N__24417\ : std_logic;
signal \N__24416\ : std_logic;
signal \N__24413\ : std_logic;
signal \N__24410\ : std_logic;
signal \N__24407\ : std_logic;
signal \N__24404\ : std_logic;
signal \N__24399\ : std_logic;
signal \N__24396\ : std_logic;
signal \N__24393\ : std_logic;
signal \N__24390\ : std_logic;
signal \N__24387\ : std_logic;
signal \N__24384\ : std_logic;
signal \N__24383\ : std_logic;
signal \N__24380\ : std_logic;
signal \N__24377\ : std_logic;
signal \N__24372\ : std_logic;
signal \N__24371\ : std_logic;
signal \N__24370\ : std_logic;
signal \N__24367\ : std_logic;
signal \N__24364\ : std_logic;
signal \N__24361\ : std_logic;
signal \N__24358\ : std_logic;
signal \N__24351\ : std_logic;
signal \N__24348\ : std_logic;
signal \N__24345\ : std_logic;
signal \N__24344\ : std_logic;
signal \N__24343\ : std_logic;
signal \N__24340\ : std_logic;
signal \N__24337\ : std_logic;
signal \N__24334\ : std_logic;
signal \N__24331\ : std_logic;
signal \N__24324\ : std_logic;
signal \N__24321\ : std_logic;
signal \N__24320\ : std_logic;
signal \N__24319\ : std_logic;
signal \N__24316\ : std_logic;
signal \N__24313\ : std_logic;
signal \N__24310\ : std_logic;
signal \N__24307\ : std_logic;
signal \N__24300\ : std_logic;
signal \N__24297\ : std_logic;
signal \N__24294\ : std_logic;
signal \N__24291\ : std_logic;
signal \N__24288\ : std_logic;
signal \N__24287\ : std_logic;
signal \N__24286\ : std_logic;
signal \N__24283\ : std_logic;
signal \N__24280\ : std_logic;
signal \N__24277\ : std_logic;
signal \N__24270\ : std_logic;
signal \N__24267\ : std_logic;
signal \N__24264\ : std_logic;
signal \N__24261\ : std_logic;
signal \N__24258\ : std_logic;
signal \N__24255\ : std_logic;
signal \N__24254\ : std_logic;
signal \N__24251\ : std_logic;
signal \N__24250\ : std_logic;
signal \N__24247\ : std_logic;
signal \N__24244\ : std_logic;
signal \N__24241\ : std_logic;
signal \N__24240\ : std_logic;
signal \N__24237\ : std_logic;
signal \N__24232\ : std_logic;
signal \N__24229\ : std_logic;
signal \N__24226\ : std_logic;
signal \N__24223\ : std_logic;
signal \N__24220\ : std_logic;
signal \N__24213\ : std_logic;
signal \N__24212\ : std_logic;
signal \N__24209\ : std_logic;
signal \N__24208\ : std_logic;
signal \N__24205\ : std_logic;
signal \N__24204\ : std_logic;
signal \N__24201\ : std_logic;
signal \N__24198\ : std_logic;
signal \N__24195\ : std_logic;
signal \N__24192\ : std_logic;
signal \N__24189\ : std_logic;
signal \N__24184\ : std_logic;
signal \N__24181\ : std_logic;
signal \N__24178\ : std_logic;
signal \N__24175\ : std_logic;
signal \N__24168\ : std_logic;
signal \N__24165\ : std_logic;
signal \N__24162\ : std_logic;
signal \N__24159\ : std_logic;
signal \N__24158\ : std_logic;
signal \N__24157\ : std_logic;
signal \N__24154\ : std_logic;
signal \N__24151\ : std_logic;
signal \N__24148\ : std_logic;
signal \N__24141\ : std_logic;
signal \N__24138\ : std_logic;
signal \N__24135\ : std_logic;
signal \N__24134\ : std_logic;
signal \N__24133\ : std_logic;
signal \N__24130\ : std_logic;
signal \N__24127\ : std_logic;
signal \N__24124\ : std_logic;
signal \N__24121\ : std_logic;
signal \N__24114\ : std_logic;
signal \N__24111\ : std_logic;
signal \N__24108\ : std_logic;
signal \N__24105\ : std_logic;
signal \N__24104\ : std_logic;
signal \N__24103\ : std_logic;
signal \N__24100\ : std_logic;
signal \N__24097\ : std_logic;
signal \N__24096\ : std_logic;
signal \N__24093\ : std_logic;
signal \N__24092\ : std_logic;
signal \N__24087\ : std_logic;
signal \N__24084\ : std_logic;
signal \N__24081\ : std_logic;
signal \N__24078\ : std_logic;
signal \N__24075\ : std_logic;
signal \N__24072\ : std_logic;
signal \N__24069\ : std_logic;
signal \N__24060\ : std_logic;
signal \N__24057\ : std_logic;
signal \N__24054\ : std_logic;
signal \N__24053\ : std_logic;
signal \N__24052\ : std_logic;
signal \N__24049\ : std_logic;
signal \N__24048\ : std_logic;
signal \N__24045\ : std_logic;
signal \N__24044\ : std_logic;
signal \N__24041\ : std_logic;
signal \N__24038\ : std_logic;
signal \N__24035\ : std_logic;
signal \N__24032\ : std_logic;
signal \N__24029\ : std_logic;
signal \N__24024\ : std_logic;
signal \N__24021\ : std_logic;
signal \N__24018\ : std_logic;
signal \N__24013\ : std_logic;
signal \N__24010\ : std_logic;
signal \N__24003\ : std_logic;
signal \N__24000\ : std_logic;
signal \N__23999\ : std_logic;
signal \N__23998\ : std_logic;
signal \N__23997\ : std_logic;
signal \N__23994\ : std_logic;
signal \N__23991\ : std_logic;
signal \N__23988\ : std_logic;
signal \N__23987\ : std_logic;
signal \N__23984\ : std_logic;
signal \N__23981\ : std_logic;
signal \N__23976\ : std_logic;
signal \N__23973\ : std_logic;
signal \N__23970\ : std_logic;
signal \N__23967\ : std_logic;
signal \N__23964\ : std_logic;
signal \N__23955\ : std_logic;
signal \N__23952\ : std_logic;
signal \N__23951\ : std_logic;
signal \N__23950\ : std_logic;
signal \N__23947\ : std_logic;
signal \N__23944\ : std_logic;
signal \N__23941\ : std_logic;
signal \N__23940\ : std_logic;
signal \N__23939\ : std_logic;
signal \N__23936\ : std_logic;
signal \N__23933\ : std_logic;
signal \N__23930\ : std_logic;
signal \N__23927\ : std_logic;
signal \N__23924\ : std_logic;
signal \N__23921\ : std_logic;
signal \N__23918\ : std_logic;
signal \N__23915\ : std_logic;
signal \N__23912\ : std_logic;
signal \N__23901\ : std_logic;
signal \N__23898\ : std_logic;
signal \N__23895\ : std_logic;
signal \N__23892\ : std_logic;
signal \N__23889\ : std_logic;
signal \N__23886\ : std_logic;
signal \N__23883\ : std_logic;
signal \N__23880\ : std_logic;
signal \N__23877\ : std_logic;
signal \N__23874\ : std_logic;
signal \N__23871\ : std_logic;
signal \N__23868\ : std_logic;
signal \N__23867\ : std_logic;
signal \N__23866\ : std_logic;
signal \N__23865\ : std_logic;
signal \N__23864\ : std_logic;
signal \N__23861\ : std_logic;
signal \N__23858\ : std_logic;
signal \N__23855\ : std_logic;
signal \N__23852\ : std_logic;
signal \N__23849\ : std_logic;
signal \N__23844\ : std_logic;
signal \N__23841\ : std_logic;
signal \N__23832\ : std_logic;
signal \N__23829\ : std_logic;
signal \N__23828\ : std_logic;
signal \N__23827\ : std_logic;
signal \N__23826\ : std_logic;
signal \N__23823\ : std_logic;
signal \N__23820\ : std_logic;
signal \N__23817\ : std_logic;
signal \N__23814\ : std_logic;
signal \N__23813\ : std_logic;
signal \N__23810\ : std_logic;
signal \N__23805\ : std_logic;
signal \N__23802\ : std_logic;
signal \N__23799\ : std_logic;
signal \N__23796\ : std_logic;
signal \N__23791\ : std_logic;
signal \N__23784\ : std_logic;
signal \N__23781\ : std_logic;
signal \N__23778\ : std_logic;
signal \N__23775\ : std_logic;
signal \N__23772\ : std_logic;
signal \N__23769\ : std_logic;
signal \N__23766\ : std_logic;
signal \N__23763\ : std_logic;
signal \N__23760\ : std_logic;
signal \N__23757\ : std_logic;
signal \N__23754\ : std_logic;
signal \N__23751\ : std_logic;
signal \N__23748\ : std_logic;
signal \N__23745\ : std_logic;
signal \N__23742\ : std_logic;
signal \N__23739\ : std_logic;
signal \N__23736\ : std_logic;
signal \N__23733\ : std_logic;
signal \N__23730\ : std_logic;
signal \N__23727\ : std_logic;
signal \N__23724\ : std_logic;
signal \N__23721\ : std_logic;
signal \N__23718\ : std_logic;
signal \N__23715\ : std_logic;
signal \N__23712\ : std_logic;
signal \N__23711\ : std_logic;
signal \N__23708\ : std_logic;
signal \N__23705\ : std_logic;
signal \N__23702\ : std_logic;
signal \N__23697\ : std_logic;
signal \N__23694\ : std_logic;
signal \N__23691\ : std_logic;
signal \N__23688\ : std_logic;
signal \N__23685\ : std_logic;
signal \N__23682\ : std_logic;
signal \N__23679\ : std_logic;
signal \N__23676\ : std_logic;
signal \N__23673\ : std_logic;
signal \N__23670\ : std_logic;
signal \N__23667\ : std_logic;
signal \N__23664\ : std_logic;
signal \N__23661\ : std_logic;
signal \N__23658\ : std_logic;
signal \N__23655\ : std_logic;
signal \N__23652\ : std_logic;
signal \N__23651\ : std_logic;
signal \N__23648\ : std_logic;
signal \N__23645\ : std_logic;
signal \N__23642\ : std_logic;
signal \N__23639\ : std_logic;
signal \N__23634\ : std_logic;
signal \N__23631\ : std_logic;
signal \N__23628\ : std_logic;
signal \N__23627\ : std_logic;
signal \N__23624\ : std_logic;
signal \N__23623\ : std_logic;
signal \N__23620\ : std_logic;
signal \N__23617\ : std_logic;
signal \N__23614\ : std_logic;
signal \N__23611\ : std_logic;
signal \N__23604\ : std_logic;
signal \N__23603\ : std_logic;
signal \N__23600\ : std_logic;
signal \N__23597\ : std_logic;
signal \N__23594\ : std_logic;
signal \N__23591\ : std_logic;
signal \N__23586\ : std_logic;
signal \N__23583\ : std_logic;
signal \N__23582\ : std_logic;
signal \N__23581\ : std_logic;
signal \N__23578\ : std_logic;
signal \N__23575\ : std_logic;
signal \N__23572\ : std_logic;
signal \N__23569\ : std_logic;
signal \N__23562\ : std_logic;
signal \N__23559\ : std_logic;
signal \N__23558\ : std_logic;
signal \N__23555\ : std_logic;
signal \N__23554\ : std_logic;
signal \N__23553\ : std_logic;
signal \N__23552\ : std_logic;
signal \N__23549\ : std_logic;
signal \N__23548\ : std_logic;
signal \N__23545\ : std_logic;
signal \N__23542\ : std_logic;
signal \N__23533\ : std_logic;
signal \N__23526\ : std_logic;
signal \N__23523\ : std_logic;
signal \N__23520\ : std_logic;
signal \N__23517\ : std_logic;
signal \N__23516\ : std_logic;
signal \N__23513\ : std_logic;
signal \N__23510\ : std_logic;
signal \N__23509\ : std_logic;
signal \N__23506\ : std_logic;
signal \N__23503\ : std_logic;
signal \N__23500\ : std_logic;
signal \N__23493\ : std_logic;
signal \N__23492\ : std_logic;
signal \N__23489\ : std_logic;
signal \N__23486\ : std_logic;
signal \N__23483\ : std_logic;
signal \N__23482\ : std_logic;
signal \N__23481\ : std_logic;
signal \N__23480\ : std_logic;
signal \N__23479\ : std_logic;
signal \N__23478\ : std_logic;
signal \N__23477\ : std_logic;
signal \N__23476\ : std_logic;
signal \N__23475\ : std_logic;
signal \N__23474\ : std_logic;
signal \N__23473\ : std_logic;
signal \N__23472\ : std_logic;
signal \N__23471\ : std_logic;
signal \N__23470\ : std_logic;
signal \N__23469\ : std_logic;
signal \N__23466\ : std_logic;
signal \N__23463\ : std_logic;
signal \N__23458\ : std_logic;
signal \N__23453\ : std_logic;
signal \N__23450\ : std_logic;
signal \N__23445\ : std_logic;
signal \N__23440\ : std_logic;
signal \N__23433\ : std_logic;
signal \N__23428\ : std_logic;
signal \N__23409\ : std_logic;
signal \N__23406\ : std_logic;
signal \N__23403\ : std_logic;
signal \N__23400\ : std_logic;
signal \N__23397\ : std_logic;
signal \N__23394\ : std_logic;
signal \N__23391\ : std_logic;
signal \N__23388\ : std_logic;
signal \N__23385\ : std_logic;
signal \N__23382\ : std_logic;
signal \N__23379\ : std_logic;
signal \N__23376\ : std_logic;
signal \N__23373\ : std_logic;
signal \N__23370\ : std_logic;
signal \N__23367\ : std_logic;
signal \N__23364\ : std_logic;
signal \N__23361\ : std_logic;
signal \N__23358\ : std_logic;
signal \N__23355\ : std_logic;
signal \N__23352\ : std_logic;
signal \N__23349\ : std_logic;
signal \N__23348\ : std_logic;
signal \N__23345\ : std_logic;
signal \N__23342\ : std_logic;
signal \N__23339\ : std_logic;
signal \N__23336\ : std_logic;
signal \N__23331\ : std_logic;
signal \N__23328\ : std_logic;
signal \N__23327\ : std_logic;
signal \N__23324\ : std_logic;
signal \N__23323\ : std_logic;
signal \N__23320\ : std_logic;
signal \N__23317\ : std_logic;
signal \N__23314\ : std_logic;
signal \N__23311\ : std_logic;
signal \N__23304\ : std_logic;
signal \N__23303\ : std_logic;
signal \N__23298\ : std_logic;
signal \N__23295\ : std_logic;
signal \N__23292\ : std_logic;
signal \N__23289\ : std_logic;
signal \N__23286\ : std_logic;
signal \N__23283\ : std_logic;
signal \N__23280\ : std_logic;
signal \N__23277\ : std_logic;
signal \N__23274\ : std_logic;
signal \N__23271\ : std_logic;
signal \N__23268\ : std_logic;
signal \N__23265\ : std_logic;
signal \N__23262\ : std_logic;
signal \N__23261\ : std_logic;
signal \N__23260\ : std_logic;
signal \N__23259\ : std_logic;
signal \N__23256\ : std_logic;
signal \N__23251\ : std_logic;
signal \N__23250\ : std_logic;
signal \N__23249\ : std_logic;
signal \N__23248\ : std_logic;
signal \N__23245\ : std_logic;
signal \N__23244\ : std_logic;
signal \N__23243\ : std_logic;
signal \N__23240\ : std_logic;
signal \N__23237\ : std_logic;
signal \N__23234\ : std_logic;
signal \N__23231\ : std_logic;
signal \N__23222\ : std_logic;
signal \N__23219\ : std_logic;
signal \N__23216\ : std_logic;
signal \N__23205\ : std_logic;
signal \N__23204\ : std_logic;
signal \N__23203\ : std_logic;
signal \N__23200\ : std_logic;
signal \N__23197\ : std_logic;
signal \N__23194\ : std_logic;
signal \N__23187\ : std_logic;
signal \N__23184\ : std_logic;
signal \N__23183\ : std_logic;
signal \N__23182\ : std_logic;
signal \N__23181\ : std_logic;
signal \N__23178\ : std_logic;
signal \N__23175\ : std_logic;
signal \N__23170\ : std_logic;
signal \N__23169\ : std_logic;
signal \N__23168\ : std_logic;
signal \N__23161\ : std_logic;
signal \N__23158\ : std_logic;
signal \N__23155\ : std_logic;
signal \N__23152\ : std_logic;
signal \N__23149\ : std_logic;
signal \N__23142\ : std_logic;
signal \N__23141\ : std_logic;
signal \N__23138\ : std_logic;
signal \N__23135\ : std_logic;
signal \N__23130\ : std_logic;
signal \N__23127\ : std_logic;
signal \N__23124\ : std_logic;
signal \N__23121\ : std_logic;
signal \N__23118\ : std_logic;
signal \N__23115\ : std_logic;
signal \N__23112\ : std_logic;
signal \N__23111\ : std_logic;
signal \N__23110\ : std_logic;
signal \N__23107\ : std_logic;
signal \N__23104\ : std_logic;
signal \N__23101\ : std_logic;
signal \N__23094\ : std_logic;
signal \N__23091\ : std_logic;
signal \N__23088\ : std_logic;
signal \N__23087\ : std_logic;
signal \N__23086\ : std_logic;
signal \N__23083\ : std_logic;
signal \N__23080\ : std_logic;
signal \N__23077\ : std_logic;
signal \N__23074\ : std_logic;
signal \N__23069\ : std_logic;
signal \N__23064\ : std_logic;
signal \N__23063\ : std_logic;
signal \N__23062\ : std_logic;
signal \N__23059\ : std_logic;
signal \N__23056\ : std_logic;
signal \N__23053\ : std_logic;
signal \N__23046\ : std_logic;
signal \N__23043\ : std_logic;
signal \N__23042\ : std_logic;
signal \N__23041\ : std_logic;
signal \N__23038\ : std_logic;
signal \N__23035\ : std_logic;
signal \N__23032\ : std_logic;
signal \N__23029\ : std_logic;
signal \N__23026\ : std_logic;
signal \N__23023\ : std_logic;
signal \N__23016\ : std_logic;
signal \N__23013\ : std_logic;
signal \N__23010\ : std_logic;
signal \N__23007\ : std_logic;
signal \N__23004\ : std_logic;
signal \N__23003\ : std_logic;
signal \N__23002\ : std_logic;
signal \N__23001\ : std_logic;
signal \N__23000\ : std_logic;
signal \N__22999\ : std_logic;
signal \N__22998\ : std_logic;
signal \N__22997\ : std_logic;
signal \N__22996\ : std_logic;
signal \N__22995\ : std_logic;
signal \N__22994\ : std_logic;
signal \N__22993\ : std_logic;
signal \N__22990\ : std_logic;
signal \N__22987\ : std_logic;
signal \N__22984\ : std_logic;
signal \N__22981\ : std_logic;
signal \N__22978\ : std_logic;
signal \N__22975\ : std_logic;
signal \N__22972\ : std_logic;
signal \N__22969\ : std_logic;
signal \N__22966\ : std_logic;
signal \N__22963\ : std_logic;
signal \N__22960\ : std_logic;
signal \N__22957\ : std_logic;
signal \N__22950\ : std_logic;
signal \N__22943\ : std_logic;
signal \N__22936\ : std_logic;
signal \N__22929\ : std_logic;
signal \N__22924\ : std_logic;
signal \N__22917\ : std_logic;
signal \N__22914\ : std_logic;
signal \N__22913\ : std_logic;
signal \N__22910\ : std_logic;
signal \N__22907\ : std_logic;
signal \N__22904\ : std_logic;
signal \N__22901\ : std_logic;
signal \N__22896\ : std_logic;
signal \N__22893\ : std_logic;
signal \N__22890\ : std_logic;
signal \N__22887\ : std_logic;
signal \N__22884\ : std_logic;
signal \N__22881\ : std_logic;
signal \N__22878\ : std_logic;
signal \N__22875\ : std_logic;
signal \N__22872\ : std_logic;
signal \N__22869\ : std_logic;
signal \N__22868\ : std_logic;
signal \N__22865\ : std_logic;
signal \N__22862\ : std_logic;
signal \N__22857\ : std_logic;
signal \N__22856\ : std_logic;
signal \N__22855\ : std_logic;
signal \N__22854\ : std_logic;
signal \N__22849\ : std_logic;
signal \N__22846\ : std_logic;
signal \N__22843\ : std_logic;
signal \N__22836\ : std_logic;
signal \N__22833\ : std_logic;
signal \N__22830\ : std_logic;
signal \N__22829\ : std_logic;
signal \N__22826\ : std_logic;
signal \N__22823\ : std_logic;
signal \N__22822\ : std_logic;
signal \N__22817\ : std_logic;
signal \N__22814\ : std_logic;
signal \N__22809\ : std_logic;
signal \N__22806\ : std_logic;
signal \N__22803\ : std_logic;
signal \N__22800\ : std_logic;
signal \N__22797\ : std_logic;
signal \N__22794\ : std_logic;
signal \N__22791\ : std_logic;
signal \N__22788\ : std_logic;
signal \N__22787\ : std_logic;
signal \N__22786\ : std_logic;
signal \N__22783\ : std_logic;
signal \N__22780\ : std_logic;
signal \N__22777\ : std_logic;
signal \N__22772\ : std_logic;
signal \N__22769\ : std_logic;
signal \N__22764\ : std_logic;
signal \N__22763\ : std_logic;
signal \N__22762\ : std_logic;
signal \N__22759\ : std_logic;
signal \N__22756\ : std_logic;
signal \N__22753\ : std_logic;
signal \N__22746\ : std_logic;
signal \N__22743\ : std_logic;
signal \N__22742\ : std_logic;
signal \N__22741\ : std_logic;
signal \N__22738\ : std_logic;
signal \N__22735\ : std_logic;
signal \N__22732\ : std_logic;
signal \N__22729\ : std_logic;
signal \N__22724\ : std_logic;
signal \N__22721\ : std_logic;
signal \N__22716\ : std_logic;
signal \N__22715\ : std_logic;
signal \N__22714\ : std_logic;
signal \N__22711\ : std_logic;
signal \N__22708\ : std_logic;
signal \N__22705\ : std_logic;
signal \N__22698\ : std_logic;
signal \N__22695\ : std_logic;
signal \N__22692\ : std_logic;
signal \N__22691\ : std_logic;
signal \N__22690\ : std_logic;
signal \N__22687\ : std_logic;
signal \N__22684\ : std_logic;
signal \N__22681\ : std_logic;
signal \N__22676\ : std_logic;
signal \N__22673\ : std_logic;
signal \N__22668\ : std_logic;
signal \N__22665\ : std_logic;
signal \N__22662\ : std_logic;
signal \N__22661\ : std_logic;
signal \N__22658\ : std_logic;
signal \N__22655\ : std_logic;
signal \N__22654\ : std_logic;
signal \N__22649\ : std_logic;
signal \N__22646\ : std_logic;
signal \N__22641\ : std_logic;
signal \N__22638\ : std_logic;
signal \N__22637\ : std_logic;
signal \N__22634\ : std_logic;
signal \N__22631\ : std_logic;
signal \N__22630\ : std_logic;
signal \N__22625\ : std_logic;
signal \N__22622\ : std_logic;
signal \N__22617\ : std_logic;
signal \N__22614\ : std_logic;
signal \N__22611\ : std_logic;
signal \N__22608\ : std_logic;
signal \N__22607\ : std_logic;
signal \N__22606\ : std_logic;
signal \N__22603\ : std_logic;
signal \N__22600\ : std_logic;
signal \N__22597\ : std_logic;
signal \N__22592\ : std_logic;
signal \N__22589\ : std_logic;
signal \N__22584\ : std_logic;
signal \N__22581\ : std_logic;
signal \N__22578\ : std_logic;
signal \N__22577\ : std_logic;
signal \N__22576\ : std_logic;
signal \N__22573\ : std_logic;
signal \N__22570\ : std_logic;
signal \N__22567\ : std_logic;
signal \N__22560\ : std_logic;
signal \N__22557\ : std_logic;
signal \N__22556\ : std_logic;
signal \N__22555\ : std_logic;
signal \N__22552\ : std_logic;
signal \N__22549\ : std_logic;
signal \N__22546\ : std_logic;
signal \N__22539\ : std_logic;
signal \N__22536\ : std_logic;
signal \N__22535\ : std_logic;
signal \N__22534\ : std_logic;
signal \N__22531\ : std_logic;
signal \N__22528\ : std_logic;
signal \N__22525\ : std_logic;
signal \N__22522\ : std_logic;
signal \N__22515\ : std_logic;
signal \N__22512\ : std_logic;
signal \N__22511\ : std_logic;
signal \N__22510\ : std_logic;
signal \N__22507\ : std_logic;
signal \N__22504\ : std_logic;
signal \N__22501\ : std_logic;
signal \N__22498\ : std_logic;
signal \N__22491\ : std_logic;
signal \N__22488\ : std_logic;
signal \N__22487\ : std_logic;
signal \N__22484\ : std_logic;
signal \N__22483\ : std_logic;
signal \N__22480\ : std_logic;
signal \N__22477\ : std_logic;
signal \N__22474\ : std_logic;
signal \N__22467\ : std_logic;
signal \N__22464\ : std_logic;
signal \N__22463\ : std_logic;
signal \N__22462\ : std_logic;
signal \N__22459\ : std_logic;
signal \N__22456\ : std_logic;
signal \N__22453\ : std_logic;
signal \N__22448\ : std_logic;
signal \N__22445\ : std_logic;
signal \N__22440\ : std_logic;
signal \N__22437\ : std_logic;
signal \N__22436\ : std_logic;
signal \N__22435\ : std_logic;
signal \N__22432\ : std_logic;
signal \N__22429\ : std_logic;
signal \N__22426\ : std_logic;
signal \N__22419\ : std_logic;
signal \N__22416\ : std_logic;
signal \N__22415\ : std_logic;
signal \N__22414\ : std_logic;
signal \N__22411\ : std_logic;
signal \N__22408\ : std_logic;
signal \N__22405\ : std_logic;
signal \N__22402\ : std_logic;
signal \N__22395\ : std_logic;
signal \N__22394\ : std_logic;
signal \N__22393\ : std_logic;
signal \N__22392\ : std_logic;
signal \N__22391\ : std_logic;
signal \N__22390\ : std_logic;
signal \N__22389\ : std_logic;
signal \N__22388\ : std_logic;
signal \N__22387\ : std_logic;
signal \N__22386\ : std_logic;
signal \N__22385\ : std_logic;
signal \N__22382\ : std_logic;
signal \N__22379\ : std_logic;
signal \N__22376\ : std_logic;
signal \N__22373\ : std_logic;
signal \N__22370\ : std_logic;
signal \N__22367\ : std_logic;
signal \N__22364\ : std_logic;
signal \N__22361\ : std_logic;
signal \N__22358\ : std_logic;
signal \N__22355\ : std_logic;
signal \N__22352\ : std_logic;
signal \N__22347\ : std_logic;
signal \N__22340\ : std_logic;
signal \N__22333\ : std_logic;
signal \N__22326\ : std_logic;
signal \N__22317\ : std_logic;
signal \N__22314\ : std_logic;
signal \N__22311\ : std_logic;
signal \N__22310\ : std_logic;
signal \N__22307\ : std_logic;
signal \N__22304\ : std_logic;
signal \N__22303\ : std_logic;
signal \N__22302\ : std_logic;
signal \N__22297\ : std_logic;
signal \N__22294\ : std_logic;
signal \N__22291\ : std_logic;
signal \N__22286\ : std_logic;
signal \N__22283\ : std_logic;
signal \N__22280\ : std_logic;
signal \N__22277\ : std_logic;
signal \N__22272\ : std_logic;
signal \N__22269\ : std_logic;
signal \N__22266\ : std_logic;
signal \N__22263\ : std_logic;
signal \N__22260\ : std_logic;
signal \N__22259\ : std_logic;
signal \N__22258\ : std_logic;
signal \N__22255\ : std_logic;
signal \N__22252\ : std_logic;
signal \N__22249\ : std_logic;
signal \N__22246\ : std_logic;
signal \N__22239\ : std_logic;
signal \N__22238\ : std_logic;
signal \N__22235\ : std_logic;
signal \N__22232\ : std_logic;
signal \N__22229\ : std_logic;
signal \N__22226\ : std_logic;
signal \N__22221\ : std_logic;
signal \N__22218\ : std_logic;
signal \N__22217\ : std_logic;
signal \N__22216\ : std_logic;
signal \N__22213\ : std_logic;
signal \N__22210\ : std_logic;
signal \N__22207\ : std_logic;
signal \N__22200\ : std_logic;
signal \N__22197\ : std_logic;
signal \N__22196\ : std_logic;
signal \N__22195\ : std_logic;
signal \N__22192\ : std_logic;
signal \N__22189\ : std_logic;
signal \N__22186\ : std_logic;
signal \N__22179\ : std_logic;
signal \N__22176\ : std_logic;
signal \N__22175\ : std_logic;
signal \N__22174\ : std_logic;
signal \N__22171\ : std_logic;
signal \N__22168\ : std_logic;
signal \N__22165\ : std_logic;
signal \N__22158\ : std_logic;
signal \N__22155\ : std_logic;
signal \N__22152\ : std_logic;
signal \N__22149\ : std_logic;
signal \N__22146\ : std_logic;
signal \N__22143\ : std_logic;
signal \N__22142\ : std_logic;
signal \N__22139\ : std_logic;
signal \N__22136\ : std_logic;
signal \N__22133\ : std_logic;
signal \N__22128\ : std_logic;
signal \N__22125\ : std_logic;
signal \N__22122\ : std_logic;
signal \N__22119\ : std_logic;
signal \N__22118\ : std_logic;
signal \N__22115\ : std_logic;
signal \N__22112\ : std_logic;
signal \N__22111\ : std_logic;
signal \N__22108\ : std_logic;
signal \N__22105\ : std_logic;
signal \N__22102\ : std_logic;
signal \N__22095\ : std_logic;
signal \N__22092\ : std_logic;
signal \N__22089\ : std_logic;
signal \N__22086\ : std_logic;
signal \N__22083\ : std_logic;
signal \N__22080\ : std_logic;
signal \N__22077\ : std_logic;
signal \N__22074\ : std_logic;
signal \N__22073\ : std_logic;
signal \N__22070\ : std_logic;
signal \N__22067\ : std_logic;
signal \N__22062\ : std_logic;
signal \N__22059\ : std_logic;
signal \N__22058\ : std_logic;
signal \N__22055\ : std_logic;
signal \N__22052\ : std_logic;
signal \N__22047\ : std_logic;
signal \N__22044\ : std_logic;
signal \N__22041\ : std_logic;
signal \N__22040\ : std_logic;
signal \N__22037\ : std_logic;
signal \N__22034\ : std_logic;
signal \N__22031\ : std_logic;
signal \N__22026\ : std_logic;
signal \N__22023\ : std_logic;
signal \N__22022\ : std_logic;
signal \N__22019\ : std_logic;
signal \N__22016\ : std_logic;
signal \N__22013\ : std_logic;
signal \N__22008\ : std_logic;
signal \N__22005\ : std_logic;
signal \N__22002\ : std_logic;
signal \N__21999\ : std_logic;
signal \N__21998\ : std_logic;
signal \N__21995\ : std_logic;
signal \N__21992\ : std_logic;
signal \N__21989\ : std_logic;
signal \N__21984\ : std_logic;
signal \N__21983\ : std_logic;
signal \N__21982\ : std_logic;
signal \N__21981\ : std_logic;
signal \N__21980\ : std_logic;
signal \N__21977\ : std_logic;
signal \N__21974\ : std_logic;
signal \N__21973\ : std_logic;
signal \N__21972\ : std_logic;
signal \N__21969\ : std_logic;
signal \N__21966\ : std_logic;
signal \N__21965\ : std_logic;
signal \N__21962\ : std_logic;
signal \N__21955\ : std_logic;
signal \N__21950\ : std_logic;
signal \N__21945\ : std_logic;
signal \N__21936\ : std_logic;
signal \N__21933\ : std_logic;
signal \N__21930\ : std_logic;
signal \N__21929\ : std_logic;
signal \N__21926\ : std_logic;
signal \N__21925\ : std_logic;
signal \N__21918\ : std_logic;
signal \N__21915\ : std_logic;
signal \N__21912\ : std_logic;
signal \N__21909\ : std_logic;
signal \N__21906\ : std_logic;
signal \N__21903\ : std_logic;
signal \N__21900\ : std_logic;
signal \N__21899\ : std_logic;
signal \N__21896\ : std_logic;
signal \N__21895\ : std_logic;
signal \N__21892\ : std_logic;
signal \N__21889\ : std_logic;
signal \N__21886\ : std_logic;
signal \N__21879\ : std_logic;
signal \N__21876\ : std_logic;
signal \N__21873\ : std_logic;
signal \N__21870\ : std_logic;
signal \N__21867\ : std_logic;
signal \N__21864\ : std_logic;
signal \N__21861\ : std_logic;
signal \N__21860\ : std_logic;
signal \N__21857\ : std_logic;
signal \N__21854\ : std_logic;
signal \N__21853\ : std_logic;
signal \N__21850\ : std_logic;
signal \N__21847\ : std_logic;
signal \N__21844\ : std_logic;
signal \N__21837\ : std_logic;
signal \N__21834\ : std_logic;
signal \N__21831\ : std_logic;
signal \N__21828\ : std_logic;
signal \N__21827\ : std_logic;
signal \N__21826\ : std_logic;
signal \N__21825\ : std_logic;
signal \N__21822\ : std_logic;
signal \N__21821\ : std_logic;
signal \N__21820\ : std_logic;
signal \N__21817\ : std_logic;
signal \N__21816\ : std_logic;
signal \N__21813\ : std_logic;
signal \N__21810\ : std_logic;
signal \N__21809\ : std_logic;
signal \N__21804\ : std_logic;
signal \N__21801\ : std_logic;
signal \N__21790\ : std_logic;
signal \N__21787\ : std_logic;
signal \N__21780\ : std_logic;
signal \N__21777\ : std_logic;
signal \N__21774\ : std_logic;
signal \N__21771\ : std_logic;
signal \N__21768\ : std_logic;
signal \N__21765\ : std_logic;
signal \N__21762\ : std_logic;
signal \N__21761\ : std_logic;
signal \N__21760\ : std_logic;
signal \N__21757\ : std_logic;
signal \N__21754\ : std_logic;
signal \N__21751\ : std_logic;
signal \N__21748\ : std_logic;
signal \N__21741\ : std_logic;
signal \N__21738\ : std_logic;
signal \N__21735\ : std_logic;
signal \N__21732\ : std_logic;
signal \N__21729\ : std_logic;
signal \N__21726\ : std_logic;
signal \N__21725\ : std_logic;
signal \N__21724\ : std_logic;
signal \N__21721\ : std_logic;
signal \N__21716\ : std_logic;
signal \N__21713\ : std_logic;
signal \N__21708\ : std_logic;
signal \N__21705\ : std_logic;
signal \N__21702\ : std_logic;
signal \N__21699\ : std_logic;
signal \N__21698\ : std_logic;
signal \N__21697\ : std_logic;
signal \N__21694\ : std_logic;
signal \N__21689\ : std_logic;
signal \N__21686\ : std_logic;
signal \N__21681\ : std_logic;
signal \N__21678\ : std_logic;
signal \N__21675\ : std_logic;
signal \N__21672\ : std_logic;
signal \N__21671\ : std_logic;
signal \N__21670\ : std_logic;
signal \N__21667\ : std_logic;
signal \N__21662\ : std_logic;
signal \N__21659\ : std_logic;
signal \N__21654\ : std_logic;
signal \N__21651\ : std_logic;
signal \N__21648\ : std_logic;
signal \N__21645\ : std_logic;
signal \N__21642\ : std_logic;
signal \N__21639\ : std_logic;
signal \N__21636\ : std_logic;
signal \N__21633\ : std_logic;
signal \N__21632\ : std_logic;
signal \N__21629\ : std_logic;
signal \N__21626\ : std_logic;
signal \N__21623\ : std_logic;
signal \N__21618\ : std_logic;
signal \N__21615\ : std_logic;
signal \N__21612\ : std_logic;
signal \N__21609\ : std_logic;
signal \N__21606\ : std_logic;
signal \N__21605\ : std_logic;
signal \N__21602\ : std_logic;
signal \N__21601\ : std_logic;
signal \N__21598\ : std_logic;
signal \N__21595\ : std_logic;
signal \N__21592\ : std_logic;
signal \N__21585\ : std_logic;
signal \N__21582\ : std_logic;
signal \N__21579\ : std_logic;
signal \N__21576\ : std_logic;
signal \N__21573\ : std_logic;
signal \N__21570\ : std_logic;
signal \N__21567\ : std_logic;
signal \N__21564\ : std_logic;
signal \N__21561\ : std_logic;
signal \N__21560\ : std_logic;
signal \N__21557\ : std_logic;
signal \N__21556\ : std_logic;
signal \N__21553\ : std_logic;
signal \N__21550\ : std_logic;
signal \N__21547\ : std_logic;
signal \N__21544\ : std_logic;
signal \N__21537\ : std_logic;
signal \N__21534\ : std_logic;
signal \N__21531\ : std_logic;
signal \N__21528\ : std_logic;
signal \N__21525\ : std_logic;
signal \N__21522\ : std_logic;
signal \N__21519\ : std_logic;
signal \N__21516\ : std_logic;
signal \N__21513\ : std_logic;
signal \N__21510\ : std_logic;
signal \N__21507\ : std_logic;
signal \N__21504\ : std_logic;
signal \N__21501\ : std_logic;
signal \N__21498\ : std_logic;
signal \N__21495\ : std_logic;
signal \N__21492\ : std_logic;
signal \N__21489\ : std_logic;
signal \N__21486\ : std_logic;
signal \N__21483\ : std_logic;
signal \N__21480\ : std_logic;
signal \N__21477\ : std_logic;
signal \N__21474\ : std_logic;
signal \N__21471\ : std_logic;
signal \N__21468\ : std_logic;
signal \N__21465\ : std_logic;
signal \N__21462\ : std_logic;
signal \N__21459\ : std_logic;
signal \N__21456\ : std_logic;
signal \N__21453\ : std_logic;
signal \N__21450\ : std_logic;
signal \N__21447\ : std_logic;
signal \N__21444\ : std_logic;
signal \N__21441\ : std_logic;
signal \N__21438\ : std_logic;
signal \N__21437\ : std_logic;
signal \N__21434\ : std_logic;
signal \N__21431\ : std_logic;
signal \N__21426\ : std_logic;
signal \N__21423\ : std_logic;
signal \N__21420\ : std_logic;
signal \N__21417\ : std_logic;
signal \N__21414\ : std_logic;
signal \N__21413\ : std_logic;
signal \N__21410\ : std_logic;
signal \N__21407\ : std_logic;
signal \N__21402\ : std_logic;
signal \N__21399\ : std_logic;
signal \N__21396\ : std_logic;
signal \N__21393\ : std_logic;
signal \N__21390\ : std_logic;
signal \N__21387\ : std_logic;
signal \N__21384\ : std_logic;
signal \N__21383\ : std_logic;
signal \N__21382\ : std_logic;
signal \N__21379\ : std_logic;
signal \N__21376\ : std_logic;
signal \N__21375\ : std_logic;
signal \N__21372\ : std_logic;
signal \N__21367\ : std_logic;
signal \N__21364\ : std_logic;
signal \N__21361\ : std_logic;
signal \N__21356\ : std_logic;
signal \N__21351\ : std_logic;
signal \N__21348\ : std_logic;
signal \N__21347\ : std_logic;
signal \N__21342\ : std_logic;
signal \N__21339\ : std_logic;
signal \N__21336\ : std_logic;
signal \N__21333\ : std_logic;
signal \N__21332\ : std_logic;
signal \N__21331\ : std_logic;
signal \N__21328\ : std_logic;
signal \N__21327\ : std_logic;
signal \N__21322\ : std_logic;
signal \N__21319\ : std_logic;
signal \N__21316\ : std_logic;
signal \N__21313\ : std_logic;
signal \N__21310\ : std_logic;
signal \N__21307\ : std_logic;
signal \N__21304\ : std_logic;
signal \N__21297\ : std_logic;
signal \N__21296\ : std_logic;
signal \N__21293\ : std_logic;
signal \N__21290\ : std_logic;
signal \N__21287\ : std_logic;
signal \N__21284\ : std_logic;
signal \N__21281\ : std_logic;
signal \N__21276\ : std_logic;
signal \N__21273\ : std_logic;
signal \N__21270\ : std_logic;
signal \N__21269\ : std_logic;
signal \N__21268\ : std_logic;
signal \N__21265\ : std_logic;
signal \N__21262\ : std_logic;
signal \N__21259\ : std_logic;
signal \N__21258\ : std_logic;
signal \N__21255\ : std_logic;
signal \N__21250\ : std_logic;
signal \N__21247\ : std_logic;
signal \N__21240\ : std_logic;
signal \N__21237\ : std_logic;
signal \N__21234\ : std_logic;
signal \N__21231\ : std_logic;
signal \N__21228\ : std_logic;
signal \N__21225\ : std_logic;
signal \N__21222\ : std_logic;
signal \N__21219\ : std_logic;
signal \N__21216\ : std_logic;
signal \N__21213\ : std_logic;
signal \N__21210\ : std_logic;
signal \N__21207\ : std_logic;
signal \N__21204\ : std_logic;
signal \N__21201\ : std_logic;
signal \N__21198\ : std_logic;
signal \N__21195\ : std_logic;
signal \N__21192\ : std_logic;
signal \N__21189\ : std_logic;
signal \N__21186\ : std_logic;
signal \N__21183\ : std_logic;
signal \N__21180\ : std_logic;
signal \N__21177\ : std_logic;
signal \N__21176\ : std_logic;
signal \N__21173\ : std_logic;
signal \N__21170\ : std_logic;
signal \N__21165\ : std_logic;
signal \N__21162\ : std_logic;
signal \N__21159\ : std_logic;
signal \N__21156\ : std_logic;
signal \N__21153\ : std_logic;
signal \N__21150\ : std_logic;
signal \N__21147\ : std_logic;
signal \N__21144\ : std_logic;
signal \N__21141\ : std_logic;
signal \N__21138\ : std_logic;
signal \N__21135\ : std_logic;
signal \N__21132\ : std_logic;
signal \N__21129\ : std_logic;
signal \N__21126\ : std_logic;
signal \N__21123\ : std_logic;
signal \N__21120\ : std_logic;
signal \N__21119\ : std_logic;
signal \N__21116\ : std_logic;
signal \N__21113\ : std_logic;
signal \N__21110\ : std_logic;
signal \N__21109\ : std_logic;
signal \N__21106\ : std_logic;
signal \N__21103\ : std_logic;
signal \N__21100\ : std_logic;
signal \N__21097\ : std_logic;
signal \N__21090\ : std_logic;
signal \N__21089\ : std_logic;
signal \N__21086\ : std_logic;
signal \N__21083\ : std_logic;
signal \N__21078\ : std_logic;
signal \N__21075\ : std_logic;
signal \N__21072\ : std_logic;
signal \N__21069\ : std_logic;
signal \N__21066\ : std_logic;
signal \N__21063\ : std_logic;
signal \N__21060\ : std_logic;
signal \N__21057\ : std_logic;
signal \N__21054\ : std_logic;
signal \N__21051\ : std_logic;
signal \N__21048\ : std_logic;
signal \N__21045\ : std_logic;
signal \N__21042\ : std_logic;
signal \N__21039\ : std_logic;
signal \N__21036\ : std_logic;
signal \N__21033\ : std_logic;
signal \N__21030\ : std_logic;
signal \N__21029\ : std_logic;
signal \N__21028\ : std_logic;
signal \N__21025\ : std_logic;
signal \N__21022\ : std_logic;
signal \N__21019\ : std_logic;
signal \N__21012\ : std_logic;
signal \N__21009\ : std_logic;
signal \N__21008\ : std_logic;
signal \N__21007\ : std_logic;
signal \N__21004\ : std_logic;
signal \N__21001\ : std_logic;
signal \N__20998\ : std_logic;
signal \N__20991\ : std_logic;
signal \N__20988\ : std_logic;
signal \N__20987\ : std_logic;
signal \N__20984\ : std_logic;
signal \N__20981\ : std_logic;
signal \N__20976\ : std_logic;
signal \N__20973\ : std_logic;
signal \N__20970\ : std_logic;
signal \N__20969\ : std_logic;
signal \N__20966\ : std_logic;
signal \N__20963\ : std_logic;
signal \N__20958\ : std_logic;
signal \N__20957\ : std_logic;
signal \N__20954\ : std_logic;
signal \N__20951\ : std_logic;
signal \N__20946\ : std_logic;
signal \N__20943\ : std_logic;
signal \N__20942\ : std_logic;
signal \N__20941\ : std_logic;
signal \N__20938\ : std_logic;
signal \N__20935\ : std_logic;
signal \N__20932\ : std_logic;
signal \N__20925\ : std_logic;
signal \N__20922\ : std_logic;
signal \N__20921\ : std_logic;
signal \N__20918\ : std_logic;
signal \N__20915\ : std_logic;
signal \N__20910\ : std_logic;
signal \N__20909\ : std_logic;
signal \N__20906\ : std_logic;
signal \N__20903\ : std_logic;
signal \N__20898\ : std_logic;
signal \N__20897\ : std_logic;
signal \N__20896\ : std_logic;
signal \N__20895\ : std_logic;
signal \N__20894\ : std_logic;
signal \N__20893\ : std_logic;
signal \N__20892\ : std_logic;
signal \N__20891\ : std_logic;
signal \N__20890\ : std_logic;
signal \N__20889\ : std_logic;
signal \N__20886\ : std_logic;
signal \N__20883\ : std_logic;
signal \N__20880\ : std_logic;
signal \N__20877\ : std_logic;
signal \N__20874\ : std_logic;
signal \N__20871\ : std_logic;
signal \N__20868\ : std_logic;
signal \N__20865\ : std_logic;
signal \N__20862\ : std_logic;
signal \N__20859\ : std_logic;
signal \N__20854\ : std_logic;
signal \N__20849\ : std_logic;
signal \N__20842\ : std_logic;
signal \N__20835\ : std_logic;
signal \N__20826\ : std_logic;
signal \N__20823\ : std_logic;
signal \N__20820\ : std_logic;
signal \N__20817\ : std_logic;
signal \N__20814\ : std_logic;
signal \N__20811\ : std_logic;
signal \N__20808\ : std_logic;
signal \N__20805\ : std_logic;
signal \N__20802\ : std_logic;
signal \N__20799\ : std_logic;
signal \N__20796\ : std_logic;
signal \N__20793\ : std_logic;
signal \N__20792\ : std_logic;
signal \N__20789\ : std_logic;
signal \N__20786\ : std_logic;
signal \N__20783\ : std_logic;
signal \N__20778\ : std_logic;
signal \N__20777\ : std_logic;
signal \N__20774\ : std_logic;
signal \N__20771\ : std_logic;
signal \N__20768\ : std_logic;
signal \N__20763\ : std_logic;
signal \N__20760\ : std_logic;
signal \N__20757\ : std_logic;
signal \N__20756\ : std_logic;
signal \N__20753\ : std_logic;
signal \N__20750\ : std_logic;
signal \N__20747\ : std_logic;
signal \N__20742\ : std_logic;
signal \N__20741\ : std_logic;
signal \N__20738\ : std_logic;
signal \N__20735\ : std_logic;
signal \N__20732\ : std_logic;
signal \N__20727\ : std_logic;
signal \N__20724\ : std_logic;
signal \N__20723\ : std_logic;
signal \N__20720\ : std_logic;
signal \N__20717\ : std_logic;
signal \N__20712\ : std_logic;
signal \N__20711\ : std_logic;
signal \N__20708\ : std_logic;
signal \N__20705\ : std_logic;
signal \N__20702\ : std_logic;
signal \N__20699\ : std_logic;
signal \N__20694\ : std_logic;
signal \N__20691\ : std_logic;
signal \N__20690\ : std_logic;
signal \N__20689\ : std_logic;
signal \N__20686\ : std_logic;
signal \N__20683\ : std_logic;
signal \N__20680\ : std_logic;
signal \N__20673\ : std_logic;
signal \N__20670\ : std_logic;
signal \N__20669\ : std_logic;
signal \N__20666\ : std_logic;
signal \N__20663\ : std_logic;
signal \N__20658\ : std_logic;
signal \N__20655\ : std_logic;
signal \N__20654\ : std_logic;
signal \N__20653\ : std_logic;
signal \N__20650\ : std_logic;
signal \N__20647\ : std_logic;
signal \N__20644\ : std_logic;
signal \N__20637\ : std_logic;
signal \N__20634\ : std_logic;
signal \N__20633\ : std_logic;
signal \N__20632\ : std_logic;
signal \N__20629\ : std_logic;
signal \N__20626\ : std_logic;
signal \N__20623\ : std_logic;
signal \N__20616\ : std_logic;
signal \N__20613\ : std_logic;
signal \N__20612\ : std_logic;
signal \N__20609\ : std_logic;
signal \N__20606\ : std_logic;
signal \N__20603\ : std_logic;
signal \N__20598\ : std_logic;
signal \N__20597\ : std_logic;
signal \N__20594\ : std_logic;
signal \N__20591\ : std_logic;
signal \N__20588\ : std_logic;
signal \N__20583\ : std_logic;
signal \N__20580\ : std_logic;
signal \N__20577\ : std_logic;
signal \N__20574\ : std_logic;
signal \N__20573\ : std_logic;
signal \N__20572\ : std_logic;
signal \N__20569\ : std_logic;
signal \N__20566\ : std_logic;
signal \N__20563\ : std_logic;
signal \N__20560\ : std_logic;
signal \N__20555\ : std_logic;
signal \N__20550\ : std_logic;
signal \N__20549\ : std_logic;
signal \N__20546\ : std_logic;
signal \N__20545\ : std_logic;
signal \N__20542\ : std_logic;
signal \N__20539\ : std_logic;
signal \N__20536\ : std_logic;
signal \N__20533\ : std_logic;
signal \N__20528\ : std_logic;
signal \N__20523\ : std_logic;
signal \N__20520\ : std_logic;
signal \N__20519\ : std_logic;
signal \N__20518\ : std_logic;
signal \N__20515\ : std_logic;
signal \N__20512\ : std_logic;
signal \N__20509\ : std_logic;
signal \N__20506\ : std_logic;
signal \N__20501\ : std_logic;
signal \N__20496\ : std_logic;
signal \N__20493\ : std_logic;
signal \N__20490\ : std_logic;
signal \N__20487\ : std_logic;
signal \N__20484\ : std_logic;
signal \N__20481\ : std_logic;
signal \N__20480\ : std_logic;
signal \N__20477\ : std_logic;
signal \N__20476\ : std_logic;
signal \N__20475\ : std_logic;
signal \N__20474\ : std_logic;
signal \N__20471\ : std_logic;
signal \N__20470\ : std_logic;
signal \N__20469\ : std_logic;
signal \N__20468\ : std_logic;
signal \N__20467\ : std_logic;
signal \N__20462\ : std_logic;
signal \N__20453\ : std_logic;
signal \N__20448\ : std_logic;
signal \N__20445\ : std_logic;
signal \N__20436\ : std_logic;
signal \N__20433\ : std_logic;
signal \N__20432\ : std_logic;
signal \N__20429\ : std_logic;
signal \N__20426\ : std_logic;
signal \N__20423\ : std_logic;
signal \N__20422\ : std_logic;
signal \N__20419\ : std_logic;
signal \N__20416\ : std_logic;
signal \N__20413\ : std_logic;
signal \N__20406\ : std_logic;
signal \N__20403\ : std_logic;
signal \N__20400\ : std_logic;
signal \N__20397\ : std_logic;
signal \N__20394\ : std_logic;
signal \N__20391\ : std_logic;
signal \N__20388\ : std_logic;
signal \N__20385\ : std_logic;
signal \N__20382\ : std_logic;
signal \N__20381\ : std_logic;
signal \N__20378\ : std_logic;
signal \N__20375\ : std_logic;
signal \N__20372\ : std_logic;
signal \N__20367\ : std_logic;
signal \N__20364\ : std_logic;
signal \N__20361\ : std_logic;
signal \N__20358\ : std_logic;
signal \N__20355\ : std_logic;
signal \N__20352\ : std_logic;
signal \N__20349\ : std_logic;
signal \N__20346\ : std_logic;
signal \N__20343\ : std_logic;
signal \N__20342\ : std_logic;
signal \N__20341\ : std_logic;
signal \N__20338\ : std_logic;
signal \N__20333\ : std_logic;
signal \N__20330\ : std_logic;
signal \N__20325\ : std_logic;
signal \N__20322\ : std_logic;
signal \N__20319\ : std_logic;
signal \N__20316\ : std_logic;
signal \N__20313\ : std_logic;
signal \N__20310\ : std_logic;
signal \N__20307\ : std_logic;
signal \N__20304\ : std_logic;
signal \N__20301\ : std_logic;
signal \N__20298\ : std_logic;
signal \N__20295\ : std_logic;
signal \N__20292\ : std_logic;
signal \N__20291\ : std_logic;
signal \N__20290\ : std_logic;
signal \N__20287\ : std_logic;
signal \N__20282\ : std_logic;
signal \N__20279\ : std_logic;
signal \N__20274\ : std_logic;
signal \N__20271\ : std_logic;
signal \N__20268\ : std_logic;
signal \N__20265\ : std_logic;
signal \N__20262\ : std_logic;
signal \N__20259\ : std_logic;
signal \N__20256\ : std_logic;
signal \N__20253\ : std_logic;
signal \N__20252\ : std_logic;
signal \N__20249\ : std_logic;
signal \N__20246\ : std_logic;
signal \N__20241\ : std_logic;
signal \N__20238\ : std_logic;
signal \N__20235\ : std_logic;
signal \N__20232\ : std_logic;
signal \N__20229\ : std_logic;
signal \N__20226\ : std_logic;
signal \N__20223\ : std_logic;
signal \N__20220\ : std_logic;
signal \N__20217\ : std_logic;
signal \N__20214\ : std_logic;
signal \N__20211\ : std_logic;
signal \N__20210\ : std_logic;
signal \N__20207\ : std_logic;
signal \N__20204\ : std_logic;
signal \N__20201\ : std_logic;
signal \N__20196\ : std_logic;
signal \N__20193\ : std_logic;
signal \N__20190\ : std_logic;
signal \N__20187\ : std_logic;
signal \N__20184\ : std_logic;
signal \N__20181\ : std_logic;
signal \N__20178\ : std_logic;
signal \N__20177\ : std_logic;
signal \N__20176\ : std_logic;
signal \N__20173\ : std_logic;
signal \N__20170\ : std_logic;
signal \N__20167\ : std_logic;
signal \N__20164\ : std_logic;
signal \N__20157\ : std_logic;
signal \N__20154\ : std_logic;
signal \N__20153\ : std_logic;
signal \N__20150\ : std_logic;
signal \N__20147\ : std_logic;
signal \N__20144\ : std_logic;
signal \N__20139\ : std_logic;
signal \N__20138\ : std_logic;
signal \N__20135\ : std_logic;
signal \N__20132\ : std_logic;
signal \N__20127\ : std_logic;
signal \N__20124\ : std_logic;
signal \N__20121\ : std_logic;
signal \N__20118\ : std_logic;
signal \N__20115\ : std_logic;
signal \N__20112\ : std_logic;
signal \N__20109\ : std_logic;
signal \N__20106\ : std_logic;
signal \N__20103\ : std_logic;
signal \N__20100\ : std_logic;
signal \N__20099\ : std_logic;
signal \N__20096\ : std_logic;
signal \N__20093\ : std_logic;
signal \N__20090\ : std_logic;
signal \N__20087\ : std_logic;
signal \N__20084\ : std_logic;
signal \N__20079\ : std_logic;
signal \N__20076\ : std_logic;
signal \N__20073\ : std_logic;
signal \N__20070\ : std_logic;
signal \N__20067\ : std_logic;
signal \N__20064\ : std_logic;
signal \N__20063\ : std_logic;
signal \N__20060\ : std_logic;
signal \N__20057\ : std_logic;
signal \N__20052\ : std_logic;
signal \N__20049\ : std_logic;
signal \N__20048\ : std_logic;
signal \N__20047\ : std_logic;
signal \N__20040\ : std_logic;
signal \N__20037\ : std_logic;
signal \N__20034\ : std_logic;
signal \N__20031\ : std_logic;
signal \N__20030\ : std_logic;
signal \N__20027\ : std_logic;
signal \N__20022\ : std_logic;
signal \N__20019\ : std_logic;
signal \N__20016\ : std_logic;
signal \N__20013\ : std_logic;
signal \N__20010\ : std_logic;
signal \N__20009\ : std_logic;
signal \N__20006\ : std_logic;
signal \N__20005\ : std_logic;
signal \N__19998\ : std_logic;
signal \N__19995\ : std_logic;
signal \N__19992\ : std_logic;
signal \N__19989\ : std_logic;
signal \N__19988\ : std_logic;
signal \N__19987\ : std_logic;
signal \N__19984\ : std_logic;
signal \N__19979\ : std_logic;
signal \N__19976\ : std_logic;
signal \N__19973\ : std_logic;
signal \N__19968\ : std_logic;
signal \N__19965\ : std_logic;
signal \N__19962\ : std_logic;
signal \N__19961\ : std_logic;
signal \N__19960\ : std_logic;
signal \N__19953\ : std_logic;
signal \N__19950\ : std_logic;
signal \N__19947\ : std_logic;
signal \N__19944\ : std_logic;
signal \N__19941\ : std_logic;
signal \N__19938\ : std_logic;
signal \N__19935\ : std_logic;
signal \N__19932\ : std_logic;
signal \N__19929\ : std_logic;
signal \N__19928\ : std_logic;
signal \N__19927\ : std_logic;
signal \N__19924\ : std_logic;
signal \N__19921\ : std_logic;
signal \N__19918\ : std_logic;
signal \N__19915\ : std_logic;
signal \N__19908\ : std_logic;
signal \N__19907\ : std_logic;
signal \N__19902\ : std_logic;
signal \N__19899\ : std_logic;
signal \N__19898\ : std_logic;
signal \N__19897\ : std_logic;
signal \N__19894\ : std_logic;
signal \N__19891\ : std_logic;
signal \N__19888\ : std_logic;
signal \N__19881\ : std_logic;
signal \N__19880\ : std_logic;
signal \N__19879\ : std_logic;
signal \N__19876\ : std_logic;
signal \N__19873\ : std_logic;
signal \N__19870\ : std_logic;
signal \N__19867\ : std_logic;
signal \N__19860\ : std_logic;
signal \N__19857\ : std_logic;
signal \N__19854\ : std_logic;
signal \N__19851\ : std_logic;
signal \N__19848\ : std_logic;
signal \N__19845\ : std_logic;
signal \N__19842\ : std_logic;
signal \N__19839\ : std_logic;
signal \N__19836\ : std_logic;
signal \N__19833\ : std_logic;
signal \N__19830\ : std_logic;
signal \N__19827\ : std_logic;
signal \N__19824\ : std_logic;
signal \N__19821\ : std_logic;
signal \N__19818\ : std_logic;
signal \N__19815\ : std_logic;
signal \N__19812\ : std_logic;
signal \N__19809\ : std_logic;
signal \N__19806\ : std_logic;
signal \N__19803\ : std_logic;
signal \N__19800\ : std_logic;
signal \N__19797\ : std_logic;
signal \N__19794\ : std_logic;
signal \N__19791\ : std_logic;
signal \N__19788\ : std_logic;
signal \N__19785\ : std_logic;
signal \N__19782\ : std_logic;
signal \N__19779\ : std_logic;
signal \N__19776\ : std_logic;
signal \N__19773\ : std_logic;
signal \N__19772\ : std_logic;
signal \N__19771\ : std_logic;
signal \N__19768\ : std_logic;
signal \N__19765\ : std_logic;
signal \N__19762\ : std_logic;
signal \N__19755\ : std_logic;
signal \N__19752\ : std_logic;
signal \N__19751\ : std_logic;
signal \N__19746\ : std_logic;
signal \N__19743\ : std_logic;
signal \N__19742\ : std_logic;
signal \N__19741\ : std_logic;
signal \N__19738\ : std_logic;
signal \N__19735\ : std_logic;
signal \N__19732\ : std_logic;
signal \N__19729\ : std_logic;
signal \N__19722\ : std_logic;
signal \N__19719\ : std_logic;
signal \N__19718\ : std_logic;
signal \N__19713\ : std_logic;
signal \N__19710\ : std_logic;
signal \N__19709\ : std_logic;
signal \N__19708\ : std_logic;
signal \N__19705\ : std_logic;
signal \N__19702\ : std_logic;
signal \N__19699\ : std_logic;
signal \N__19696\ : std_logic;
signal \N__19689\ : std_logic;
signal \N__19688\ : std_logic;
signal \N__19685\ : std_logic;
signal \N__19682\ : std_logic;
signal \N__19677\ : std_logic;
signal \N__19674\ : std_logic;
signal \N__19671\ : std_logic;
signal \N__19670\ : std_logic;
signal \N__19667\ : std_logic;
signal \N__19664\ : std_logic;
signal \N__19661\ : std_logic;
signal \N__19658\ : std_logic;
signal \N__19655\ : std_logic;
signal \N__19652\ : std_logic;
signal \N__19647\ : std_logic;
signal \N__19644\ : std_logic;
signal \N__19641\ : std_logic;
signal \N__19638\ : std_logic;
signal \N__19635\ : std_logic;
signal \N__19632\ : std_logic;
signal \N__19629\ : std_logic;
signal \N__19626\ : std_logic;
signal \N__19623\ : std_logic;
signal \N__19620\ : std_logic;
signal \N__19617\ : std_logic;
signal \N__19614\ : std_logic;
signal \N__19611\ : std_logic;
signal \N__19608\ : std_logic;
signal \N__19607\ : std_logic;
signal \N__19604\ : std_logic;
signal \N__19603\ : std_logic;
signal \N__19600\ : std_logic;
signal \N__19597\ : std_logic;
signal \N__19594\ : std_logic;
signal \N__19587\ : std_logic;
signal \N__19584\ : std_logic;
signal \N__19581\ : std_logic;
signal \N__19578\ : std_logic;
signal \N__19575\ : std_logic;
signal \N__19572\ : std_logic;
signal \N__19571\ : std_logic;
signal \N__19568\ : std_logic;
signal \N__19565\ : std_logic;
signal \N__19564\ : std_logic;
signal \N__19561\ : std_logic;
signal \N__19558\ : std_logic;
signal \N__19555\ : std_logic;
signal \N__19548\ : std_logic;
signal \N__19545\ : std_logic;
signal \N__19542\ : std_logic;
signal \N__19539\ : std_logic;
signal \N__19536\ : std_logic;
signal \N__19533\ : std_logic;
signal \N__19530\ : std_logic;
signal \N__19527\ : std_logic;
signal \N__19524\ : std_logic;
signal \N__19521\ : std_logic;
signal \N__19520\ : std_logic;
signal \N__19519\ : std_logic;
signal \N__19518\ : std_logic;
signal \N__19515\ : std_logic;
signal \N__19514\ : std_logic;
signal \N__19513\ : std_logic;
signal \N__19510\ : std_logic;
signal \N__19509\ : std_logic;
signal \N__19506\ : std_logic;
signal \N__19505\ : std_logic;
signal \N__19502\ : std_logic;
signal \N__19501\ : std_logic;
signal \N__19500\ : std_logic;
signal \N__19495\ : std_logic;
signal \N__19484\ : std_logic;
signal \N__19477\ : std_logic;
signal \N__19470\ : std_logic;
signal \N__19467\ : std_logic;
signal \N__19464\ : std_logic;
signal \N__19461\ : std_logic;
signal \N__19458\ : std_logic;
signal \N__19455\ : std_logic;
signal \N__19452\ : std_logic;
signal \N__19449\ : std_logic;
signal \N__19446\ : std_logic;
signal \N__19443\ : std_logic;
signal \N__19442\ : std_logic;
signal \N__19439\ : std_logic;
signal \N__19438\ : std_logic;
signal \N__19435\ : std_logic;
signal \N__19432\ : std_logic;
signal \N__19429\ : std_logic;
signal \N__19422\ : std_logic;
signal \N__19419\ : std_logic;
signal \N__19418\ : std_logic;
signal \N__19417\ : std_logic;
signal \N__19414\ : std_logic;
signal \N__19409\ : std_logic;
signal \N__19404\ : std_logic;
signal \N__19401\ : std_logic;
signal \N__19398\ : std_logic;
signal \N__19395\ : std_logic;
signal \N__19392\ : std_logic;
signal \N__19389\ : std_logic;
signal \N__19388\ : std_logic;
signal \N__19387\ : std_logic;
signal \N__19384\ : std_logic;
signal \N__19381\ : std_logic;
signal \N__19378\ : std_logic;
signal \N__19373\ : std_logic;
signal \N__19370\ : std_logic;
signal \N__19365\ : std_logic;
signal \N__19362\ : std_logic;
signal \N__19359\ : std_logic;
signal \N__19356\ : std_logic;
signal \N__19353\ : std_logic;
signal \N__19350\ : std_logic;
signal \N__19349\ : std_logic;
signal \N__19346\ : std_logic;
signal \N__19343\ : std_logic;
signal \N__19340\ : std_logic;
signal \N__19337\ : std_logic;
signal \N__19332\ : std_logic;
signal \N__19329\ : std_logic;
signal \N__19326\ : std_logic;
signal \N__19323\ : std_logic;
signal \N__19322\ : std_logic;
signal \N__19319\ : std_logic;
signal \N__19318\ : std_logic;
signal \N__19315\ : std_logic;
signal \N__19310\ : std_logic;
signal \N__19307\ : std_logic;
signal \N__19302\ : std_logic;
signal \N__19299\ : std_logic;
signal \N__19298\ : std_logic;
signal \N__19295\ : std_logic;
signal \N__19292\ : std_logic;
signal \N__19289\ : std_logic;
signal \N__19284\ : std_logic;
signal \N__19281\ : std_logic;
signal \N__19278\ : std_logic;
signal \N__19277\ : std_logic;
signal \N__19274\ : std_logic;
signal \N__19271\ : std_logic;
signal \N__19268\ : std_logic;
signal \N__19263\ : std_logic;
signal \N__19260\ : std_logic;
signal \N__19257\ : std_logic;
signal \N__19254\ : std_logic;
signal \N__19251\ : std_logic;
signal \N__19248\ : std_logic;
signal \N__19245\ : std_logic;
signal \N__19242\ : std_logic;
signal \N__19239\ : std_logic;
signal \N__19238\ : std_logic;
signal \N__19233\ : std_logic;
signal \N__19232\ : std_logic;
signal \N__19229\ : std_logic;
signal \N__19226\ : std_logic;
signal \N__19221\ : std_logic;
signal \N__19218\ : std_logic;
signal \N__19217\ : std_logic;
signal \N__19214\ : std_logic;
signal \N__19211\ : std_logic;
signal \N__19208\ : std_logic;
signal \N__19203\ : std_logic;
signal \N__19200\ : std_logic;
signal \N__19197\ : std_logic;
signal \N__19196\ : std_logic;
signal \N__19193\ : std_logic;
signal \N__19190\ : std_logic;
signal \N__19187\ : std_logic;
signal \N__19182\ : std_logic;
signal \N__19179\ : std_logic;
signal \N__19176\ : std_logic;
signal \N__19173\ : std_logic;
signal \N__19170\ : std_logic;
signal \N__19167\ : std_logic;
signal \N__19164\ : std_logic;
signal \N__19161\ : std_logic;
signal \N__19158\ : std_logic;
signal \N__19155\ : std_logic;
signal \N__19154\ : std_logic;
signal \N__19151\ : std_logic;
signal \N__19148\ : std_logic;
signal \N__19143\ : std_logic;
signal \N__19140\ : std_logic;
signal \N__19139\ : std_logic;
signal \N__19138\ : std_logic;
signal \N__19135\ : std_logic;
signal \N__19132\ : std_logic;
signal \N__19129\ : std_logic;
signal \N__19122\ : std_logic;
signal \N__19121\ : std_logic;
signal \N__19118\ : std_logic;
signal \N__19115\ : std_logic;
signal \N__19110\ : std_logic;
signal \N__19107\ : std_logic;
signal \N__19104\ : std_logic;
signal \N__19101\ : std_logic;
signal \N__19098\ : std_logic;
signal \N__19095\ : std_logic;
signal \N__19092\ : std_logic;
signal \N__19089\ : std_logic;
signal \N__19088\ : std_logic;
signal \N__19085\ : std_logic;
signal \N__19084\ : std_logic;
signal \N__19081\ : std_logic;
signal \N__19078\ : std_logic;
signal \N__19075\ : std_logic;
signal \N__19070\ : std_logic;
signal \N__19065\ : std_logic;
signal \N__19062\ : std_logic;
signal \N__19059\ : std_logic;
signal \N__19056\ : std_logic;
signal \N__19053\ : std_logic;
signal \N__19050\ : std_logic;
signal \N__19047\ : std_logic;
signal \N__19046\ : std_logic;
signal \N__19045\ : std_logic;
signal \N__19042\ : std_logic;
signal \N__19039\ : std_logic;
signal \N__19036\ : std_logic;
signal \N__19033\ : std_logic;
signal \N__19030\ : std_logic;
signal \N__19023\ : std_logic;
signal \N__19020\ : std_logic;
signal \N__19017\ : std_logic;
signal \N__19014\ : std_logic;
signal \N__19011\ : std_logic;
signal \N__19008\ : std_logic;
signal \N__19007\ : std_logic;
signal \N__19004\ : std_logic;
signal \N__19001\ : std_logic;
signal \N__18996\ : std_logic;
signal \N__18993\ : std_logic;
signal \N__18992\ : std_logic;
signal \N__18989\ : std_logic;
signal \N__18988\ : std_logic;
signal \N__18985\ : std_logic;
signal \N__18982\ : std_logic;
signal \N__18979\ : std_logic;
signal \N__18976\ : std_logic;
signal \N__18969\ : std_logic;
signal \N__18966\ : std_logic;
signal \N__18965\ : std_logic;
signal \N__18962\ : std_logic;
signal \N__18959\ : std_logic;
signal \N__18958\ : std_logic;
signal \N__18955\ : std_logic;
signal \N__18952\ : std_logic;
signal \N__18949\ : std_logic;
signal \N__18944\ : std_logic;
signal \N__18939\ : std_logic;
signal \N__18936\ : std_logic;
signal \N__18933\ : std_logic;
signal \N__18930\ : std_logic;
signal \N__18927\ : std_logic;
signal \N__18926\ : std_logic;
signal \N__18925\ : std_logic;
signal \N__18922\ : std_logic;
signal \N__18919\ : std_logic;
signal \N__18916\ : std_logic;
signal \N__18909\ : std_logic;
signal \N__18906\ : std_logic;
signal \N__18903\ : std_logic;
signal \N__18902\ : std_logic;
signal \N__18899\ : std_logic;
signal \N__18898\ : std_logic;
signal \N__18895\ : std_logic;
signal \N__18892\ : std_logic;
signal \N__18889\ : std_logic;
signal \N__18886\ : std_logic;
signal \N__18879\ : std_logic;
signal \N__18876\ : std_logic;
signal \N__18875\ : std_logic;
signal \N__18872\ : std_logic;
signal \N__18869\ : std_logic;
signal \N__18868\ : std_logic;
signal \N__18865\ : std_logic;
signal \N__18862\ : std_logic;
signal \N__18859\ : std_logic;
signal \N__18854\ : std_logic;
signal \N__18849\ : std_logic;
signal \N__18846\ : std_logic;
signal \N__18843\ : std_logic;
signal \N__18842\ : std_logic;
signal \N__18841\ : std_logic;
signal \N__18838\ : std_logic;
signal \N__18835\ : std_logic;
signal \N__18832\ : std_logic;
signal \N__18827\ : std_logic;
signal \N__18822\ : std_logic;
signal \N__18819\ : std_logic;
signal \N__18818\ : std_logic;
signal \N__18815\ : std_logic;
signal \N__18814\ : std_logic;
signal \N__18811\ : std_logic;
signal \N__18808\ : std_logic;
signal \N__18805\ : std_logic;
signal \N__18802\ : std_logic;
signal \N__18795\ : std_logic;
signal \N__18792\ : std_logic;
signal \N__18789\ : std_logic;
signal \N__18788\ : std_logic;
signal \N__18787\ : std_logic;
signal \N__18784\ : std_logic;
signal \N__18781\ : std_logic;
signal \N__18778\ : std_logic;
signal \N__18771\ : std_logic;
signal \N__18768\ : std_logic;
signal \N__18765\ : std_logic;
signal \N__18764\ : std_logic;
signal \N__18763\ : std_logic;
signal \N__18760\ : std_logic;
signal \N__18757\ : std_logic;
signal \N__18754\ : std_logic;
signal \N__18747\ : std_logic;
signal \N__18744\ : std_logic;
signal \N__18743\ : std_logic;
signal \N__18740\ : std_logic;
signal \N__18739\ : std_logic;
signal \N__18736\ : std_logic;
signal \N__18733\ : std_logic;
signal \N__18730\ : std_logic;
signal \N__18727\ : std_logic;
signal \N__18720\ : std_logic;
signal \N__18717\ : std_logic;
signal \N__18714\ : std_logic;
signal \N__18711\ : std_logic;
signal \N__18710\ : std_logic;
signal \N__18707\ : std_logic;
signal \N__18706\ : std_logic;
signal \N__18703\ : std_logic;
signal \N__18700\ : std_logic;
signal \N__18697\ : std_logic;
signal \N__18694\ : std_logic;
signal \N__18687\ : std_logic;
signal \N__18684\ : std_logic;
signal \N__18681\ : std_logic;
signal \N__18680\ : std_logic;
signal \N__18677\ : std_logic;
signal \N__18676\ : std_logic;
signal \N__18673\ : std_logic;
signal \N__18670\ : std_logic;
signal \N__18667\ : std_logic;
signal \N__18664\ : std_logic;
signal \N__18657\ : std_logic;
signal \N__18654\ : std_logic;
signal \N__18651\ : std_logic;
signal \N__18650\ : std_logic;
signal \N__18649\ : std_logic;
signal \N__18646\ : std_logic;
signal \N__18643\ : std_logic;
signal \N__18640\ : std_logic;
signal \N__18635\ : std_logic;
signal \N__18630\ : std_logic;
signal \N__18627\ : std_logic;
signal \N__18624\ : std_logic;
signal \N__18621\ : std_logic;
signal \N__18620\ : std_logic;
signal \N__18617\ : std_logic;
signal \N__18616\ : std_logic;
signal \N__18613\ : std_logic;
signal \N__18610\ : std_logic;
signal \N__18607\ : std_logic;
signal \N__18604\ : std_logic;
signal \N__18597\ : std_logic;
signal \N__18594\ : std_logic;
signal \N__18591\ : std_logic;
signal \N__18590\ : std_logic;
signal \N__18589\ : std_logic;
signal \N__18586\ : std_logic;
signal \N__18583\ : std_logic;
signal \N__18580\ : std_logic;
signal \N__18577\ : std_logic;
signal \N__18570\ : std_logic;
signal \N__18567\ : std_logic;
signal \N__18564\ : std_logic;
signal \N__18563\ : std_logic;
signal \N__18560\ : std_logic;
signal \N__18559\ : std_logic;
signal \N__18556\ : std_logic;
signal \N__18553\ : std_logic;
signal \N__18550\ : std_logic;
signal \N__18547\ : std_logic;
signal \N__18540\ : std_logic;
signal \N__18537\ : std_logic;
signal \N__18534\ : std_logic;
signal \N__18533\ : std_logic;
signal \N__18532\ : std_logic;
signal \N__18529\ : std_logic;
signal \N__18526\ : std_logic;
signal \N__18523\ : std_logic;
signal \N__18520\ : std_logic;
signal \N__18513\ : std_logic;
signal \N__18510\ : std_logic;
signal \N__18509\ : std_logic;
signal \N__18506\ : std_logic;
signal \N__18505\ : std_logic;
signal \N__18502\ : std_logic;
signal \N__18499\ : std_logic;
signal \N__18496\ : std_logic;
signal \N__18493\ : std_logic;
signal \N__18486\ : std_logic;
signal \N__18483\ : std_logic;
signal \N__18480\ : std_logic;
signal \N__18477\ : std_logic;
signal \N__18474\ : std_logic;
signal \N__18471\ : std_logic;
signal \N__18468\ : std_logic;
signal \N__18467\ : std_logic;
signal \N__18462\ : std_logic;
signal \N__18459\ : std_logic;
signal \N__18456\ : std_logic;
signal \N__18453\ : std_logic;
signal \N__18450\ : std_logic;
signal \N__18447\ : std_logic;
signal \N__18444\ : std_logic;
signal \N__18441\ : std_logic;
signal \N__18438\ : std_logic;
signal \N__18435\ : std_logic;
signal \N__18432\ : std_logic;
signal \N__18429\ : std_logic;
signal \N__18426\ : std_logic;
signal \N__18423\ : std_logic;
signal \N__18420\ : std_logic;
signal \N__18417\ : std_logic;
signal \N__18414\ : std_logic;
signal \N__18411\ : std_logic;
signal \N__18408\ : std_logic;
signal \N__18405\ : std_logic;
signal \N__18402\ : std_logic;
signal \N__18399\ : std_logic;
signal \N__18396\ : std_logic;
signal \N__18393\ : std_logic;
signal \N__18390\ : std_logic;
signal \N__18387\ : std_logic;
signal \N__18384\ : std_logic;
signal \N__18381\ : std_logic;
signal \N__18378\ : std_logic;
signal \N__18375\ : std_logic;
signal \N__18372\ : std_logic;
signal \N__18369\ : std_logic;
signal \N__18366\ : std_logic;
signal \N__18363\ : std_logic;
signal \N__18360\ : std_logic;
signal \N__18357\ : std_logic;
signal \N__18354\ : std_logic;
signal \N__18351\ : std_logic;
signal \N__18348\ : std_logic;
signal \N__18347\ : std_logic;
signal \N__18342\ : std_logic;
signal \N__18339\ : std_logic;
signal \N__18336\ : std_logic;
signal \N__18333\ : std_logic;
signal \N__18330\ : std_logic;
signal \N__18327\ : std_logic;
signal \N__18324\ : std_logic;
signal \N__18321\ : std_logic;
signal \N__18318\ : std_logic;
signal \N__18315\ : std_logic;
signal \N__18312\ : std_logic;
signal \N__18309\ : std_logic;
signal \N__18306\ : std_logic;
signal \N__18303\ : std_logic;
signal \N__18300\ : std_logic;
signal \N__18297\ : std_logic;
signal \N__18294\ : std_logic;
signal \N__18291\ : std_logic;
signal \N__18288\ : std_logic;
signal \N__18285\ : std_logic;
signal \N__18282\ : std_logic;
signal \N__18279\ : std_logic;
signal \N__18276\ : std_logic;
signal \N__18273\ : std_logic;
signal \N__18270\ : std_logic;
signal \N__18267\ : std_logic;
signal \N__18264\ : std_logic;
signal \N__18261\ : std_logic;
signal \N__18258\ : std_logic;
signal \N__18255\ : std_logic;
signal \N__18252\ : std_logic;
signal \N__18249\ : std_logic;
signal \N__18246\ : std_logic;
signal \N__18243\ : std_logic;
signal \N__18240\ : std_logic;
signal \N__18237\ : std_logic;
signal \N__18234\ : std_logic;
signal \N__18231\ : std_logic;
signal \N__18228\ : std_logic;
signal \N__18225\ : std_logic;
signal \N__18222\ : std_logic;
signal \N__18219\ : std_logic;
signal \N__18216\ : std_logic;
signal \N__18213\ : std_logic;
signal \N__18210\ : std_logic;
signal \N__18207\ : std_logic;
signal \N__18204\ : std_logic;
signal \N__18201\ : std_logic;
signal \N__18198\ : std_logic;
signal \N__18195\ : std_logic;
signal \N__18192\ : std_logic;
signal \N__18189\ : std_logic;
signal \N__18186\ : std_logic;
signal \N__18183\ : std_logic;
signal \N__18180\ : std_logic;
signal \N__18177\ : std_logic;
signal \N__18174\ : std_logic;
signal \N__18171\ : std_logic;
signal \N__18168\ : std_logic;
signal \N__18165\ : std_logic;
signal \N__18162\ : std_logic;
signal \N__18159\ : std_logic;
signal \N__18156\ : std_logic;
signal \N__18153\ : std_logic;
signal \N__18150\ : std_logic;
signal \N__18147\ : std_logic;
signal \N__18144\ : std_logic;
signal \N__18141\ : std_logic;
signal \N__18138\ : std_logic;
signal \N__18135\ : std_logic;
signal \N__18132\ : std_logic;
signal \N__18129\ : std_logic;
signal \N__18126\ : std_logic;
signal \N__18123\ : std_logic;
signal \N__18120\ : std_logic;
signal \N__18117\ : std_logic;
signal \N__18114\ : std_logic;
signal \N__18111\ : std_logic;
signal \N__18108\ : std_logic;
signal \N__18105\ : std_logic;
signal \N__18102\ : std_logic;
signal \N__18099\ : std_logic;
signal \N__18096\ : std_logic;
signal \N__18093\ : std_logic;
signal \N__18090\ : std_logic;
signal \N__18087\ : std_logic;
signal \N__18084\ : std_logic;
signal \N__18081\ : std_logic;
signal \N__18078\ : std_logic;
signal \N__18075\ : std_logic;
signal \N__18072\ : std_logic;
signal \N__18069\ : std_logic;
signal \N__18066\ : std_logic;
signal \N__18063\ : std_logic;
signal \N__18060\ : std_logic;
signal \N__18057\ : std_logic;
signal \N__18054\ : std_logic;
signal \N__18051\ : std_logic;
signal \N__18048\ : std_logic;
signal \N__18047\ : std_logic;
signal \N__18042\ : std_logic;
signal \N__18039\ : std_logic;
signal \N__18038\ : std_logic;
signal \N__18033\ : std_logic;
signal \N__18030\ : std_logic;
signal \N__18027\ : std_logic;
signal \N__18024\ : std_logic;
signal \N__18021\ : std_logic;
signal \N__18018\ : std_logic;
signal \N__18015\ : std_logic;
signal \N__18012\ : std_logic;
signal \N__18009\ : std_logic;
signal \N__18006\ : std_logic;
signal \N__18003\ : std_logic;
signal \N__18000\ : std_logic;
signal \N__17997\ : std_logic;
signal \N__17994\ : std_logic;
signal \N__17991\ : std_logic;
signal \N__17988\ : std_logic;
signal \N__17985\ : std_logic;
signal \N__17982\ : std_logic;
signal \N__17981\ : std_logic;
signal \N__17976\ : std_logic;
signal \N__17973\ : std_logic;
signal \N__17972\ : std_logic;
signal \N__17967\ : std_logic;
signal \N__17964\ : std_logic;
signal \N__17963\ : std_logic;
signal \N__17958\ : std_logic;
signal \N__17955\ : std_logic;
signal \N__17954\ : std_logic;
signal \N__17949\ : std_logic;
signal \N__17946\ : std_logic;
signal \N__17945\ : std_logic;
signal \N__17942\ : std_logic;
signal \N__17939\ : std_logic;
signal \N__17934\ : std_logic;
signal \N__17933\ : std_logic;
signal \N__17928\ : std_logic;
signal \N__17925\ : std_logic;
signal \N__17924\ : std_logic;
signal \N__17921\ : std_logic;
signal \N__17918\ : std_logic;
signal \N__17915\ : std_logic;
signal \N__17910\ : std_logic;
signal \N__17907\ : std_logic;
signal \N__17904\ : std_logic;
signal \N__17901\ : std_logic;
signal \N__17900\ : std_logic;
signal \N__17897\ : std_logic;
signal \N__17894\ : std_logic;
signal \N__17891\ : std_logic;
signal \N__17886\ : std_logic;
signal \N__17883\ : std_logic;
signal \N__17880\ : std_logic;
signal \N__17877\ : std_logic;
signal \N__17874\ : std_logic;
signal \N__17871\ : std_logic;
signal \N__17868\ : std_logic;
signal \N__17865\ : std_logic;
signal \N__17862\ : std_logic;
signal \N__17861\ : std_logic;
signal \N__17858\ : std_logic;
signal \N__17855\ : std_logic;
signal \N__17852\ : std_logic;
signal \N__17847\ : std_logic;
signal \N__17844\ : std_logic;
signal \N__17841\ : std_logic;
signal \N__17840\ : std_logic;
signal \N__17837\ : std_logic;
signal \N__17834\ : std_logic;
signal \N__17831\ : std_logic;
signal \N__17826\ : std_logic;
signal \N__17823\ : std_logic;
signal \N__17820\ : std_logic;
signal \N__17817\ : std_logic;
signal \N__17816\ : std_logic;
signal \N__17813\ : std_logic;
signal \N__17810\ : std_logic;
signal \N__17807\ : std_logic;
signal \N__17802\ : std_logic;
signal \N__17799\ : std_logic;
signal \N__17798\ : std_logic;
signal \N__17795\ : std_logic;
signal \N__17792\ : std_logic;
signal \N__17789\ : std_logic;
signal \N__17784\ : std_logic;
signal \N__17781\ : std_logic;
signal \N__17780\ : std_logic;
signal \N__17777\ : std_logic;
signal \N__17774\ : std_logic;
signal \N__17771\ : std_logic;
signal \N__17766\ : std_logic;
signal \N__17763\ : std_logic;
signal \N__17762\ : std_logic;
signal \N__17759\ : std_logic;
signal \N__17756\ : std_logic;
signal \N__17753\ : std_logic;
signal \N__17748\ : std_logic;
signal \N__17745\ : std_logic;
signal \N__17744\ : std_logic;
signal \N__17741\ : std_logic;
signal \N__17738\ : std_logic;
signal \N__17735\ : std_logic;
signal \N__17730\ : std_logic;
signal \N__17727\ : std_logic;
signal \N__17726\ : std_logic;
signal \N__17723\ : std_logic;
signal \N__17720\ : std_logic;
signal \N__17717\ : std_logic;
signal \N__17712\ : std_logic;
signal \N__17709\ : std_logic;
signal \N__17706\ : std_logic;
signal \N__17703\ : std_logic;
signal \N__17700\ : std_logic;
signal \N__17699\ : std_logic;
signal \N__17696\ : std_logic;
signal \N__17693\ : std_logic;
signal \N__17688\ : std_logic;
signal \N__17685\ : std_logic;
signal \N__17684\ : std_logic;
signal \N__17681\ : std_logic;
signal \N__17678\ : std_logic;
signal \N__17675\ : std_logic;
signal \N__17670\ : std_logic;
signal \N__17667\ : std_logic;
signal \N__17666\ : std_logic;
signal \N__17663\ : std_logic;
signal \N__17660\ : std_logic;
signal \N__17655\ : std_logic;
signal \N__17652\ : std_logic;
signal \N__17651\ : std_logic;
signal \N__17648\ : std_logic;
signal \N__17645\ : std_logic;
signal \N__17640\ : std_logic;
signal \N__17637\ : std_logic;
signal \N__17636\ : std_logic;
signal \N__17633\ : std_logic;
signal \N__17630\ : std_logic;
signal \N__17625\ : std_logic;
signal \N__17622\ : std_logic;
signal \N__17621\ : std_logic;
signal \N__17618\ : std_logic;
signal \N__17615\ : std_logic;
signal \N__17610\ : std_logic;
signal \N__17607\ : std_logic;
signal \N__17604\ : std_logic;
signal \N__17603\ : std_logic;
signal \N__17600\ : std_logic;
signal \N__17597\ : std_logic;
signal \N__17594\ : std_logic;
signal \N__17589\ : std_logic;
signal \N__17586\ : std_logic;
signal \N__17585\ : std_logic;
signal \N__17582\ : std_logic;
signal \N__17579\ : std_logic;
signal \N__17576\ : std_logic;
signal \N__17571\ : std_logic;
signal \N__17568\ : std_logic;
signal \N__17567\ : std_logic;
signal \N__17564\ : std_logic;
signal \N__17561\ : std_logic;
signal \N__17556\ : std_logic;
signal \N__17555\ : std_logic;
signal \N__17552\ : std_logic;
signal \N__17549\ : std_logic;
signal \N__17544\ : std_logic;
signal \N__17543\ : std_logic;
signal \N__17538\ : std_logic;
signal \N__17535\ : std_logic;
signal \N__17534\ : std_logic;
signal \N__17529\ : std_logic;
signal \N__17526\ : std_logic;
signal \N__17523\ : std_logic;
signal \N__17520\ : std_logic;
signal \N__17517\ : std_logic;
signal \N__17514\ : std_logic;
signal \N__17513\ : std_logic;
signal \N__17510\ : std_logic;
signal \N__17507\ : std_logic;
signal \N__17504\ : std_logic;
signal \N__17499\ : std_logic;
signal \N__17496\ : std_logic;
signal \N__17495\ : std_logic;
signal \N__17490\ : std_logic;
signal \N__17487\ : std_logic;
signal \N__17484\ : std_logic;
signal \N__17481\ : std_logic;
signal \N__17478\ : std_logic;
signal \N__17475\ : std_logic;
signal \N__17472\ : std_logic;
signal \N__17469\ : std_logic;
signal \N__17466\ : std_logic;
signal \N__17463\ : std_logic;
signal \N__17462\ : std_logic;
signal \N__17457\ : std_logic;
signal \N__17454\ : std_logic;
signal \N__17453\ : std_logic;
signal \N__17448\ : std_logic;
signal \N__17445\ : std_logic;
signal \N__17444\ : std_logic;
signal \N__17439\ : std_logic;
signal \N__17436\ : std_logic;
signal \N__17435\ : std_logic;
signal \N__17430\ : std_logic;
signal \N__17427\ : std_logic;
signal \N__17426\ : std_logic;
signal \N__17421\ : std_logic;
signal \N__17418\ : std_logic;
signal \N__17415\ : std_logic;
signal \N__17412\ : std_logic;
signal \N__17409\ : std_logic;
signal \N__17406\ : std_logic;
signal \N__17403\ : std_logic;
signal \CLK_pad_gb_input\ : std_logic;
signal \VCCG0\ : std_logic;
signal neo_pixel_transmitter_t0_0 : std_logic;
signal neo_pixel_transmitter_t0_21 : std_logic;
signal neo_pixel_transmitter_t0_7 : std_logic;
signal neo_pixel_transmitter_t0_12 : std_logic;
signal neo_pixel_transmitter_t0_4 : std_logic;
signal neo_pixel_transmitter_t0_9 : std_logic;
signal neopxl_color_prev_12 : std_logic;
signal \n24_adj_801_cascade_\ : std_logic;
signal n12414 : std_logic;
signal neopxl_color_prev_6 : std_logic;
signal neo_pixel_transmitter_t0_18 : std_logic;
signal neo_pixel_transmitter_t0_20 : std_logic;
signal neo_pixel_transmitter_t0_24 : std_logic;
signal neo_pixel_transmitter_t0_31 : std_logic;
signal n15_adj_841 : std_logic;
signal n14_adj_842 : std_logic;
signal delay_counter_0 : std_logic;
signal \bfn_1_22_0_\ : std_logic;
signal delay_counter_1 : std_logic;
signal n10582 : std_logic;
signal delay_counter_2 : std_logic;
signal n10583 : std_logic;
signal delay_counter_3 : std_logic;
signal n10584 : std_logic;
signal delay_counter_4 : std_logic;
signal n10585 : std_logic;
signal delay_counter_5 : std_logic;
signal n10586 : std_logic;
signal delay_counter_6 : std_logic;
signal n10587 : std_logic;
signal delay_counter_7 : std_logic;
signal n10588 : std_logic;
signal n10589 : std_logic;
signal delay_counter_8 : std_logic;
signal \bfn_1_23_0_\ : std_logic;
signal delay_counter_9 : std_logic;
signal n10590 : std_logic;
signal delay_counter_10 : std_logic;
signal n10591 : std_logic;
signal delay_counter_11 : std_logic;
signal n10592 : std_logic;
signal delay_counter_12 : std_logic;
signal n10593 : std_logic;
signal delay_counter_13 : std_logic;
signal n10594 : std_logic;
signal delay_counter_14 : std_logic;
signal n10595 : std_logic;
signal n10596 : std_logic;
signal n10597 : std_logic;
signal \bfn_1_24_0_\ : std_logic;
signal n10598 : std_logic;
signal n10599 : std_logic;
signal n10600 : std_logic;
signal n10601 : std_logic;
signal n10602 : std_logic;
signal n10603 : std_logic;
signal delay_counter_23 : std_logic;
signal n10604 : std_logic;
signal n10605 : std_logic;
signal \bfn_1_25_0_\ : std_logic;
signal delay_counter_25 : std_logic;
signal n10606 : std_logic;
signal n10607 : std_logic;
signal delay_counter_27 : std_logic;
signal n10608 : std_logic;
signal n10609 : std_logic;
signal n10610 : std_logic;
signal delay_counter_30 : std_logic;
signal n10611 : std_logic;
signal n10612 : std_logic;
signal neo_pixel_transmitter_t0_23 : std_logic;
signal neo_pixel_transmitter_t0_15 : std_logic;
signal neo_pixel_transmitter_t0_8 : std_logic;
signal neo_pixel_transmitter_t0_2 : std_logic;
signal neo_pixel_transmitter_t0_6 : std_logic;
signal neo_pixel_transmitter_t0_17 : std_logic;
signal neo_pixel_transmitter_t0_22 : std_logic;
signal neo_pixel_transmitter_t0_10 : std_logic;
signal \nx.n33\ : std_logic;
signal \bfn_2_19_0_\ : std_logic;
signal \nx.n10669\ : std_logic;
signal \nx.n31_adj_711\ : std_logic;
signal \nx.n10670\ : std_logic;
signal \nx.n10671\ : std_logic;
signal \nx.n29_adj_714\ : std_logic;
signal \nx.n10672\ : std_logic;
signal \nx.n10673\ : std_logic;
signal \nx.n27_adj_720\ : std_logic;
signal \nx.n10674\ : std_logic;
signal \nx.n26_adj_722\ : std_logic;
signal \nx.n10675\ : std_logic;
signal \nx.n10676\ : std_logic;
signal \nx.n25_adj_724\ : std_logic;
signal \bfn_2_20_0_\ : std_logic;
signal \nx.n24_adj_734\ : std_logic;
signal \nx.n10677\ : std_logic;
signal \nx.n23\ : std_logic;
signal \nx.n10678\ : std_logic;
signal \nx.n10679\ : std_logic;
signal \nx.one_wire_N_599_11\ : std_logic;
signal \nx.n21_adj_737\ : std_logic;
signal \nx.n10680\ : std_logic;
signal \nx.n13173\ : std_logic;
signal \nx.n10681\ : std_logic;
signal \nx.n13175\ : std_logic;
signal \nx.n10682\ : std_logic;
signal \nx.n10683\ : std_logic;
signal \nx.n10683_THRU_CRY_0_THRU_CO\ : std_logic;
signal \nx.n13177\ : std_logic;
signal \nx.n18_adj_723\ : std_logic;
signal \bfn_2_21_0_\ : std_logic;
signal \nx.n13179\ : std_logic;
signal \nx.n10684\ : std_logic;
signal \nx.n13181\ : std_logic;
signal \nx.n16_adj_672\ : std_logic;
signal \nx.n10685\ : std_logic;
signal \nx.n13183\ : std_logic;
signal \nx.n15\ : std_logic;
signal \nx.n10686\ : std_logic;
signal \nx.n13185\ : std_logic;
signal \nx.n10687\ : std_logic;
signal \nx.n13187\ : std_logic;
signal \nx.n13\ : std_logic;
signal \nx.n10688\ : std_logic;
signal \nx.n10689\ : std_logic;
signal \nx.n10689_THRU_CRY_0_THRU_CO\ : std_logic;
signal \nx.n10689_THRU_CRY_1_THRU_CO\ : std_logic;
signal \nx.n13189\ : std_logic;
signal \nx.n12\ : std_logic;
signal \bfn_2_22_0_\ : std_logic;
signal \nx.n13191\ : std_logic;
signal \nx.n11\ : std_logic;
signal \nx.n10690\ : std_logic;
signal \nx.n13193\ : std_logic;
signal \nx.n10\ : std_logic;
signal \nx.n10691\ : std_logic;
signal \nx.n13195\ : std_logic;
signal \nx.n9\ : std_logic;
signal \nx.n10692\ : std_logic;
signal \nx.n13197\ : std_logic;
signal \nx.n10693\ : std_logic;
signal \nx.n13199\ : std_logic;
signal \nx.n10694\ : std_logic;
signal \nx.n10695\ : std_logic;
signal \GNDG0\ : std_logic;
signal \nx.n10695_THRU_CRY_0_THRU_CO\ : std_logic;
signal \nx.n10695_THRU_CRY_1_THRU_CO\ : std_logic;
signal \nx.n13201\ : std_logic;
signal \bfn_2_23_0_\ : std_logic;
signal \nx.n13203\ : std_logic;
signal \nx.n10696\ : std_logic;
signal \nx.n13205\ : std_logic;
signal \nx.n4_adj_710\ : std_logic;
signal \nx.n10697\ : std_logic;
signal \nx.n13207\ : std_logic;
signal \nx.n10698\ : std_logic;
signal \nx.n2\ : std_logic;
signal \nx.n13209\ : std_logic;
signal \nx.n10699\ : std_logic;
signal \nx.n6\ : std_logic;
signal neo_pixel_transmitter_t0_27 : std_logic;
signal \bfn_2_25_0_\ : std_logic;
signal \nx.n10773\ : std_logic;
signal \nx.n10774\ : std_logic;
signal \nx.n10775\ : std_logic;
signal \nx.n10776\ : std_logic;
signal \nx.n10777\ : std_logic;
signal \nx.n10778\ : std_logic;
signal \nx.n10779\ : std_logic;
signal \nx.n10780\ : std_logic;
signal \bfn_2_26_0_\ : std_logic;
signal \nx.n10781\ : std_logic;
signal \nx.n10782\ : std_logic;
signal \nx.n1469\ : std_logic;
signal neo_pixel_transmitter_t0_14 : std_logic;
signal \nx.n19_adj_725\ : std_logic;
signal \nx.n11834_cascade_\ : std_logic;
signal timer_0 : std_logic;
signal \bfn_3_18_0_\ : std_logic;
signal \nx.n10707\ : std_logic;
signal timer_2 : std_logic;
signal \nx.n10708\ : std_logic;
signal \nx.n10709\ : std_logic;
signal timer_4 : std_logic;
signal \nx.n10710\ : std_logic;
signal \nx.n10711\ : std_logic;
signal timer_6 : std_logic;
signal \nx.n10712\ : std_logic;
signal timer_7 : std_logic;
signal \nx.n10713\ : std_logic;
signal \nx.n10714\ : std_logic;
signal timer_8 : std_logic;
signal \bfn_3_19_0_\ : std_logic;
signal timer_9 : std_logic;
signal \nx.n10715\ : std_logic;
signal timer_10 : std_logic;
signal \nx.n10716\ : std_logic;
signal \nx.n10717\ : std_logic;
signal timer_12 : std_logic;
signal \nx.n10718\ : std_logic;
signal \nx.n10719\ : std_logic;
signal timer_14 : std_logic;
signal \nx.n10720\ : std_logic;
signal timer_15 : std_logic;
signal \nx.n10721\ : std_logic;
signal \nx.n10722\ : std_logic;
signal \bfn_3_20_0_\ : std_logic;
signal timer_17 : std_logic;
signal \nx.n10723\ : std_logic;
signal timer_18 : std_logic;
signal \nx.n10724\ : std_logic;
signal \nx.n10725\ : std_logic;
signal timer_20 : std_logic;
signal \nx.n10726\ : std_logic;
signal timer_21 : std_logic;
signal \nx.n10727\ : std_logic;
signal timer_22 : std_logic;
signal \nx.n10728\ : std_logic;
signal timer_23 : std_logic;
signal \nx.n10729\ : std_logic;
signal \nx.n10730\ : std_logic;
signal timer_24 : std_logic;
signal \bfn_3_21_0_\ : std_logic;
signal \nx.n10731\ : std_logic;
signal \nx.n10732\ : std_logic;
signal timer_27 : std_logic;
signal \nx.n10733\ : std_logic;
signal \nx.n10734\ : std_logic;
signal \nx.n10735\ : std_logic;
signal \nx.n10736\ : std_logic;
signal \nx.n10737\ : std_logic;
signal timer_31 : std_logic;
signal \n11826_cascade_\ : std_logic;
signal pin_oe_1 : std_logic;
signal delay_counter_17 : std_logic;
signal delay_counter_15 : std_logic;
signal n12382 : std_logic;
signal \n11828_cascade_\ : std_logic;
signal pin_oe_5 : std_logic;
signal timer_16 : std_logic;
signal neo_pixel_transmitter_t0_16 : std_logic;
signal \nx.n17\ : std_logic;
signal \nx.n1309_cascade_\ : std_logic;
signal delay_counter_21 : std_logic;
signal delay_counter_29 : std_logic;
signal n12379 : std_logic;
signal \nx.n12_adj_669\ : std_logic;
signal \nx.n1308_cascade_\ : std_logic;
signal \nx.n1334_cascade_\ : std_logic;
signal \nx.n1403_cascade_\ : std_logic;
signal \nx.n1402\ : std_logic;
signal \nx.n16_adj_727_cascade_\ : std_logic;
signal \nx.n1471\ : std_logic;
signal \nx.n1473\ : std_logic;
signal \nx.n1406\ : std_logic;
signal \nx.n1404\ : std_logic;
signal \nx.n13_adj_729\ : std_logic;
signal \nx.n18_adj_728\ : std_logic;
signal \nx.n1405\ : std_logic;
signal \nx.n1433_cascade_\ : std_logic;
signal \nx.n1472\ : std_logic;
signal \nx.n1470\ : std_logic;
signal \nx.n1403\ : std_logic;
signal \nx.n1502_cascade_\ : std_logic;
signal \nx.n1474\ : std_logic;
signal \nx.n1407\ : std_logic;
signal \nx.n1476\ : std_logic;
signal \nx.n1409\ : std_logic;
signal \nx.n1468\ : std_logic;
signal \nx.n1475\ : std_logic;
signal \nx.n1408\ : std_logic;
signal \nx.n1507_cascade_\ : std_logic;
signal \nx.n18_adj_731_cascade_\ : std_logic;
signal \nx.n20_adj_733_cascade_\ : std_logic;
signal \nx.n16_adj_732\ : std_logic;
signal \nx.n1532_cascade_\ : std_logic;
signal \nx.n1477\ : std_logic;
signal \nx.n1433\ : std_logic;
signal \nx.n1509_cascade_\ : std_logic;
signal \nx.n9729\ : std_logic;
signal \nx.n46_adj_779\ : std_logic;
signal \nx.n3\ : std_logic;
signal \nx.n7_adj_764_cascade_\ : std_logic;
signal \nx.n11864_cascade_\ : std_logic;
signal \nx.n7_adj_667\ : std_logic;
signal \nx.n103\ : std_logic;
signal \nx.n11892\ : std_logic;
signal \nx.n30_adj_712\ : std_logic;
signal \nx.n32\ : std_logic;
signal \nx.n28_adj_715\ : std_logic;
signal timer_5 : std_logic;
signal neo_pixel_transmitter_t0_5 : std_logic;
signal timer_1 : std_logic;
signal neo_pixel_transmitter_t0_1 : std_logic;
signal timer_3 : std_logic;
signal neo_pixel_transmitter_t0_3 : std_logic;
signal \nx.n16_adj_785\ : std_logic;
signal \nx.one_wire_N_599_4\ : std_logic;
signal \nx.n6_adj_786_cascade_\ : std_logic;
signal \nx.one_wire_N_599_5\ : std_logic;
signal \nx.n13659\ : std_logic;
signal \nx.one_wire_N_599_7\ : std_logic;
signal \nx.one_wire_N_599_8\ : std_logic;
signal \nx.one_wire_N_599_6\ : std_logic;
signal \nx.n13211\ : std_logic;
signal \nx.one_wire_N_599_10\ : std_logic;
signal \nx.one_wire_N_599_9\ : std_logic;
signal \nx.n13217_cascade_\ : std_logic;
signal \nx.n7608\ : std_logic;
signal \nx.n20_adj_726\ : std_logic;
signal timer_13 : std_logic;
signal neo_pixel_transmitter_t0_13 : std_logic;
signal timer_25 : std_logic;
signal timer_19 : std_logic;
signal pin_in_7 : std_logic;
signal pin_in_6 : std_logic;
signal timer_29 : std_logic;
signal neo_pixel_transmitter_t0_29 : std_logic;
signal neo_pixel_transmitter_t0_25 : std_logic;
signal \nx.n8\ : std_logic;
signal \nx.n1205_cascade_\ : std_logic;
signal \nx.n11_adj_674\ : std_logic;
signal \nx.n1235_cascade_\ : std_logic;
signal \nx.n1203_cascade_\ : std_logic;
signal \nx.n13_adj_675\ : std_logic;
signal \nx.n1377\ : std_logic;
signal \bfn_4_23_0_\ : std_logic;
signal \nx.n1309\ : std_logic;
signal \nx.n1376\ : std_logic;
signal \nx.n10764\ : std_logic;
signal \nx.n1308\ : std_logic;
signal \nx.n1375\ : std_logic;
signal \nx.n10765\ : std_logic;
signal \nx.n1374\ : std_logic;
signal \nx.n10766\ : std_logic;
signal \nx.n1306\ : std_logic;
signal \nx.n1373\ : std_logic;
signal \nx.n10767\ : std_logic;
signal \nx.n1372\ : std_logic;
signal \nx.n10768\ : std_logic;
signal \nx.n1371\ : std_logic;
signal \nx.n10769\ : std_logic;
signal \nx.n1303\ : std_logic;
signal \nx.n1370\ : std_logic;
signal \nx.n10770\ : std_logic;
signal \nx.n10771\ : std_logic;
signal \bfn_4_24_0_\ : std_logic;
signal \nx.n10772\ : std_logic;
signal \nx.n1400\ : std_logic;
signal delay_counter_18 : std_logic;
signal delay_counter_16 : std_logic;
signal n6_adj_843 : std_logic;
signal \nx.n1304\ : std_logic;
signal \nx.n1305\ : std_logic;
signal \nx.n10_adj_668_cascade_\ : std_logic;
signal \nx.n1307\ : std_logic;
signal \nx.n16\ : std_logic;
signal \nx.n1369\ : std_logic;
signal \nx.n1334\ : std_logic;
signal \nx.n1401\ : std_logic;
signal n22_adj_795 : std_logic;
signal \nx.n1631_cascade_\ : std_logic;
signal \nx.n15_adj_676_cascade_\ : std_logic;
signal \nx.n22\ : std_logic;
signal \nx.n47_adj_780\ : std_logic;
signal \nx.n18\ : std_logic;
signal delay_counter_28 : std_logic;
signal delay_counter_24 : std_logic;
signal delay_counter_22 : std_logic;
signal delay_counter_26 : std_logic;
signal \bfn_4_26_0_\ : std_logic;
signal \nx.n1509\ : std_logic;
signal \nx.n13604\ : std_logic;
signal \nx.n10783\ : std_logic;
signal \nx.n1508\ : std_logic;
signal \nx.n10784\ : std_logic;
signal \nx.n1507\ : std_logic;
signal \nx.n10785\ : std_logic;
signal \nx.n1506\ : std_logic;
signal \nx.n10786\ : std_logic;
signal \nx.n1505\ : std_logic;
signal \nx.n10787\ : std_logic;
signal \nx.n1504\ : std_logic;
signal \nx.n10788\ : std_logic;
signal \nx.n1503\ : std_logic;
signal \nx.n10789\ : std_logic;
signal \nx.n10790\ : std_logic;
signal \nx.n1502\ : std_logic;
signal \bfn_4_27_0_\ : std_logic;
signal \nx.n1501\ : std_logic;
signal \nx.n10791\ : std_logic;
signal \nx.n1500\ : std_logic;
signal \nx.n10792\ : std_logic;
signal \nx.n1499\ : std_logic;
signal \nx.n1532\ : std_logic;
signal \nx.n10793\ : std_logic;
signal \nx.n45_adj_781\ : std_logic;
signal \nx.n19\ : std_logic;
signal pin_in_10 : std_logic;
signal pin_in_11 : std_logic;
signal pin_oe_6 : std_logic;
signal pin_in_9 : std_logic;
signal pin_in_8 : std_logic;
signal n13649 : std_logic;
signal timer_30 : std_logic;
signal neo_pixel_transmitter_t0_30 : std_logic;
signal \nx.n11946\ : std_logic;
signal \nx.n13445\ : std_logic;
signal \nx.n11948_cascade_\ : std_logic;
signal pin_in_2 : std_logic;
signal pin_in_3 : std_logic;
signal \n13379_cascade_\ : std_logic;
signal \nx.n13438\ : std_logic;
signal \nx.one_wire_N_599_3\ : std_logic;
signal \nx.n11908_cascade_\ : std_logic;
signal \nx.n11926\ : std_logic;
signal \nx.n11926_cascade_\ : std_logic;
signal \n7671_cascade_\ : std_logic;
signal \nx.one_wire_N_599_2\ : std_logic;
signal \nx.n4_adj_771\ : std_logic;
signal \nx.n9747\ : std_logic;
signal \nx.n12381\ : std_logic;
signal timer_11 : std_logic;
signal pin_in_0 : std_logic;
signal pin_in_1 : std_logic;
signal n13378 : std_logic;
signal pin_in_4 : std_logic;
signal pin_in_5 : std_logic;
signal n13382 : std_logic;
signal \n13381_cascade_\ : std_logic;
signal n13613 : std_logic;
signal neo_pixel_transmitter_t0_11 : std_logic;
signal \nx.n22_adj_749\ : std_logic;
signal neo_pixel_transmitter_t0_19 : std_logic;
signal \nx.n14\ : std_logic;
signal \nx.n1109_cascade_\ : std_logic;
signal \nx.n9737_cascade_\ : std_logic;
signal \nx.n12_adj_673_cascade_\ : std_logic;
signal \nx.n1177\ : std_logic;
signal \bfn_5_21_0_\ : std_logic;
signal \nx.n1109\ : std_logic;
signal \nx.n1176\ : std_logic;
signal \nx.n10749\ : std_logic;
signal \nx.n1108\ : std_logic;
signal \nx.n1175\ : std_logic;
signal \nx.n10750\ : std_logic;
signal \nx.n1174\ : std_logic;
signal \nx.n10751\ : std_logic;
signal \nx.n1106\ : std_logic;
signal \nx.n1173\ : std_logic;
signal \nx.n10752\ : std_logic;
signal \nx.n1172\ : std_logic;
signal \nx.n10753\ : std_logic;
signal \nx.n1104\ : std_logic;
signal \nx.n1171\ : std_logic;
signal \nx.n10754\ : std_logic;
signal \nx.n1136\ : std_logic;
signal \nx.n10755\ : std_logic;
signal \nx.n1277\ : std_logic;
signal \bfn_5_22_0_\ : std_logic;
signal \nx.n1209\ : std_logic;
signal \nx.n1276\ : std_logic;
signal \nx.n10756\ : std_logic;
signal \nx.n1208\ : std_logic;
signal \nx.n1275\ : std_logic;
signal \nx.n10757\ : std_logic;
signal \nx.n1207\ : std_logic;
signal \nx.n1274\ : std_logic;
signal \nx.n10758\ : std_logic;
signal \nx.n1206\ : std_logic;
signal \nx.n1273\ : std_logic;
signal \nx.n10759\ : std_logic;
signal \nx.n1205\ : std_logic;
signal \nx.n1272\ : std_logic;
signal \nx.n10760\ : std_logic;
signal \nx.n1204\ : std_logic;
signal \nx.n1271\ : std_logic;
signal \nx.n10761\ : std_logic;
signal \nx.n10762\ : std_logic;
signal \nx.n10763\ : std_logic;
signal \nx.n1202\ : std_logic;
signal \bfn_5_23_0_\ : std_logic;
signal \nx.n1301\ : std_logic;
signal delay_counter_19 : std_logic;
signal delay_counter_20 : std_logic;
signal n4 : std_logic;
signal \nx.n1203\ : std_logic;
signal \nx.n1235\ : std_logic;
signal \nx.n1270\ : std_logic;
signal \nx.n1302\ : std_logic;
signal \nx.n49_adj_784_cascade_\ : std_logic;
signal \nx.n54\ : std_logic;
signal n7664 : std_logic;
signal \nx.n30_adj_777_cascade_\ : std_logic;
signal \nx.n43_adj_783\ : std_logic;
signal \bfn_5_25_0_\ : std_logic;
signal \nx.n1609\ : std_logic;
signal \nx.n13602\ : std_logic;
signal \nx.n10794\ : std_logic;
signal \nx.n1608\ : std_logic;
signal \nx.n10795\ : std_logic;
signal \nx.n1607\ : std_logic;
signal \nx.n10796\ : std_logic;
signal \nx.n1606\ : std_logic;
signal \nx.n10797\ : std_logic;
signal \nx.n1605\ : std_logic;
signal \nx.n10798\ : std_logic;
signal \nx.n1604\ : std_logic;
signal \nx.n10799\ : std_logic;
signal \nx.n1603\ : std_logic;
signal \nx.n10800\ : std_logic;
signal \nx.n10801\ : std_logic;
signal \nx.n1602\ : std_logic;
signal \bfn_5_26_0_\ : std_logic;
signal \nx.n1601\ : std_logic;
signal \nx.n10802\ : std_logic;
signal \nx.n1600\ : std_logic;
signal \nx.n10803\ : std_logic;
signal \nx.n1599\ : std_logic;
signal \nx.n10804\ : std_logic;
signal \nx.n1598\ : std_logic;
signal \nx.n1631\ : std_logic;
signal \nx.n10805\ : std_logic;
signal \bfn_5_27_0_\ : std_logic;
signal \nx.n1709\ : std_logic;
signal \nx.n10806\ : std_logic;
signal \nx.n1708\ : std_logic;
signal \nx.n10807\ : std_logic;
signal \nx.n1707\ : std_logic;
signal \nx.n10808\ : std_logic;
signal \nx.n10809\ : std_logic;
signal \nx.n10810\ : std_logic;
signal \nx.n1704\ : std_logic;
signal \nx.n10811\ : std_logic;
signal \nx.n10812\ : std_logic;
signal \nx.n10813\ : std_logic;
signal \bfn_5_28_0_\ : std_logic;
signal \nx.n1701\ : std_logic;
signal \nx.n10814\ : std_logic;
signal \nx.n10815\ : std_logic;
signal \nx.n10816\ : std_logic;
signal \nx.n10817\ : std_logic;
signal \nx.n10818\ : std_logic;
signal \nx.n1703\ : std_logic;
signal \nx.n1706\ : std_logic;
signal \nx.n1705\ : std_logic;
signal \nx.n1700\ : std_logic;
signal \nx.n16_adj_766\ : std_logic;
signal \nx.n1702\ : std_logic;
signal \nx.n22_adj_774_cascade_\ : std_logic;
signal \nx.n1698\ : std_logic;
signal \nx.n1699\ : std_logic;
signal \nx.n1697\ : std_logic;
signal \nx.n24_adj_776_cascade_\ : std_logic;
signal \nx.n20_adj_775\ : std_logic;
signal \nx.n1730\ : std_logic;
signal \nx.n1730_cascade_\ : std_logic;
signal \nx.n13601\ : std_logic;
signal n11972 : std_logic;
signal \nx.n13514\ : std_logic;
signal \nx.n13513\ : std_logic;
signal \nx.n7598\ : std_logic;
signal \nx.n11113\ : std_logic;
signal \nx.n7598_cascade_\ : std_logic;
signal timer_26 : std_logic;
signal neo_pixel_transmitter_t0_26 : std_logic;
signal \nx.n7\ : std_logic;
signal \nx.n10_adj_760\ : std_logic;
signal n12_adj_844 : std_logic;
signal \nx.start\ : std_logic;
signal \nx.n11908\ : std_logic;
signal \nx.n7564\ : std_logic;
signal update_color : std_logic;
signal \nx.n13436_cascade_\ : std_logic;
signal \nx.n3901\ : std_logic;
signal state_1_adj_791 : std_logic;
signal \nx.n3901_cascade_\ : std_logic;
signal \nx.n13435\ : std_logic;
signal \nx.n1077\ : std_logic;
signal \bfn_6_20_0_\ : std_logic;
signal \nx.n1076\ : std_logic;
signal \nx.n10743\ : std_logic;
signal \nx.n10744\ : std_logic;
signal \nx.n1074\ : std_logic;
signal \nx.n10745\ : std_logic;
signal \nx.n10746\ : std_logic;
signal \nx.n1072\ : std_logic;
signal \nx.n10747\ : std_logic;
signal \nx.n10748\ : std_logic;
signal \nx.n1103\ : std_logic;
signal \nx.n5\ : std_logic;
signal \nx.n1007\ : std_logic;
signal \nx.n1075\ : std_logic;
signal \nx.n1107\ : std_logic;
signal \nx.n1005\ : std_logic;
signal \nx.n1005_cascade_\ : std_logic;
signal \nx.n1009\ : std_logic;
signal \nx.n7_adj_690_cascade_\ : std_logic;
signal \nx.n1037\ : std_logic;
signal \nx.n1037_cascade_\ : std_logic;
signal \nx.n1073\ : std_logic;
signal \nx.n1105\ : std_logic;
signal \nx.n7899_cascade_\ : std_logic;
signal \nx.n740\ : std_logic;
signal \nx.n740_cascade_\ : std_logic;
signal \nx.n11866_cascade_\ : std_logic;
signal \nx.n838_cascade_\ : std_logic;
signal n18_adj_815 : std_logic;
signal delay_counter_31 : std_logic;
signal n19_adj_814 : std_logic;
signal n17_adj_816 : std_logic;
signal \bfn_6_23_0_\ : std_logic;
signal \nx.n10613\ : std_logic;
signal \nx.n10614\ : std_logic;
signal \nx.n10615\ : std_logic;
signal \nx.n10616\ : std_logic;
signal \nx.n10617\ : std_logic;
signal \nx.n10618\ : std_logic;
signal \nx.n10619\ : std_logic;
signal \nx.n10620\ : std_logic;
signal \bfn_6_24_0_\ : std_logic;
signal \nx.n10621\ : std_logic;
signal \nx.n10622\ : std_logic;
signal \nx.n10623\ : std_logic;
signal \nx.n10624\ : std_logic;
signal \nx.n10625\ : std_logic;
signal \nx.n10626\ : std_logic;
signal \nx.n10627\ : std_logic;
signal \nx.n10628\ : std_logic;
signal \bfn_6_25_0_\ : std_logic;
signal \nx.n10629\ : std_logic;
signal \nx.n10630\ : std_logic;
signal \nx.bit_ctr_19\ : std_logic;
signal \nx.n10631\ : std_logic;
signal \nx.bit_ctr_20\ : std_logic;
signal \nx.n10632\ : std_logic;
signal \nx.bit_ctr_21\ : std_logic;
signal \nx.n10633\ : std_logic;
signal \nx.n10634\ : std_logic;
signal \nx.bit_ctr_23\ : std_logic;
signal \nx.n10635\ : std_logic;
signal \nx.n10636\ : std_logic;
signal \nx.bit_ctr_24\ : std_logic;
signal \bfn_6_26_0_\ : std_logic;
signal \nx.bit_ctr_25\ : std_logic;
signal \nx.n10637\ : std_logic;
signal \nx.n10638\ : std_logic;
signal \nx.n10639\ : std_logic;
signal \nx.n10640\ : std_logic;
signal \nx.n10641\ : std_logic;
signal \nx.n10642\ : std_logic;
signal \nx.n10643\ : std_logic;
signal \nx.n7657\ : std_logic;
signal \nx.n7994\ : std_logic;
signal \bfn_6_27_0_\ : std_logic;
signal \nx.n10819\ : std_logic;
signal \nx.n10820\ : std_logic;
signal \nx.n1807\ : std_logic;
signal \nx.n10821\ : std_logic;
signal \nx.n1806\ : std_logic;
signal \nx.n10822\ : std_logic;
signal \nx.n10823\ : std_logic;
signal \nx.n1804\ : std_logic;
signal \nx.n10824\ : std_logic;
signal \nx.n10825\ : std_logic;
signal \nx.n10826\ : std_logic;
signal \nx.n1802\ : std_logic;
signal \bfn_6_28_0_\ : std_logic;
signal \nx.n1801\ : std_logic;
signal \nx.n10827\ : std_logic;
signal \nx.n10828\ : std_logic;
signal \nx.n10829\ : std_logic;
signal \nx.n10830\ : std_logic;
signal \nx.n1797\ : std_logic;
signal \nx.n10831\ : std_logic;
signal \nx.n10832\ : std_logic;
signal \nx.bit_ctr_18\ : std_logic;
signal \nx.n48_adj_778\ : std_logic;
signal \nx.n18_adj_716\ : std_logic;
signal \nx.n1799\ : std_logic;
signal \nx.n1805\ : std_logic;
signal \nx.n24_adj_717\ : std_logic;
signal \nx.n1798\ : std_logic;
signal \nx.n1808\ : std_logic;
signal \nx.n26_adj_719_cascade_\ : std_logic;
signal \nx.n1809\ : std_logic;
signal \nx.n1803\ : std_logic;
signal \nx.n1800\ : std_logic;
signal \nx.n9717_cascade_\ : std_logic;
signal \nx.n1796\ : std_logic;
signal \nx.n22_adj_718\ : std_logic;
signal \nx.n1829\ : std_logic;
signal \nx.n13605\ : std_logic;
signal pin_oe_7 : std_logic;
signal \nx.neo_pixel_transmitter_done\ : std_logic;
signal \NEOPXL_c\ : std_logic;
signal \nx.n11988\ : std_logic;
signal \nx.n12451\ : std_logic;
signal \nx.bit_ctr_1\ : std_logic;
signal \nx.n13364\ : std_logic;
signal \nx.n11156_cascade_\ : std_logic;
signal \nx.n13363\ : std_logic;
signal \nx.n13619_cascade_\ : std_logic;
signal \nx.n11156\ : std_logic;
signal n11966 : std_logic;
signal pin_oe_2 : std_logic;
signal \nx.n13372\ : std_logic;
signal timer_28 : std_logic;
signal n11353 : std_logic;
signal neo_pixel_transmitter_t0_28 : std_logic;
signal n9_adj_847 : std_logic;
signal \current_pin_7__N_153\ : std_logic;
signal neopxl_color_prev_14 : std_logic;
signal neopxl_color_13 : std_logic;
signal neopxl_color_prev_13 : std_logic;
signal n11_adj_845 : std_logic;
signal neopxl_color_prev_4 : std_logic;
signal neopxl_color_14 : std_logic;
signal \nx.n11941\ : std_logic;
signal \nx.n1008\ : std_logic;
signal \nx.n1006\ : std_logic;
signal \nx.n12837_cascade_\ : std_logic;
signal \nx.n905_cascade_\ : std_logic;
signal \nx.n12839\ : std_logic;
signal \nx.n11174\ : std_logic;
signal \nx.n11174_cascade_\ : std_logic;
signal \nx.bit_ctr_26\ : std_logic;
signal \nx.n977\ : std_logic;
signal \bfn_7_22_0_\ : std_logic;
signal \nx.n7497\ : std_logic;
signal \nx.n976\ : std_logic;
signal \nx.n10738\ : std_logic;
signal \nx.n7899\ : std_logic;
signal \nx.n975\ : std_logic;
signal \nx.n10739\ : std_logic;
signal \nx.n974\ : std_logic;
signal \nx.n10740\ : std_logic;
signal \nx.n906\ : std_logic;
signal \nx.n973\ : std_logic;
signal \nx.n10741\ : std_logic;
signal \nx.n13594\ : std_logic;
signal \nx.n905\ : std_logic;
signal \nx.n10742\ : std_logic;
signal \nx.n4\ : std_logic;
signal \nx.n807\ : std_logic;
signal \nx.n11866\ : std_logic;
signal \nx.n838\ : std_logic;
signal \nx.n11868\ : std_logic;
signal \nx.bit_ctr_17\ : std_logic;
signal \nx.bit_ctr_22\ : std_logic;
signal \nx.n44_adj_782\ : std_logic;
signal \nx.n11912_cascade_\ : std_logic;
signal \nx.n58\ : std_logic;
signal \nx.bit_ctr_29\ : std_logic;
signal \nx.bit_ctr_30\ : std_logic;
signal \nx.bit_ctr_31\ : std_logic;
signal \nx.n9803\ : std_logic;
signal \nx.bit_ctr_27\ : std_logic;
signal \nx.bit_ctr_28\ : std_logic;
signal \nx.n11912\ : std_logic;
signal \nx.n708\ : std_logic;
signal \nx.n5703\ : std_logic;
signal n10_adj_846 : std_logic;
signal neopxl_color_prev_7 : std_logic;
signal neopxl_color_15 : std_logic;
signal neopxl_color_prev_15 : std_logic;
signal neopxl_color_6 : std_logic;
signal \nx.bit_ctr_0\ : std_logic;
signal \nx.n13373\ : std_logic;
signal neopxl_color_7 : std_logic;
signal n22_adj_793 : std_logic;
signal \nx.n26_cascade_\ : std_logic;
signal \nx.n20\ : std_logic;
signal \nx.n28_adj_679_cascade_\ : std_logic;
signal \nx.n16_adj_678\ : std_logic;
signal \nx.n1928_cascade_\ : std_logic;
signal \nx.bit_ctr_16\ : std_logic;
signal \nx.n1977\ : std_logic;
signal \bfn_7_27_0_\ : std_logic;
signal \nx.n1909\ : std_logic;
signal \nx.n1976\ : std_logic;
signal \nx.n10833\ : std_logic;
signal \nx.n1908\ : std_logic;
signal \nx.n1975\ : std_logic;
signal \nx.n10834\ : std_logic;
signal \nx.n1907\ : std_logic;
signal \nx.n1974\ : std_logic;
signal \nx.n10835\ : std_logic;
signal \nx.n1906\ : std_logic;
signal \nx.n1973\ : std_logic;
signal \nx.n10836\ : std_logic;
signal \nx.n10837\ : std_logic;
signal \nx.n10838\ : std_logic;
signal \nx.n10839\ : std_logic;
signal \nx.n10840\ : std_logic;
signal \bfn_7_28_0_\ : std_logic;
signal \nx.n10841\ : std_logic;
signal \nx.n10842\ : std_logic;
signal \nx.n10843\ : std_logic;
signal \nx.n10844\ : std_logic;
signal \nx.n10845\ : std_logic;
signal \nx.n10846\ : std_logic;
signal \nx.n1895\ : std_logic;
signal \nx.n10847\ : std_logic;
signal \nx.n24\ : std_logic;
signal \nx.n1963\ : std_logic;
signal \nx.n1896\ : std_logic;
signal \nx.n1995_cascade_\ : std_logic;
signal \nx.n1965\ : std_logic;
signal \nx.n1898\ : std_logic;
signal \nx.n1964\ : std_logic;
signal \nx.n1897\ : std_logic;
signal \nx.n1971\ : std_logic;
signal \nx.n1904\ : std_logic;
signal n13360 : std_logic;
signal \n13361_cascade_\ : std_logic;
signal \LED_c\ : std_logic;
signal neopxl_color_12 : std_logic;
signal \nx.n59\ : std_logic;
signal \nx.n61_cascade_\ : std_logic;
signal \nx.n11153\ : std_logic;
signal \nx.bit_ctr_2\ : std_logic;
signal \state_3_N_448_1\ : std_logic;
signal \nx.color_bit_N_642_4\ : std_logic;
signal \nx.n13622\ : std_logic;
signal state_0_adj_792 : std_logic;
signal n7671 : std_logic;
signal \nx.n7983\ : std_logic;
signal \nx.n12817\ : std_logic;
signal \nx.n12819_cascade_\ : std_logic;
signal \nx.n12821\ : std_logic;
signal \nx.n3009_cascade_\ : std_logic;
signal \nx.n2791_cascade_\ : std_logic;
signal \bfn_9_21_0_\ : std_logic;
signal \nx.n2876\ : std_logic;
signal \nx.n11004\ : std_logic;
signal \nx.n2875\ : std_logic;
signal \nx.n11005\ : std_logic;
signal \nx.n11006\ : std_logic;
signal \nx.n11007\ : std_logic;
signal \nx.n11008\ : std_logic;
signal \nx.n11009\ : std_logic;
signal \nx.n11010\ : std_logic;
signal \nx.n11011\ : std_logic;
signal \bfn_9_22_0_\ : std_logic;
signal \nx.n11012\ : std_logic;
signal \nx.n11013\ : std_logic;
signal \nx.n11014\ : std_logic;
signal \nx.n11015\ : std_logic;
signal \nx.n11016\ : std_logic;
signal \nx.n11017\ : std_logic;
signal \nx.n11018\ : std_logic;
signal \nx.n11019\ : std_logic;
signal \bfn_9_23_0_\ : std_logic;
signal \nx.n11020\ : std_logic;
signal \nx.n2859\ : std_logic;
signal \nx.n11021\ : std_logic;
signal \nx.n2791\ : std_logic;
signal \nx.n2858\ : std_logic;
signal \nx.n11022\ : std_logic;
signal \nx.n11023\ : std_logic;
signal \nx.n2856\ : std_logic;
signal \nx.n11024\ : std_logic;
signal \nx.n11025\ : std_logic;
signal \nx.n11026\ : std_logic;
signal \nx.n11027\ : std_logic;
signal \bfn_9_24_0_\ : std_logic;
signal \nx.n2792\ : std_logic;
signal neopxl_color_prev_5 : std_logic;
signal neopxl_color_5 : std_logic;
signal n22 : std_logic;
signal \nx.n1966\ : std_logic;
signal \nx.n1899\ : std_logic;
signal \nx.n1967\ : std_logic;
signal \nx.n1900\ : std_logic;
signal \nx.n1970\ : std_logic;
signal \nx.n1903\ : std_logic;
signal \nx.n1972\ : std_logic;
signal \nx.n1905\ : std_logic;
signal \bfn_9_26_0_\ : std_logic;
signal \nx.n10848\ : std_logic;
signal \nx.n10849\ : std_logic;
signal \nx.n10850\ : std_logic;
signal \nx.n10851\ : std_logic;
signal \nx.n10852\ : std_logic;
signal \nx.n10853\ : std_logic;
signal \nx.n10854\ : std_logic;
signal \nx.n10855\ : std_logic;
signal \bfn_9_27_0_\ : std_logic;
signal \nx.n10856\ : std_logic;
signal \nx.n10857\ : std_logic;
signal \nx.n10858\ : std_logic;
signal \nx.n10859\ : std_logic;
signal \nx.n10860\ : std_logic;
signal \nx.n10861\ : std_logic;
signal \nx.n10862\ : std_logic;
signal \nx.n10863\ : std_logic;
signal \nx.n1994\ : std_logic;
signal \bfn_9_28_0_\ : std_logic;
signal \nx.n1995\ : std_logic;
signal \nx.n2062\ : std_logic;
signal \nx.n2094_cascade_\ : std_logic;
signal \nx.n1901\ : std_logic;
signal \nx.n1968\ : std_logic;
signal \nx.n1969\ : std_logic;
signal \nx.n1902\ : std_logic;
signal \nx.n1928\ : std_logic;
signal \nx.n2068\ : std_logic;
signal \nx.n2001_cascade_\ : std_logic;
signal \nx.n2067\ : std_logic;
signal \nx.n2099_cascade_\ : std_logic;
signal n26_adj_798 : std_logic;
signal \bfn_9_29_0_\ : std_logic;
signal n25 : std_logic;
signal n10644 : std_logic;
signal n24 : std_logic;
signal n10645 : std_logic;
signal n23 : std_logic;
signal n10646 : std_logic;
signal n22_adj_799 : std_logic;
signal n10647 : std_logic;
signal n21 : std_logic;
signal n10648 : std_logic;
signal n20 : std_logic;
signal n10649 : std_logic;
signal n19_adj_800 : std_logic;
signal n10650 : std_logic;
signal n10651 : std_logic;
signal n18 : std_logic;
signal \bfn_9_30_0_\ : std_logic;
signal n17 : std_logic;
signal n10652 : std_logic;
signal n16 : std_logic;
signal n10653 : std_logic;
signal n15 : std_logic;
signal n10654 : std_logic;
signal n14_adj_802 : std_logic;
signal n10655 : std_logic;
signal n13 : std_logic;
signal n10656 : std_logic;
signal n12 : std_logic;
signal n10657 : std_logic;
signal n11 : std_logic;
signal n10658 : std_logic;
signal n10659 : std_logic;
signal n10_adj_806 : std_logic;
signal \bfn_9_31_0_\ : std_logic;
signal n9_adj_807 : std_logic;
signal n10660 : std_logic;
signal n8 : std_logic;
signal n10661 : std_logic;
signal n7_adj_808 : std_logic;
signal n10662 : std_logic;
signal n6_adj_809 : std_logic;
signal n10663 : std_logic;
signal blink_counter_21 : std_logic;
signal n10664 : std_logic;
signal blink_counter_22 : std_logic;
signal n10665 : std_logic;
signal blink_counter_23 : std_logic;
signal n10666 : std_logic;
signal n10667 : std_logic;
signal blink_counter_24 : std_logic;
signal \bfn_9_32_0_\ : std_logic;
signal n10668 : std_logic;
signal blink_counter_25 : std_logic;
signal \nx.n45_adj_754_cascade_\ : std_logic;
signal \nx.n12809_cascade_\ : std_logic;
signal \nx.n12811_cascade_\ : std_logic;
signal \nx.n12813_cascade_\ : std_logic;
signal \nx.n12815\ : std_logic;
signal \nx.n43_adj_753\ : std_logic;
signal \nx.n46_cascade_\ : std_logic;
signal \nx.n13_adj_743_cascade_\ : std_logic;
signal \nx.n12775\ : std_logic;
signal \nx.n12787_cascade_\ : std_logic;
signal \nx.n12803\ : std_logic;
signal \nx.n35_adj_738\ : std_logic;
signal \nx.n2987_cascade_\ : std_logic;
signal \nx.n41_cascade_\ : std_logic;
signal \nx.n39_adj_671\ : std_logic;
signal \nx.n50_cascade_\ : std_logic;
signal \nx.n2877\ : std_logic;
signal \nx.n2857\ : std_logic;
signal \nx.n2790\ : std_logic;
signal \nx.n2889_cascade_\ : std_logic;
signal \nx.n2868\ : std_logic;
signal \nx.n2801\ : std_logic;
signal \nx.n2808\ : std_logic;
signal \nx.n40_adj_705_cascade_\ : std_logic;
signal \nx.n44_adj_721_cascade_\ : std_logic;
signal \nx.n2862\ : std_logic;
signal \nx.n2819_cascade_\ : std_logic;
signal \nx.n2874\ : std_logic;
signal \nx.n42_adj_730\ : std_logic;
signal \nx.n2807\ : std_logic;
signal \nx.n2809\ : std_logic;
signal \nx.n2809_cascade_\ : std_logic;
signal \nx.bit_ctr_7\ : std_logic;
signal \nx.n30_adj_704\ : std_logic;
signal \nx.n2802\ : std_logic;
signal \nx.n2869\ : std_logic;
signal \nx.n2802_cascade_\ : std_logic;
signal \nx.n2795\ : std_logic;
signal \nx.n2720_cascade_\ : std_logic;
signal \nx.n2788_cascade_\ : std_logic;
signal \nx.n2789\ : std_logic;
signal \nx.n26_adj_706_cascade_\ : std_logic;
signal \nx.n38_adj_713\ : std_logic;
signal \nx.n43_adj_735\ : std_logic;
signal \nx.n2777\ : std_logic;
signal \bfn_10_23_0_\ : std_logic;
signal \nx.n2776\ : std_logic;
signal \nx.n10981\ : std_logic;
signal \nx.n2775\ : std_logic;
signal \nx.n10982\ : std_logic;
signal \nx.n10983\ : std_logic;
signal \nx.n2773\ : std_logic;
signal \nx.n10984\ : std_logic;
signal \nx.n2772\ : std_logic;
signal \nx.n10985\ : std_logic;
signal \nx.n2771\ : std_logic;
signal \nx.n10986\ : std_logic;
signal \nx.n2770\ : std_logic;
signal \nx.n10987\ : std_logic;
signal \nx.n10988\ : std_logic;
signal \nx.n2769\ : std_logic;
signal \bfn_10_24_0_\ : std_logic;
signal \nx.n2768\ : std_logic;
signal \nx.n10989\ : std_logic;
signal \nx.n10990\ : std_logic;
signal \nx.n10991\ : std_logic;
signal \nx.n10992\ : std_logic;
signal \nx.n10993\ : std_logic;
signal \nx.n2763\ : std_logic;
signal \nx.n10994\ : std_logic;
signal \nx.n2762\ : std_logic;
signal \nx.n10995\ : std_logic;
signal \nx.n10996\ : std_logic;
signal \nx.n2761\ : std_logic;
signal \bfn_10_25_0_\ : std_logic;
signal \nx.n2760\ : std_logic;
signal \nx.n10997\ : std_logic;
signal \nx.n2759\ : std_logic;
signal \nx.n10998\ : std_logic;
signal \nx.n2758\ : std_logic;
signal \nx.n10999\ : std_logic;
signal \nx.n2757\ : std_logic;
signal \nx.n11000\ : std_logic;
signal \nx.n2756\ : std_logic;
signal \nx.n11001\ : std_logic;
signal \nx.n11002\ : std_logic;
signal \nx.n11003\ : std_logic;
signal \nx.n2786\ : std_logic;
signal \nx.n2070\ : std_logic;
signal \nx.n9709_cascade_\ : std_logic;
signal \nx.n25\ : std_logic;
signal \nx.n26_adj_681_cascade_\ : std_logic;
signal \nx.n2027_cascade_\ : std_logic;
signal \nx.n2074\ : std_logic;
signal \nx.n2001\ : std_logic;
signal \nx.n28_adj_680\ : std_logic;
signal \nx.n1999\ : std_logic;
signal \nx.n2066\ : std_logic;
signal \nx.n2007\ : std_logic;
signal \nx.n2003\ : std_logic;
signal \nx.n2000\ : std_logic;
signal \nx.n27\ : std_logic;
signal \nx.n2004\ : std_logic;
signal \nx.n2071\ : std_logic;
signal \nx.n2103_cascade_\ : std_logic;
signal \nx.n1998\ : std_logic;
signal \nx.n2065\ : std_logic;
signal \nx.n2073\ : std_logic;
signal \nx.n2006\ : std_logic;
signal \nx.n2105_cascade_\ : std_logic;
signal \nx.n2005\ : std_logic;
signal \nx.n2072\ : std_logic;
signal \nx.n2002\ : std_logic;
signal \nx.n2069\ : std_logic;
signal \nx.n2075\ : std_logic;
signal \nx.n2008\ : std_logic;
signal \nx.n2107_cascade_\ : std_logic;
signal \nx.n24_adj_684\ : std_logic;
signal \nx.n1997\ : std_logic;
signal \nx.n2064\ : std_logic;
signal \nx.n2096_cascade_\ : std_logic;
signal \nx.bit_ctr_15\ : std_logic;
signal \nx.n2077\ : std_logic;
signal \nx.n2109_cascade_\ : std_logic;
signal \nx.n2202_cascade_\ : std_logic;
signal \nx.n18_adj_682\ : std_logic;
signal \nx.n2193_cascade_\ : std_logic;
signal \nx.n2009\ : std_logic;
signal \nx.n2076\ : std_logic;
signal \nx.n2108_cascade_\ : std_logic;
signal \nx.n1996\ : std_logic;
signal \nx.n2027\ : std_logic;
signal \nx.n2063\ : std_logic;
signal \nx.n42_adj_739_cascade_\ : std_logic;
signal \nx.n32_adj_740_cascade_\ : std_logic;
signal \nx.n44_adj_741\ : std_logic;
signal \nx.n50_adj_742\ : std_logic;
signal \nx.n47\ : std_logic;
signal \nx.n49_cascade_\ : std_logic;
signal \nx.n48\ : std_logic;
signal \nx.n3116_cascade_\ : std_logic;
signal \nx.bit_ctr_5\ : std_logic;
signal \bfn_11_18_0_\ : std_logic;
signal \nx.n3009\ : std_logic;
signal \nx.n13600\ : std_logic;
signal \nx.n11053\ : std_logic;
signal \nx.n3008\ : std_logic;
signal \nx.n11054\ : std_logic;
signal \nx.n3007\ : std_logic;
signal \nx.n11055\ : std_logic;
signal \nx.n11056\ : std_logic;
signal \nx.n11057\ : std_logic;
signal \nx.n11058\ : std_logic;
signal \nx.n11059\ : std_logic;
signal \nx.n11060\ : std_logic;
signal \bfn_11_19_0_\ : std_logic;
signal \nx.n11061\ : std_logic;
signal \nx.n11062\ : std_logic;
signal \nx.n11063\ : std_logic;
signal \nx.n11064\ : std_logic;
signal \nx.n11065\ : std_logic;
signal \nx.n11066\ : std_logic;
signal \nx.n11067\ : std_logic;
signal \nx.n11068\ : std_logic;
signal \bfn_11_20_0_\ : std_logic;
signal \nx.n11069\ : std_logic;
signal \nx.n11070\ : std_logic;
signal \nx.n11071\ : std_logic;
signal \nx.n11072\ : std_logic;
signal \nx.n11073\ : std_logic;
signal \nx.n11074\ : std_logic;
signal \nx.n2987\ : std_logic;
signal \nx.n11075\ : std_logic;
signal \nx.n11076\ : std_logic;
signal \bfn_11_21_0_\ : std_logic;
signal \nx.n11077\ : std_logic;
signal \nx.n3017\ : std_logic;
signal \nx.n11078\ : std_logic;
signal \nx.n40_adj_670\ : std_logic;
signal \nx.n2996\ : std_logic;
signal \nx.n41_adj_736\ : std_logic;
signal \nx.n2998\ : std_logic;
signal \nx.n2765\ : std_logic;
signal \nx.n41_adj_688\ : std_logic;
signal \nx.n2767\ : std_logic;
signal \nx.n2854\ : std_logic;
signal \nx.n2886_cascade_\ : std_logic;
signal \nx.n2985\ : std_logic;
signal \nx.n2774\ : std_logic;
signal \nx.n2800\ : std_logic;
signal \nx.n2867\ : std_logic;
signal \nx.n2706\ : std_logic;
signal \nx.n2706_cascade_\ : std_logic;
signal \nx.n40_adj_687\ : std_logic;
signal \nx.n2755\ : std_logic;
signal \nx.n2787\ : std_logic;
signal \nx.n2699\ : std_logic;
signal \nx.n2766\ : std_logic;
signal \nx.n2699_cascade_\ : std_logic;
signal \nx.n2701\ : std_logic;
signal \nx.n2701_cascade_\ : std_logic;
signal \nx.n42_adj_683\ : std_logic;
signal \nx.n2698\ : std_logic;
signal \nx.bit_ctr_8\ : std_logic;
signal \nx.n2698_cascade_\ : std_logic;
signal \nx.n30\ : std_logic;
signal \nx.n2693\ : std_logic;
signal \nx.n2694\ : std_logic;
signal \nx.n2693_cascade_\ : std_logic;
signal \nx.n2696\ : std_logic;
signal \nx.n37_adj_677\ : std_logic;
signal \nx.n2709\ : std_logic;
signal \bfn_11_25_0_\ : std_logic;
signal \nx.n10881\ : std_logic;
signal \nx.n10882\ : std_logic;
signal \nx.n10883\ : std_logic;
signal \nx.n10884\ : std_logic;
signal \nx.n10885\ : std_logic;
signal \nx.n10886\ : std_logic;
signal \nx.n10887\ : std_logic;
signal \nx.n10888\ : std_logic;
signal \bfn_11_26_0_\ : std_logic;
signal \nx.n10889\ : std_logic;
signal \nx.n10890\ : std_logic;
signal \nx.n10891\ : std_logic;
signal \nx.n10892\ : std_logic;
signal \nx.n2264\ : std_logic;
signal \nx.n10893\ : std_logic;
signal \nx.n10894\ : std_logic;
signal \nx.n10895\ : std_logic;
signal \nx.n10896\ : std_logic;
signal \bfn_11_27_0_\ : std_logic;
signal \nx.n10897\ : std_logic;
signal \nx.n10898\ : std_logic;
signal \nx.n2263\ : std_logic;
signal \nx.n2196_cascade_\ : std_logic;
signal \nx.n2193\ : std_logic;
signal \nx.n2260\ : std_logic;
signal \nx.n29\ : std_logic;
signal \nx.n28_adj_686\ : std_logic;
signal \nx.n27_adj_691\ : std_logic;
signal \nx.n30_adj_685\ : std_logic;
signal \nx.n2126_cascade_\ : std_logic;
signal \nx.n2199_cascade_\ : std_logic;
signal \nx.n31_cascade_\ : std_logic;
signal \nx.n28_adj_692\ : std_logic;
signal \nx.bit_ctr_14\ : std_logic;
signal \nx.n2177\ : std_logic;
signal \bfn_11_29_0_\ : std_logic;
signal \nx.n2109\ : std_logic;
signal \nx.n2176\ : std_logic;
signal \nx.n10864\ : std_logic;
signal \nx.n2108\ : std_logic;
signal \nx.n2175\ : std_logic;
signal \nx.n10865\ : std_logic;
signal \nx.n2107\ : std_logic;
signal \nx.n2174\ : std_logic;
signal \nx.n10866\ : std_logic;
signal \nx.n2106\ : std_logic;
signal \nx.n2173\ : std_logic;
signal \nx.n10867\ : std_logic;
signal \nx.n2105\ : std_logic;
signal \nx.n2172\ : std_logic;
signal \nx.n10868\ : std_logic;
signal \nx.n2104\ : std_logic;
signal \nx.n2171\ : std_logic;
signal \nx.n10869\ : std_logic;
signal \nx.n2103\ : std_logic;
signal \nx.n2170\ : std_logic;
signal \nx.n10870\ : std_logic;
signal \nx.n10871\ : std_logic;
signal \bfn_11_30_0_\ : std_logic;
signal \nx.n10872\ : std_logic;
signal \nx.n2100\ : std_logic;
signal \nx.n2167\ : std_logic;
signal \nx.n10873\ : std_logic;
signal \nx.n10874\ : std_logic;
signal \nx.n2098\ : std_logic;
signal \nx.n2165\ : std_logic;
signal \nx.n10875\ : std_logic;
signal \nx.n2097\ : std_logic;
signal \nx.n2164\ : std_logic;
signal \nx.n10876\ : std_logic;
signal \nx.n2096\ : std_logic;
signal \nx.n2163\ : std_logic;
signal \nx.n10877\ : std_logic;
signal \nx.n2095\ : std_logic;
signal \nx.n2162\ : std_logic;
signal \nx.n10878\ : std_logic;
signal \nx.n10879\ : std_logic;
signal \nx.n2094\ : std_logic;
signal \nx.n2161\ : std_logic;
signal \bfn_11_31_0_\ : std_logic;
signal \nx.n2093\ : std_logic;
signal \nx.n10880\ : std_logic;
signal \nx.n2192\ : std_logic;
signal \nx.n21_adj_750_cascade_\ : std_logic;
signal \nx.bit_ctr_3\ : std_logic;
signal \nx.n12781_cascade_\ : std_logic;
signal \nx.n12801\ : std_logic;
signal \nx.n27_adj_744_cascade_\ : std_logic;
signal \nx.n3209\ : std_logic;
signal \nx.n25_adj_748_cascade_\ : std_logic;
signal \nx.n12785\ : std_logic;
signal \nx.n19_adj_745\ : std_logic;
signal \nx.n12777_cascade_\ : std_logic;
signal \nx.n12779\ : std_logic;
signal \nx.n39_adj_747_cascade_\ : std_logic;
signal \nx.n12789\ : std_logic;
signal \nx.n12799\ : std_logic;
signal \nx.n29_adj_746\ : std_logic;
signal \nx.n11_adj_751\ : std_logic;
signal \nx.n41_adj_752\ : std_logic;
signal \nx.n2989\ : std_logic;
signal \nx.n3000\ : std_logic;
signal \nx.n3001\ : std_logic;
signal \nx.n3001_cascade_\ : std_logic;
signal \nx.n44\ : std_logic;
signal \nx.n3003\ : std_logic;
signal \nx.n3005\ : std_logic;
signal \nx.n2863\ : std_logic;
signal \nx.n2895_cascade_\ : std_logic;
signal \nx.n2994\ : std_logic;
signal \nx.n2799\ : std_logic;
signal \nx.n2866\ : std_logic;
signal \nx.n2898_cascade_\ : std_logic;
signal \nx.n2997\ : std_logic;
signal \nx.n2997_cascade_\ : std_logic;
signal \nx.n45\ : std_logic;
signal \nx.n2988\ : std_logic;
signal \nx.n2855\ : std_logic;
signal \nx.n2788\ : std_logic;
signal \nx.n2764\ : std_logic;
signal \nx.n2697\ : std_logic;
signal \nx.n2720\ : std_logic;
signal \nx.n2796\ : std_logic;
signal \nx.n2597_cascade_\ : std_logic;
signal \nx.n2691\ : std_logic;
signal \nx.n2690\ : std_logic;
signal \nx.n2691_cascade_\ : std_logic;
signal \nx.n2692\ : std_logic;
signal \nx.n36\ : std_logic;
signal \nx.n2700\ : std_logic;
signal \nx.n2688\ : std_logic;
signal \nx.n2689\ : std_logic;
signal \nx.n34_cascade_\ : std_logic;
signal \nx.n38\ : std_logic;
signal \nx.n37\ : std_logic;
signal \nx.n39_cascade_\ : std_logic;
signal \nx.n2621_cascade_\ : std_logic;
signal \nx.n2707\ : std_logic;
signal \nx.bit_ctr_13\ : std_logic;
signal \nx.n2277\ : std_logic;
signal \nx.n2309_cascade_\ : std_logic;
signal \nx.n9697_cascade_\ : std_logic;
signal \nx.n2273\ : std_logic;
signal \nx.n2206\ : std_logic;
signal \nx.n2209\ : std_logic;
signal \nx.n2276\ : std_logic;
signal \nx.n2695\ : std_logic;
signal \nx.n2204\ : std_logic;
signal \nx.n2271\ : std_logic;
signal \nx.n2303_cascade_\ : std_logic;
signal \nx.n2269\ : std_logic;
signal \nx.n2202\ : std_logic;
signal \nx.n2203\ : std_logic;
signal \nx.n2270\ : std_logic;
signal \nx.n2302_cascade_\ : std_logic;
signal \nx.n2401_cascade_\ : std_logic;
signal \nx.n2274\ : std_logic;
signal \nx.n2207\ : std_logic;
signal \nx.n2208\ : std_logic;
signal \nx.n2275\ : std_logic;
signal \nx.n2272\ : std_logic;
signal \nx.n2205\ : std_logic;
signal \nx.n2391_cascade_\ : std_logic;
signal \nx.n30_adj_696_cascade_\ : std_logic;
signal \nx.n2266\ : std_logic;
signal \nx.n2199\ : std_logic;
signal \nx.n2267\ : std_logic;
signal \nx.n2299_cascade_\ : std_logic;
signal \nx.n2265\ : std_logic;
signal \nx.n2197\ : std_logic;
signal \nx.n2196\ : std_logic;
signal \nx.n30_adj_694\ : std_logic;
signal \nx.n22_adj_693\ : std_logic;
signal \nx.n21_cascade_\ : std_logic;
signal \nx.n34_adj_695\ : std_logic;
signal \nx.n2268\ : std_logic;
signal \nx.n2225_cascade_\ : std_logic;
signal neopxl_color_4 : std_logic;
signal n22_adj_787 : std_logic;
signal \nx.n2099\ : std_logic;
signal \nx.n2166\ : std_logic;
signal \nx.n2198\ : std_logic;
signal \nx.n2169\ : std_logic;
signal \nx.n2102\ : std_logic;
signal \nx.n2201\ : std_logic;
signal \nx.n2261\ : std_logic;
signal \nx.n2194\ : std_logic;
signal \nx.n2262\ : std_logic;
signal \nx.n2195\ : std_logic;
signal \nx.n2225\ : std_logic;
signal pin_oe_4 : std_logic;
signal \n11970_cascade_\ : std_logic;
signal pin_oe_0 : std_logic;
signal n11968 : std_logic;
signal \nx.bit_ctr_4\ : std_logic;
signal \nx.n3177\ : std_logic;
signal \bfn_13_17_0_\ : std_logic;
signal \nx.n3109\ : std_logic;
signal \nx.n3176\ : std_logic;
signal \nx.n11079\ : std_logic;
signal \nx.n3108\ : std_logic;
signal \nx.n3175\ : std_logic;
signal \nx.n11080\ : std_logic;
signal \nx.n3107\ : std_logic;
signal \nx.n3174\ : std_logic;
signal \nx.n11081\ : std_logic;
signal \nx.n3106\ : std_logic;
signal \nx.n3173\ : std_logic;
signal \nx.n11082\ : std_logic;
signal \nx.n3105\ : std_logic;
signal \nx.n3172\ : std_logic;
signal \nx.n11083\ : std_logic;
signal \nx.n3104\ : std_logic;
signal \nx.n3171\ : std_logic;
signal \nx.n11084\ : std_logic;
signal \nx.n3103\ : std_logic;
signal \nx.n3170\ : std_logic;
signal \nx.n11085\ : std_logic;
signal \nx.n11086\ : std_logic;
signal \nx.n3102\ : std_logic;
signal \nx.n3169\ : std_logic;
signal \bfn_13_18_0_\ : std_logic;
signal \nx.n3101\ : std_logic;
signal \nx.n3168\ : std_logic;
signal \nx.n11087\ : std_logic;
signal \nx.n3100\ : std_logic;
signal \nx.n3167\ : std_logic;
signal \nx.n11088\ : std_logic;
signal \nx.n3099\ : std_logic;
signal \nx.n3166\ : std_logic;
signal \nx.n11089\ : std_logic;
signal \nx.n3098\ : std_logic;
signal \nx.n3165\ : std_logic;
signal \nx.n11090\ : std_logic;
signal \nx.n3097\ : std_logic;
signal \nx.n3164\ : std_logic;
signal \nx.n11091\ : std_logic;
signal \nx.n3096\ : std_logic;
signal \nx.n3163\ : std_logic;
signal \nx.n11092\ : std_logic;
signal \nx.n3095\ : std_logic;
signal \nx.n3162\ : std_logic;
signal \nx.n11093\ : std_logic;
signal \nx.n11094\ : std_logic;
signal \nx.n3094\ : std_logic;
signal \nx.n3161\ : std_logic;
signal \bfn_13_19_0_\ : std_logic;
signal \nx.n3093\ : std_logic;
signal \nx.n3160\ : std_logic;
signal \nx.n11095\ : std_logic;
signal \nx.n3092\ : std_logic;
signal \nx.n3159\ : std_logic;
signal \nx.n11096\ : std_logic;
signal \nx.n3091\ : std_logic;
signal \nx.n3158\ : std_logic;
signal \nx.n11097\ : std_logic;
signal \nx.n3090\ : std_logic;
signal \nx.n3157\ : std_logic;
signal \nx.n11098\ : std_logic;
signal \nx.n3089\ : std_logic;
signal \nx.n3156\ : std_logic;
signal \nx.n11099\ : std_logic;
signal \nx.n3088\ : std_logic;
signal \nx.n3155\ : std_logic;
signal \nx.n11100\ : std_logic;
signal \nx.n3087\ : std_logic;
signal \nx.n3154\ : std_logic;
signal \nx.n11101\ : std_logic;
signal \nx.n11102\ : std_logic;
signal \nx.n3086\ : std_logic;
signal \nx.n3153\ : std_logic;
signal \bfn_13_20_0_\ : std_logic;
signal \nx.n3085\ : std_logic;
signal \nx.n3152\ : std_logic;
signal \nx.n11103\ : std_logic;
signal \nx.n3084\ : std_logic;
signal \nx.n3151\ : std_logic;
signal \nx.n11104\ : std_logic;
signal \nx.n3116\ : std_logic;
signal \nx.n3083\ : std_logic;
signal \nx.n11105\ : std_logic;
signal \nx.n13280\ : std_logic;
signal \nx.n2805\ : std_logic;
signal \nx.n2872\ : std_logic;
signal \nx.n2798\ : std_logic;
signal \nx.n2865\ : std_logic;
signal \nx.n2986\ : std_logic;
signal \nx.n2991\ : std_logic;
signal \nx.n2603_cascade_\ : std_logic;
signal \nx.n2702\ : std_logic;
signal \nx.n2803\ : std_logic;
signal \nx.n2870\ : std_logic;
signal \nx.n2501_cascade_\ : std_logic;
signal \nx.n2507_cascade_\ : std_logic;
signal \nx.n2398_cascade_\ : std_logic;
signal \nx.n31_adj_700\ : std_logic;
signal \nx.n32_adj_698\ : std_logic;
signal \nx.n33_adj_699\ : std_logic;
signal \nx.n34_adj_697\ : std_logic;
signal \nx.n2324_cascade_\ : std_logic;
signal \nx.bit_ctr_12\ : std_logic;
signal \nx.n2377\ : std_logic;
signal \bfn_13_26_0_\ : std_logic;
signal \nx.n2309\ : std_logic;
signal \nx.n2376\ : std_logic;
signal \nx.n10899\ : std_logic;
signal \nx.n2308\ : std_logic;
signal \nx.n2375\ : std_logic;
signal \nx.n10900\ : std_logic;
signal \nx.n10901\ : std_logic;
signal \nx.n2306\ : std_logic;
signal \nx.n2373\ : std_logic;
signal \nx.n10902\ : std_logic;
signal \nx.n2305\ : std_logic;
signal \nx.n2372\ : std_logic;
signal \nx.n10903\ : std_logic;
signal \nx.n2304\ : std_logic;
signal \nx.n2371\ : std_logic;
signal \nx.n10904\ : std_logic;
signal \nx.n2303\ : std_logic;
signal \nx.n2370\ : std_logic;
signal \nx.n10905\ : std_logic;
signal \nx.n10906\ : std_logic;
signal \nx.n2302\ : std_logic;
signal \nx.n2369\ : std_logic;
signal \bfn_13_27_0_\ : std_logic;
signal \nx.n10907\ : std_logic;
signal \nx.n2300\ : std_logic;
signal \nx.n2367\ : std_logic;
signal \nx.n10908\ : std_logic;
signal \nx.n2299\ : std_logic;
signal \nx.n2366\ : std_logic;
signal \nx.n10909\ : std_logic;
signal \nx.n10910\ : std_logic;
signal \nx.n10911\ : std_logic;
signal \nx.n2296\ : std_logic;
signal \nx.n2363\ : std_logic;
signal \nx.n10912\ : std_logic;
signal \nx.n10913\ : std_logic;
signal \nx.n10914\ : std_logic;
signal \nx.n2294\ : std_logic;
signal \nx.n2361\ : std_logic;
signal \bfn_13_28_0_\ : std_logic;
signal \nx.n2293\ : std_logic;
signal \nx.n2360\ : std_logic;
signal \nx.n10915\ : std_logic;
signal \nx.n2292\ : std_logic;
signal \nx.n2359\ : std_logic;
signal \nx.n10916\ : std_logic;
signal \nx.n2291\ : std_logic;
signal \nx.n10917\ : std_logic;
signal \nx.n3006\ : std_logic;
signal \nx.n3004\ : std_logic;
signal \nx.n3006_cascade_\ : std_logic;
signal \nx.n43\ : std_logic;
signal \nx.n2999\ : std_logic;
signal \nx.n2797\ : std_logic;
signal \nx.n2864\ : std_logic;
signal \nx.n2896_cascade_\ : std_logic;
signal \nx.n43_adj_763_cascade_\ : std_logic;
signal \nx.n38_adj_762\ : std_logic;
signal \nx.n2806\ : std_logic;
signal \nx.n2873\ : std_logic;
signal \nx.bit_ctr_6\ : std_logic;
signal \nx.n2977\ : std_logic;
signal \bfn_14_19_0_\ : std_logic;
signal \nx.n2909\ : std_logic;
signal \nx.n2976\ : std_logic;
signal \nx.n11028\ : std_logic;
signal \nx.n2908\ : std_logic;
signal \nx.n2975\ : std_logic;
signal \nx.n11029\ : std_logic;
signal \nx.n2907\ : std_logic;
signal \nx.n2974\ : std_logic;
signal \nx.n11030\ : std_logic;
signal \nx.n2906\ : std_logic;
signal \nx.n2973\ : std_logic;
signal \nx.n11031\ : std_logic;
signal \nx.n2905\ : std_logic;
signal \nx.n2972\ : std_logic;
signal \nx.n11032\ : std_logic;
signal \nx.n2971\ : std_logic;
signal \nx.n11033\ : std_logic;
signal \nx.n11034\ : std_logic;
signal \nx.n11035\ : std_logic;
signal \nx.n2902\ : std_logic;
signal \nx.n2969\ : std_logic;
signal \bfn_14_20_0_\ : std_logic;
signal \nx.n2901\ : std_logic;
signal \nx.n2968\ : std_logic;
signal \nx.n11036\ : std_logic;
signal \nx.n2900\ : std_logic;
signal \nx.n2967\ : std_logic;
signal \nx.n11037\ : std_logic;
signal \nx.n2899\ : std_logic;
signal \nx.n2966\ : std_logic;
signal \nx.n11038\ : std_logic;
signal \nx.n2965\ : std_logic;
signal \nx.n11039\ : std_logic;
signal \nx.n2964\ : std_logic;
signal \nx.n11040\ : std_logic;
signal \nx.n11041\ : std_logic;
signal \nx.n2895\ : std_logic;
signal \nx.n2962\ : std_logic;
signal \nx.n11042\ : std_logic;
signal \nx.n11043\ : std_logic;
signal \bfn_14_21_0_\ : std_logic;
signal \nx.n11044\ : std_logic;
signal \nx.n2959\ : std_logic;
signal \nx.n11045\ : std_logic;
signal \nx.n11046\ : std_logic;
signal \nx.n2957\ : std_logic;
signal \nx.n11047\ : std_logic;
signal \nx.n2889\ : std_logic;
signal \nx.n2956\ : std_logic;
signal \nx.n11048\ : std_logic;
signal \nx.n2888\ : std_logic;
signal \nx.n2955\ : std_logic;
signal \nx.n11049\ : std_logic;
signal \nx.n2887\ : std_logic;
signal \nx.n2954\ : std_logic;
signal \nx.n11050\ : std_logic;
signal \nx.n11051\ : std_logic;
signal \nx.n2886\ : std_logic;
signal \nx.n2953\ : std_logic;
signal \bfn_14_22_0_\ : std_logic;
signal \nx.n2885\ : std_logic;
signal \nx.n11052\ : std_logic;
signal \nx.n2984\ : std_logic;
signal \nx.n27_adj_757\ : std_logic;
signal \nx.n36_adj_756\ : std_logic;
signal \nx.n2708\ : std_logic;
signal \nx.n2703\ : std_logic;
signal \nx.n39_adj_689\ : std_logic;
signal \nx.n25_adj_702_cascade_\ : std_logic;
signal \nx.n34_adj_701\ : std_logic;
signal \nx.n35_adj_708\ : std_logic;
signal \nx.n32_adj_703\ : std_logic;
signal \nx.n37_adj_709_cascade_\ : std_logic;
signal \nx.n31_adj_707\ : std_logic;
signal \nx.n2423_cascade_\ : std_logic;
signal \nx.n2374\ : std_logic;
signal \nx.bit_ctr_11\ : std_logic;
signal \nx.n2477\ : std_logic;
signal \bfn_14_24_0_\ : std_logic;
signal \nx.n10918\ : std_logic;
signal \nx.n2408\ : std_logic;
signal \nx.n2475\ : std_logic;
signal \nx.n10919\ : std_logic;
signal \nx.n2407\ : std_logic;
signal \nx.n2474\ : std_logic;
signal \nx.n10920\ : std_logic;
signal \nx.n2406\ : std_logic;
signal \nx.n2473\ : std_logic;
signal \nx.n10921\ : std_logic;
signal \nx.n2405\ : std_logic;
signal \nx.n2472\ : std_logic;
signal \nx.n10922\ : std_logic;
signal \nx.n2404\ : std_logic;
signal \nx.n2471\ : std_logic;
signal \nx.n10923\ : std_logic;
signal \nx.n2403\ : std_logic;
signal \nx.n2470\ : std_logic;
signal \nx.n10924\ : std_logic;
signal \nx.n10925\ : std_logic;
signal \nx.n2402\ : std_logic;
signal \nx.n2469\ : std_logic;
signal \bfn_14_25_0_\ : std_logic;
signal \nx.n2401\ : std_logic;
signal \nx.n2468\ : std_logic;
signal \nx.n10926\ : std_logic;
signal \nx.n10927\ : std_logic;
signal \nx.n2399\ : std_logic;
signal \nx.n2466\ : std_logic;
signal \nx.n10928\ : std_logic;
signal \nx.n10929\ : std_logic;
signal \nx.n10930\ : std_logic;
signal \nx.n10931\ : std_logic;
signal \nx.n10932\ : std_logic;
signal \nx.n10933\ : std_logic;
signal \bfn_14_26_0_\ : std_logic;
signal \nx.n10934\ : std_logic;
signal \nx.n10935\ : std_logic;
signal \nx.n10936\ : std_logic;
signal \nx.n2390\ : std_logic;
signal \nx.n10937\ : std_logic;
signal pin_oe_18 : std_logic;
signal \nx.n2295\ : std_logic;
signal \nx.n2362\ : std_logic;
signal \nx.n2297\ : std_logic;
signal \nx.n2364\ : std_logic;
signal \nx.n2298\ : std_logic;
signal \nx.n2365\ : std_logic;
signal \nx.n2168\ : std_logic;
signal \nx.n2101\ : std_logic;
signal \nx.n2126\ : std_logic;
signal \nx.n2200\ : std_logic;
signal \nx.n2301\ : std_logic;
signal \nx.n2368\ : std_logic;
signal \n7602_cascade_\ : std_logic;
signal \n7730_cascade_\ : std_logic;
signal pin_oe_9 : std_logic;
signal pin_oe_10 : std_logic;
signal n11960 : std_logic;
signal n2618 : std_logic;
signal pin_oe_3 : std_logic;
signal \n8_adj_825_cascade_\ : std_logic;
signal pin_out_9 : std_logic;
signal \n6_adj_813_cascade_\ : std_logic;
signal n11974 : std_logic;
signal \nx.n2890\ : std_logic;
signal \nx.n30_adj_759\ : std_logic;
signal \nx.n39_adj_761\ : std_logic;
signal \nx.n42_adj_765\ : std_logic;
signal \nx.n45_adj_769_cascade_\ : std_logic;
signal \nx.n47_adj_770\ : std_logic;
signal \nx.n2896\ : std_logic;
signal \nx.n2918_cascade_\ : std_logic;
signal \nx.n2963\ : std_logic;
signal \nx.n2970\ : std_logic;
signal \nx.n3002\ : std_logic;
signal \nx.n2995\ : std_logic;
signal \nx.n3002_cascade_\ : std_logic;
signal \nx.n42\ : std_logic;
signal \nx.n2958\ : std_logic;
signal \nx.n2891\ : std_logic;
signal \nx.n2990\ : std_logic;
signal \nx.n2804\ : std_logic;
signal \nx.n2871\ : std_logic;
signal \nx.n2903\ : std_logic;
signal \nx.n2793\ : std_logic;
signal \nx.n2860\ : std_logic;
signal \nx.n2892\ : std_logic;
signal \nx.n2960\ : std_logic;
signal \nx.n2992\ : std_logic;
signal \nx.n2794\ : std_logic;
signal \nx.n2861\ : std_logic;
signal \nx.n2819\ : std_logic;
signal \nx.n2893\ : std_logic;
signal \nx.n2898\ : std_logic;
signal \nx.n2904\ : std_logic;
signal \nx.n2893_cascade_\ : std_logic;
signal \nx.n2897\ : std_logic;
signal \nx.n41_adj_768\ : std_logic;
signal \nx.n2894\ : std_logic;
signal \nx.n2918\ : std_logic;
signal \nx.n2961\ : std_logic;
signal \nx.n2993\ : std_logic;
signal \nx.n40\ : std_logic;
signal \nx.n2609_cascade_\ : std_logic;
signal \nx.n28\ : std_logic;
signal \nx.n2606_cascade_\ : std_logic;
signal \nx.n2705\ : std_logic;
signal \nx.n2704\ : std_logic;
signal \nx.n37_adj_772_cascade_\ : std_logic;
signal \nx.n39_adj_773\ : std_logic;
signal \nx.n2522_cascade_\ : std_logic;
signal \nx.n2592_cascade_\ : std_logic;
signal \nx.n35\ : std_logic;
signal \nx.n2391\ : std_logic;
signal \nx.n2458\ : std_logic;
signal \nx.n2490_cascade_\ : std_logic;
signal \nx.n22_adj_755\ : std_logic;
signal \nx.n2324\ : std_logic;
signal \nx.n2307\ : std_logic;
signal \nx.n13321\ : std_logic;
signal \nx.n2505_cascade_\ : std_logic;
signal \nx.n2476\ : std_logic;
signal \nx.n2409\ : std_logic;
signal \nx.n2400\ : std_logic;
signal \nx.n2467\ : std_logic;
signal \nx.n2396\ : std_logic;
signal \nx.n2463\ : std_logic;
signal \nx.n2495_cascade_\ : std_logic;
signal \nx.n34_adj_758\ : std_logic;
signal \nx.n2398\ : std_logic;
signal \nx.n2465\ : std_logic;
signal \nx.n2395\ : std_logic;
signal \nx.n2462\ : std_logic;
signal \nx.n2397\ : std_logic;
signal \nx.n2464\ : std_logic;
signal \nx.n2496_cascade_\ : std_logic;
signal \nx.n2394\ : std_logic;
signal \nx.n2461\ : std_logic;
signal pin_oe_22 : std_logic;
signal \nx.n2392\ : std_logic;
signal \nx.n2459\ : std_logic;
signal \nx.n2491_cascade_\ : std_logic;
signal \nx.n33_adj_767\ : std_logic;
signal \nx.n2460\ : std_logic;
signal \nx.n2393\ : std_logic;
signal \nx.n2423\ : std_logic;
signal n7992 : std_logic;
signal n7602 : std_logic;
signal pin_oe_11 : std_logic;
signal n9 : std_logic;
signal \n9_cascade_\ : std_logic;
signal \n8_adj_820_cascade_\ : std_logic;
signal \n6_adj_805_cascade_\ : std_logic;
signal n1788 : std_logic;
signal \n9488_cascade_\ : std_logic;
signal \n7_adj_818_cascade_\ : std_logic;
signal n7_adj_821 : std_logic;
signal pin_out_3 : std_logic;
signal pin_out_2 : std_logic;
signal \n13355_cascade_\ : std_logic;
signal n13354 : std_logic;
signal \n7_adj_840_cascade_\ : std_logic;
signal pin_out_0 : std_logic;
signal n8_adj_817 : std_logic;
signal pin_out_1 : std_logic;
signal n11952 : std_logic;
signal pin_oe_8 : std_logic;
signal \nx.bit_ctr_9\ : std_logic;
signal \nx.n2677\ : std_logic;
signal \bfn_16_21_0_\ : std_logic;
signal \nx.n2609\ : std_logic;
signal \nx.n2676\ : std_logic;
signal \nx.n10959\ : std_logic;
signal \nx.n2608\ : std_logic;
signal \nx.n2675\ : std_logic;
signal \nx.n10960\ : std_logic;
signal \nx.n2607\ : std_logic;
signal \nx.n2674\ : std_logic;
signal \nx.n10961\ : std_logic;
signal \nx.n2606\ : std_logic;
signal \nx.n2673\ : std_logic;
signal \nx.n10962\ : std_logic;
signal \nx.n2605\ : std_logic;
signal \nx.n2672\ : std_logic;
signal \nx.n10963\ : std_logic;
signal \nx.n2604\ : std_logic;
signal \nx.n2671\ : std_logic;
signal \nx.n10964\ : std_logic;
signal \nx.n2603\ : std_logic;
signal \nx.n2670\ : std_logic;
signal \nx.n10965\ : std_logic;
signal \nx.n10966\ : std_logic;
signal \nx.n2602\ : std_logic;
signal \nx.n2669\ : std_logic;
signal \bfn_16_22_0_\ : std_logic;
signal \nx.n2601\ : std_logic;
signal \nx.n2668\ : std_logic;
signal \nx.n10967\ : std_logic;
signal \nx.n2600\ : std_logic;
signal \nx.n2667\ : std_logic;
signal \nx.n10968\ : std_logic;
signal \nx.n2599\ : std_logic;
signal \nx.n2666\ : std_logic;
signal \nx.n10969\ : std_logic;
signal \nx.n2598\ : std_logic;
signal \nx.n2665\ : std_logic;
signal \nx.n10970\ : std_logic;
signal \nx.n2597\ : std_logic;
signal \nx.n2664\ : std_logic;
signal \nx.n10971\ : std_logic;
signal \nx.n2596\ : std_logic;
signal \nx.n2663\ : std_logic;
signal \nx.n10972\ : std_logic;
signal \nx.n2595\ : std_logic;
signal \nx.n2662\ : std_logic;
signal \nx.n10973\ : std_logic;
signal \nx.n10974\ : std_logic;
signal \nx.n2594\ : std_logic;
signal \nx.n2661\ : std_logic;
signal \bfn_16_23_0_\ : std_logic;
signal \nx.n2593\ : std_logic;
signal \nx.n2660\ : std_logic;
signal \nx.n10975\ : std_logic;
signal \nx.n2592\ : std_logic;
signal \nx.n2659\ : std_logic;
signal \nx.n10976\ : std_logic;
signal \nx.n2591\ : std_logic;
signal \nx.n2658\ : std_logic;
signal \nx.n10977\ : std_logic;
signal \nx.n2590\ : std_logic;
signal \nx.n2657\ : std_logic;
signal \nx.n10978\ : std_logic;
signal \nx.n2656\ : std_logic;
signal \nx.n10979\ : std_logic;
signal \nx.n2621\ : std_logic;
signal \nx.n10980\ : std_logic;
signal \nx.n2687\ : std_logic;
signal \nx.n2589\ : std_logic;
signal \nx.bit_ctr_10\ : std_logic;
signal \nx.n2577\ : std_logic;
signal \bfn_16_24_0_\ : std_logic;
signal \nx.n2509\ : std_logic;
signal \nx.n2576\ : std_logic;
signal \nx.n10938\ : std_logic;
signal \nx.n2508\ : std_logic;
signal \nx.n2575\ : std_logic;
signal \nx.n10939\ : std_logic;
signal \nx.n2507\ : std_logic;
signal \nx.n2574\ : std_logic;
signal \nx.n10940\ : std_logic;
signal \nx.n2506\ : std_logic;
signal \nx.n2573\ : std_logic;
signal \nx.n10941\ : std_logic;
signal \nx.n2505\ : std_logic;
signal \nx.n2572\ : std_logic;
signal \nx.n10942\ : std_logic;
signal \nx.n2504\ : std_logic;
signal \nx.n2571\ : std_logic;
signal \nx.n10943\ : std_logic;
signal \nx.n2503\ : std_logic;
signal \nx.n2570\ : std_logic;
signal \nx.n10944\ : std_logic;
signal \nx.n10945\ : std_logic;
signal \nx.n2502\ : std_logic;
signal \nx.n2569\ : std_logic;
signal \bfn_16_25_0_\ : std_logic;
signal \nx.n2501\ : std_logic;
signal \nx.n2568\ : std_logic;
signal \nx.n10946\ : std_logic;
signal \nx.n2500\ : std_logic;
signal \nx.n2567\ : std_logic;
signal \nx.n10947\ : std_logic;
signal \nx.n2499\ : std_logic;
signal \nx.n2566\ : std_logic;
signal \nx.n10948\ : std_logic;
signal \nx.n2498\ : std_logic;
signal \nx.n2565\ : std_logic;
signal \nx.n10949\ : std_logic;
signal \nx.n2497\ : std_logic;
signal \nx.n2564\ : std_logic;
signal \nx.n10950\ : std_logic;
signal \nx.n2496\ : std_logic;
signal \nx.n2563\ : std_logic;
signal \nx.n10951\ : std_logic;
signal \nx.n2495\ : std_logic;
signal \nx.n2562\ : std_logic;
signal \nx.n10952\ : std_logic;
signal \nx.n10953\ : std_logic;
signal \nx.n2494\ : std_logic;
signal \nx.n2561\ : std_logic;
signal \bfn_16_26_0_\ : std_logic;
signal \nx.n2493\ : std_logic;
signal \nx.n2560\ : std_logic;
signal \nx.n10954\ : std_logic;
signal \nx.n2492\ : std_logic;
signal \nx.n2559\ : std_logic;
signal \nx.n10955\ : std_logic;
signal \nx.n2491\ : std_logic;
signal \nx.n2558\ : std_logic;
signal \nx.n10956\ : std_logic;
signal \nx.n2490\ : std_logic;
signal \nx.n2557\ : std_logic;
signal \nx.n10957\ : std_logic;
signal \CONSTANT_ONE_NET\ : std_logic;
signal \nx.n2489\ : std_logic;
signal \nx.n2522\ : std_logic;
signal \nx.n10958\ : std_logic;
signal \nx.n2588\ : std_logic;
signal pin_oe_12 : std_logic;
signal n45 : std_logic;
signal \bfn_17_15_0_\ : std_logic;
signal n10700 : std_logic;
signal n10701 : std_logic;
signal n10702 : std_logic;
signal n10703 : std_logic;
signal n10704 : std_logic;
signal n10705 : std_logic;
signal n13603 : std_logic;
signal n10706 : std_logic;
signal n7681 : std_logic;
signal n11824 : std_logic;
signal \bfn_17_17_0_\ : std_logic;
signal n10575 : std_logic;
signal n10576 : std_logic;
signal n10577 : std_logic;
signal n10578 : std_logic;
signal current_pin_5 : std_logic;
signal n10579 : std_logic;
signal current_pin_6 : std_logic;
signal n10580 : std_logic;
signal n10581 : std_logic;
signal current_pin_7 : std_logic;
signal n7985 : std_logic;
signal n7635 : std_logic;
signal \n9_adj_824_cascade_\ : std_logic;
signal \n8_adj_822_cascade_\ : std_logic;
signal pin_out_5 : std_logic;
signal pin_out_4 : std_logic;
signal \n13357_cascade_\ : std_logic;
signal n13625 : std_logic;
signal \n6_adj_810_cascade_\ : std_logic;
signal n11874 : std_logic;
signal n11823 : std_logic;
signal n7 : std_logic;
signal \n7_adj_823_cascade_\ : std_logic;
signal pin_oe_19 : std_logic;
signal pin_out_7 : std_logic;
signal pin_out_6 : std_logic;
signal n13358 : std_logic;
signal n3762 : std_logic;
signal n11964 : std_logic;
signal pin_oe_16 : std_logic;
signal n11820 : std_logic;
signal counter_7 : std_logic;
signal counter_0 : std_logic;
signal counter_6 : std_logic;
signal counter_1 : std_logic;
signal \n10_cascade_\ : std_logic;
signal counter_4 : std_logic;
signal counter_5 : std_logic;
signal counter_2 : std_logic;
signal counter_3 : std_logic;
signal n14 : std_logic;
signal pin_out_11 : std_logic;
signal \n7_adj_827_cascade_\ : std_logic;
signal pin_out_10 : std_logic;
signal \n9675_cascade_\ : std_logic;
signal n8_adj_832 : std_logic;
signal \pin_out_22__N_216\ : std_logic;
signal \pin_out_22__N_216_cascade_\ : std_logic;
signal n13370 : std_logic;
signal n13369 : std_logic;
signal \n13640_cascade_\ : std_logic;
signal n13628 : std_logic;
signal n13540 : std_logic;
signal current_pin_4 : std_logic;
signal \n7_adj_797_cascade_\ : std_logic;
signal n13551 : std_logic;
signal \state_7_N_167_2\ : std_logic;
signal n26 : std_logic;
signal \n11825_cascade_\ : std_logic;
signal pin_oe_15 : std_logic;
signal n1907 : std_logic;
signal state_1 : std_logic;
signal state_2 : std_logic;
signal n8025 : std_logic;
signal \n11954_cascade_\ : std_logic;
signal pin_oe_20 : std_logic;
signal n9488 : std_logic;
signal n11821 : std_logic;
signal n8_adj_826 : std_logic;
signal pin_out_8 : std_logic;
signal \n11962_cascade_\ : std_logic;
signal pin_oe_14 : std_logic;
signal n9_adj_812 : std_logic;
signal n8_adj_828 : std_logic;
signal \n11958_cascade_\ : std_logic;
signal pin_oe_21 : std_logic;
signal n13652 : std_logic;
signal \n13536_cascade_\ : std_logic;
signal n13616 : std_logic;
signal n13542 : std_logic;
signal \n7_adj_831_cascade_\ : std_logic;
signal n6_adj_813 : std_logic;
signal \n7_adj_833_cascade_\ : std_logic;
signal n8_adj_836 : std_logic;
signal n7_adj_811 : std_logic;
signal \n7_adj_835_cascade_\ : std_logic;
signal n6_adj_810 : std_logic;
signal \n7_adj_839_cascade_\ : std_logic;
signal pin_out_18 : std_logic;
signal pin_out_19 : std_logic;
signal n7_adj_797 : std_logic;
signal n6 : std_logic;
signal n6_adj_819 : std_logic;
signal \n8_adj_834_cascade_\ : std_logic;
signal pin_out_17 : std_logic;
signal n13631 : std_logic;
signal pin_out_16 : std_logic;
signal \n13634_cascade_\ : std_logic;
signal n13389 : std_logic;
signal n7_adj_838 : std_logic;
signal n7_adj_837 : std_logic;
signal pin_out_21 : std_logic;
signal pin_out_20 : std_logic;
signal pin_out_22 : std_logic;
signal \n19_adj_790_cascade_\ : std_logic;
signal n13388 : std_logic;
signal \n13375_cascade_\ : std_logic;
signal n13637 : std_logic;
signal n8_adj_829 : std_logic;
signal pin_out_12 : std_logic;
signal n9675 : std_logic;
signal n7_adj_830 : std_logic;
signal n11789 : std_logic;
signal pin_out_13 : std_logic;
signal pin_out_15 : std_logic;
signal pin_out_14 : std_logic;
signal n13376 : std_logic;
signal n11956 : std_logic;
signal pin_oe_13 : std_logic;
signal current_pin_2 : std_logic;
signal current_pin_3 : std_logic;
signal n13465 : std_logic;
signal pin_in_15 : std_logic;
signal pin_in_14 : std_logic;
signal pin_in_13 : std_logic;
signal \n13643_cascade_\ : std_logic;
signal pin_in_12 : std_logic;
signal n13646 : std_logic;
signal n11822 : std_logic;
signal state_0 : std_logic;
signal n7730 : std_logic;
signal pin_oe_17 : std_logic;
signal \CLK_c\ : std_logic;
signal pin_in_22 : std_logic;
signal n13352 : std_logic;
signal pin_in_17 : std_logic;
signal pin_in_16 : std_logic;
signal n13610 : std_logic;
signal pin_in_19 : std_logic;
signal pin_in_18 : std_logic;
signal current_pin_1 : std_logic;
signal n13607 : std_logic;
signal current_pin_0 : std_logic;
signal pin_in_21 : std_logic;
signal pin_in_20 : std_logic;
signal n19_adj_789 : std_logic;
signal \_gnd_net_\ : std_logic;

signal \LED_wire\ : std_logic;
signal \NEOPXL_wire\ : std_logic;
signal \CLK_wire\ : std_logic;

begin
    LED <= \LED_wire\;
    NEOPXL <= \NEOPXL_wire\;
    \CLK_wire\ <= CLK;

    \LED_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__47950\,
            DIN => \N__47949\,
            DOUT => \N__47948\,
            PACKAGEPIN => \LED_wire\
        );

    \LED_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__47950\,
            PADOUT => \N__47949\,
            PADIN => \N__47948\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__26619\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \NEOPXL_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__47941\,
            DIN => \N__47940\,
            DOUT => \N__47939\,
            PACKAGEPIN => \NEOPXL_wire\
        );

    \NEOPXL_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__47941\,
            PADOUT => \N__47940\,
            PADIN => \N__47939\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__24873\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \pin0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '1'
        )
    port map (
            OE => \N__47932\,
            DIN => \N__47931\,
            DOUT => \N__47930\,
            PACKAGEPIN => USBPU
        );

    \pin0_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "101001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__47932\,
            PADOUT => \N__47931\,
            PADIN => \N__47930\,
            CLOCKENABLE => 'H',
            DIN0 => pin_in_0,
            DIN1 => OPEN,
            DOUT0 => \N__39036\,
            DOUT1 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => \N__32448\
        );

    \pin1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '1'
        )
    port map (
            OE => \N__47923\,
            DIN => \N__47922\,
            DOUT => \N__47921\,
            PACKAGEPIN => ENCODER0_A
        );

    \pin1_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "101001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__47923\,
            PADOUT => \N__47922\,
            PADIN => \N__47921\,
            CLOCKENABLE => 'H',
            DIN0 => pin_in_1,
            DIN1 => OPEN,
            DOUT0 => \N__38997\,
            DOUT1 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => \N__19020\
        );

    \pin10_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '1'
        )
    port map (
            OE => \N__47914\,
            DIN => \N__47913\,
            DOUT => \N__47912\,
            PACKAGEPIN => TX
        );

    \pin10_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "101001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__47914\,
            PADOUT => \N__47913\,
            PADIN => \N__47912\,
            CLOCKENABLE => 'H',
            DIN0 => pin_in_10,
            DIN1 => OPEN,
            DOUT0 => \N__43026\,
            DOUT1 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => \N__36756\
        );

    \pin11_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '1'
        )
    port map (
            OE => \N__47905\,
            DIN => \N__47904\,
            DOUT => \N__47903\,
            PACKAGEPIN => RX
        );

    \pin11_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "101001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__47905\,
            PADOUT => \N__47904\,
            PADIN => \N__47903\,
            CLOCKENABLE => 'H',
            DIN0 => pin_in_11,
            DIN1 => OPEN,
            DOUT0 => \N__43056\,
            DOUT1 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => \N__38364\
        );

    \pin12_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '1'
        )
    port map (
            OE => \N__47896\,
            DIN => \N__47895\,
            DOUT => \N__47894\,
            PACKAGEPIN => CS_CLK
        );

    \pin12_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "101001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__47896\,
            PADOUT => \N__47895\,
            PADIN => \N__47894\,
            CLOCKENABLE => 'H',
            DIN0 => pin_in_12,
            DIN1 => OPEN,
            DOUT0 => \N__46185\,
            DOUT1 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => \N__40779\
        );

    \pin13_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '1'
        )
    port map (
            OE => \N__47887\,
            DIN => \N__47886\,
            DOUT => \N__47885\,
            PACKAGEPIN => CS
        );

    \pin13_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "101001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__47887\,
            PADOUT => \N__47886\,
            PADIN => \N__47885\,
            CLOCKENABLE => 'H',
            DIN0 => pin_in_13,
            DIN1 => OPEN,
            DOUT0 => \N__45819\,
            DOUT1 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => \N__45723\
        );

    \pin14_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '1'
        )
    port map (
            OE => \N__47878\,
            DIN => \N__47877\,
            DOUT => \N__47876\,
            PACKAGEPIN => CS_MISO
        );

    \pin14_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "101001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__47878\,
            PADOUT => \N__47877\,
            PADIN => \N__47876\,
            CLOCKENABLE => 'H',
            DIN0 => pin_in_14,
            DIN1 => OPEN,
            DOUT0 => \N__45768\,
            DOUT1 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => \N__44247\
        );

    \pin15_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '1'
        )
    port map (
            OE => \N__47869\,
            DIN => \N__47868\,
            DOUT => \N__47867\,
            PACKAGEPIN => SCL
        );

    \pin15_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "101001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__47869\,
            PADOUT => \N__47868\,
            PADIN => \N__47867\,
            CLOCKENABLE => 'H',
            DIN0 => pin_in_15,
            DIN1 => OPEN,
            DOUT0 => \N__45798\,
            DOUT1 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => \N__44004\
        );

    \pin16_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '1'
        )
    port map (
            OE => \N__47860\,
            DIN => \N__47859\,
            DOUT => \N__47858\,
            PACKAGEPIN => SDA
        );

    \pin16_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "101001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__47860\,
            PADOUT => \N__47859\,
            PADIN => \N__47858\,
            CLOCKENABLE => 'H',
            DIN0 => pin_in_16,
            DIN1 => OPEN,
            DOUT0 => \N__44718\,
            DOUT1 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => \N__42834\
        );

    \pin17_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '1'
        )
    port map (
            OE => \N__47851\,
            DIN => \N__47850\,
            DOUT => \N__47849\,
            PACKAGEPIN => INLC
        );

    \pin17_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "101001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__47851\,
            PADOUT => \N__47850\,
            PADIN => \N__47849\,
            CLOCKENABLE => 'H',
            DIN0 => pin_in_17,
            DIN1 => OPEN,
            DOUT0 => \N__44751\,
            DOUT1 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => \N__46950\
        );

    \pin18_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '1'
        )
    port map (
            OE => \N__47842\,
            DIN => \N__47841\,
            DOUT => \N__47840\,
            PACKAGEPIN => INHC
        );

    \pin18_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "101001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__47842\,
            PADOUT => \N__47841\,
            PADIN => \N__47840\,
            CLOCKENABLE => 'H',
            DIN0 => pin_in_18,
            DIN1 => OPEN,
            DOUT0 => \N__44325\,
            DOUT1 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => \N__36339\
        );

    \pin19_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '1'
        )
    port map (
            OE => \N__47833\,
            DIN => \N__47832\,
            DOUT => \N__47831\,
            PACKAGEPIN => INLB
        );

    \pin19_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "101001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__47833\,
            PADOUT => \N__47832\,
            PADIN => \N__47831\,
            CLOCKENABLE => 'H',
            DIN0 => pin_in_19,
            DIN1 => OPEN,
            DOUT0 => \N__44292\,
            DOUT1 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => \N__42990\
        );

    \pin2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '1'
        )
    port map (
            OE => \N__47824\,
            DIN => \N__47823\,
            DOUT => \N__47822\,
            PACKAGEPIN => ENCODER0_B
        );

    \pin2_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "101001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__47824\,
            PADOUT => \N__47823\,
            PADIN => \N__47822\,
            CLOCKENABLE => 'H',
            DIN0 => pin_in_2,
            DIN1 => OPEN,
            DOUT0 => \N__38688\,
            DOUT1 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => \N__24792\
        );

    \pin20_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '1'
        )
    port map (
            OE => \N__47815\,
            DIN => \N__47814\,
            DOUT => \N__47813\,
            PACKAGEPIN => INHB
        );

    \pin20_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "101001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__47815\,
            PADOUT => \N__47814\,
            PADIN => \N__47813\,
            CLOCKENABLE => 'H',
            DIN0 => pin_in_20,
            DIN1 => OPEN,
            DOUT0 => \N__44619\,
            DOUT1 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => \N__43455\
        );

    \pin21_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '1'
        )
    port map (
            OE => \N__47806\,
            DIN => \N__47805\,
            DOUT => \N__47804\,
            PACKAGEPIN => INLA
        );

    \pin21_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "101001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__47806\,
            PADOUT => \N__47805\,
            PADIN => \N__47804\,
            CLOCKENABLE => 'H',
            DIN0 => pin_in_21,
            DIN1 => OPEN,
            DOUT0 => \N__44655\,
            DOUT1 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => \N__44187\
        );

    \pin22_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '1'
        )
    port map (
            OE => \N__47797\,
            DIN => \N__47796\,
            DOUT => \N__47795\,
            PACKAGEPIN => INHA
        );

    \pin22_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "101001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__47797\,
            PADOUT => \N__47796\,
            PADIN => \N__47795\,
            CLOCKENABLE => 'H',
            DIN0 => pin_in_22,
            DIN1 => OPEN,
            DOUT0 => \N__44595\,
            DOUT1 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => \N__38616\
        );

    \pin3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '1'
        )
    port map (
            OE => \N__47788\,
            DIN => \N__47787\,
            DOUT => \N__47786\,
            PACKAGEPIN => ENCODER1_A
        );

    \pin3_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "101001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__47788\,
            PADOUT => \N__47787\,
            PADIN => \N__47786\,
            CLOCKENABLE => 'H',
            DIN0 => pin_in_3,
            DIN1 => OPEN,
            DOUT0 => \N__38721\,
            DOUT1 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => \N__36723\
        );

    \pin4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '1'
        )
    port map (
            OE => \N__47779\,
            DIN => \N__47778\,
            DOUT => \N__47777\,
            PACKAGEPIN => ENCODER1_B
        );

    \pin4_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "101001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__47779\,
            PADOUT => \N__47778\,
            PADIN => \N__47777\,
            CLOCKENABLE => 'H',
            DIN0 => pin_in_4,
            DIN1 => OPEN,
            DOUT0 => \N__42705\,
            DOUT1 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => \N__32475\
        );

    \pin5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '1'
        )
    port map (
            OE => \N__47770\,
            DIN => \N__47769\,
            DOUT => \N__47768\,
            PACKAGEPIN => HALL1
        );

    \pin5_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "101001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__47770\,
            PADOUT => \N__47769\,
            PADIN => \N__47768\,
            CLOCKENABLE => 'H',
            DIN0 => pin_in_5,
            DIN1 => OPEN,
            DOUT0 => \N__42735\,
            DOUT1 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => \N__19167\
        );

    \pin6_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '1'
        )
    port map (
            OE => \N__47761\,
            DIN => \N__47760\,
            DOUT => \N__47759\,
            PACKAGEPIN => HALL2
        );

    \pin6_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "101001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__47761\,
            PADOUT => \N__47760\,
            PADIN => \N__47759\,
            CLOCKENABLE => 'H',
            DIN0 => pin_in_6,
            DIN1 => OPEN,
            DOUT0 => \N__42927\,
            DOUT1 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => \N__21192\
        );

    \pin7_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '1'
        )
    port map (
            OE => \N__47752\,
            DIN => \N__47751\,
            DOUT => \N__47750\,
            PACKAGEPIN => HALL3
        );

    \pin7_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "101001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__47752\,
            PADOUT => \N__47751\,
            PADIN => \N__47750\,
            CLOCKENABLE => 'H',
            DIN0 => pin_in_7,
            DIN1 => OPEN,
            DOUT0 => \N__42966\,
            DOUT1 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => \N__24396\
        );

    \pin8_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '1'
        )
    port map (
            OE => \N__47743\,
            DIN => \N__47742\,
            DOUT => \N__47741\,
            PACKAGEPIN => FAULT_N
        );

    \pin8_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "101001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__47743\,
            PADOUT => \N__47742\,
            PADIN => \N__47741\,
            CLOCKENABLE => 'H',
            DIN0 => pin_in_8,
            DIN1 => OPEN,
            DOUT0 => \N__43353\,
            DOUT1 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => \N__38952\
        );

    \pin9_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '1'
        )
    port map (
            OE => \N__47734\,
            DIN => \N__47733\,
            DOUT => \N__47732\,
            PACKAGEPIN => DE
        );

    \pin9_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "101001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__47734\,
            PADOUT => \N__47733\,
            PADIN => \N__47732\,
            CLOCKENABLE => 'H',
            DIN0 => pin_in_9,
            DIN1 => OPEN,
            DOUT0 => \N__36699\,
            DOUT1 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => \N__36777\
        );

    \CLK_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__47725\,
            DIN => \N__47724\,
            DOUT => \N__47723\,
            PACKAGEPIN => \CLK_wire\
        );

    \CLK_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__47725\,
            PADOUT => \N__47724\,
            PADIN => \N__47723\,
            CLOCKENABLE => 'H',
            DIN0 => \CLK_pad_gb_input\,
            DIN1 => OPEN,
            DOUT0 => '0',
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \I__11563\ : InMux
    port map (
            O => \N__47706\,
            I => \N__47703\
        );

    \I__11562\ : LocalMux
    port map (
            O => \N__47703\,
            I => \N__47700\
        );

    \I__11561\ : Odrv12
    port map (
            O => \N__47700\,
            I => n11822
        );

    \I__11560\ : CascadeMux
    port map (
            O => \N__47697\,
            I => \N__47690\
        );

    \I__11559\ : CascadeMux
    port map (
            O => \N__47696\,
            I => \N__47687\
        );

    \I__11558\ : CascadeMux
    port map (
            O => \N__47695\,
            I => \N__47684\
        );

    \I__11557\ : CascadeMux
    port map (
            O => \N__47694\,
            I => \N__47681\
        );

    \I__11556\ : InMux
    port map (
            O => \N__47693\,
            I => \N__47678\
        );

    \I__11555\ : InMux
    port map (
            O => \N__47690\,
            I => \N__47669\
        );

    \I__11554\ : InMux
    port map (
            O => \N__47687\,
            I => \N__47660\
        );

    \I__11553\ : InMux
    port map (
            O => \N__47684\,
            I => \N__47654\
        );

    \I__11552\ : InMux
    port map (
            O => \N__47681\,
            I => \N__47651\
        );

    \I__11551\ : LocalMux
    port map (
            O => \N__47678\,
            I => \N__47648\
        );

    \I__11550\ : CascadeMux
    port map (
            O => \N__47677\,
            I => \N__47643\
        );

    \I__11549\ : CascadeMux
    port map (
            O => \N__47676\,
            I => \N__47638\
        );

    \I__11548\ : CascadeMux
    port map (
            O => \N__47675\,
            I => \N__47632\
        );

    \I__11547\ : CascadeMux
    port map (
            O => \N__47674\,
            I => \N__47628\
        );

    \I__11546\ : InMux
    port map (
            O => \N__47673\,
            I => \N__47625\
        );

    \I__11545\ : InMux
    port map (
            O => \N__47672\,
            I => \N__47621\
        );

    \I__11544\ : LocalMux
    port map (
            O => \N__47669\,
            I => \N__47618\
        );

    \I__11543\ : InMux
    port map (
            O => \N__47668\,
            I => \N__47611\
        );

    \I__11542\ : InMux
    port map (
            O => \N__47667\,
            I => \N__47611\
        );

    \I__11541\ : InMux
    port map (
            O => \N__47666\,
            I => \N__47611\
        );

    \I__11540\ : InMux
    port map (
            O => \N__47665\,
            I => \N__47607\
        );

    \I__11539\ : InMux
    port map (
            O => \N__47664\,
            I => \N__47604\
        );

    \I__11538\ : CascadeMux
    port map (
            O => \N__47663\,
            I => \N__47601\
        );

    \I__11537\ : LocalMux
    port map (
            O => \N__47660\,
            I => \N__47595\
        );

    \I__11536\ : CascadeMux
    port map (
            O => \N__47659\,
            I => \N__47591\
        );

    \I__11535\ : CascadeMux
    port map (
            O => \N__47658\,
            I => \N__47587\
        );

    \I__11534\ : CascadeMux
    port map (
            O => \N__47657\,
            I => \N__47578\
        );

    \I__11533\ : LocalMux
    port map (
            O => \N__47654\,
            I => \N__47570\
        );

    \I__11532\ : LocalMux
    port map (
            O => \N__47651\,
            I => \N__47570\
        );

    \I__11531\ : Span4Mux_h
    port map (
            O => \N__47648\,
            I => \N__47570\
        );

    \I__11530\ : InMux
    port map (
            O => \N__47647\,
            I => \N__47563\
        );

    \I__11529\ : InMux
    port map (
            O => \N__47646\,
            I => \N__47563\
        );

    \I__11528\ : InMux
    port map (
            O => \N__47643\,
            I => \N__47563\
        );

    \I__11527\ : InMux
    port map (
            O => \N__47642\,
            I => \N__47560\
        );

    \I__11526\ : InMux
    port map (
            O => \N__47641\,
            I => \N__47555\
        );

    \I__11525\ : InMux
    port map (
            O => \N__47638\,
            I => \N__47555\
        );

    \I__11524\ : InMux
    port map (
            O => \N__47637\,
            I => \N__47550\
        );

    \I__11523\ : InMux
    port map (
            O => \N__47636\,
            I => \N__47550\
        );

    \I__11522\ : CascadeMux
    port map (
            O => \N__47635\,
            I => \N__47546\
        );

    \I__11521\ : InMux
    port map (
            O => \N__47632\,
            I => \N__47543\
        );

    \I__11520\ : CascadeMux
    port map (
            O => \N__47631\,
            I => \N__47540\
        );

    \I__11519\ : InMux
    port map (
            O => \N__47628\,
            I => \N__47536\
        );

    \I__11518\ : LocalMux
    port map (
            O => \N__47625\,
            I => \N__47533\
        );

    \I__11517\ : InMux
    port map (
            O => \N__47624\,
            I => \N__47530\
        );

    \I__11516\ : LocalMux
    port map (
            O => \N__47621\,
            I => \N__47523\
        );

    \I__11515\ : Span4Mux_v
    port map (
            O => \N__47618\,
            I => \N__47523\
        );

    \I__11514\ : LocalMux
    port map (
            O => \N__47611\,
            I => \N__47523\
        );

    \I__11513\ : CascadeMux
    port map (
            O => \N__47610\,
            I => \N__47520\
        );

    \I__11512\ : LocalMux
    port map (
            O => \N__47607\,
            I => \N__47509\
        );

    \I__11511\ : LocalMux
    port map (
            O => \N__47604\,
            I => \N__47509\
        );

    \I__11510\ : InMux
    port map (
            O => \N__47601\,
            I => \N__47506\
        );

    \I__11509\ : CascadeMux
    port map (
            O => \N__47600\,
            I => \N__47503\
        );

    \I__11508\ : CascadeMux
    port map (
            O => \N__47599\,
            I => \N__47499\
        );

    \I__11507\ : InMux
    port map (
            O => \N__47598\,
            I => \N__47496\
        );

    \I__11506\ : Span4Mux_h
    port map (
            O => \N__47595\,
            I => \N__47493\
        );

    \I__11505\ : InMux
    port map (
            O => \N__47594\,
            I => \N__47490\
        );

    \I__11504\ : InMux
    port map (
            O => \N__47591\,
            I => \N__47485\
        );

    \I__11503\ : InMux
    port map (
            O => \N__47590\,
            I => \N__47475\
        );

    \I__11502\ : InMux
    port map (
            O => \N__47587\,
            I => \N__47470\
        );

    \I__11501\ : InMux
    port map (
            O => \N__47586\,
            I => \N__47470\
        );

    \I__11500\ : InMux
    port map (
            O => \N__47585\,
            I => \N__47461\
        );

    \I__11499\ : InMux
    port map (
            O => \N__47584\,
            I => \N__47461\
        );

    \I__11498\ : InMux
    port map (
            O => \N__47583\,
            I => \N__47461\
        );

    \I__11497\ : InMux
    port map (
            O => \N__47582\,
            I => \N__47461\
        );

    \I__11496\ : InMux
    port map (
            O => \N__47581\,
            I => \N__47456\
        );

    \I__11495\ : InMux
    port map (
            O => \N__47578\,
            I => \N__47453\
        );

    \I__11494\ : CascadeMux
    port map (
            O => \N__47577\,
            I => \N__47450\
        );

    \I__11493\ : Span4Mux_v
    port map (
            O => \N__47570\,
            I => \N__47447\
        );

    \I__11492\ : LocalMux
    port map (
            O => \N__47563\,
            I => \N__47444\
        );

    \I__11491\ : LocalMux
    port map (
            O => \N__47560\,
            I => \N__47437\
        );

    \I__11490\ : LocalMux
    port map (
            O => \N__47555\,
            I => \N__47437\
        );

    \I__11489\ : LocalMux
    port map (
            O => \N__47550\,
            I => \N__47437\
        );

    \I__11488\ : InMux
    port map (
            O => \N__47549\,
            I => \N__47432\
        );

    \I__11487\ : InMux
    port map (
            O => \N__47546\,
            I => \N__47432\
        );

    \I__11486\ : LocalMux
    port map (
            O => \N__47543\,
            I => \N__47428\
        );

    \I__11485\ : InMux
    port map (
            O => \N__47540\,
            I => \N__47425\
        );

    \I__11484\ : InMux
    port map (
            O => \N__47539\,
            I => \N__47422\
        );

    \I__11483\ : LocalMux
    port map (
            O => \N__47536\,
            I => \N__47415\
        );

    \I__11482\ : Span4Mux_h
    port map (
            O => \N__47533\,
            I => \N__47415\
        );

    \I__11481\ : LocalMux
    port map (
            O => \N__47530\,
            I => \N__47415\
        );

    \I__11480\ : Span4Mux_h
    port map (
            O => \N__47523\,
            I => \N__47412\
        );

    \I__11479\ : InMux
    port map (
            O => \N__47520\,
            I => \N__47407\
        );

    \I__11478\ : InMux
    port map (
            O => \N__47519\,
            I => \N__47407\
        );

    \I__11477\ : InMux
    port map (
            O => \N__47518\,
            I => \N__47402\
        );

    \I__11476\ : InMux
    port map (
            O => \N__47517\,
            I => \N__47402\
        );

    \I__11475\ : InMux
    port map (
            O => \N__47516\,
            I => \N__47397\
        );

    \I__11474\ : InMux
    port map (
            O => \N__47515\,
            I => \N__47397\
        );

    \I__11473\ : InMux
    port map (
            O => \N__47514\,
            I => \N__47394\
        );

    \I__11472\ : Span4Mux_h
    port map (
            O => \N__47509\,
            I => \N__47391\
        );

    \I__11471\ : LocalMux
    port map (
            O => \N__47506\,
            I => \N__47388\
        );

    \I__11470\ : InMux
    port map (
            O => \N__47503\,
            I => \N__47385\
        );

    \I__11469\ : InMux
    port map (
            O => \N__47502\,
            I => \N__47380\
        );

    \I__11468\ : InMux
    port map (
            O => \N__47499\,
            I => \N__47380\
        );

    \I__11467\ : LocalMux
    port map (
            O => \N__47496\,
            I => \N__47377\
        );

    \I__11466\ : Span4Mux_v
    port map (
            O => \N__47493\,
            I => \N__47372\
        );

    \I__11465\ : LocalMux
    port map (
            O => \N__47490\,
            I => \N__47372\
        );

    \I__11464\ : CascadeMux
    port map (
            O => \N__47489\,
            I => \N__47369\
        );

    \I__11463\ : CascadeMux
    port map (
            O => \N__47488\,
            I => \N__47364\
        );

    \I__11462\ : LocalMux
    port map (
            O => \N__47485\,
            I => \N__47360\
        );

    \I__11461\ : InMux
    port map (
            O => \N__47484\,
            I => \N__47355\
        );

    \I__11460\ : InMux
    port map (
            O => \N__47483\,
            I => \N__47355\
        );

    \I__11459\ : InMux
    port map (
            O => \N__47482\,
            I => \N__47350\
        );

    \I__11458\ : InMux
    port map (
            O => \N__47481\,
            I => \N__47350\
        );

    \I__11457\ : InMux
    port map (
            O => \N__47480\,
            I => \N__47347\
        );

    \I__11456\ : InMux
    port map (
            O => \N__47479\,
            I => \N__47344\
        );

    \I__11455\ : InMux
    port map (
            O => \N__47478\,
            I => \N__47341\
        );

    \I__11454\ : LocalMux
    port map (
            O => \N__47475\,
            I => \N__47336\
        );

    \I__11453\ : LocalMux
    port map (
            O => \N__47470\,
            I => \N__47336\
        );

    \I__11452\ : LocalMux
    port map (
            O => \N__47461\,
            I => \N__47333\
        );

    \I__11451\ : CascadeMux
    port map (
            O => \N__47460\,
            I => \N__47330\
        );

    \I__11450\ : CascadeMux
    port map (
            O => \N__47459\,
            I => \N__47326\
        );

    \I__11449\ : LocalMux
    port map (
            O => \N__47456\,
            I => \N__47318\
        );

    \I__11448\ : LocalMux
    port map (
            O => \N__47453\,
            I => \N__47318\
        );

    \I__11447\ : InMux
    port map (
            O => \N__47450\,
            I => \N__47315\
        );

    \I__11446\ : Span4Mux_v
    port map (
            O => \N__47447\,
            I => \N__47308\
        );

    \I__11445\ : Span4Mux_h
    port map (
            O => \N__47444\,
            I => \N__47308\
        );

    \I__11444\ : Span4Mux_h
    port map (
            O => \N__47437\,
            I => \N__47308\
        );

    \I__11443\ : LocalMux
    port map (
            O => \N__47432\,
            I => \N__47305\
        );

    \I__11442\ : CascadeMux
    port map (
            O => \N__47431\,
            I => \N__47302\
        );

    \I__11441\ : Span4Mux_v
    port map (
            O => \N__47428\,
            I => \N__47296\
        );

    \I__11440\ : LocalMux
    port map (
            O => \N__47425\,
            I => \N__47277\
        );

    \I__11439\ : LocalMux
    port map (
            O => \N__47422\,
            I => \N__47277\
        );

    \I__11438\ : Sp12to4
    port map (
            O => \N__47415\,
            I => \N__47277\
        );

    \I__11437\ : Sp12to4
    port map (
            O => \N__47412\,
            I => \N__47277\
        );

    \I__11436\ : LocalMux
    port map (
            O => \N__47407\,
            I => \N__47277\
        );

    \I__11435\ : LocalMux
    port map (
            O => \N__47402\,
            I => \N__47277\
        );

    \I__11434\ : LocalMux
    port map (
            O => \N__47397\,
            I => \N__47277\
        );

    \I__11433\ : LocalMux
    port map (
            O => \N__47394\,
            I => \N__47277\
        );

    \I__11432\ : Sp12to4
    port map (
            O => \N__47391\,
            I => \N__47277\
        );

    \I__11431\ : Span4Mux_h
    port map (
            O => \N__47388\,
            I => \N__47272\
        );

    \I__11430\ : LocalMux
    port map (
            O => \N__47385\,
            I => \N__47272\
        );

    \I__11429\ : LocalMux
    port map (
            O => \N__47380\,
            I => \N__47269\
        );

    \I__11428\ : Span4Mux_h
    port map (
            O => \N__47377\,
            I => \N__47264\
        );

    \I__11427\ : Span4Mux_v
    port map (
            O => \N__47372\,
            I => \N__47264\
        );

    \I__11426\ : InMux
    port map (
            O => \N__47369\,
            I => \N__47259\
        );

    \I__11425\ : InMux
    port map (
            O => \N__47368\,
            I => \N__47259\
        );

    \I__11424\ : InMux
    port map (
            O => \N__47367\,
            I => \N__47256\
        );

    \I__11423\ : InMux
    port map (
            O => \N__47364\,
            I => \N__47251\
        );

    \I__11422\ : InMux
    port map (
            O => \N__47363\,
            I => \N__47251\
        );

    \I__11421\ : Span4Mux_h
    port map (
            O => \N__47360\,
            I => \N__47234\
        );

    \I__11420\ : LocalMux
    port map (
            O => \N__47355\,
            I => \N__47234\
        );

    \I__11419\ : LocalMux
    port map (
            O => \N__47350\,
            I => \N__47234\
        );

    \I__11418\ : LocalMux
    port map (
            O => \N__47347\,
            I => \N__47234\
        );

    \I__11417\ : LocalMux
    port map (
            O => \N__47344\,
            I => \N__47234\
        );

    \I__11416\ : LocalMux
    port map (
            O => \N__47341\,
            I => \N__47234\
        );

    \I__11415\ : Span4Mux_h
    port map (
            O => \N__47336\,
            I => \N__47234\
        );

    \I__11414\ : Span4Mux_v
    port map (
            O => \N__47333\,
            I => \N__47234\
        );

    \I__11413\ : InMux
    port map (
            O => \N__47330\,
            I => \N__47229\
        );

    \I__11412\ : InMux
    port map (
            O => \N__47329\,
            I => \N__47229\
        );

    \I__11411\ : InMux
    port map (
            O => \N__47326\,
            I => \N__47226\
        );

    \I__11410\ : InMux
    port map (
            O => \N__47325\,
            I => \N__47221\
        );

    \I__11409\ : InMux
    port map (
            O => \N__47324\,
            I => \N__47221\
        );

    \I__11408\ : InMux
    port map (
            O => \N__47323\,
            I => \N__47218\
        );

    \I__11407\ : Span4Mux_v
    port map (
            O => \N__47318\,
            I => \N__47215\
        );

    \I__11406\ : LocalMux
    port map (
            O => \N__47315\,
            I => \N__47208\
        );

    \I__11405\ : Span4Mux_v
    port map (
            O => \N__47308\,
            I => \N__47208\
        );

    \I__11404\ : Span4Mux_h
    port map (
            O => \N__47305\,
            I => \N__47208\
        );

    \I__11403\ : InMux
    port map (
            O => \N__47302\,
            I => \N__47199\
        );

    \I__11402\ : InMux
    port map (
            O => \N__47301\,
            I => \N__47199\
        );

    \I__11401\ : InMux
    port map (
            O => \N__47300\,
            I => \N__47199\
        );

    \I__11400\ : InMux
    port map (
            O => \N__47299\,
            I => \N__47199\
        );

    \I__11399\ : Sp12to4
    port map (
            O => \N__47296\,
            I => \N__47194\
        );

    \I__11398\ : Span12Mux_v
    port map (
            O => \N__47277\,
            I => \N__47194\
        );

    \I__11397\ : Span4Mux_h
    port map (
            O => \N__47272\,
            I => \N__47183\
        );

    \I__11396\ : Span4Mux_v
    port map (
            O => \N__47269\,
            I => \N__47183\
        );

    \I__11395\ : Span4Mux_h
    port map (
            O => \N__47264\,
            I => \N__47183\
        );

    \I__11394\ : LocalMux
    port map (
            O => \N__47259\,
            I => \N__47183\
        );

    \I__11393\ : LocalMux
    port map (
            O => \N__47256\,
            I => \N__47183\
        );

    \I__11392\ : LocalMux
    port map (
            O => \N__47251\,
            I => \N__47176\
        );

    \I__11391\ : Span4Mux_v
    port map (
            O => \N__47234\,
            I => \N__47176\
        );

    \I__11390\ : LocalMux
    port map (
            O => \N__47229\,
            I => \N__47176\
        );

    \I__11389\ : LocalMux
    port map (
            O => \N__47226\,
            I => state_0
        );

    \I__11388\ : LocalMux
    port map (
            O => \N__47221\,
            I => state_0
        );

    \I__11387\ : LocalMux
    port map (
            O => \N__47218\,
            I => state_0
        );

    \I__11386\ : Odrv4
    port map (
            O => \N__47215\,
            I => state_0
        );

    \I__11385\ : Odrv4
    port map (
            O => \N__47208\,
            I => state_0
        );

    \I__11384\ : LocalMux
    port map (
            O => \N__47199\,
            I => state_0
        );

    \I__11383\ : Odrv12
    port map (
            O => \N__47194\,
            I => state_0
        );

    \I__11382\ : Odrv4
    port map (
            O => \N__47183\,
            I => state_0
        );

    \I__11381\ : Odrv4
    port map (
            O => \N__47176\,
            I => state_0
        );

    \I__11380\ : InMux
    port map (
            O => \N__47157\,
            I => \N__47150\
        );

    \I__11379\ : InMux
    port map (
            O => \N__47156\,
            I => \N__47143\
        );

    \I__11378\ : InMux
    port map (
            O => \N__47155\,
            I => \N__47140\
        );

    \I__11377\ : InMux
    port map (
            O => \N__47154\,
            I => \N__47137\
        );

    \I__11376\ : InMux
    port map (
            O => \N__47153\,
            I => \N__47134\
        );

    \I__11375\ : LocalMux
    port map (
            O => \N__47150\,
            I => \N__47131\
        );

    \I__11374\ : CascadeMux
    port map (
            O => \N__47149\,
            I => \N__47127\
        );

    \I__11373\ : InMux
    port map (
            O => \N__47148\,
            I => \N__47116\
        );

    \I__11372\ : InMux
    port map (
            O => \N__47147\,
            I => \N__47113\
        );

    \I__11371\ : InMux
    port map (
            O => \N__47146\,
            I => \N__47110\
        );

    \I__11370\ : LocalMux
    port map (
            O => \N__47143\,
            I => \N__47107\
        );

    \I__11369\ : LocalMux
    port map (
            O => \N__47140\,
            I => \N__47102\
        );

    \I__11368\ : LocalMux
    port map (
            O => \N__47137\,
            I => \N__47102\
        );

    \I__11367\ : LocalMux
    port map (
            O => \N__47134\,
            I => \N__47099\
        );

    \I__11366\ : Span4Mux_v
    port map (
            O => \N__47131\,
            I => \N__47096\
        );

    \I__11365\ : InMux
    port map (
            O => \N__47130\,
            I => \N__47093\
        );

    \I__11364\ : InMux
    port map (
            O => \N__47127\,
            I => \N__47090\
        );

    \I__11363\ : InMux
    port map (
            O => \N__47126\,
            I => \N__47085\
        );

    \I__11362\ : InMux
    port map (
            O => \N__47125\,
            I => \N__47085\
        );

    \I__11361\ : InMux
    port map (
            O => \N__47124\,
            I => \N__47082\
        );

    \I__11360\ : InMux
    port map (
            O => \N__47123\,
            I => \N__47079\
        );

    \I__11359\ : InMux
    port map (
            O => \N__47122\,
            I => \N__47076\
        );

    \I__11358\ : InMux
    port map (
            O => \N__47121\,
            I => \N__47073\
        );

    \I__11357\ : InMux
    port map (
            O => \N__47120\,
            I => \N__47069\
        );

    \I__11356\ : InMux
    port map (
            O => \N__47119\,
            I => \N__47066\
        );

    \I__11355\ : LocalMux
    port map (
            O => \N__47116\,
            I => \N__47061\
        );

    \I__11354\ : LocalMux
    port map (
            O => \N__47113\,
            I => \N__47061\
        );

    \I__11353\ : LocalMux
    port map (
            O => \N__47110\,
            I => \N__47058\
        );

    \I__11352\ : Span4Mux_h
    port map (
            O => \N__47107\,
            I => \N__47053\
        );

    \I__11351\ : Span4Mux_v
    port map (
            O => \N__47102\,
            I => \N__47053\
        );

    \I__11350\ : Span4Mux_h
    port map (
            O => \N__47099\,
            I => \N__47048\
        );

    \I__11349\ : Span4Mux_h
    port map (
            O => \N__47096\,
            I => \N__47048\
        );

    \I__11348\ : LocalMux
    port map (
            O => \N__47093\,
            I => \N__47043\
        );

    \I__11347\ : LocalMux
    port map (
            O => \N__47090\,
            I => \N__47043\
        );

    \I__11346\ : LocalMux
    port map (
            O => \N__47085\,
            I => \N__47040\
        );

    \I__11345\ : LocalMux
    port map (
            O => \N__47082\,
            I => \N__47034\
        );

    \I__11344\ : LocalMux
    port map (
            O => \N__47079\,
            I => \N__47031\
        );

    \I__11343\ : LocalMux
    port map (
            O => \N__47076\,
            I => \N__47028\
        );

    \I__11342\ : LocalMux
    port map (
            O => \N__47073\,
            I => \N__47025\
        );

    \I__11341\ : InMux
    port map (
            O => \N__47072\,
            I => \N__47022\
        );

    \I__11340\ : LocalMux
    port map (
            O => \N__47069\,
            I => \N__47019\
        );

    \I__11339\ : LocalMux
    port map (
            O => \N__47066\,
            I => \N__47014\
        );

    \I__11338\ : Span4Mux_v
    port map (
            O => \N__47061\,
            I => \N__47014\
        );

    \I__11337\ : Span4Mux_h
    port map (
            O => \N__47058\,
            I => \N__47005\
        );

    \I__11336\ : Span4Mux_v
    port map (
            O => \N__47053\,
            I => \N__47005\
        );

    \I__11335\ : Span4Mux_h
    port map (
            O => \N__47048\,
            I => \N__47005\
        );

    \I__11334\ : Span4Mux_h
    port map (
            O => \N__47043\,
            I => \N__47005\
        );

    \I__11333\ : Span12Mux_v
    port map (
            O => \N__47040\,
            I => \N__47002\
        );

    \I__11332\ : InMux
    port map (
            O => \N__47039\,
            I => \N__46999\
        );

    \I__11331\ : InMux
    port map (
            O => \N__47038\,
            I => \N__46996\
        );

    \I__11330\ : InMux
    port map (
            O => \N__47037\,
            I => \N__46993\
        );

    \I__11329\ : Span4Mux_h
    port map (
            O => \N__47034\,
            I => \N__46990\
        );

    \I__11328\ : Span4Mux_v
    port map (
            O => \N__47031\,
            I => \N__46985\
        );

    \I__11327\ : Span4Mux_v
    port map (
            O => \N__47028\,
            I => \N__46985\
        );

    \I__11326\ : Span12Mux_s9_h
    port map (
            O => \N__47025\,
            I => \N__46982\
        );

    \I__11325\ : LocalMux
    port map (
            O => \N__47022\,
            I => \N__46975\
        );

    \I__11324\ : Span4Mux_v
    port map (
            O => \N__47019\,
            I => \N__46975\
        );

    \I__11323\ : Span4Mux_h
    port map (
            O => \N__47014\,
            I => \N__46975\
        );

    \I__11322\ : Span4Mux_v
    port map (
            O => \N__47005\,
            I => \N__46972\
        );

    \I__11321\ : Span12Mux_h
    port map (
            O => \N__47002\,
            I => \N__46969\
        );

    \I__11320\ : LocalMux
    port map (
            O => \N__46999\,
            I => n7730
        );

    \I__11319\ : LocalMux
    port map (
            O => \N__46996\,
            I => n7730
        );

    \I__11318\ : LocalMux
    port map (
            O => \N__46993\,
            I => n7730
        );

    \I__11317\ : Odrv4
    port map (
            O => \N__46990\,
            I => n7730
        );

    \I__11316\ : Odrv4
    port map (
            O => \N__46985\,
            I => n7730
        );

    \I__11315\ : Odrv12
    port map (
            O => \N__46982\,
            I => n7730
        );

    \I__11314\ : Odrv4
    port map (
            O => \N__46975\,
            I => n7730
        );

    \I__11313\ : Odrv4
    port map (
            O => \N__46972\,
            I => n7730
        );

    \I__11312\ : Odrv12
    port map (
            O => \N__46969\,
            I => n7730
        );

    \I__11311\ : IoInMux
    port map (
            O => \N__46950\,
            I => \N__46947\
        );

    \I__11310\ : LocalMux
    port map (
            O => \N__46947\,
            I => \N__46944\
        );

    \I__11309\ : Span4Mux_s3_v
    port map (
            O => \N__46944\,
            I => \N__46941\
        );

    \I__11308\ : Sp12to4
    port map (
            O => \N__46941\,
            I => \N__46938\
        );

    \I__11307\ : Span12Mux_s11_h
    port map (
            O => \N__46938\,
            I => \N__46935\
        );

    \I__11306\ : Span12Mux_v
    port map (
            O => \N__46935\,
            I => \N__46931\
        );

    \I__11305\ : InMux
    port map (
            O => \N__46934\,
            I => \N__46928\
        );

    \I__11304\ : Odrv12
    port map (
            O => \N__46931\,
            I => pin_oe_17
        );

    \I__11303\ : LocalMux
    port map (
            O => \N__46928\,
            I => pin_oe_17
        );

    \I__11302\ : ClkMux
    port map (
            O => \N__46923\,
            I => \N__46668\
        );

    \I__11301\ : ClkMux
    port map (
            O => \N__46922\,
            I => \N__46668\
        );

    \I__11300\ : ClkMux
    port map (
            O => \N__46921\,
            I => \N__46668\
        );

    \I__11299\ : ClkMux
    port map (
            O => \N__46920\,
            I => \N__46668\
        );

    \I__11298\ : ClkMux
    port map (
            O => \N__46919\,
            I => \N__46668\
        );

    \I__11297\ : ClkMux
    port map (
            O => \N__46918\,
            I => \N__46668\
        );

    \I__11296\ : ClkMux
    port map (
            O => \N__46917\,
            I => \N__46668\
        );

    \I__11295\ : ClkMux
    port map (
            O => \N__46916\,
            I => \N__46668\
        );

    \I__11294\ : ClkMux
    port map (
            O => \N__46915\,
            I => \N__46668\
        );

    \I__11293\ : ClkMux
    port map (
            O => \N__46914\,
            I => \N__46668\
        );

    \I__11292\ : ClkMux
    port map (
            O => \N__46913\,
            I => \N__46668\
        );

    \I__11291\ : ClkMux
    port map (
            O => \N__46912\,
            I => \N__46668\
        );

    \I__11290\ : ClkMux
    port map (
            O => \N__46911\,
            I => \N__46668\
        );

    \I__11289\ : ClkMux
    port map (
            O => \N__46910\,
            I => \N__46668\
        );

    \I__11288\ : ClkMux
    port map (
            O => \N__46909\,
            I => \N__46668\
        );

    \I__11287\ : ClkMux
    port map (
            O => \N__46908\,
            I => \N__46668\
        );

    \I__11286\ : ClkMux
    port map (
            O => \N__46907\,
            I => \N__46668\
        );

    \I__11285\ : ClkMux
    port map (
            O => \N__46906\,
            I => \N__46668\
        );

    \I__11284\ : ClkMux
    port map (
            O => \N__46905\,
            I => \N__46668\
        );

    \I__11283\ : ClkMux
    port map (
            O => \N__46904\,
            I => \N__46668\
        );

    \I__11282\ : ClkMux
    port map (
            O => \N__46903\,
            I => \N__46668\
        );

    \I__11281\ : ClkMux
    port map (
            O => \N__46902\,
            I => \N__46668\
        );

    \I__11280\ : ClkMux
    port map (
            O => \N__46901\,
            I => \N__46668\
        );

    \I__11279\ : ClkMux
    port map (
            O => \N__46900\,
            I => \N__46668\
        );

    \I__11278\ : ClkMux
    port map (
            O => \N__46899\,
            I => \N__46668\
        );

    \I__11277\ : ClkMux
    port map (
            O => \N__46898\,
            I => \N__46668\
        );

    \I__11276\ : ClkMux
    port map (
            O => \N__46897\,
            I => \N__46668\
        );

    \I__11275\ : ClkMux
    port map (
            O => \N__46896\,
            I => \N__46668\
        );

    \I__11274\ : ClkMux
    port map (
            O => \N__46895\,
            I => \N__46668\
        );

    \I__11273\ : ClkMux
    port map (
            O => \N__46894\,
            I => \N__46668\
        );

    \I__11272\ : ClkMux
    port map (
            O => \N__46893\,
            I => \N__46668\
        );

    \I__11271\ : ClkMux
    port map (
            O => \N__46892\,
            I => \N__46668\
        );

    \I__11270\ : ClkMux
    port map (
            O => \N__46891\,
            I => \N__46668\
        );

    \I__11269\ : ClkMux
    port map (
            O => \N__46890\,
            I => \N__46668\
        );

    \I__11268\ : ClkMux
    port map (
            O => \N__46889\,
            I => \N__46668\
        );

    \I__11267\ : ClkMux
    port map (
            O => \N__46888\,
            I => \N__46668\
        );

    \I__11266\ : ClkMux
    port map (
            O => \N__46887\,
            I => \N__46668\
        );

    \I__11265\ : ClkMux
    port map (
            O => \N__46886\,
            I => \N__46668\
        );

    \I__11264\ : ClkMux
    port map (
            O => \N__46885\,
            I => \N__46668\
        );

    \I__11263\ : ClkMux
    port map (
            O => \N__46884\,
            I => \N__46668\
        );

    \I__11262\ : ClkMux
    port map (
            O => \N__46883\,
            I => \N__46668\
        );

    \I__11261\ : ClkMux
    port map (
            O => \N__46882\,
            I => \N__46668\
        );

    \I__11260\ : ClkMux
    port map (
            O => \N__46881\,
            I => \N__46668\
        );

    \I__11259\ : ClkMux
    port map (
            O => \N__46880\,
            I => \N__46668\
        );

    \I__11258\ : ClkMux
    port map (
            O => \N__46879\,
            I => \N__46668\
        );

    \I__11257\ : ClkMux
    port map (
            O => \N__46878\,
            I => \N__46668\
        );

    \I__11256\ : ClkMux
    port map (
            O => \N__46877\,
            I => \N__46668\
        );

    \I__11255\ : ClkMux
    port map (
            O => \N__46876\,
            I => \N__46668\
        );

    \I__11254\ : ClkMux
    port map (
            O => \N__46875\,
            I => \N__46668\
        );

    \I__11253\ : ClkMux
    port map (
            O => \N__46874\,
            I => \N__46668\
        );

    \I__11252\ : ClkMux
    port map (
            O => \N__46873\,
            I => \N__46668\
        );

    \I__11251\ : ClkMux
    port map (
            O => \N__46872\,
            I => \N__46668\
        );

    \I__11250\ : ClkMux
    port map (
            O => \N__46871\,
            I => \N__46668\
        );

    \I__11249\ : ClkMux
    port map (
            O => \N__46870\,
            I => \N__46668\
        );

    \I__11248\ : ClkMux
    port map (
            O => \N__46869\,
            I => \N__46668\
        );

    \I__11247\ : ClkMux
    port map (
            O => \N__46868\,
            I => \N__46668\
        );

    \I__11246\ : ClkMux
    port map (
            O => \N__46867\,
            I => \N__46668\
        );

    \I__11245\ : ClkMux
    port map (
            O => \N__46866\,
            I => \N__46668\
        );

    \I__11244\ : ClkMux
    port map (
            O => \N__46865\,
            I => \N__46668\
        );

    \I__11243\ : ClkMux
    port map (
            O => \N__46864\,
            I => \N__46668\
        );

    \I__11242\ : ClkMux
    port map (
            O => \N__46863\,
            I => \N__46668\
        );

    \I__11241\ : ClkMux
    port map (
            O => \N__46862\,
            I => \N__46668\
        );

    \I__11240\ : ClkMux
    port map (
            O => \N__46861\,
            I => \N__46668\
        );

    \I__11239\ : ClkMux
    port map (
            O => \N__46860\,
            I => \N__46668\
        );

    \I__11238\ : ClkMux
    port map (
            O => \N__46859\,
            I => \N__46668\
        );

    \I__11237\ : ClkMux
    port map (
            O => \N__46858\,
            I => \N__46668\
        );

    \I__11236\ : ClkMux
    port map (
            O => \N__46857\,
            I => \N__46668\
        );

    \I__11235\ : ClkMux
    port map (
            O => \N__46856\,
            I => \N__46668\
        );

    \I__11234\ : ClkMux
    port map (
            O => \N__46855\,
            I => \N__46668\
        );

    \I__11233\ : ClkMux
    port map (
            O => \N__46854\,
            I => \N__46668\
        );

    \I__11232\ : ClkMux
    port map (
            O => \N__46853\,
            I => \N__46668\
        );

    \I__11231\ : ClkMux
    port map (
            O => \N__46852\,
            I => \N__46668\
        );

    \I__11230\ : ClkMux
    port map (
            O => \N__46851\,
            I => \N__46668\
        );

    \I__11229\ : ClkMux
    port map (
            O => \N__46850\,
            I => \N__46668\
        );

    \I__11228\ : ClkMux
    port map (
            O => \N__46849\,
            I => \N__46668\
        );

    \I__11227\ : ClkMux
    port map (
            O => \N__46848\,
            I => \N__46668\
        );

    \I__11226\ : ClkMux
    port map (
            O => \N__46847\,
            I => \N__46668\
        );

    \I__11225\ : ClkMux
    port map (
            O => \N__46846\,
            I => \N__46668\
        );

    \I__11224\ : ClkMux
    port map (
            O => \N__46845\,
            I => \N__46668\
        );

    \I__11223\ : ClkMux
    port map (
            O => \N__46844\,
            I => \N__46668\
        );

    \I__11222\ : ClkMux
    port map (
            O => \N__46843\,
            I => \N__46668\
        );

    \I__11221\ : ClkMux
    port map (
            O => \N__46842\,
            I => \N__46668\
        );

    \I__11220\ : ClkMux
    port map (
            O => \N__46841\,
            I => \N__46668\
        );

    \I__11219\ : ClkMux
    port map (
            O => \N__46840\,
            I => \N__46668\
        );

    \I__11218\ : ClkMux
    port map (
            O => \N__46839\,
            I => \N__46668\
        );

    \I__11217\ : GlobalMux
    port map (
            O => \N__46668\,
            I => \N__46665\
        );

    \I__11216\ : gio2CtrlBuf
    port map (
            O => \N__46665\,
            I => \CLK_c\
        );

    \I__11215\ : InMux
    port map (
            O => \N__46662\,
            I => \N__46659\
        );

    \I__11214\ : LocalMux
    port map (
            O => \N__46659\,
            I => pin_in_22
        );

    \I__11213\ : InMux
    port map (
            O => \N__46656\,
            I => \N__46653\
        );

    \I__11212\ : LocalMux
    port map (
            O => \N__46653\,
            I => \N__46650\
        );

    \I__11211\ : Span12Mux_h
    port map (
            O => \N__46650\,
            I => \N__46647\
        );

    \I__11210\ : Odrv12
    port map (
            O => \N__46647\,
            I => n13352
        );

    \I__11209\ : InMux
    port map (
            O => \N__46644\,
            I => \N__46641\
        );

    \I__11208\ : LocalMux
    port map (
            O => \N__46641\,
            I => \N__46638\
        );

    \I__11207\ : Span12Mux_h
    port map (
            O => \N__46638\,
            I => \N__46635\
        );

    \I__11206\ : Odrv12
    port map (
            O => \N__46635\,
            I => pin_in_17
        );

    \I__11205\ : CascadeMux
    port map (
            O => \N__46632\,
            I => \N__46629\
        );

    \I__11204\ : InMux
    port map (
            O => \N__46629\,
            I => \N__46626\
        );

    \I__11203\ : LocalMux
    port map (
            O => \N__46626\,
            I => \N__46623\
        );

    \I__11202\ : Span4Mux_v
    port map (
            O => \N__46623\,
            I => \N__46620\
        );

    \I__11201\ : Sp12to4
    port map (
            O => \N__46620\,
            I => \N__46617\
        );

    \I__11200\ : Span12Mux_s6_h
    port map (
            O => \N__46617\,
            I => \N__46614\
        );

    \I__11199\ : Span12Mux_v
    port map (
            O => \N__46614\,
            I => \N__46611\
        );

    \I__11198\ : Span12Mux_v
    port map (
            O => \N__46611\,
            I => \N__46608\
        );

    \I__11197\ : Odrv12
    port map (
            O => \N__46608\,
            I => pin_in_16
        );

    \I__11196\ : InMux
    port map (
            O => \N__46605\,
            I => \N__46602\
        );

    \I__11195\ : LocalMux
    port map (
            O => \N__46602\,
            I => \N__46599\
        );

    \I__11194\ : Span12Mux_h
    port map (
            O => \N__46599\,
            I => \N__46596\
        );

    \I__11193\ : Odrv12
    port map (
            O => \N__46596\,
            I => n13610
        );

    \I__11192\ : InMux
    port map (
            O => \N__46593\,
            I => \N__46590\
        );

    \I__11191\ : LocalMux
    port map (
            O => \N__46590\,
            I => pin_in_19
        );

    \I__11190\ : CascadeMux
    port map (
            O => \N__46587\,
            I => \N__46584\
        );

    \I__11189\ : InMux
    port map (
            O => \N__46584\,
            I => \N__46581\
        );

    \I__11188\ : LocalMux
    port map (
            O => \N__46581\,
            I => \N__46578\
        );

    \I__11187\ : Span4Mux_h
    port map (
            O => \N__46578\,
            I => \N__46575\
        );

    \I__11186\ : Odrv4
    port map (
            O => \N__46575\,
            I => pin_in_18
        );

    \I__11185\ : InMux
    port map (
            O => \N__46572\,
            I => \N__46568\
        );

    \I__11184\ : InMux
    port map (
            O => \N__46571\,
            I => \N__46560\
        );

    \I__11183\ : LocalMux
    port map (
            O => \N__46568\,
            I => \N__46556\
        );

    \I__11182\ : InMux
    port map (
            O => \N__46567\,
            I => \N__46552\
        );

    \I__11181\ : InMux
    port map (
            O => \N__46566\,
            I => \N__46549\
        );

    \I__11180\ : InMux
    port map (
            O => \N__46565\,
            I => \N__46546\
        );

    \I__11179\ : InMux
    port map (
            O => \N__46564\,
            I => \N__46542\
        );

    \I__11178\ : InMux
    port map (
            O => \N__46563\,
            I => \N__46539\
        );

    \I__11177\ : LocalMux
    port map (
            O => \N__46560\,
            I => \N__46536\
        );

    \I__11176\ : InMux
    port map (
            O => \N__46559\,
            I => \N__46533\
        );

    \I__11175\ : Span4Mux_s2_v
    port map (
            O => \N__46556\,
            I => \N__46530\
        );

    \I__11174\ : InMux
    port map (
            O => \N__46555\,
            I => \N__46527\
        );

    \I__11173\ : LocalMux
    port map (
            O => \N__46552\,
            I => \N__46524\
        );

    \I__11172\ : LocalMux
    port map (
            O => \N__46549\,
            I => \N__46517\
        );

    \I__11171\ : LocalMux
    port map (
            O => \N__46546\,
            I => \N__46517\
        );

    \I__11170\ : InMux
    port map (
            O => \N__46545\,
            I => \N__46514\
        );

    \I__11169\ : LocalMux
    port map (
            O => \N__46542\,
            I => \N__46505\
        );

    \I__11168\ : LocalMux
    port map (
            O => \N__46539\,
            I => \N__46498\
        );

    \I__11167\ : Span4Mux_v
    port map (
            O => \N__46536\,
            I => \N__46498\
        );

    \I__11166\ : LocalMux
    port map (
            O => \N__46533\,
            I => \N__46498\
        );

    \I__11165\ : Sp12to4
    port map (
            O => \N__46530\,
            I => \N__46491\
        );

    \I__11164\ : LocalMux
    port map (
            O => \N__46527\,
            I => \N__46491\
        );

    \I__11163\ : Span12Mux_s3_v
    port map (
            O => \N__46524\,
            I => \N__46491\
        );

    \I__11162\ : InMux
    port map (
            O => \N__46523\,
            I => \N__46486\
        );

    \I__11161\ : InMux
    port map (
            O => \N__46522\,
            I => \N__46486\
        );

    \I__11160\ : Span12Mux_v
    port map (
            O => \N__46517\,
            I => \N__46481\
        );

    \I__11159\ : LocalMux
    port map (
            O => \N__46514\,
            I => \N__46481\
        );

    \I__11158\ : InMux
    port map (
            O => \N__46513\,
            I => \N__46478\
        );

    \I__11157\ : InMux
    port map (
            O => \N__46512\,
            I => \N__46473\
        );

    \I__11156\ : InMux
    port map (
            O => \N__46511\,
            I => \N__46473\
        );

    \I__11155\ : InMux
    port map (
            O => \N__46510\,
            I => \N__46470\
        );

    \I__11154\ : InMux
    port map (
            O => \N__46509\,
            I => \N__46467\
        );

    \I__11153\ : InMux
    port map (
            O => \N__46508\,
            I => \N__46464\
        );

    \I__11152\ : Span4Mux_v
    port map (
            O => \N__46505\,
            I => \N__46459\
        );

    \I__11151\ : Span4Mux_v
    port map (
            O => \N__46498\,
            I => \N__46459\
        );

    \I__11150\ : Span12Mux_v
    port map (
            O => \N__46491\,
            I => \N__46454\
        );

    \I__11149\ : LocalMux
    port map (
            O => \N__46486\,
            I => \N__46454\
        );

    \I__11148\ : Span12Mux_h
    port map (
            O => \N__46481\,
            I => \N__46451\
        );

    \I__11147\ : LocalMux
    port map (
            O => \N__46478\,
            I => \N__46448\
        );

    \I__11146\ : LocalMux
    port map (
            O => \N__46473\,
            I => \N__46445\
        );

    \I__11145\ : LocalMux
    port map (
            O => \N__46470\,
            I => current_pin_1
        );

    \I__11144\ : LocalMux
    port map (
            O => \N__46467\,
            I => current_pin_1
        );

    \I__11143\ : LocalMux
    port map (
            O => \N__46464\,
            I => current_pin_1
        );

    \I__11142\ : Odrv4
    port map (
            O => \N__46459\,
            I => current_pin_1
        );

    \I__11141\ : Odrv12
    port map (
            O => \N__46454\,
            I => current_pin_1
        );

    \I__11140\ : Odrv12
    port map (
            O => \N__46451\,
            I => current_pin_1
        );

    \I__11139\ : Odrv4
    port map (
            O => \N__46448\,
            I => current_pin_1
        );

    \I__11138\ : Odrv4
    port map (
            O => \N__46445\,
            I => current_pin_1
        );

    \I__11137\ : InMux
    port map (
            O => \N__46428\,
            I => \N__46425\
        );

    \I__11136\ : LocalMux
    port map (
            O => \N__46425\,
            I => \N__46422\
        );

    \I__11135\ : Odrv12
    port map (
            O => \N__46422\,
            I => n13607
        );

    \I__11134\ : CascadeMux
    port map (
            O => \N__46419\,
            I => \N__46416\
        );

    \I__11133\ : InMux
    port map (
            O => \N__46416\,
            I => \N__46413\
        );

    \I__11132\ : LocalMux
    port map (
            O => \N__46413\,
            I => \N__46402\
        );

    \I__11131\ : InMux
    port map (
            O => \N__46412\,
            I => \N__46397\
        );

    \I__11130\ : InMux
    port map (
            O => \N__46411\,
            I => \N__46397\
        );

    \I__11129\ : InMux
    port map (
            O => \N__46410\,
            I => \N__46393\
        );

    \I__11128\ : InMux
    port map (
            O => \N__46409\,
            I => \N__46387\
        );

    \I__11127\ : InMux
    port map (
            O => \N__46408\,
            I => \N__46387\
        );

    \I__11126\ : InMux
    port map (
            O => \N__46407\,
            I => \N__46378\
        );

    \I__11125\ : InMux
    port map (
            O => \N__46406\,
            I => \N__46378\
        );

    \I__11124\ : InMux
    port map (
            O => \N__46405\,
            I => \N__46375\
        );

    \I__11123\ : Span4Mux_s3_v
    port map (
            O => \N__46402\,
            I => \N__46372\
        );

    \I__11122\ : LocalMux
    port map (
            O => \N__46397\,
            I => \N__46369\
        );

    \I__11121\ : InMux
    port map (
            O => \N__46396\,
            I => \N__46366\
        );

    \I__11120\ : LocalMux
    port map (
            O => \N__46393\,
            I => \N__46363\
        );

    \I__11119\ : InMux
    port map (
            O => \N__46392\,
            I => \N__46360\
        );

    \I__11118\ : LocalMux
    port map (
            O => \N__46387\,
            I => \N__46357\
        );

    \I__11117\ : InMux
    port map (
            O => \N__46386\,
            I => \N__46352\
        );

    \I__11116\ : InMux
    port map (
            O => \N__46385\,
            I => \N__46352\
        );

    \I__11115\ : InMux
    port map (
            O => \N__46384\,
            I => \N__46349\
        );

    \I__11114\ : InMux
    port map (
            O => \N__46383\,
            I => \N__46346\
        );

    \I__11113\ : LocalMux
    port map (
            O => \N__46378\,
            I => \N__46338\
        );

    \I__11112\ : LocalMux
    port map (
            O => \N__46375\,
            I => \N__46338\
        );

    \I__11111\ : Sp12to4
    port map (
            O => \N__46372\,
            I => \N__46332\
        );

    \I__11110\ : Sp12to4
    port map (
            O => \N__46369\,
            I => \N__46329\
        );

    \I__11109\ : LocalMux
    port map (
            O => \N__46366\,
            I => \N__46324\
        );

    \I__11108\ : Span4Mux_v
    port map (
            O => \N__46363\,
            I => \N__46324\
        );

    \I__11107\ : LocalMux
    port map (
            O => \N__46360\,
            I => \N__46315\
        );

    \I__11106\ : Span4Mux_v
    port map (
            O => \N__46357\,
            I => \N__46315\
        );

    \I__11105\ : LocalMux
    port map (
            O => \N__46352\,
            I => \N__46308\
        );

    \I__11104\ : LocalMux
    port map (
            O => \N__46349\,
            I => \N__46308\
        );

    \I__11103\ : LocalMux
    port map (
            O => \N__46346\,
            I => \N__46308\
        );

    \I__11102\ : InMux
    port map (
            O => \N__46345\,
            I => \N__46303\
        );

    \I__11101\ : InMux
    port map (
            O => \N__46344\,
            I => \N__46303\
        );

    \I__11100\ : InMux
    port map (
            O => \N__46343\,
            I => \N__46300\
        );

    \I__11099\ : Span12Mux_v
    port map (
            O => \N__46338\,
            I => \N__46297\
        );

    \I__11098\ : InMux
    port map (
            O => \N__46337\,
            I => \N__46294\
        );

    \I__11097\ : InMux
    port map (
            O => \N__46336\,
            I => \N__46289\
        );

    \I__11096\ : InMux
    port map (
            O => \N__46335\,
            I => \N__46289\
        );

    \I__11095\ : Span12Mux_h
    port map (
            O => \N__46332\,
            I => \N__46284\
        );

    \I__11094\ : Span12Mux_s3_v
    port map (
            O => \N__46329\,
            I => \N__46284\
        );

    \I__11093\ : Sp12to4
    port map (
            O => \N__46324\,
            I => \N__46281\
        );

    \I__11092\ : InMux
    port map (
            O => \N__46323\,
            I => \N__46278\
        );

    \I__11091\ : InMux
    port map (
            O => \N__46322\,
            I => \N__46275\
        );

    \I__11090\ : InMux
    port map (
            O => \N__46321\,
            I => \N__46272\
        );

    \I__11089\ : InMux
    port map (
            O => \N__46320\,
            I => \N__46269\
        );

    \I__11088\ : Span4Mux_v
    port map (
            O => \N__46315\,
            I => \N__46264\
        );

    \I__11087\ : Span4Mux_v
    port map (
            O => \N__46308\,
            I => \N__46264\
        );

    \I__11086\ : LocalMux
    port map (
            O => \N__46303\,
            I => \N__46257\
        );

    \I__11085\ : LocalMux
    port map (
            O => \N__46300\,
            I => \N__46257\
        );

    \I__11084\ : Span12Mux_h
    port map (
            O => \N__46297\,
            I => \N__46257\
        );

    \I__11083\ : LocalMux
    port map (
            O => \N__46294\,
            I => \N__46248\
        );

    \I__11082\ : LocalMux
    port map (
            O => \N__46289\,
            I => \N__46248\
        );

    \I__11081\ : Span12Mux_v
    port map (
            O => \N__46284\,
            I => \N__46248\
        );

    \I__11080\ : Span12Mux_h
    port map (
            O => \N__46281\,
            I => \N__46248\
        );

    \I__11079\ : LocalMux
    port map (
            O => \N__46278\,
            I => current_pin_0
        );

    \I__11078\ : LocalMux
    port map (
            O => \N__46275\,
            I => current_pin_0
        );

    \I__11077\ : LocalMux
    port map (
            O => \N__46272\,
            I => current_pin_0
        );

    \I__11076\ : LocalMux
    port map (
            O => \N__46269\,
            I => current_pin_0
        );

    \I__11075\ : Odrv4
    port map (
            O => \N__46264\,
            I => current_pin_0
        );

    \I__11074\ : Odrv12
    port map (
            O => \N__46257\,
            I => current_pin_0
        );

    \I__11073\ : Odrv12
    port map (
            O => \N__46248\,
            I => current_pin_0
        );

    \I__11072\ : InMux
    port map (
            O => \N__46233\,
            I => \N__46230\
        );

    \I__11071\ : LocalMux
    port map (
            O => \N__46230\,
            I => pin_in_21
        );

    \I__11070\ : InMux
    port map (
            O => \N__46227\,
            I => \N__46224\
        );

    \I__11069\ : LocalMux
    port map (
            O => \N__46224\,
            I => \N__46221\
        );

    \I__11068\ : Span4Mux_h
    port map (
            O => \N__46221\,
            I => \N__46218\
        );

    \I__11067\ : Odrv4
    port map (
            O => \N__46218\,
            I => pin_in_20
        );

    \I__11066\ : InMux
    port map (
            O => \N__46215\,
            I => \N__46212\
        );

    \I__11065\ : LocalMux
    port map (
            O => \N__46212\,
            I => n19_adj_789
        );

    \I__11064\ : CascadeMux
    port map (
            O => \N__46209\,
            I => \n13375_cascade_\
        );

    \I__11063\ : InMux
    port map (
            O => \N__46206\,
            I => \N__46203\
        );

    \I__11062\ : LocalMux
    port map (
            O => \N__46203\,
            I => \N__46200\
        );

    \I__11061\ : Span4Mux_h
    port map (
            O => \N__46200\,
            I => \N__46197\
        );

    \I__11060\ : Odrv4
    port map (
            O => \N__46197\,
            I => n13637
        );

    \I__11059\ : InMux
    port map (
            O => \N__46194\,
            I => \N__46191\
        );

    \I__11058\ : LocalMux
    port map (
            O => \N__46191\,
            I => \N__46188\
        );

    \I__11057\ : Odrv4
    port map (
            O => \N__46188\,
            I => n8_adj_829
        );

    \I__11056\ : IoInMux
    port map (
            O => \N__46185\,
            I => \N__46182\
        );

    \I__11055\ : LocalMux
    port map (
            O => \N__46182\,
            I => \N__46179\
        );

    \I__11054\ : IoSpan4Mux
    port map (
            O => \N__46179\,
            I => \N__46176\
        );

    \I__11053\ : Span4Mux_s2_v
    port map (
            O => \N__46176\,
            I => \N__46173\
        );

    \I__11052\ : Sp12to4
    port map (
            O => \N__46173\,
            I => \N__46170\
        );

    \I__11051\ : Span12Mux_h
    port map (
            O => \N__46170\,
            I => \N__46167\
        );

    \I__11050\ : Span12Mux_v
    port map (
            O => \N__46167\,
            I => \N__46162\
        );

    \I__11049\ : InMux
    port map (
            O => \N__46166\,
            I => \N__46157\
        );

    \I__11048\ : InMux
    port map (
            O => \N__46165\,
            I => \N__46157\
        );

    \I__11047\ : Odrv12
    port map (
            O => \N__46162\,
            I => pin_out_12
        );

    \I__11046\ : LocalMux
    port map (
            O => \N__46157\,
            I => pin_out_12
        );

    \I__11045\ : CascadeMux
    port map (
            O => \N__46152\,
            I => \N__46148\
        );

    \I__11044\ : CascadeMux
    port map (
            O => \N__46151\,
            I => \N__46133\
        );

    \I__11043\ : InMux
    port map (
            O => \N__46148\,
            I => \N__46129\
        );

    \I__11042\ : InMux
    port map (
            O => \N__46147\,
            I => \N__46126\
        );

    \I__11041\ : InMux
    port map (
            O => \N__46146\,
            I => \N__46121\
        );

    \I__11040\ : InMux
    port map (
            O => \N__46145\,
            I => \N__46121\
        );

    \I__11039\ : InMux
    port map (
            O => \N__46144\,
            I => \N__46118\
        );

    \I__11038\ : InMux
    port map (
            O => \N__46143\,
            I => \N__46115\
        );

    \I__11037\ : InMux
    port map (
            O => \N__46142\,
            I => \N__46112\
        );

    \I__11036\ : InMux
    port map (
            O => \N__46141\,
            I => \N__46107\
        );

    \I__11035\ : InMux
    port map (
            O => \N__46140\,
            I => \N__46104\
        );

    \I__11034\ : InMux
    port map (
            O => \N__46139\,
            I => \N__46099\
        );

    \I__11033\ : InMux
    port map (
            O => \N__46138\,
            I => \N__46099\
        );

    \I__11032\ : InMux
    port map (
            O => \N__46137\,
            I => \N__46089\
        );

    \I__11031\ : InMux
    port map (
            O => \N__46136\,
            I => \N__46089\
        );

    \I__11030\ : InMux
    port map (
            O => \N__46133\,
            I => \N__46086\
        );

    \I__11029\ : InMux
    port map (
            O => \N__46132\,
            I => \N__46083\
        );

    \I__11028\ : LocalMux
    port map (
            O => \N__46129\,
            I => \N__46080\
        );

    \I__11027\ : LocalMux
    port map (
            O => \N__46126\,
            I => \N__46077\
        );

    \I__11026\ : LocalMux
    port map (
            O => \N__46121\,
            I => \N__46074\
        );

    \I__11025\ : LocalMux
    port map (
            O => \N__46118\,
            I => \N__46067\
        );

    \I__11024\ : LocalMux
    port map (
            O => \N__46115\,
            I => \N__46067\
        );

    \I__11023\ : LocalMux
    port map (
            O => \N__46112\,
            I => \N__46067\
        );

    \I__11022\ : InMux
    port map (
            O => \N__46111\,
            I => \N__46064\
        );

    \I__11021\ : InMux
    port map (
            O => \N__46110\,
            I => \N__46061\
        );

    \I__11020\ : LocalMux
    port map (
            O => \N__46107\,
            I => \N__46054\
        );

    \I__11019\ : LocalMux
    port map (
            O => \N__46104\,
            I => \N__46054\
        );

    \I__11018\ : LocalMux
    port map (
            O => \N__46099\,
            I => \N__46054\
        );

    \I__11017\ : InMux
    port map (
            O => \N__46098\,
            I => \N__46049\
        );

    \I__11016\ : InMux
    port map (
            O => \N__46097\,
            I => \N__46049\
        );

    \I__11015\ : InMux
    port map (
            O => \N__46096\,
            I => \N__46046\
        );

    \I__11014\ : InMux
    port map (
            O => \N__46095\,
            I => \N__46041\
        );

    \I__11013\ : InMux
    port map (
            O => \N__46094\,
            I => \N__46041\
        );

    \I__11012\ : LocalMux
    port map (
            O => \N__46089\,
            I => \N__46026\
        );

    \I__11011\ : LocalMux
    port map (
            O => \N__46086\,
            I => \N__46026\
        );

    \I__11010\ : LocalMux
    port map (
            O => \N__46083\,
            I => \N__46026\
        );

    \I__11009\ : Span4Mux_v
    port map (
            O => \N__46080\,
            I => \N__46026\
        );

    \I__11008\ : Span4Mux_h
    port map (
            O => \N__46077\,
            I => \N__46026\
        );

    \I__11007\ : Span4Mux_h
    port map (
            O => \N__46074\,
            I => \N__46026\
        );

    \I__11006\ : Span4Mux_v
    port map (
            O => \N__46067\,
            I => \N__46026\
        );

    \I__11005\ : LocalMux
    port map (
            O => \N__46064\,
            I => \N__46019\
        );

    \I__11004\ : LocalMux
    port map (
            O => \N__46061\,
            I => \N__46019\
        );

    \I__11003\ : Span4Mux_v
    port map (
            O => \N__46054\,
            I => \N__46019\
        );

    \I__11002\ : LocalMux
    port map (
            O => \N__46049\,
            I => n9675
        );

    \I__11001\ : LocalMux
    port map (
            O => \N__46046\,
            I => n9675
        );

    \I__11000\ : LocalMux
    port map (
            O => \N__46041\,
            I => n9675
        );

    \I__10999\ : Odrv4
    port map (
            O => \N__46026\,
            I => n9675
        );

    \I__10998\ : Odrv4
    port map (
            O => \N__46019\,
            I => n9675
        );

    \I__10997\ : InMux
    port map (
            O => \N__46008\,
            I => \N__46005\
        );

    \I__10996\ : LocalMux
    port map (
            O => \N__46005\,
            I => \N__46002\
        );

    \I__10995\ : Span4Mux_h
    port map (
            O => \N__46002\,
            I => \N__45999\
        );

    \I__10994\ : Odrv4
    port map (
            O => \N__45999\,
            I => n7_adj_830
        );

    \I__10993\ : InMux
    port map (
            O => \N__45996\,
            I => \N__45987\
        );

    \I__10992\ : InMux
    port map (
            O => \N__45995\,
            I => \N__45987\
        );

    \I__10991\ : InMux
    port map (
            O => \N__45994\,
            I => \N__45982\
        );

    \I__10990\ : InMux
    port map (
            O => \N__45993\,
            I => \N__45982\
        );

    \I__10989\ : CascadeMux
    port map (
            O => \N__45992\,
            I => \N__45975\
        );

    \I__10988\ : LocalMux
    port map (
            O => \N__45987\,
            I => \N__45965\
        );

    \I__10987\ : LocalMux
    port map (
            O => \N__45982\,
            I => \N__45965\
        );

    \I__10986\ : CEMux
    port map (
            O => \N__45981\,
            I => \N__45962\
        );

    \I__10985\ : InMux
    port map (
            O => \N__45980\,
            I => \N__45953\
        );

    \I__10984\ : InMux
    port map (
            O => \N__45979\,
            I => \N__45949\
        );

    \I__10983\ : InMux
    port map (
            O => \N__45978\,
            I => \N__45944\
        );

    \I__10982\ : InMux
    port map (
            O => \N__45975\,
            I => \N__45944\
        );

    \I__10981\ : InMux
    port map (
            O => \N__45974\,
            I => \N__45941\
        );

    \I__10980\ : InMux
    port map (
            O => \N__45973\,
            I => \N__45936\
        );

    \I__10979\ : InMux
    port map (
            O => \N__45972\,
            I => \N__45936\
        );

    \I__10978\ : InMux
    port map (
            O => \N__45971\,
            I => \N__45931\
        );

    \I__10977\ : InMux
    port map (
            O => \N__45970\,
            I => \N__45931\
        );

    \I__10976\ : Span4Mux_v
    port map (
            O => \N__45965\,
            I => \N__45926\
        );

    \I__10975\ : LocalMux
    port map (
            O => \N__45962\,
            I => \N__45926\
        );

    \I__10974\ : CEMux
    port map (
            O => \N__45961\,
            I => \N__45923\
        );

    \I__10973\ : InMux
    port map (
            O => \N__45960\,
            I => \N__45920\
        );

    \I__10972\ : InMux
    port map (
            O => \N__45959\,
            I => \N__45917\
        );

    \I__10971\ : InMux
    port map (
            O => \N__45958\,
            I => \N__45912\
        );

    \I__10970\ : InMux
    port map (
            O => \N__45957\,
            I => \N__45912\
        );

    \I__10969\ : InMux
    port map (
            O => \N__45956\,
            I => \N__45909\
        );

    \I__10968\ : LocalMux
    port map (
            O => \N__45953\,
            I => \N__45906\
        );

    \I__10967\ : InMux
    port map (
            O => \N__45952\,
            I => \N__45903\
        );

    \I__10966\ : LocalMux
    port map (
            O => \N__45949\,
            I => \N__45893\
        );

    \I__10965\ : LocalMux
    port map (
            O => \N__45944\,
            I => \N__45893\
        );

    \I__10964\ : LocalMux
    port map (
            O => \N__45941\,
            I => \N__45886\
        );

    \I__10963\ : LocalMux
    port map (
            O => \N__45936\,
            I => \N__45886\
        );

    \I__10962\ : LocalMux
    port map (
            O => \N__45931\,
            I => \N__45886\
        );

    \I__10961\ : Span4Mux_h
    port map (
            O => \N__45926\,
            I => \N__45883\
        );

    \I__10960\ : LocalMux
    port map (
            O => \N__45923\,
            I => \N__45880\
        );

    \I__10959\ : LocalMux
    port map (
            O => \N__45920\,
            I => \N__45867\
        );

    \I__10958\ : LocalMux
    port map (
            O => \N__45917\,
            I => \N__45867\
        );

    \I__10957\ : LocalMux
    port map (
            O => \N__45912\,
            I => \N__45867\
        );

    \I__10956\ : LocalMux
    port map (
            O => \N__45909\,
            I => \N__45867\
        );

    \I__10955\ : Sp12to4
    port map (
            O => \N__45906\,
            I => \N__45867\
        );

    \I__10954\ : LocalMux
    port map (
            O => \N__45903\,
            I => \N__45867\
        );

    \I__10953\ : InMux
    port map (
            O => \N__45902\,
            I => \N__45864\
        );

    \I__10952\ : InMux
    port map (
            O => \N__45901\,
            I => \N__45861\
        );

    \I__10951\ : InMux
    port map (
            O => \N__45900\,
            I => \N__45856\
        );

    \I__10950\ : InMux
    port map (
            O => \N__45899\,
            I => \N__45856\
        );

    \I__10949\ : InMux
    port map (
            O => \N__45898\,
            I => \N__45853\
        );

    \I__10948\ : Span4Mux_h
    port map (
            O => \N__45893\,
            I => \N__45848\
        );

    \I__10947\ : Span4Mux_v
    port map (
            O => \N__45886\,
            I => \N__45848\
        );

    \I__10946\ : Span4Mux_h
    port map (
            O => \N__45883\,
            I => \N__45845\
        );

    \I__10945\ : Span4Mux_v
    port map (
            O => \N__45880\,
            I => \N__45842\
        );

    \I__10944\ : Span12Mux_v
    port map (
            O => \N__45867\,
            I => \N__45839\
        );

    \I__10943\ : LocalMux
    port map (
            O => \N__45864\,
            I => \N__45836\
        );

    \I__10942\ : LocalMux
    port map (
            O => \N__45861\,
            I => n11789
        );

    \I__10941\ : LocalMux
    port map (
            O => \N__45856\,
            I => n11789
        );

    \I__10940\ : LocalMux
    port map (
            O => \N__45853\,
            I => n11789
        );

    \I__10939\ : Odrv4
    port map (
            O => \N__45848\,
            I => n11789
        );

    \I__10938\ : Odrv4
    port map (
            O => \N__45845\,
            I => n11789
        );

    \I__10937\ : Odrv4
    port map (
            O => \N__45842\,
            I => n11789
        );

    \I__10936\ : Odrv12
    port map (
            O => \N__45839\,
            I => n11789
        );

    \I__10935\ : Odrv4
    port map (
            O => \N__45836\,
            I => n11789
        );

    \I__10934\ : IoInMux
    port map (
            O => \N__45819\,
            I => \N__45816\
        );

    \I__10933\ : LocalMux
    port map (
            O => \N__45816\,
            I => \N__45813\
        );

    \I__10932\ : Span12Mux_s7_h
    port map (
            O => \N__45813\,
            I => \N__45808\
        );

    \I__10931\ : InMux
    port map (
            O => \N__45812\,
            I => \N__45803\
        );

    \I__10930\ : InMux
    port map (
            O => \N__45811\,
            I => \N__45803\
        );

    \I__10929\ : Odrv12
    port map (
            O => \N__45808\,
            I => pin_out_13
        );

    \I__10928\ : LocalMux
    port map (
            O => \N__45803\,
            I => pin_out_13
        );

    \I__10927\ : IoInMux
    port map (
            O => \N__45798\,
            I => \N__45795\
        );

    \I__10926\ : LocalMux
    port map (
            O => \N__45795\,
            I => \N__45792\
        );

    \I__10925\ : IoSpan4Mux
    port map (
            O => \N__45792\,
            I => \N__45789\
        );

    \I__10924\ : Sp12to4
    port map (
            O => \N__45789\,
            I => \N__45784\
        );

    \I__10923\ : InMux
    port map (
            O => \N__45788\,
            I => \N__45781\
        );

    \I__10922\ : InMux
    port map (
            O => \N__45787\,
            I => \N__45778\
        );

    \I__10921\ : Span12Mux_s9_h
    port map (
            O => \N__45784\,
            I => \N__45773\
        );

    \I__10920\ : LocalMux
    port map (
            O => \N__45781\,
            I => \N__45773\
        );

    \I__10919\ : LocalMux
    port map (
            O => \N__45778\,
            I => pin_out_15
        );

    \I__10918\ : Odrv12
    port map (
            O => \N__45773\,
            I => pin_out_15
        );

    \I__10917\ : IoInMux
    port map (
            O => \N__45768\,
            I => \N__45765\
        );

    \I__10916\ : LocalMux
    port map (
            O => \N__45765\,
            I => \N__45762\
        );

    \I__10915\ : IoSpan4Mux
    port map (
            O => \N__45762\,
            I => \N__45759\
        );

    \I__10914\ : Span4Mux_s0_h
    port map (
            O => \N__45759\,
            I => \N__45756\
        );

    \I__10913\ : Sp12to4
    port map (
            O => \N__45756\,
            I => \N__45753\
        );

    \I__10912\ : Span12Mux_h
    port map (
            O => \N__45753\,
            I => \N__45748\
        );

    \I__10911\ : InMux
    port map (
            O => \N__45752\,
            I => \N__45745\
        );

    \I__10910\ : InMux
    port map (
            O => \N__45751\,
            I => \N__45742\
        );

    \I__10909\ : Odrv12
    port map (
            O => \N__45748\,
            I => pin_out_14
        );

    \I__10908\ : LocalMux
    port map (
            O => \N__45745\,
            I => pin_out_14
        );

    \I__10907\ : LocalMux
    port map (
            O => \N__45742\,
            I => pin_out_14
        );

    \I__10906\ : InMux
    port map (
            O => \N__45735\,
            I => \N__45732\
        );

    \I__10905\ : LocalMux
    port map (
            O => \N__45732\,
            I => n13376
        );

    \I__10904\ : InMux
    port map (
            O => \N__45729\,
            I => \N__45726\
        );

    \I__10903\ : LocalMux
    port map (
            O => \N__45726\,
            I => n11956
        );

    \I__10902\ : IoInMux
    port map (
            O => \N__45723\,
            I => \N__45720\
        );

    \I__10901\ : LocalMux
    port map (
            O => \N__45720\,
            I => \N__45717\
        );

    \I__10900\ : IoSpan4Mux
    port map (
            O => \N__45717\,
            I => \N__45714\
        );

    \I__10899\ : Span4Mux_s1_h
    port map (
            O => \N__45714\,
            I => \N__45711\
        );

    \I__10898\ : Span4Mux_h
    port map (
            O => \N__45711\,
            I => \N__45708\
        );

    \I__10897\ : Span4Mux_h
    port map (
            O => \N__45708\,
            I => \N__45704\
        );

    \I__10896\ : InMux
    port map (
            O => \N__45707\,
            I => \N__45701\
        );

    \I__10895\ : Odrv4
    port map (
            O => \N__45704\,
            I => pin_oe_13
        );

    \I__10894\ : LocalMux
    port map (
            O => \N__45701\,
            I => pin_oe_13
        );

    \I__10893\ : CascadeMux
    port map (
            O => \N__45696\,
            I => \N__45692\
        );

    \I__10892\ : CascadeMux
    port map (
            O => \N__45695\,
            I => \N__45689\
        );

    \I__10891\ : InMux
    port map (
            O => \N__45692\,
            I => \N__45686\
        );

    \I__10890\ : InMux
    port map (
            O => \N__45689\,
            I => \N__45683\
        );

    \I__10889\ : LocalMux
    port map (
            O => \N__45686\,
            I => \N__45678\
        );

    \I__10888\ : LocalMux
    port map (
            O => \N__45683\,
            I => \N__45675\
        );

    \I__10887\ : CascadeMux
    port map (
            O => \N__45682\,
            I => \N__45672\
        );

    \I__10886\ : CascadeMux
    port map (
            O => \N__45681\,
            I => \N__45665\
        );

    \I__10885\ : Span4Mux_v
    port map (
            O => \N__45678\,
            I => \N__45661\
        );

    \I__10884\ : Span4Mux_v
    port map (
            O => \N__45675\,
            I => \N__45658\
        );

    \I__10883\ : InMux
    port map (
            O => \N__45672\,
            I => \N__45655\
        );

    \I__10882\ : InMux
    port map (
            O => \N__45671\,
            I => \N__45646\
        );

    \I__10881\ : CascadeMux
    port map (
            O => \N__45670\,
            I => \N__45638\
        );

    \I__10880\ : CascadeMux
    port map (
            O => \N__45669\,
            I => \N__45635\
        );

    \I__10879\ : InMux
    port map (
            O => \N__45668\,
            I => \N__45631\
        );

    \I__10878\ : InMux
    port map (
            O => \N__45665\,
            I => \N__45628\
        );

    \I__10877\ : CascadeMux
    port map (
            O => \N__45664\,
            I => \N__45624\
        );

    \I__10876\ : Span4Mux_h
    port map (
            O => \N__45661\,
            I => \N__45619\
        );

    \I__10875\ : Span4Mux_h
    port map (
            O => \N__45658\,
            I => \N__45619\
        );

    \I__10874\ : LocalMux
    port map (
            O => \N__45655\,
            I => \N__45616\
        );

    \I__10873\ : CascadeMux
    port map (
            O => \N__45654\,
            I => \N__45612\
        );

    \I__10872\ : CascadeMux
    port map (
            O => \N__45653\,
            I => \N__45608\
        );

    \I__10871\ : CascadeMux
    port map (
            O => \N__45652\,
            I => \N__45605\
        );

    \I__10870\ : CascadeMux
    port map (
            O => \N__45651\,
            I => \N__45602\
        );

    \I__10869\ : CascadeMux
    port map (
            O => \N__45650\,
            I => \N__45599\
        );

    \I__10868\ : CascadeMux
    port map (
            O => \N__45649\,
            I => \N__45593\
        );

    \I__10867\ : LocalMux
    port map (
            O => \N__45646\,
            I => \N__45589\
        );

    \I__10866\ : InMux
    port map (
            O => \N__45645\,
            I => \N__45584\
        );

    \I__10865\ : InMux
    port map (
            O => \N__45644\,
            I => \N__45581\
        );

    \I__10864\ : CascadeMux
    port map (
            O => \N__45643\,
            I => \N__45578\
        );

    \I__10863\ : CascadeMux
    port map (
            O => \N__45642\,
            I => \N__45575\
        );

    \I__10862\ : CascadeMux
    port map (
            O => \N__45641\,
            I => \N__45571\
        );

    \I__10861\ : InMux
    port map (
            O => \N__45638\,
            I => \N__45564\
        );

    \I__10860\ : InMux
    port map (
            O => \N__45635\,
            I => \N__45561\
        );

    \I__10859\ : CascadeMux
    port map (
            O => \N__45634\,
            I => \N__45557\
        );

    \I__10858\ : LocalMux
    port map (
            O => \N__45631\,
            I => \N__45553\
        );

    \I__10857\ : LocalMux
    port map (
            O => \N__45628\,
            I => \N__45550\
        );

    \I__10856\ : InMux
    port map (
            O => \N__45627\,
            I => \N__45547\
        );

    \I__10855\ : InMux
    port map (
            O => \N__45624\,
            I => \N__45544\
        );

    \I__10854\ : Span4Mux_v
    port map (
            O => \N__45619\,
            I => \N__45539\
        );

    \I__10853\ : Span4Mux_v
    port map (
            O => \N__45616\,
            I => \N__45539\
        );

    \I__10852\ : CascadeMux
    port map (
            O => \N__45615\,
            I => \N__45535\
        );

    \I__10851\ : InMux
    port map (
            O => \N__45612\,
            I => \N__45531\
        );

    \I__10850\ : InMux
    port map (
            O => \N__45611\,
            I => \N__45526\
        );

    \I__10849\ : InMux
    port map (
            O => \N__45608\,
            I => \N__45526\
        );

    \I__10848\ : InMux
    port map (
            O => \N__45605\,
            I => \N__45523\
        );

    \I__10847\ : InMux
    port map (
            O => \N__45602\,
            I => \N__45520\
        );

    \I__10846\ : InMux
    port map (
            O => \N__45599\,
            I => \N__45515\
        );

    \I__10845\ : InMux
    port map (
            O => \N__45598\,
            I => \N__45515\
        );

    \I__10844\ : CascadeMux
    port map (
            O => \N__45597\,
            I => \N__45512\
        );

    \I__10843\ : CascadeMux
    port map (
            O => \N__45596\,
            I => \N__45509\
        );

    \I__10842\ : InMux
    port map (
            O => \N__45593\,
            I => \N__45502\
        );

    \I__10841\ : InMux
    port map (
            O => \N__45592\,
            I => \N__45502\
        );

    \I__10840\ : Span4Mux_h
    port map (
            O => \N__45589\,
            I => \N__45499\
        );

    \I__10839\ : CascadeMux
    port map (
            O => \N__45588\,
            I => \N__45494\
        );

    \I__10838\ : CascadeMux
    port map (
            O => \N__45587\,
            I => \N__45489\
        );

    \I__10837\ : LocalMux
    port map (
            O => \N__45584\,
            I => \N__45482\
        );

    \I__10836\ : LocalMux
    port map (
            O => \N__45581\,
            I => \N__45482\
        );

    \I__10835\ : InMux
    port map (
            O => \N__45578\,
            I => \N__45478\
        );

    \I__10834\ : InMux
    port map (
            O => \N__45575\,
            I => \N__45475\
        );

    \I__10833\ : InMux
    port map (
            O => \N__45574\,
            I => \N__45472\
        );

    \I__10832\ : InMux
    port map (
            O => \N__45571\,
            I => \N__45467\
        );

    \I__10831\ : InMux
    port map (
            O => \N__45570\,
            I => \N__45467\
        );

    \I__10830\ : CascadeMux
    port map (
            O => \N__45569\,
            I => \N__45463\
        );

    \I__10829\ : CascadeMux
    port map (
            O => \N__45568\,
            I => \N__45458\
        );

    \I__10828\ : CascadeMux
    port map (
            O => \N__45567\,
            I => \N__45455\
        );

    \I__10827\ : LocalMux
    port map (
            O => \N__45564\,
            I => \N__45449\
        );

    \I__10826\ : LocalMux
    port map (
            O => \N__45561\,
            I => \N__45446\
        );

    \I__10825\ : InMux
    port map (
            O => \N__45560\,
            I => \N__45443\
        );

    \I__10824\ : InMux
    port map (
            O => \N__45557\,
            I => \N__45438\
        );

    \I__10823\ : InMux
    port map (
            O => \N__45556\,
            I => \N__45438\
        );

    \I__10822\ : Span4Mux_h
    port map (
            O => \N__45553\,
            I => \N__45431\
        );

    \I__10821\ : Span4Mux_v
    port map (
            O => \N__45550\,
            I => \N__45431\
        );

    \I__10820\ : LocalMux
    port map (
            O => \N__45547\,
            I => \N__45431\
        );

    \I__10819\ : LocalMux
    port map (
            O => \N__45544\,
            I => \N__45426\
        );

    \I__10818\ : Span4Mux_h
    port map (
            O => \N__45539\,
            I => \N__45426\
        );

    \I__10817\ : InMux
    port map (
            O => \N__45538\,
            I => \N__45419\
        );

    \I__10816\ : InMux
    port map (
            O => \N__45535\,
            I => \N__45419\
        );

    \I__10815\ : InMux
    port map (
            O => \N__45534\,
            I => \N__45419\
        );

    \I__10814\ : LocalMux
    port map (
            O => \N__45531\,
            I => \N__45408\
        );

    \I__10813\ : LocalMux
    port map (
            O => \N__45526\,
            I => \N__45408\
        );

    \I__10812\ : LocalMux
    port map (
            O => \N__45523\,
            I => \N__45408\
        );

    \I__10811\ : LocalMux
    port map (
            O => \N__45520\,
            I => \N__45408\
        );

    \I__10810\ : LocalMux
    port map (
            O => \N__45515\,
            I => \N__45408\
        );

    \I__10809\ : InMux
    port map (
            O => \N__45512\,
            I => \N__45403\
        );

    \I__10808\ : InMux
    port map (
            O => \N__45509\,
            I => \N__45403\
        );

    \I__10807\ : InMux
    port map (
            O => \N__45508\,
            I => \N__45398\
        );

    \I__10806\ : InMux
    port map (
            O => \N__45507\,
            I => \N__45398\
        );

    \I__10805\ : LocalMux
    port map (
            O => \N__45502\,
            I => \N__45393\
        );

    \I__10804\ : Span4Mux_h
    port map (
            O => \N__45499\,
            I => \N__45393\
        );

    \I__10803\ : InMux
    port map (
            O => \N__45498\,
            I => \N__45388\
        );

    \I__10802\ : InMux
    port map (
            O => \N__45497\,
            I => \N__45388\
        );

    \I__10801\ : InMux
    port map (
            O => \N__45494\,
            I => \N__45383\
        );

    \I__10800\ : InMux
    port map (
            O => \N__45493\,
            I => \N__45383\
        );

    \I__10799\ : InMux
    port map (
            O => \N__45492\,
            I => \N__45380\
        );

    \I__10798\ : InMux
    port map (
            O => \N__45489\,
            I => \N__45377\
        );

    \I__10797\ : InMux
    port map (
            O => \N__45488\,
            I => \N__45372\
        );

    \I__10796\ : InMux
    port map (
            O => \N__45487\,
            I => \N__45372\
        );

    \I__10795\ : Span12Mux_v
    port map (
            O => \N__45482\,
            I => \N__45369\
        );

    \I__10794\ : InMux
    port map (
            O => \N__45481\,
            I => \N__45366\
        );

    \I__10793\ : LocalMux
    port map (
            O => \N__45478\,
            I => \N__45361\
        );

    \I__10792\ : LocalMux
    port map (
            O => \N__45475\,
            I => \N__45361\
        );

    \I__10791\ : LocalMux
    port map (
            O => \N__45472\,
            I => \N__45356\
        );

    \I__10790\ : LocalMux
    port map (
            O => \N__45467\,
            I => \N__45356\
        );

    \I__10789\ : InMux
    port map (
            O => \N__45466\,
            I => \N__45351\
        );

    \I__10788\ : InMux
    port map (
            O => \N__45463\,
            I => \N__45351\
        );

    \I__10787\ : InMux
    port map (
            O => \N__45462\,
            I => \N__45348\
        );

    \I__10786\ : InMux
    port map (
            O => \N__45461\,
            I => \N__45345\
        );

    \I__10785\ : InMux
    port map (
            O => \N__45458\,
            I => \N__45338\
        );

    \I__10784\ : InMux
    port map (
            O => \N__45455\,
            I => \N__45338\
        );

    \I__10783\ : InMux
    port map (
            O => \N__45454\,
            I => \N__45338\
        );

    \I__10782\ : InMux
    port map (
            O => \N__45453\,
            I => \N__45333\
        );

    \I__10781\ : InMux
    port map (
            O => \N__45452\,
            I => \N__45333\
        );

    \I__10780\ : Span4Mux_v
    port map (
            O => \N__45449\,
            I => \N__45316\
        );

    \I__10779\ : Span4Mux_v
    port map (
            O => \N__45446\,
            I => \N__45316\
        );

    \I__10778\ : LocalMux
    port map (
            O => \N__45443\,
            I => \N__45316\
        );

    \I__10777\ : LocalMux
    port map (
            O => \N__45438\,
            I => \N__45316\
        );

    \I__10776\ : Span4Mux_v
    port map (
            O => \N__45431\,
            I => \N__45316\
        );

    \I__10775\ : Span4Mux_h
    port map (
            O => \N__45426\,
            I => \N__45316\
        );

    \I__10774\ : LocalMux
    port map (
            O => \N__45419\,
            I => \N__45316\
        );

    \I__10773\ : Span4Mux_v
    port map (
            O => \N__45408\,
            I => \N__45316\
        );

    \I__10772\ : LocalMux
    port map (
            O => \N__45403\,
            I => \N__45305\
        );

    \I__10771\ : LocalMux
    port map (
            O => \N__45398\,
            I => \N__45305\
        );

    \I__10770\ : Span4Mux_h
    port map (
            O => \N__45393\,
            I => \N__45305\
        );

    \I__10769\ : LocalMux
    port map (
            O => \N__45388\,
            I => \N__45305\
        );

    \I__10768\ : LocalMux
    port map (
            O => \N__45383\,
            I => \N__45305\
        );

    \I__10767\ : LocalMux
    port map (
            O => \N__45380\,
            I => \N__45302\
        );

    \I__10766\ : LocalMux
    port map (
            O => \N__45377\,
            I => \N__45295\
        );

    \I__10765\ : LocalMux
    port map (
            O => \N__45372\,
            I => \N__45295\
        );

    \I__10764\ : Span12Mux_h
    port map (
            O => \N__45369\,
            I => \N__45295\
        );

    \I__10763\ : LocalMux
    port map (
            O => \N__45366\,
            I => current_pin_2
        );

    \I__10762\ : Odrv4
    port map (
            O => \N__45361\,
            I => current_pin_2
        );

    \I__10761\ : Odrv4
    port map (
            O => \N__45356\,
            I => current_pin_2
        );

    \I__10760\ : LocalMux
    port map (
            O => \N__45351\,
            I => current_pin_2
        );

    \I__10759\ : LocalMux
    port map (
            O => \N__45348\,
            I => current_pin_2
        );

    \I__10758\ : LocalMux
    port map (
            O => \N__45345\,
            I => current_pin_2
        );

    \I__10757\ : LocalMux
    port map (
            O => \N__45338\,
            I => current_pin_2
        );

    \I__10756\ : LocalMux
    port map (
            O => \N__45333\,
            I => current_pin_2
        );

    \I__10755\ : Odrv4
    port map (
            O => \N__45316\,
            I => current_pin_2
        );

    \I__10754\ : Odrv4
    port map (
            O => \N__45305\,
            I => current_pin_2
        );

    \I__10753\ : Odrv4
    port map (
            O => \N__45302\,
            I => current_pin_2
        );

    \I__10752\ : Odrv12
    port map (
            O => \N__45295\,
            I => current_pin_2
        );

    \I__10751\ : CascadeMux
    port map (
            O => \N__45270\,
            I => \N__45264\
        );

    \I__10750\ : InMux
    port map (
            O => \N__45269\,
            I => \N__45258\
        );

    \I__10749\ : InMux
    port map (
            O => \N__45268\,
            I => \N__45255\
        );

    \I__10748\ : InMux
    port map (
            O => \N__45267\,
            I => \N__45247\
        );

    \I__10747\ : InMux
    port map (
            O => \N__45264\,
            I => \N__45240\
        );

    \I__10746\ : InMux
    port map (
            O => \N__45263\,
            I => \N__45240\
        );

    \I__10745\ : InMux
    port map (
            O => \N__45262\,
            I => \N__45240\
        );

    \I__10744\ : InMux
    port map (
            O => \N__45261\,
            I => \N__45237\
        );

    \I__10743\ : LocalMux
    port map (
            O => \N__45258\,
            I => \N__45234\
        );

    \I__10742\ : LocalMux
    port map (
            O => \N__45255\,
            I => \N__45231\
        );

    \I__10741\ : InMux
    port map (
            O => \N__45254\,
            I => \N__45226\
        );

    \I__10740\ : InMux
    port map (
            O => \N__45253\,
            I => \N__45226\
        );

    \I__10739\ : InMux
    port map (
            O => \N__45252\,
            I => \N__45219\
        );

    \I__10738\ : InMux
    port map (
            O => \N__45251\,
            I => \N__45219\
        );

    \I__10737\ : InMux
    port map (
            O => \N__45250\,
            I => \N__45219\
        );

    \I__10736\ : LocalMux
    port map (
            O => \N__45247\,
            I => \N__45210\
        );

    \I__10735\ : LocalMux
    port map (
            O => \N__45240\,
            I => \N__45210\
        );

    \I__10734\ : LocalMux
    port map (
            O => \N__45237\,
            I => \N__45210\
        );

    \I__10733\ : Span4Mux_v
    port map (
            O => \N__45234\,
            I => \N__45210\
        );

    \I__10732\ : Odrv4
    port map (
            O => \N__45231\,
            I => current_pin_3
        );

    \I__10731\ : LocalMux
    port map (
            O => \N__45226\,
            I => current_pin_3
        );

    \I__10730\ : LocalMux
    port map (
            O => \N__45219\,
            I => current_pin_3
        );

    \I__10729\ : Odrv4
    port map (
            O => \N__45210\,
            I => current_pin_3
        );

    \I__10728\ : InMux
    port map (
            O => \N__45201\,
            I => \N__45198\
        );

    \I__10727\ : LocalMux
    port map (
            O => \N__45198\,
            I => \N__45195\
        );

    \I__10726\ : Span4Mux_h
    port map (
            O => \N__45195\,
            I => \N__45192\
        );

    \I__10725\ : Odrv4
    port map (
            O => \N__45192\,
            I => n13465
        );

    \I__10724\ : InMux
    port map (
            O => \N__45189\,
            I => \N__45186\
        );

    \I__10723\ : LocalMux
    port map (
            O => \N__45186\,
            I => \N__45183\
        );

    \I__10722\ : Sp12to4
    port map (
            O => \N__45183\,
            I => \N__45180\
        );

    \I__10721\ : Span12Mux_v
    port map (
            O => \N__45180\,
            I => \N__45177\
        );

    \I__10720\ : Odrv12
    port map (
            O => \N__45177\,
            I => pin_in_15
        );

    \I__10719\ : CascadeMux
    port map (
            O => \N__45174\,
            I => \N__45171\
        );

    \I__10718\ : InMux
    port map (
            O => \N__45171\,
            I => \N__45168\
        );

    \I__10717\ : LocalMux
    port map (
            O => \N__45168\,
            I => \N__45165\
        );

    \I__10716\ : Span4Mux_v
    port map (
            O => \N__45165\,
            I => \N__45162\
        );

    \I__10715\ : Sp12to4
    port map (
            O => \N__45162\,
            I => \N__45159\
        );

    \I__10714\ : Span12Mux_h
    port map (
            O => \N__45159\,
            I => \N__45156\
        );

    \I__10713\ : Span12Mux_v
    port map (
            O => \N__45156\,
            I => \N__45153\
        );

    \I__10712\ : Odrv12
    port map (
            O => \N__45153\,
            I => pin_in_14
        );

    \I__10711\ : InMux
    port map (
            O => \N__45150\,
            I => \N__45147\
        );

    \I__10710\ : LocalMux
    port map (
            O => \N__45147\,
            I => \N__45144\
        );

    \I__10709\ : Span12Mux_h
    port map (
            O => \N__45144\,
            I => \N__45141\
        );

    \I__10708\ : Odrv12
    port map (
            O => \N__45141\,
            I => pin_in_13
        );

    \I__10707\ : CascadeMux
    port map (
            O => \N__45138\,
            I => \n13643_cascade_\
        );

    \I__10706\ : InMux
    port map (
            O => \N__45135\,
            I => \N__45132\
        );

    \I__10705\ : LocalMux
    port map (
            O => \N__45132\,
            I => \N__45129\
        );

    \I__10704\ : Span4Mux_v
    port map (
            O => \N__45129\,
            I => \N__45126\
        );

    \I__10703\ : Sp12to4
    port map (
            O => \N__45126\,
            I => \N__45123\
        );

    \I__10702\ : Span12Mux_v
    port map (
            O => \N__45123\,
            I => \N__45120\
        );

    \I__10701\ : Odrv12
    port map (
            O => \N__45120\,
            I => pin_in_12
        );

    \I__10700\ : InMux
    port map (
            O => \N__45117\,
            I => \N__45114\
        );

    \I__10699\ : LocalMux
    port map (
            O => \N__45114\,
            I => \N__45111\
        );

    \I__10698\ : Odrv12
    port map (
            O => \N__45111\,
            I => n13646
        );

    \I__10697\ : InMux
    port map (
            O => \N__45108\,
            I => \N__45102\
        );

    \I__10696\ : InMux
    port map (
            O => \N__45107\,
            I => \N__45095\
        );

    \I__10695\ : InMux
    port map (
            O => \N__45106\,
            I => \N__45092\
        );

    \I__10694\ : InMux
    port map (
            O => \N__45105\,
            I => \N__45086\
        );

    \I__10693\ : LocalMux
    port map (
            O => \N__45102\,
            I => \N__45083\
        );

    \I__10692\ : InMux
    port map (
            O => \N__45101\,
            I => \N__45080\
        );

    \I__10691\ : InMux
    port map (
            O => \N__45100\,
            I => \N__45077\
        );

    \I__10690\ : InMux
    port map (
            O => \N__45099\,
            I => \N__45072\
        );

    \I__10689\ : InMux
    port map (
            O => \N__45098\,
            I => \N__45072\
        );

    \I__10688\ : LocalMux
    port map (
            O => \N__45095\,
            I => \N__45069\
        );

    \I__10687\ : LocalMux
    port map (
            O => \N__45092\,
            I => \N__45066\
        );

    \I__10686\ : InMux
    port map (
            O => \N__45091\,
            I => \N__45063\
        );

    \I__10685\ : InMux
    port map (
            O => \N__45090\,
            I => \N__45059\
        );

    \I__10684\ : InMux
    port map (
            O => \N__45089\,
            I => \N__45056\
        );

    \I__10683\ : LocalMux
    port map (
            O => \N__45086\,
            I => \N__45053\
        );

    \I__10682\ : Span4Mux_h
    port map (
            O => \N__45083\,
            I => \N__45046\
        );

    \I__10681\ : LocalMux
    port map (
            O => \N__45080\,
            I => \N__45046\
        );

    \I__10680\ : LocalMux
    port map (
            O => \N__45077\,
            I => \N__45046\
        );

    \I__10679\ : LocalMux
    port map (
            O => \N__45072\,
            I => \N__45037\
        );

    \I__10678\ : Span4Mux_h
    port map (
            O => \N__45069\,
            I => \N__45037\
        );

    \I__10677\ : Span4Mux_h
    port map (
            O => \N__45066\,
            I => \N__45037\
        );

    \I__10676\ : LocalMux
    port map (
            O => \N__45063\,
            I => \N__45037\
        );

    \I__10675\ : InMux
    port map (
            O => \N__45062\,
            I => \N__45034\
        );

    \I__10674\ : LocalMux
    port map (
            O => \N__45059\,
            I => n7_adj_797
        );

    \I__10673\ : LocalMux
    port map (
            O => \N__45056\,
            I => n7_adj_797
        );

    \I__10672\ : Odrv4
    port map (
            O => \N__45053\,
            I => n7_adj_797
        );

    \I__10671\ : Odrv4
    port map (
            O => \N__45046\,
            I => n7_adj_797
        );

    \I__10670\ : Odrv4
    port map (
            O => \N__45037\,
            I => n7_adj_797
        );

    \I__10669\ : LocalMux
    port map (
            O => \N__45034\,
            I => n7_adj_797
        );

    \I__10668\ : InMux
    port map (
            O => \N__45021\,
            I => \N__45014\
        );

    \I__10667\ : InMux
    port map (
            O => \N__45020\,
            I => \N__45014\
        );

    \I__10666\ : InMux
    port map (
            O => \N__45019\,
            I => \N__45011\
        );

    \I__10665\ : LocalMux
    port map (
            O => \N__45014\,
            I => \N__45007\
        );

    \I__10664\ : LocalMux
    port map (
            O => \N__45011\,
            I => \N__45003\
        );

    \I__10663\ : InMux
    port map (
            O => \N__45010\,
            I => \N__45000\
        );

    \I__10662\ : Span4Mux_v
    port map (
            O => \N__45007\,
            I => \N__44997\
        );

    \I__10661\ : InMux
    port map (
            O => \N__45006\,
            I => \N__44992\
        );

    \I__10660\ : Span4Mux_v
    port map (
            O => \N__45003\,
            I => \N__44985\
        );

    \I__10659\ : LocalMux
    port map (
            O => \N__45000\,
            I => \N__44985\
        );

    \I__10658\ : Span4Mux_h
    port map (
            O => \N__44997\,
            I => \N__44982\
        );

    \I__10657\ : CascadeMux
    port map (
            O => \N__44996\,
            I => \N__44978\
        );

    \I__10656\ : InMux
    port map (
            O => \N__44995\,
            I => \N__44975\
        );

    \I__10655\ : LocalMux
    port map (
            O => \N__44992\,
            I => \N__44972\
        );

    \I__10654\ : InMux
    port map (
            O => \N__44991\,
            I => \N__44969\
        );

    \I__10653\ : InMux
    port map (
            O => \N__44990\,
            I => \N__44965\
        );

    \I__10652\ : Span4Mux_h
    port map (
            O => \N__44985\,
            I => \N__44959\
        );

    \I__10651\ : Span4Mux_h
    port map (
            O => \N__44982\,
            I => \N__44959\
        );

    \I__10650\ : InMux
    port map (
            O => \N__44981\,
            I => \N__44956\
        );

    \I__10649\ : InMux
    port map (
            O => \N__44978\,
            I => \N__44953\
        );

    \I__10648\ : LocalMux
    port map (
            O => \N__44975\,
            I => \N__44946\
        );

    \I__10647\ : Span4Mux_h
    port map (
            O => \N__44972\,
            I => \N__44946\
        );

    \I__10646\ : LocalMux
    port map (
            O => \N__44969\,
            I => \N__44946\
        );

    \I__10645\ : InMux
    port map (
            O => \N__44968\,
            I => \N__44943\
        );

    \I__10644\ : LocalMux
    port map (
            O => \N__44965\,
            I => \N__44940\
        );

    \I__10643\ : InMux
    port map (
            O => \N__44964\,
            I => \N__44937\
        );

    \I__10642\ : Span4Mux_h
    port map (
            O => \N__44959\,
            I => \N__44934\
        );

    \I__10641\ : LocalMux
    port map (
            O => \N__44956\,
            I => \N__44929\
        );

    \I__10640\ : LocalMux
    port map (
            O => \N__44953\,
            I => \N__44929\
        );

    \I__10639\ : Span4Mux_v
    port map (
            O => \N__44946\,
            I => \N__44926\
        );

    \I__10638\ : LocalMux
    port map (
            O => \N__44943\,
            I => n6
        );

    \I__10637\ : Odrv4
    port map (
            O => \N__44940\,
            I => n6
        );

    \I__10636\ : LocalMux
    port map (
            O => \N__44937\,
            I => n6
        );

    \I__10635\ : Odrv4
    port map (
            O => \N__44934\,
            I => n6
        );

    \I__10634\ : Odrv12
    port map (
            O => \N__44929\,
            I => n6
        );

    \I__10633\ : Odrv4
    port map (
            O => \N__44926\,
            I => n6
        );

    \I__10632\ : CascadeMux
    port map (
            O => \N__44913\,
            I => \N__44904\
        );

    \I__10631\ : CascadeMux
    port map (
            O => \N__44912\,
            I => \N__44899\
        );

    \I__10630\ : InMux
    port map (
            O => \N__44911\,
            I => \N__44896\
        );

    \I__10629\ : CascadeMux
    port map (
            O => \N__44910\,
            I => \N__44893\
        );

    \I__10628\ : CascadeMux
    port map (
            O => \N__44909\,
            I => \N__44887\
        );

    \I__10627\ : InMux
    port map (
            O => \N__44908\,
            I => \N__44883\
        );

    \I__10626\ : InMux
    port map (
            O => \N__44907\,
            I => \N__44880\
        );

    \I__10625\ : InMux
    port map (
            O => \N__44904\,
            I => \N__44875\
        );

    \I__10624\ : InMux
    port map (
            O => \N__44903\,
            I => \N__44868\
        );

    \I__10623\ : InMux
    port map (
            O => \N__44902\,
            I => \N__44863\
        );

    \I__10622\ : InMux
    port map (
            O => \N__44899\,
            I => \N__44863\
        );

    \I__10621\ : LocalMux
    port map (
            O => \N__44896\,
            I => \N__44860\
        );

    \I__10620\ : InMux
    port map (
            O => \N__44893\,
            I => \N__44855\
        );

    \I__10619\ : InMux
    port map (
            O => \N__44892\,
            I => \N__44855\
        );

    \I__10618\ : InMux
    port map (
            O => \N__44891\,
            I => \N__44848\
        );

    \I__10617\ : InMux
    port map (
            O => \N__44890\,
            I => \N__44848\
        );

    \I__10616\ : InMux
    port map (
            O => \N__44887\,
            I => \N__44845\
        );

    \I__10615\ : InMux
    port map (
            O => \N__44886\,
            I => \N__44842\
        );

    \I__10614\ : LocalMux
    port map (
            O => \N__44883\,
            I => \N__44837\
        );

    \I__10613\ : LocalMux
    port map (
            O => \N__44880\,
            I => \N__44837\
        );

    \I__10612\ : InMux
    port map (
            O => \N__44879\,
            I => \N__44832\
        );

    \I__10611\ : InMux
    port map (
            O => \N__44878\,
            I => \N__44832\
        );

    \I__10610\ : LocalMux
    port map (
            O => \N__44875\,
            I => \N__44827\
        );

    \I__10609\ : InMux
    port map (
            O => \N__44874\,
            I => \N__44824\
        );

    \I__10608\ : InMux
    port map (
            O => \N__44873\,
            I => \N__44819\
        );

    \I__10607\ : InMux
    port map (
            O => \N__44872\,
            I => \N__44819\
        );

    \I__10606\ : InMux
    port map (
            O => \N__44871\,
            I => \N__44816\
        );

    \I__10605\ : LocalMux
    port map (
            O => \N__44868\,
            I => \N__44807\
        );

    \I__10604\ : LocalMux
    port map (
            O => \N__44863\,
            I => \N__44807\
        );

    \I__10603\ : Span4Mux_v
    port map (
            O => \N__44860\,
            I => \N__44807\
        );

    \I__10602\ : LocalMux
    port map (
            O => \N__44855\,
            I => \N__44807\
        );

    \I__10601\ : InMux
    port map (
            O => \N__44854\,
            I => \N__44802\
        );

    \I__10600\ : InMux
    port map (
            O => \N__44853\,
            I => \N__44802\
        );

    \I__10599\ : LocalMux
    port map (
            O => \N__44848\,
            I => \N__44799\
        );

    \I__10598\ : LocalMux
    port map (
            O => \N__44845\,
            I => \N__44790\
        );

    \I__10597\ : LocalMux
    port map (
            O => \N__44842\,
            I => \N__44790\
        );

    \I__10596\ : Span4Mux_v
    port map (
            O => \N__44837\,
            I => \N__44790\
        );

    \I__10595\ : LocalMux
    port map (
            O => \N__44832\,
            I => \N__44790\
        );

    \I__10594\ : InMux
    port map (
            O => \N__44831\,
            I => \N__44787\
        );

    \I__10593\ : InMux
    port map (
            O => \N__44830\,
            I => \N__44784\
        );

    \I__10592\ : Span4Mux_v
    port map (
            O => \N__44827\,
            I => \N__44777\
        );

    \I__10591\ : LocalMux
    port map (
            O => \N__44824\,
            I => \N__44777\
        );

    \I__10590\ : LocalMux
    port map (
            O => \N__44819\,
            I => \N__44777\
        );

    \I__10589\ : LocalMux
    port map (
            O => \N__44816\,
            I => \N__44770\
        );

    \I__10588\ : Span4Mux_v
    port map (
            O => \N__44807\,
            I => \N__44770\
        );

    \I__10587\ : LocalMux
    port map (
            O => \N__44802\,
            I => \N__44770\
        );

    \I__10586\ : Span4Mux_v
    port map (
            O => \N__44799\,
            I => \N__44765\
        );

    \I__10585\ : Span4Mux_v
    port map (
            O => \N__44790\,
            I => \N__44765\
        );

    \I__10584\ : LocalMux
    port map (
            O => \N__44787\,
            I => n6_adj_819
        );

    \I__10583\ : LocalMux
    port map (
            O => \N__44784\,
            I => n6_adj_819
        );

    \I__10582\ : Odrv4
    port map (
            O => \N__44777\,
            I => n6_adj_819
        );

    \I__10581\ : Odrv4
    port map (
            O => \N__44770\,
            I => n6_adj_819
        );

    \I__10580\ : Odrv4
    port map (
            O => \N__44765\,
            I => n6_adj_819
        );

    \I__10579\ : CascadeMux
    port map (
            O => \N__44754\,
            I => \n8_adj_834_cascade_\
        );

    \I__10578\ : IoInMux
    port map (
            O => \N__44751\,
            I => \N__44748\
        );

    \I__10577\ : LocalMux
    port map (
            O => \N__44748\,
            I => \N__44745\
        );

    \I__10576\ : Span4Mux_s1_v
    port map (
            O => \N__44745\,
            I => \N__44742\
        );

    \I__10575\ : Sp12to4
    port map (
            O => \N__44742\,
            I => \N__44739\
        );

    \I__10574\ : Span12Mux_h
    port map (
            O => \N__44739\,
            I => \N__44734\
        );

    \I__10573\ : InMux
    port map (
            O => \N__44738\,
            I => \N__44729\
        );

    \I__10572\ : InMux
    port map (
            O => \N__44737\,
            I => \N__44729\
        );

    \I__10571\ : Odrv12
    port map (
            O => \N__44734\,
            I => pin_out_17
        );

    \I__10570\ : LocalMux
    port map (
            O => \N__44729\,
            I => pin_out_17
        );

    \I__10569\ : InMux
    port map (
            O => \N__44724\,
            I => \N__44721\
        );

    \I__10568\ : LocalMux
    port map (
            O => \N__44721\,
            I => n13631
        );

    \I__10567\ : IoInMux
    port map (
            O => \N__44718\,
            I => \N__44715\
        );

    \I__10566\ : LocalMux
    port map (
            O => \N__44715\,
            I => \N__44712\
        );

    \I__10565\ : Span4Mux_s0_h
    port map (
            O => \N__44712\,
            I => \N__44709\
        );

    \I__10564\ : Sp12to4
    port map (
            O => \N__44709\,
            I => \N__44705\
        );

    \I__10563\ : CascadeMux
    port map (
            O => \N__44708\,
            I => \N__44702\
        );

    \I__10562\ : Span12Mux_v
    port map (
            O => \N__44705\,
            I => \N__44699\
        );

    \I__10561\ : InMux
    port map (
            O => \N__44702\,
            I => \N__44695\
        );

    \I__10560\ : Span12Mux_h
    port map (
            O => \N__44699\,
            I => \N__44692\
        );

    \I__10559\ : InMux
    port map (
            O => \N__44698\,
            I => \N__44689\
        );

    \I__10558\ : LocalMux
    port map (
            O => \N__44695\,
            I => \N__44686\
        );

    \I__10557\ : Odrv12
    port map (
            O => \N__44692\,
            I => pin_out_16
        );

    \I__10556\ : LocalMux
    port map (
            O => \N__44689\,
            I => pin_out_16
        );

    \I__10555\ : Odrv12
    port map (
            O => \N__44686\,
            I => pin_out_16
        );

    \I__10554\ : CascadeMux
    port map (
            O => \N__44679\,
            I => \n13634_cascade_\
        );

    \I__10553\ : InMux
    port map (
            O => \N__44676\,
            I => \N__44673\
        );

    \I__10552\ : LocalMux
    port map (
            O => \N__44673\,
            I => \N__44670\
        );

    \I__10551\ : Odrv4
    port map (
            O => \N__44670\,
            I => n13389
        );

    \I__10550\ : InMux
    port map (
            O => \N__44667\,
            I => \N__44664\
        );

    \I__10549\ : LocalMux
    port map (
            O => \N__44664\,
            I => n7_adj_838
        );

    \I__10548\ : InMux
    port map (
            O => \N__44661\,
            I => \N__44658\
        );

    \I__10547\ : LocalMux
    port map (
            O => \N__44658\,
            I => n7_adj_837
        );

    \I__10546\ : IoInMux
    port map (
            O => \N__44655\,
            I => \N__44652\
        );

    \I__10545\ : LocalMux
    port map (
            O => \N__44652\,
            I => \N__44649\
        );

    \I__10544\ : IoSpan4Mux
    port map (
            O => \N__44649\,
            I => \N__44646\
        );

    \I__10543\ : Span4Mux_s3_v
    port map (
            O => \N__44646\,
            I => \N__44643\
        );

    \I__10542\ : Span4Mux_v
    port map (
            O => \N__44643\,
            I => \N__44639\
        );

    \I__10541\ : CascadeMux
    port map (
            O => \N__44642\,
            I => \N__44636\
        );

    \I__10540\ : Span4Mux_v
    port map (
            O => \N__44639\,
            I => \N__44632\
        );

    \I__10539\ : InMux
    port map (
            O => \N__44636\,
            I => \N__44629\
        );

    \I__10538\ : InMux
    port map (
            O => \N__44635\,
            I => \N__44626\
        );

    \I__10537\ : Odrv4
    port map (
            O => \N__44632\,
            I => pin_out_21
        );

    \I__10536\ : LocalMux
    port map (
            O => \N__44629\,
            I => pin_out_21
        );

    \I__10535\ : LocalMux
    port map (
            O => \N__44626\,
            I => pin_out_21
        );

    \I__10534\ : IoInMux
    port map (
            O => \N__44619\,
            I => \N__44616\
        );

    \I__10533\ : LocalMux
    port map (
            O => \N__44616\,
            I => \N__44612\
        );

    \I__10532\ : CascadeMux
    port map (
            O => \N__44615\,
            I => \N__44609\
        );

    \I__10531\ : Span12Mux_s10_v
    port map (
            O => \N__44612\,
            I => \N__44605\
        );

    \I__10530\ : InMux
    port map (
            O => \N__44609\,
            I => \N__44600\
        );

    \I__10529\ : InMux
    port map (
            O => \N__44608\,
            I => \N__44600\
        );

    \I__10528\ : Odrv12
    port map (
            O => \N__44605\,
            I => pin_out_20
        );

    \I__10527\ : LocalMux
    port map (
            O => \N__44600\,
            I => pin_out_20
        );

    \I__10526\ : IoInMux
    port map (
            O => \N__44595\,
            I => \N__44592\
        );

    \I__10525\ : LocalMux
    port map (
            O => \N__44592\,
            I => \N__44589\
        );

    \I__10524\ : Span4Mux_s2_v
    port map (
            O => \N__44589\,
            I => \N__44586\
        );

    \I__10523\ : Span4Mux_h
    port map (
            O => \N__44586\,
            I => \N__44582\
        );

    \I__10522\ : InMux
    port map (
            O => \N__44585\,
            I => \N__44578\
        );

    \I__10521\ : Sp12to4
    port map (
            O => \N__44582\,
            I => \N__44575\
        );

    \I__10520\ : InMux
    port map (
            O => \N__44581\,
            I => \N__44572\
        );

    \I__10519\ : LocalMux
    port map (
            O => \N__44578\,
            I => \N__44569\
        );

    \I__10518\ : Odrv12
    port map (
            O => \N__44575\,
            I => pin_out_22
        );

    \I__10517\ : LocalMux
    port map (
            O => \N__44572\,
            I => pin_out_22
        );

    \I__10516\ : Odrv4
    port map (
            O => \N__44569\,
            I => pin_out_22
        );

    \I__10515\ : CascadeMux
    port map (
            O => \N__44562\,
            I => \n19_adj_790_cascade_\
        );

    \I__10514\ : InMux
    port map (
            O => \N__44559\,
            I => \N__44556\
        );

    \I__10513\ : LocalMux
    port map (
            O => \N__44556\,
            I => n13388
        );

    \I__10512\ : CascadeMux
    port map (
            O => \N__44553\,
            I => \n7_adj_833_cascade_\
        );

    \I__10511\ : InMux
    port map (
            O => \N__44550\,
            I => \N__44547\
        );

    \I__10510\ : LocalMux
    port map (
            O => \N__44547\,
            I => n8_adj_836
        );

    \I__10509\ : CascadeMux
    port map (
            O => \N__44544\,
            I => \N__44541\
        );

    \I__10508\ : InMux
    port map (
            O => \N__44541\,
            I => \N__44526\
        );

    \I__10507\ : InMux
    port map (
            O => \N__44540\,
            I => \N__44523\
        );

    \I__10506\ : InMux
    port map (
            O => \N__44539\,
            I => \N__44520\
        );

    \I__10505\ : InMux
    port map (
            O => \N__44538\,
            I => \N__44517\
        );

    \I__10504\ : InMux
    port map (
            O => \N__44537\,
            I => \N__44514\
        );

    \I__10503\ : InMux
    port map (
            O => \N__44536\,
            I => \N__44509\
        );

    \I__10502\ : InMux
    port map (
            O => \N__44535\,
            I => \N__44509\
        );

    \I__10501\ : InMux
    port map (
            O => \N__44534\,
            I => \N__44504\
        );

    \I__10500\ : InMux
    port map (
            O => \N__44533\,
            I => \N__44504\
        );

    \I__10499\ : InMux
    port map (
            O => \N__44532\,
            I => \N__44500\
        );

    \I__10498\ : InMux
    port map (
            O => \N__44531\,
            I => \N__44497\
        );

    \I__10497\ : InMux
    port map (
            O => \N__44530\,
            I => \N__44494\
        );

    \I__10496\ : InMux
    port map (
            O => \N__44529\,
            I => \N__44491\
        );

    \I__10495\ : LocalMux
    port map (
            O => \N__44526\,
            I => \N__44488\
        );

    \I__10494\ : LocalMux
    port map (
            O => \N__44523\,
            I => \N__44485\
        );

    \I__10493\ : LocalMux
    port map (
            O => \N__44520\,
            I => \N__44474\
        );

    \I__10492\ : LocalMux
    port map (
            O => \N__44517\,
            I => \N__44474\
        );

    \I__10491\ : LocalMux
    port map (
            O => \N__44514\,
            I => \N__44474\
        );

    \I__10490\ : LocalMux
    port map (
            O => \N__44509\,
            I => \N__44474\
        );

    \I__10489\ : LocalMux
    port map (
            O => \N__44504\,
            I => \N__44474\
        );

    \I__10488\ : InMux
    port map (
            O => \N__44503\,
            I => \N__44471\
        );

    \I__10487\ : LocalMux
    port map (
            O => \N__44500\,
            I => \N__44468\
        );

    \I__10486\ : LocalMux
    port map (
            O => \N__44497\,
            I => \N__44463\
        );

    \I__10485\ : LocalMux
    port map (
            O => \N__44494\,
            I => \N__44463\
        );

    \I__10484\ : LocalMux
    port map (
            O => \N__44491\,
            I => \N__44460\
        );

    \I__10483\ : Span4Mux_v
    port map (
            O => \N__44488\,
            I => \N__44453\
        );

    \I__10482\ : Span4Mux_h
    port map (
            O => \N__44485\,
            I => \N__44453\
        );

    \I__10481\ : Span4Mux_v
    port map (
            O => \N__44474\,
            I => \N__44453\
        );

    \I__10480\ : LocalMux
    port map (
            O => \N__44471\,
            I => n7_adj_811
        );

    \I__10479\ : Odrv4
    port map (
            O => \N__44468\,
            I => n7_adj_811
        );

    \I__10478\ : Odrv4
    port map (
            O => \N__44463\,
            I => n7_adj_811
        );

    \I__10477\ : Odrv4
    port map (
            O => \N__44460\,
            I => n7_adj_811
        );

    \I__10476\ : Odrv4
    port map (
            O => \N__44453\,
            I => n7_adj_811
        );

    \I__10475\ : CascadeMux
    port map (
            O => \N__44442\,
            I => \n7_adj_835_cascade_\
        );

    \I__10474\ : CascadeMux
    port map (
            O => \N__44439\,
            I => \N__44436\
        );

    \I__10473\ : InMux
    port map (
            O => \N__44436\,
            I => \N__44432\
        );

    \I__10472\ : InMux
    port map (
            O => \N__44435\,
            I => \N__44427\
        );

    \I__10471\ : LocalMux
    port map (
            O => \N__44432\,
            I => \N__44423\
        );

    \I__10470\ : InMux
    port map (
            O => \N__44431\,
            I => \N__44418\
        );

    \I__10469\ : InMux
    port map (
            O => \N__44430\,
            I => \N__44415\
        );

    \I__10468\ : LocalMux
    port map (
            O => \N__44427\,
            I => \N__44412\
        );

    \I__10467\ : InMux
    port map (
            O => \N__44426\,
            I => \N__44409\
        );

    \I__10466\ : Span4Mux_v
    port map (
            O => \N__44423\,
            I => \N__44406\
        );

    \I__10465\ : InMux
    port map (
            O => \N__44422\,
            I => \N__44402\
        );

    \I__10464\ : InMux
    port map (
            O => \N__44421\,
            I => \N__44399\
        );

    \I__10463\ : LocalMux
    port map (
            O => \N__44418\,
            I => \N__44396\
        );

    \I__10462\ : LocalMux
    port map (
            O => \N__44415\,
            I => \N__44393\
        );

    \I__10461\ : Span4Mux_v
    port map (
            O => \N__44412\,
            I => \N__44390\
        );

    \I__10460\ : LocalMux
    port map (
            O => \N__44409\,
            I => \N__44384\
        );

    \I__10459\ : Span4Mux_h
    port map (
            O => \N__44406\,
            I => \N__44381\
        );

    \I__10458\ : InMux
    port map (
            O => \N__44405\,
            I => \N__44378\
        );

    \I__10457\ : LocalMux
    port map (
            O => \N__44402\,
            I => \N__44375\
        );

    \I__10456\ : LocalMux
    port map (
            O => \N__44399\,
            I => \N__44372\
        );

    \I__10455\ : Span4Mux_h
    port map (
            O => \N__44396\,
            I => \N__44367\
        );

    \I__10454\ : Span4Mux_h
    port map (
            O => \N__44393\,
            I => \N__44367\
        );

    \I__10453\ : Span4Mux_h
    port map (
            O => \N__44390\,
            I => \N__44364\
        );

    \I__10452\ : InMux
    port map (
            O => \N__44389\,
            I => \N__44361\
        );

    \I__10451\ : InMux
    port map (
            O => \N__44388\,
            I => \N__44358\
        );

    \I__10450\ : InMux
    port map (
            O => \N__44387\,
            I => \N__44355\
        );

    \I__10449\ : Span4Mux_v
    port map (
            O => \N__44384\,
            I => \N__44350\
        );

    \I__10448\ : Span4Mux_h
    port map (
            O => \N__44381\,
            I => \N__44350\
        );

    \I__10447\ : LocalMux
    port map (
            O => \N__44378\,
            I => \N__44339\
        );

    \I__10446\ : Span4Mux_v
    port map (
            O => \N__44375\,
            I => \N__44339\
        );

    \I__10445\ : Span4Mux_v
    port map (
            O => \N__44372\,
            I => \N__44339\
        );

    \I__10444\ : Span4Mux_v
    port map (
            O => \N__44367\,
            I => \N__44339\
        );

    \I__10443\ : Span4Mux_h
    port map (
            O => \N__44364\,
            I => \N__44339\
        );

    \I__10442\ : LocalMux
    port map (
            O => \N__44361\,
            I => n6_adj_810
        );

    \I__10441\ : LocalMux
    port map (
            O => \N__44358\,
            I => n6_adj_810
        );

    \I__10440\ : LocalMux
    port map (
            O => \N__44355\,
            I => n6_adj_810
        );

    \I__10439\ : Odrv4
    port map (
            O => \N__44350\,
            I => n6_adj_810
        );

    \I__10438\ : Odrv4
    port map (
            O => \N__44339\,
            I => n6_adj_810
        );

    \I__10437\ : CascadeMux
    port map (
            O => \N__44328\,
            I => \n7_adj_839_cascade_\
        );

    \I__10436\ : IoInMux
    port map (
            O => \N__44325\,
            I => \N__44322\
        );

    \I__10435\ : LocalMux
    port map (
            O => \N__44322\,
            I => \N__44319\
        );

    \I__10434\ : IoSpan4Mux
    port map (
            O => \N__44319\,
            I => \N__44316\
        );

    \I__10433\ : Sp12to4
    port map (
            O => \N__44316\,
            I => \N__44313\
        );

    \I__10432\ : Span12Mux_s6_v
    port map (
            O => \N__44313\,
            I => \N__44310\
        );

    \I__10431\ : Span12Mux_h
    port map (
            O => \N__44310\,
            I => \N__44305\
        );

    \I__10430\ : InMux
    port map (
            O => \N__44309\,
            I => \N__44302\
        );

    \I__10429\ : InMux
    port map (
            O => \N__44308\,
            I => \N__44299\
        );

    \I__10428\ : Odrv12
    port map (
            O => \N__44305\,
            I => pin_out_18
        );

    \I__10427\ : LocalMux
    port map (
            O => \N__44302\,
            I => pin_out_18
        );

    \I__10426\ : LocalMux
    port map (
            O => \N__44299\,
            I => pin_out_18
        );

    \I__10425\ : IoInMux
    port map (
            O => \N__44292\,
            I => \N__44289\
        );

    \I__10424\ : LocalMux
    port map (
            O => \N__44289\,
            I => \N__44286\
        );

    \I__10423\ : IoSpan4Mux
    port map (
            O => \N__44286\,
            I => \N__44283\
        );

    \I__10422\ : Span4Mux_s1_v
    port map (
            O => \N__44283\,
            I => \N__44279\
        );

    \I__10421\ : CascadeMux
    port map (
            O => \N__44282\,
            I => \N__44275\
        );

    \I__10420\ : Sp12to4
    port map (
            O => \N__44279\,
            I => \N__44272\
        );

    \I__10419\ : CascadeMux
    port map (
            O => \N__44278\,
            I => \N__44269\
        );

    \I__10418\ : InMux
    port map (
            O => \N__44275\,
            I => \N__44266\
        );

    \I__10417\ : Span12Mux_v
    port map (
            O => \N__44272\,
            I => \N__44263\
        );

    \I__10416\ : InMux
    port map (
            O => \N__44269\,
            I => \N__44260\
        );

    \I__10415\ : LocalMux
    port map (
            O => \N__44266\,
            I => \N__44257\
        );

    \I__10414\ : Odrv12
    port map (
            O => \N__44263\,
            I => pin_out_19
        );

    \I__10413\ : LocalMux
    port map (
            O => \N__44260\,
            I => pin_out_19
        );

    \I__10412\ : Odrv4
    port map (
            O => \N__44257\,
            I => pin_out_19
        );

    \I__10411\ : CascadeMux
    port map (
            O => \N__44250\,
            I => \n11962_cascade_\
        );

    \I__10410\ : IoInMux
    port map (
            O => \N__44247\,
            I => \N__44244\
        );

    \I__10409\ : LocalMux
    port map (
            O => \N__44244\,
            I => \N__44241\
        );

    \I__10408\ : Span4Mux_s3_h
    port map (
            O => \N__44241\,
            I => \N__44238\
        );

    \I__10407\ : Span4Mux_v
    port map (
            O => \N__44238\,
            I => \N__44235\
        );

    \I__10406\ : Sp12to4
    port map (
            O => \N__44235\,
            I => \N__44232\
        );

    \I__10405\ : Span12Mux_h
    port map (
            O => \N__44232\,
            I => \N__44228\
        );

    \I__10404\ : InMux
    port map (
            O => \N__44231\,
            I => \N__44225\
        );

    \I__10403\ : Odrv12
    port map (
            O => \N__44228\,
            I => pin_oe_14
        );

    \I__10402\ : LocalMux
    port map (
            O => \N__44225\,
            I => pin_oe_14
        );

    \I__10401\ : InMux
    port map (
            O => \N__44220\,
            I => \N__44216\
        );

    \I__10400\ : InMux
    port map (
            O => \N__44219\,
            I => \N__44213\
        );

    \I__10399\ : LocalMux
    port map (
            O => \N__44216\,
            I => \N__44210\
        );

    \I__10398\ : LocalMux
    port map (
            O => \N__44213\,
            I => \N__44207\
        );

    \I__10397\ : Span4Mux_v
    port map (
            O => \N__44210\,
            I => \N__44204\
        );

    \I__10396\ : Odrv4
    port map (
            O => \N__44207\,
            I => n9_adj_812
        );

    \I__10395\ : Odrv4
    port map (
            O => \N__44204\,
            I => n9_adj_812
        );

    \I__10394\ : CascadeMux
    port map (
            O => \N__44199\,
            I => \N__44196\
        );

    \I__10393\ : InMux
    port map (
            O => \N__44196\,
            I => \N__44193\
        );

    \I__10392\ : LocalMux
    port map (
            O => \N__44193\,
            I => n8_adj_828
        );

    \I__10391\ : CascadeMux
    port map (
            O => \N__44190\,
            I => \n11958_cascade_\
        );

    \I__10390\ : IoInMux
    port map (
            O => \N__44187\,
            I => \N__44184\
        );

    \I__10389\ : LocalMux
    port map (
            O => \N__44184\,
            I => \N__44181\
        );

    \I__10388\ : Span4Mux_s0_v
    port map (
            O => \N__44181\,
            I => \N__44178\
        );

    \I__10387\ : Span4Mux_v
    port map (
            O => \N__44178\,
            I => \N__44175\
        );

    \I__10386\ : Sp12to4
    port map (
            O => \N__44175\,
            I => \N__44172\
        );

    \I__10385\ : Span12Mux_h
    port map (
            O => \N__44172\,
            I => \N__44169\
        );

    \I__10384\ : Span12Mux_v
    port map (
            O => \N__44169\,
            I => \N__44165\
        );

    \I__10383\ : InMux
    port map (
            O => \N__44168\,
            I => \N__44162\
        );

    \I__10382\ : Odrv12
    port map (
            O => \N__44165\,
            I => pin_oe_21
        );

    \I__10381\ : LocalMux
    port map (
            O => \N__44162\,
            I => pin_oe_21
        );

    \I__10380\ : InMux
    port map (
            O => \N__44157\,
            I => \N__44154\
        );

    \I__10379\ : LocalMux
    port map (
            O => \N__44154\,
            I => \N__44151\
        );

    \I__10378\ : Span4Mux_v
    port map (
            O => \N__44151\,
            I => \N__44148\
        );

    \I__10377\ : Sp12to4
    port map (
            O => \N__44148\,
            I => \N__44145\
        );

    \I__10376\ : Span12Mux_h
    port map (
            O => \N__44145\,
            I => \N__44142\
        );

    \I__10375\ : Odrv12
    port map (
            O => \N__44142\,
            I => n13652
        );

    \I__10374\ : CascadeMux
    port map (
            O => \N__44139\,
            I => \n13536_cascade_\
        );

    \I__10373\ : InMux
    port map (
            O => \N__44136\,
            I => \N__44133\
        );

    \I__10372\ : LocalMux
    port map (
            O => \N__44133\,
            I => \N__44130\
        );

    \I__10371\ : Span12Mux_h
    port map (
            O => \N__44130\,
            I => \N__44127\
        );

    \I__10370\ : Odrv12
    port map (
            O => \N__44127\,
            I => n13616
        );

    \I__10369\ : InMux
    port map (
            O => \N__44124\,
            I => \N__44121\
        );

    \I__10368\ : LocalMux
    port map (
            O => \N__44121\,
            I => n13542
        );

    \I__10367\ : CascadeMux
    port map (
            O => \N__44118\,
            I => \n7_adj_831_cascade_\
        );

    \I__10366\ : CascadeMux
    port map (
            O => \N__44115\,
            I => \N__44108\
        );

    \I__10365\ : CascadeMux
    port map (
            O => \N__44114\,
            I => \N__44102\
        );

    \I__10364\ : CascadeMux
    port map (
            O => \N__44113\,
            I => \N__44099\
        );

    \I__10363\ : InMux
    port map (
            O => \N__44112\,
            I => \N__44096\
        );

    \I__10362\ : CascadeMux
    port map (
            O => \N__44111\,
            I => \N__44092\
        );

    \I__10361\ : InMux
    port map (
            O => \N__44108\,
            I => \N__44088\
        );

    \I__10360\ : InMux
    port map (
            O => \N__44107\,
            I => \N__44085\
        );

    \I__10359\ : InMux
    port map (
            O => \N__44106\,
            I => \N__44082\
        );

    \I__10358\ : InMux
    port map (
            O => \N__44105\,
            I => \N__44079\
        );

    \I__10357\ : InMux
    port map (
            O => \N__44102\,
            I => \N__44076\
        );

    \I__10356\ : InMux
    port map (
            O => \N__44099\,
            I => \N__44073\
        );

    \I__10355\ : LocalMux
    port map (
            O => \N__44096\,
            I => \N__44070\
        );

    \I__10354\ : InMux
    port map (
            O => \N__44095\,
            I => \N__44067\
        );

    \I__10353\ : InMux
    port map (
            O => \N__44092\,
            I => \N__44064\
        );

    \I__10352\ : InMux
    port map (
            O => \N__44091\,
            I => \N__44060\
        );

    \I__10351\ : LocalMux
    port map (
            O => \N__44088\,
            I => \N__44055\
        );

    \I__10350\ : LocalMux
    port map (
            O => \N__44085\,
            I => \N__44055\
        );

    \I__10349\ : LocalMux
    port map (
            O => \N__44082\,
            I => \N__44052\
        );

    \I__10348\ : LocalMux
    port map (
            O => \N__44079\,
            I => \N__44047\
        );

    \I__10347\ : LocalMux
    port map (
            O => \N__44076\,
            I => \N__44047\
        );

    \I__10346\ : LocalMux
    port map (
            O => \N__44073\,
            I => \N__44044\
        );

    \I__10345\ : Span4Mux_v
    port map (
            O => \N__44070\,
            I => \N__44041\
        );

    \I__10344\ : LocalMux
    port map (
            O => \N__44067\,
            I => \N__44036\
        );

    \I__10343\ : LocalMux
    port map (
            O => \N__44064\,
            I => \N__44036\
        );

    \I__10342\ : InMux
    port map (
            O => \N__44063\,
            I => \N__44033\
        );

    \I__10341\ : LocalMux
    port map (
            O => \N__44060\,
            I => \N__44028\
        );

    \I__10340\ : Span4Mux_h
    port map (
            O => \N__44055\,
            I => \N__44028\
        );

    \I__10339\ : Span4Mux_h
    port map (
            O => \N__44052\,
            I => \N__44021\
        );

    \I__10338\ : Span4Mux_h
    port map (
            O => \N__44047\,
            I => \N__44021\
        );

    \I__10337\ : Span4Mux_h
    port map (
            O => \N__44044\,
            I => \N__44021\
        );

    \I__10336\ : Span4Mux_h
    port map (
            O => \N__44041\,
            I => \N__44016\
        );

    \I__10335\ : Span4Mux_v
    port map (
            O => \N__44036\,
            I => \N__44016\
        );

    \I__10334\ : LocalMux
    port map (
            O => \N__44033\,
            I => n6_adj_813
        );

    \I__10333\ : Odrv4
    port map (
            O => \N__44028\,
            I => n6_adj_813
        );

    \I__10332\ : Odrv4
    port map (
            O => \N__44021\,
            I => n6_adj_813
        );

    \I__10331\ : Odrv4
    port map (
            O => \N__44016\,
            I => n6_adj_813
        );

    \I__10330\ : CascadeMux
    port map (
            O => \N__44007\,
            I => \n11825_cascade_\
        );

    \I__10329\ : IoInMux
    port map (
            O => \N__44004\,
            I => \N__44001\
        );

    \I__10328\ : LocalMux
    port map (
            O => \N__44001\,
            I => \N__43998\
        );

    \I__10327\ : IoSpan4Mux
    port map (
            O => \N__43998\,
            I => \N__43995\
        );

    \I__10326\ : Span4Mux_s3_h
    port map (
            O => \N__43995\,
            I => \N__43992\
        );

    \I__10325\ : Span4Mux_h
    port map (
            O => \N__43992\,
            I => \N__43989\
        );

    \I__10324\ : Span4Mux_h
    port map (
            O => \N__43989\,
            I => \N__43985\
        );

    \I__10323\ : InMux
    port map (
            O => \N__43988\,
            I => \N__43982\
        );

    \I__10322\ : Odrv4
    port map (
            O => \N__43985\,
            I => pin_oe_15
        );

    \I__10321\ : LocalMux
    port map (
            O => \N__43982\,
            I => pin_oe_15
        );

    \I__10320\ : InMux
    port map (
            O => \N__43977\,
            I => \N__43971\
        );

    \I__10319\ : InMux
    port map (
            O => \N__43976\,
            I => \N__43971\
        );

    \I__10318\ : LocalMux
    port map (
            O => \N__43971\,
            I => \N__43968\
        );

    \I__10317\ : Span4Mux_h
    port map (
            O => \N__43968\,
            I => \N__43965\
        );

    \I__10316\ : Span4Mux_h
    port map (
            O => \N__43965\,
            I => \N__43962\
        );

    \I__10315\ : Span4Mux_h
    port map (
            O => \N__43962\,
            I => \N__43959\
        );

    \I__10314\ : Odrv4
    port map (
            O => \N__43959\,
            I => n1907
        );

    \I__10313\ : CascadeMux
    port map (
            O => \N__43956\,
            I => \N__43952\
        );

    \I__10312\ : InMux
    port map (
            O => \N__43955\,
            I => \N__43948\
        );

    \I__10311\ : InMux
    port map (
            O => \N__43952\,
            I => \N__43944\
        );

    \I__10310\ : InMux
    port map (
            O => \N__43951\,
            I => \N__43941\
        );

    \I__10309\ : LocalMux
    port map (
            O => \N__43948\,
            I => \N__43936\
        );

    \I__10308\ : InMux
    port map (
            O => \N__43947\,
            I => \N__43933\
        );

    \I__10307\ : LocalMux
    port map (
            O => \N__43944\,
            I => \N__43929\
        );

    \I__10306\ : LocalMux
    port map (
            O => \N__43941\,
            I => \N__43926\
        );

    \I__10305\ : CascadeMux
    port map (
            O => \N__43940\,
            I => \N__43922\
        );

    \I__10304\ : InMux
    port map (
            O => \N__43939\,
            I => \N__43919\
        );

    \I__10303\ : Span4Mux_v
    port map (
            O => \N__43936\,
            I => \N__43916\
        );

    \I__10302\ : LocalMux
    port map (
            O => \N__43933\,
            I => \N__43913\
        );

    \I__10301\ : InMux
    port map (
            O => \N__43932\,
            I => \N__43907\
        );

    \I__10300\ : Span4Mux_v
    port map (
            O => \N__43929\,
            I => \N__43902\
        );

    \I__10299\ : Span4Mux_h
    port map (
            O => \N__43926\,
            I => \N__43902\
        );

    \I__10298\ : InMux
    port map (
            O => \N__43925\,
            I => \N__43899\
        );

    \I__10297\ : InMux
    port map (
            O => \N__43922\,
            I => \N__43887\
        );

    \I__10296\ : LocalMux
    port map (
            O => \N__43919\,
            I => \N__43884\
        );

    \I__10295\ : Span4Mux_h
    port map (
            O => \N__43916\,
            I => \N__43879\
        );

    \I__10294\ : Span4Mux_v
    port map (
            O => \N__43913\,
            I => \N__43879\
        );

    \I__10293\ : CascadeMux
    port map (
            O => \N__43912\,
            I => \N__43876\
        );

    \I__10292\ : InMux
    port map (
            O => \N__43911\,
            I => \N__43869\
        );

    \I__10291\ : InMux
    port map (
            O => \N__43910\,
            I => \N__43869\
        );

    \I__10290\ : LocalMux
    port map (
            O => \N__43907\,
            I => \N__43866\
        );

    \I__10289\ : Span4Mux_v
    port map (
            O => \N__43902\,
            I => \N__43861\
        );

    \I__10288\ : LocalMux
    port map (
            O => \N__43899\,
            I => \N__43861\
        );

    \I__10287\ : InMux
    port map (
            O => \N__43898\,
            I => \N__43858\
        );

    \I__10286\ : InMux
    port map (
            O => \N__43897\,
            I => \N__43853\
        );

    \I__10285\ : InMux
    port map (
            O => \N__43896\,
            I => \N__43853\
        );

    \I__10284\ : InMux
    port map (
            O => \N__43895\,
            I => \N__43846\
        );

    \I__10283\ : InMux
    port map (
            O => \N__43894\,
            I => \N__43846\
        );

    \I__10282\ : InMux
    port map (
            O => \N__43893\,
            I => \N__43846\
        );

    \I__10281\ : InMux
    port map (
            O => \N__43892\,
            I => \N__43843\
        );

    \I__10280\ : InMux
    port map (
            O => \N__43891\,
            I => \N__43840\
        );

    \I__10279\ : CascadeMux
    port map (
            O => \N__43890\,
            I => \N__43837\
        );

    \I__10278\ : LocalMux
    port map (
            O => \N__43887\,
            I => \N__43833\
        );

    \I__10277\ : Span4Mux_v
    port map (
            O => \N__43884\,
            I => \N__43828\
        );

    \I__10276\ : Span4Mux_v
    port map (
            O => \N__43879\,
            I => \N__43828\
        );

    \I__10275\ : InMux
    port map (
            O => \N__43876\,
            I => \N__43825\
        );

    \I__10274\ : CascadeMux
    port map (
            O => \N__43875\,
            I => \N__43819\
        );

    \I__10273\ : InMux
    port map (
            O => \N__43874\,
            I => \N__43814\
        );

    \I__10272\ : LocalMux
    port map (
            O => \N__43869\,
            I => \N__43811\
        );

    \I__10271\ : Span4Mux_h
    port map (
            O => \N__43866\,
            I => \N__43806\
        );

    \I__10270\ : Span4Mux_v
    port map (
            O => \N__43861\,
            I => \N__43806\
        );

    \I__10269\ : LocalMux
    port map (
            O => \N__43858\,
            I => \N__43797\
        );

    \I__10268\ : LocalMux
    port map (
            O => \N__43853\,
            I => \N__43797\
        );

    \I__10267\ : LocalMux
    port map (
            O => \N__43846\,
            I => \N__43797\
        );

    \I__10266\ : LocalMux
    port map (
            O => \N__43843\,
            I => \N__43797\
        );

    \I__10265\ : LocalMux
    port map (
            O => \N__43840\,
            I => \N__43794\
        );

    \I__10264\ : InMux
    port map (
            O => \N__43837\,
            I => \N__43791\
        );

    \I__10263\ : InMux
    port map (
            O => \N__43836\,
            I => \N__43788\
        );

    \I__10262\ : Span12Mux_v
    port map (
            O => \N__43833\,
            I => \N__43783\
        );

    \I__10261\ : Sp12to4
    port map (
            O => \N__43828\,
            I => \N__43783\
        );

    \I__10260\ : LocalMux
    port map (
            O => \N__43825\,
            I => \N__43780\
        );

    \I__10259\ : InMux
    port map (
            O => \N__43824\,
            I => \N__43777\
        );

    \I__10258\ : InMux
    port map (
            O => \N__43823\,
            I => \N__43774\
        );

    \I__10257\ : InMux
    port map (
            O => \N__43822\,
            I => \N__43771\
        );

    \I__10256\ : InMux
    port map (
            O => \N__43819\,
            I => \N__43768\
        );

    \I__10255\ : InMux
    port map (
            O => \N__43818\,
            I => \N__43765\
        );

    \I__10254\ : InMux
    port map (
            O => \N__43817\,
            I => \N__43762\
        );

    \I__10253\ : LocalMux
    port map (
            O => \N__43814\,
            I => \N__43755\
        );

    \I__10252\ : Span4Mux_v
    port map (
            O => \N__43811\,
            I => \N__43755\
        );

    \I__10251\ : Span4Mux_h
    port map (
            O => \N__43806\,
            I => \N__43755\
        );

    \I__10250\ : Span12Mux_v
    port map (
            O => \N__43797\,
            I => \N__43752\
        );

    \I__10249\ : Span4Mux_h
    port map (
            O => \N__43794\,
            I => \N__43745\
        );

    \I__10248\ : LocalMux
    port map (
            O => \N__43791\,
            I => \N__43745\
        );

    \I__10247\ : LocalMux
    port map (
            O => \N__43788\,
            I => \N__43745\
        );

    \I__10246\ : Span12Mux_h
    port map (
            O => \N__43783\,
            I => \N__43740\
        );

    \I__10245\ : Span12Mux_h
    port map (
            O => \N__43780\,
            I => \N__43740\
        );

    \I__10244\ : LocalMux
    port map (
            O => \N__43777\,
            I => \N__43737\
        );

    \I__10243\ : LocalMux
    port map (
            O => \N__43774\,
            I => state_1
        );

    \I__10242\ : LocalMux
    port map (
            O => \N__43771\,
            I => state_1
        );

    \I__10241\ : LocalMux
    port map (
            O => \N__43768\,
            I => state_1
        );

    \I__10240\ : LocalMux
    port map (
            O => \N__43765\,
            I => state_1
        );

    \I__10239\ : LocalMux
    port map (
            O => \N__43762\,
            I => state_1
        );

    \I__10238\ : Odrv4
    port map (
            O => \N__43755\,
            I => state_1
        );

    \I__10237\ : Odrv12
    port map (
            O => \N__43752\,
            I => state_1
        );

    \I__10236\ : Odrv4
    port map (
            O => \N__43745\,
            I => state_1
        );

    \I__10235\ : Odrv12
    port map (
            O => \N__43740\,
            I => state_1
        );

    \I__10234\ : Odrv4
    port map (
            O => \N__43737\,
            I => state_1
        );

    \I__10233\ : InMux
    port map (
            O => \N__43716\,
            I => \N__43712\
        );

    \I__10232\ : CascadeMux
    port map (
            O => \N__43715\,
            I => \N__43708\
        );

    \I__10231\ : LocalMux
    port map (
            O => \N__43712\,
            I => \N__43705\
        );

    \I__10230\ : InMux
    port map (
            O => \N__43711\,
            I => \N__43702\
        );

    \I__10229\ : InMux
    port map (
            O => \N__43708\,
            I => \N__43698\
        );

    \I__10228\ : Span4Mux_h
    port map (
            O => \N__43705\,
            I => \N__43693\
        );

    \I__10227\ : LocalMux
    port map (
            O => \N__43702\,
            I => \N__43693\
        );

    \I__10226\ : CascadeMux
    port map (
            O => \N__43701\,
            I => \N__43688\
        );

    \I__10225\ : LocalMux
    port map (
            O => \N__43698\,
            I => \N__43685\
        );

    \I__10224\ : Span4Mux_v
    port map (
            O => \N__43693\,
            I => \N__43682\
        );

    \I__10223\ : CascadeMux
    port map (
            O => \N__43692\,
            I => \N__43677\
        );

    \I__10222\ : CascadeMux
    port map (
            O => \N__43691\,
            I => \N__43672\
        );

    \I__10221\ : InMux
    port map (
            O => \N__43688\,
            I => \N__43669\
        );

    \I__10220\ : Span4Mux_v
    port map (
            O => \N__43685\,
            I => \N__43663\
        );

    \I__10219\ : Span4Mux_v
    port map (
            O => \N__43682\,
            I => \N__43663\
        );

    \I__10218\ : InMux
    port map (
            O => \N__43681\,
            I => \N__43660\
        );

    \I__10217\ : InMux
    port map (
            O => \N__43680\,
            I => \N__43653\
        );

    \I__10216\ : InMux
    port map (
            O => \N__43677\,
            I => \N__43653\
        );

    \I__10215\ : InMux
    port map (
            O => \N__43676\,
            I => \N__43653\
        );

    \I__10214\ : InMux
    port map (
            O => \N__43675\,
            I => \N__43648\
        );

    \I__10213\ : InMux
    port map (
            O => \N__43672\,
            I => \N__43645\
        );

    \I__10212\ : LocalMux
    port map (
            O => \N__43669\,
            I => \N__43642\
        );

    \I__10211\ : CascadeMux
    port map (
            O => \N__43668\,
            I => \N__43637\
        );

    \I__10210\ : Span4Mux_h
    port map (
            O => \N__43663\,
            I => \N__43632\
        );

    \I__10209\ : LocalMux
    port map (
            O => \N__43660\,
            I => \N__43632\
        );

    \I__10208\ : LocalMux
    port map (
            O => \N__43653\,
            I => \N__43629\
        );

    \I__10207\ : InMux
    port map (
            O => \N__43652\,
            I => \N__43626\
        );

    \I__10206\ : CascadeMux
    port map (
            O => \N__43651\,
            I => \N__43622\
        );

    \I__10205\ : LocalMux
    port map (
            O => \N__43648\,
            I => \N__43619\
        );

    \I__10204\ : LocalMux
    port map (
            O => \N__43645\,
            I => \N__43614\
        );

    \I__10203\ : Span4Mux_h
    port map (
            O => \N__43642\,
            I => \N__43614\
        );

    \I__10202\ : InMux
    port map (
            O => \N__43641\,
            I => \N__43611\
        );

    \I__10201\ : InMux
    port map (
            O => \N__43640\,
            I => \N__43606\
        );

    \I__10200\ : InMux
    port map (
            O => \N__43637\,
            I => \N__43606\
        );

    \I__10199\ : Span4Mux_v
    port map (
            O => \N__43632\,
            I => \N__43601\
        );

    \I__10198\ : Span4Mux_v
    port map (
            O => \N__43629\,
            I => \N__43601\
        );

    \I__10197\ : LocalMux
    port map (
            O => \N__43626\,
            I => \N__43597\
        );

    \I__10196\ : InMux
    port map (
            O => \N__43625\,
            I => \N__43593\
        );

    \I__10195\ : InMux
    port map (
            O => \N__43622\,
            I => \N__43589\
        );

    \I__10194\ : Span12Mux_v
    port map (
            O => \N__43619\,
            I => \N__43585\
        );

    \I__10193\ : Span4Mux_v
    port map (
            O => \N__43614\,
            I => \N__43581\
        );

    \I__10192\ : LocalMux
    port map (
            O => \N__43611\,
            I => \N__43576\
        );

    \I__10191\ : LocalMux
    port map (
            O => \N__43606\,
            I => \N__43576\
        );

    \I__10190\ : Span4Mux_h
    port map (
            O => \N__43601\,
            I => \N__43573\
        );

    \I__10189\ : InMux
    port map (
            O => \N__43600\,
            I => \N__43570\
        );

    \I__10188\ : Sp12to4
    port map (
            O => \N__43597\,
            I => \N__43567\
        );

    \I__10187\ : InMux
    port map (
            O => \N__43596\,
            I => \N__43564\
        );

    \I__10186\ : LocalMux
    port map (
            O => \N__43593\,
            I => \N__43561\
        );

    \I__10185\ : InMux
    port map (
            O => \N__43592\,
            I => \N__43558\
        );

    \I__10184\ : LocalMux
    port map (
            O => \N__43589\,
            I => \N__43555\
        );

    \I__10183\ : InMux
    port map (
            O => \N__43588\,
            I => \N__43552\
        );

    \I__10182\ : Span12Mux_h
    port map (
            O => \N__43585\,
            I => \N__43549\
        );

    \I__10181\ : InMux
    port map (
            O => \N__43584\,
            I => \N__43546\
        );

    \I__10180\ : Span4Mux_h
    port map (
            O => \N__43581\,
            I => \N__43541\
        );

    \I__10179\ : Span4Mux_v
    port map (
            O => \N__43576\,
            I => \N__43541\
        );

    \I__10178\ : Span4Mux_h
    port map (
            O => \N__43573\,
            I => \N__43536\
        );

    \I__10177\ : LocalMux
    port map (
            O => \N__43570\,
            I => \N__43536\
        );

    \I__10176\ : Span12Mux_v
    port map (
            O => \N__43567\,
            I => \N__43533\
        );

    \I__10175\ : LocalMux
    port map (
            O => \N__43564\,
            I => \N__43528\
        );

    \I__10174\ : Span12Mux_h
    port map (
            O => \N__43561\,
            I => \N__43528\
        );

    \I__10173\ : LocalMux
    port map (
            O => \N__43558\,
            I => \N__43521\
        );

    \I__10172\ : Span4Mux_v
    port map (
            O => \N__43555\,
            I => \N__43521\
        );

    \I__10171\ : LocalMux
    port map (
            O => \N__43552\,
            I => \N__43521\
        );

    \I__10170\ : Odrv12
    port map (
            O => \N__43549\,
            I => state_2
        );

    \I__10169\ : LocalMux
    port map (
            O => \N__43546\,
            I => state_2
        );

    \I__10168\ : Odrv4
    port map (
            O => \N__43541\,
            I => state_2
        );

    \I__10167\ : Odrv4
    port map (
            O => \N__43536\,
            I => state_2
        );

    \I__10166\ : Odrv12
    port map (
            O => \N__43533\,
            I => state_2
        );

    \I__10165\ : Odrv12
    port map (
            O => \N__43528\,
            I => state_2
        );

    \I__10164\ : Odrv4
    port map (
            O => \N__43521\,
            I => state_2
        );

    \I__10163\ : SRMux
    port map (
            O => \N__43506\,
            I => \N__43502\
        );

    \I__10162\ : SRMux
    port map (
            O => \N__43505\,
            I => \N__43499\
        );

    \I__10161\ : LocalMux
    port map (
            O => \N__43502\,
            I => \N__43496\
        );

    \I__10160\ : LocalMux
    port map (
            O => \N__43499\,
            I => \N__43493\
        );

    \I__10159\ : Span4Mux_s1_h
    port map (
            O => \N__43496\,
            I => \N__43486\
        );

    \I__10158\ : Span4Mux_v
    port map (
            O => \N__43493\,
            I => \N__43486\
        );

    \I__10157\ : SRMux
    port map (
            O => \N__43492\,
            I => \N__43483\
        );

    \I__10156\ : SRMux
    port map (
            O => \N__43491\,
            I => \N__43480\
        );

    \I__10155\ : Span4Mux_v
    port map (
            O => \N__43486\,
            I => \N__43473\
        );

    \I__10154\ : LocalMux
    port map (
            O => \N__43483\,
            I => \N__43473\
        );

    \I__10153\ : LocalMux
    port map (
            O => \N__43480\,
            I => \N__43473\
        );

    \I__10152\ : Span4Mux_v
    port map (
            O => \N__43473\,
            I => \N__43470\
        );

    \I__10151\ : Sp12to4
    port map (
            O => \N__43470\,
            I => \N__43467\
        );

    \I__10150\ : Span12Mux_s5_h
    port map (
            O => \N__43467\,
            I => \N__43464\
        );

    \I__10149\ : Span12Mux_h
    port map (
            O => \N__43464\,
            I => \N__43461\
        );

    \I__10148\ : Odrv12
    port map (
            O => \N__43461\,
            I => n8025
        );

    \I__10147\ : CascadeMux
    port map (
            O => \N__43458\,
            I => \n11954_cascade_\
        );

    \I__10146\ : IoInMux
    port map (
            O => \N__43455\,
            I => \N__43452\
        );

    \I__10145\ : LocalMux
    port map (
            O => \N__43452\,
            I => \N__43449\
        );

    \I__10144\ : IoSpan4Mux
    port map (
            O => \N__43449\,
            I => \N__43446\
        );

    \I__10143\ : Sp12to4
    port map (
            O => \N__43446\,
            I => \N__43443\
        );

    \I__10142\ : Span12Mux_v
    port map (
            O => \N__43443\,
            I => \N__43439\
        );

    \I__10141\ : InMux
    port map (
            O => \N__43442\,
            I => \N__43436\
        );

    \I__10140\ : Odrv12
    port map (
            O => \N__43439\,
            I => pin_oe_20
        );

    \I__10139\ : LocalMux
    port map (
            O => \N__43436\,
            I => pin_oe_20
        );

    \I__10138\ : InMux
    port map (
            O => \N__43431\,
            I => \N__43425\
        );

    \I__10137\ : InMux
    port map (
            O => \N__43430\,
            I => \N__43421\
        );

    \I__10136\ : InMux
    port map (
            O => \N__43429\,
            I => \N__43418\
        );

    \I__10135\ : InMux
    port map (
            O => \N__43428\,
            I => \N__43415\
        );

    \I__10134\ : LocalMux
    port map (
            O => \N__43425\,
            I => \N__43411\
        );

    \I__10133\ : InMux
    port map (
            O => \N__43424\,
            I => \N__43408\
        );

    \I__10132\ : LocalMux
    port map (
            O => \N__43421\,
            I => \N__43405\
        );

    \I__10131\ : LocalMux
    port map (
            O => \N__43418\,
            I => \N__43402\
        );

    \I__10130\ : LocalMux
    port map (
            O => \N__43415\,
            I => \N__43399\
        );

    \I__10129\ : InMux
    port map (
            O => \N__43414\,
            I => \N__43395\
        );

    \I__10128\ : Span4Mux_v
    port map (
            O => \N__43411\,
            I => \N__43392\
        );

    \I__10127\ : LocalMux
    port map (
            O => \N__43408\,
            I => \N__43389\
        );

    \I__10126\ : Span4Mux_h
    port map (
            O => \N__43405\,
            I => \N__43386\
        );

    \I__10125\ : Span4Mux_h
    port map (
            O => \N__43402\,
            I => \N__43381\
        );

    \I__10124\ : Span4Mux_h
    port map (
            O => \N__43399\,
            I => \N__43381\
        );

    \I__10123\ : InMux
    port map (
            O => \N__43398\,
            I => \N__43378\
        );

    \I__10122\ : LocalMux
    port map (
            O => \N__43395\,
            I => n9488
        );

    \I__10121\ : Odrv4
    port map (
            O => \N__43392\,
            I => n9488
        );

    \I__10120\ : Odrv12
    port map (
            O => \N__43389\,
            I => n9488
        );

    \I__10119\ : Odrv4
    port map (
            O => \N__43386\,
            I => n9488
        );

    \I__10118\ : Odrv4
    port map (
            O => \N__43381\,
            I => n9488
        );

    \I__10117\ : LocalMux
    port map (
            O => \N__43378\,
            I => n9488
        );

    \I__10116\ : InMux
    port map (
            O => \N__43365\,
            I => \N__43362\
        );

    \I__10115\ : LocalMux
    port map (
            O => \N__43362\,
            I => n11821
        );

    \I__10114\ : InMux
    port map (
            O => \N__43359\,
            I => \N__43356\
        );

    \I__10113\ : LocalMux
    port map (
            O => \N__43356\,
            I => n8_adj_826
        );

    \I__10112\ : IoInMux
    port map (
            O => \N__43353\,
            I => \N__43350\
        );

    \I__10111\ : LocalMux
    port map (
            O => \N__43350\,
            I => \N__43347\
        );

    \I__10110\ : IoSpan4Mux
    port map (
            O => \N__43347\,
            I => \N__43344\
        );

    \I__10109\ : IoSpan4Mux
    port map (
            O => \N__43344\,
            I => \N__43341\
        );

    \I__10108\ : Span4Mux_s3_v
    port map (
            O => \N__43341\,
            I => \N__43337\
        );

    \I__10107\ : InMux
    port map (
            O => \N__43340\,
            I => \N__43333\
        );

    \I__10106\ : Sp12to4
    port map (
            O => \N__43337\,
            I => \N__43330\
        );

    \I__10105\ : CascadeMux
    port map (
            O => \N__43336\,
            I => \N__43327\
        );

    \I__10104\ : LocalMux
    port map (
            O => \N__43333\,
            I => \N__43324\
        );

    \I__10103\ : Span12Mux_s10_v
    port map (
            O => \N__43330\,
            I => \N__43321\
        );

    \I__10102\ : InMux
    port map (
            O => \N__43327\,
            I => \N__43318\
        );

    \I__10101\ : Span4Mux_h
    port map (
            O => \N__43324\,
            I => \N__43315\
        );

    \I__10100\ : Odrv12
    port map (
            O => \N__43321\,
            I => pin_out_8
        );

    \I__10099\ : LocalMux
    port map (
            O => \N__43318\,
            I => pin_out_8
        );

    \I__10098\ : Odrv4
    port map (
            O => \N__43315\,
            I => pin_out_8
        );

    \I__10097\ : InMux
    port map (
            O => \N__43308\,
            I => \N__43305\
        );

    \I__10096\ : LocalMux
    port map (
            O => \N__43305\,
            I => n8_adj_832
        );

    \I__10095\ : InMux
    port map (
            O => \N__43302\,
            I => \N__43299\
        );

    \I__10094\ : LocalMux
    port map (
            O => \N__43299\,
            I => \pin_out_22__N_216\
        );

    \I__10093\ : CascadeMux
    port map (
            O => \N__43296\,
            I => \pin_out_22__N_216_cascade_\
        );

    \I__10092\ : InMux
    port map (
            O => \N__43293\,
            I => \N__43290\
        );

    \I__10091\ : LocalMux
    port map (
            O => \N__43290\,
            I => \N__43287\
        );

    \I__10090\ : Odrv4
    port map (
            O => \N__43287\,
            I => n13370
        );

    \I__10089\ : CascadeMux
    port map (
            O => \N__43284\,
            I => \N__43281\
        );

    \I__10088\ : InMux
    port map (
            O => \N__43281\,
            I => \N__43278\
        );

    \I__10087\ : LocalMux
    port map (
            O => \N__43278\,
            I => \N__43275\
        );

    \I__10086\ : Odrv4
    port map (
            O => \N__43275\,
            I => n13369
        );

    \I__10085\ : CascadeMux
    port map (
            O => \N__43272\,
            I => \n13640_cascade_\
        );

    \I__10084\ : InMux
    port map (
            O => \N__43269\,
            I => \N__43266\
        );

    \I__10083\ : LocalMux
    port map (
            O => \N__43266\,
            I => \N__43263\
        );

    \I__10082\ : Span4Mux_h
    port map (
            O => \N__43263\,
            I => \N__43260\
        );

    \I__10081\ : Odrv4
    port map (
            O => \N__43260\,
            I => n13628
        );

    \I__10080\ : CascadeMux
    port map (
            O => \N__43257\,
            I => \N__43254\
        );

    \I__10079\ : InMux
    port map (
            O => \N__43254\,
            I => \N__43251\
        );

    \I__10078\ : LocalMux
    port map (
            O => \N__43251\,
            I => n13540
        );

    \I__10077\ : InMux
    port map (
            O => \N__43248\,
            I => \N__43245\
        );

    \I__10076\ : LocalMux
    port map (
            O => \N__43245\,
            I => \N__43233\
        );

    \I__10075\ : InMux
    port map (
            O => \N__43244\,
            I => \N__43230\
        );

    \I__10074\ : InMux
    port map (
            O => \N__43243\,
            I => \N__43225\
        );

    \I__10073\ : InMux
    port map (
            O => \N__43242\,
            I => \N__43225\
        );

    \I__10072\ : InMux
    port map (
            O => \N__43241\,
            I => \N__43218\
        );

    \I__10071\ : InMux
    port map (
            O => \N__43240\,
            I => \N__43218\
        );

    \I__10070\ : InMux
    port map (
            O => \N__43239\,
            I => \N__43218\
        );

    \I__10069\ : InMux
    port map (
            O => \N__43238\,
            I => \N__43211\
        );

    \I__10068\ : InMux
    port map (
            O => \N__43237\,
            I => \N__43211\
        );

    \I__10067\ : InMux
    port map (
            O => \N__43236\,
            I => \N__43211\
        );

    \I__10066\ : Odrv4
    port map (
            O => \N__43233\,
            I => current_pin_4
        );

    \I__10065\ : LocalMux
    port map (
            O => \N__43230\,
            I => current_pin_4
        );

    \I__10064\ : LocalMux
    port map (
            O => \N__43225\,
            I => current_pin_4
        );

    \I__10063\ : LocalMux
    port map (
            O => \N__43218\,
            I => current_pin_4
        );

    \I__10062\ : LocalMux
    port map (
            O => \N__43211\,
            I => current_pin_4
        );

    \I__10061\ : CascadeMux
    port map (
            O => \N__43200\,
            I => \n7_adj_797_cascade_\
        );

    \I__10060\ : InMux
    port map (
            O => \N__43197\,
            I => \N__43194\
        );

    \I__10059\ : LocalMux
    port map (
            O => \N__43194\,
            I => n13551
        );

    \I__10058\ : CascadeMux
    port map (
            O => \N__43191\,
            I => \N__43187\
        );

    \I__10057\ : InMux
    port map (
            O => \N__43190\,
            I => \N__43180\
        );

    \I__10056\ : InMux
    port map (
            O => \N__43187\,
            I => \N__43175\
        );

    \I__10055\ : InMux
    port map (
            O => \N__43186\,
            I => \N__43175\
        );

    \I__10054\ : CascadeMux
    port map (
            O => \N__43185\,
            I => \N__43171\
        );

    \I__10053\ : InMux
    port map (
            O => \N__43184\,
            I => \N__43168\
        );

    \I__10052\ : CascadeMux
    port map (
            O => \N__43183\,
            I => \N__43165\
        );

    \I__10051\ : LocalMux
    port map (
            O => \N__43180\,
            I => \N__43160\
        );

    \I__10050\ : LocalMux
    port map (
            O => \N__43175\,
            I => \N__43160\
        );

    \I__10049\ : InMux
    port map (
            O => \N__43174\,
            I => \N__43157\
        );

    \I__10048\ : InMux
    port map (
            O => \N__43171\,
            I => \N__43154\
        );

    \I__10047\ : LocalMux
    port map (
            O => \N__43168\,
            I => \N__43151\
        );

    \I__10046\ : InMux
    port map (
            O => \N__43165\,
            I => \N__43148\
        );

    \I__10045\ : Span4Mux_h
    port map (
            O => \N__43160\,
            I => \N__43143\
        );

    \I__10044\ : LocalMux
    port map (
            O => \N__43157\,
            I => \N__43143\
        );

    \I__10043\ : LocalMux
    port map (
            O => \N__43154\,
            I => \N__43140\
        );

    \I__10042\ : Span4Mux_h
    port map (
            O => \N__43151\,
            I => \N__43137\
        );

    \I__10041\ : LocalMux
    port map (
            O => \N__43148\,
            I => \state_7_N_167_2\
        );

    \I__10040\ : Odrv4
    port map (
            O => \N__43143\,
            I => \state_7_N_167_2\
        );

    \I__10039\ : Odrv12
    port map (
            O => \N__43140\,
            I => \state_7_N_167_2\
        );

    \I__10038\ : Odrv4
    port map (
            O => \N__43137\,
            I => \state_7_N_167_2\
        );

    \I__10037\ : InMux
    port map (
            O => \N__43128\,
            I => \N__43125\
        );

    \I__10036\ : LocalMux
    port map (
            O => \N__43125\,
            I => \N__43122\
        );

    \I__10035\ : Odrv4
    port map (
            O => \N__43122\,
            I => n26
        );

    \I__10034\ : CascadeMux
    port map (
            O => \N__43119\,
            I => \N__43116\
        );

    \I__10033\ : InMux
    port map (
            O => \N__43116\,
            I => \N__43112\
        );

    \I__10032\ : InMux
    port map (
            O => \N__43115\,
            I => \N__43109\
        );

    \I__10031\ : LocalMux
    port map (
            O => \N__43112\,
            I => counter_4
        );

    \I__10030\ : LocalMux
    port map (
            O => \N__43109\,
            I => counter_4
        );

    \I__10029\ : InMux
    port map (
            O => \N__43104\,
            I => \N__43100\
        );

    \I__10028\ : InMux
    port map (
            O => \N__43103\,
            I => \N__43097\
        );

    \I__10027\ : LocalMux
    port map (
            O => \N__43100\,
            I => counter_5
        );

    \I__10026\ : LocalMux
    port map (
            O => \N__43097\,
            I => counter_5
        );

    \I__10025\ : CascadeMux
    port map (
            O => \N__43092\,
            I => \N__43088\
        );

    \I__10024\ : CascadeMux
    port map (
            O => \N__43091\,
            I => \N__43085\
        );

    \I__10023\ : InMux
    port map (
            O => \N__43088\,
            I => \N__43082\
        );

    \I__10022\ : InMux
    port map (
            O => \N__43085\,
            I => \N__43079\
        );

    \I__10021\ : LocalMux
    port map (
            O => \N__43082\,
            I => counter_2
        );

    \I__10020\ : LocalMux
    port map (
            O => \N__43079\,
            I => counter_2
        );

    \I__10019\ : InMux
    port map (
            O => \N__43074\,
            I => \N__43070\
        );

    \I__10018\ : InMux
    port map (
            O => \N__43073\,
            I => \N__43067\
        );

    \I__10017\ : LocalMux
    port map (
            O => \N__43070\,
            I => counter_3
        );

    \I__10016\ : LocalMux
    port map (
            O => \N__43067\,
            I => counter_3
        );

    \I__10015\ : InMux
    port map (
            O => \N__43062\,
            I => \N__43059\
        );

    \I__10014\ : LocalMux
    port map (
            O => \N__43059\,
            I => n14
        );

    \I__10013\ : IoInMux
    port map (
            O => \N__43056\,
            I => \N__43053\
        );

    \I__10012\ : LocalMux
    port map (
            O => \N__43053\,
            I => \N__43050\
        );

    \I__10011\ : Span12Mux_s5_h
    port map (
            O => \N__43050\,
            I => \N__43047\
        );

    \I__10010\ : Span12Mux_h
    port map (
            O => \N__43047\,
            I => \N__43044\
        );

    \I__10009\ : Span12Mux_v
    port map (
            O => \N__43044\,
            I => \N__43039\
        );

    \I__10008\ : InMux
    port map (
            O => \N__43043\,
            I => \N__43034\
        );

    \I__10007\ : InMux
    port map (
            O => \N__43042\,
            I => \N__43034\
        );

    \I__10006\ : Odrv12
    port map (
            O => \N__43039\,
            I => pin_out_11
        );

    \I__10005\ : LocalMux
    port map (
            O => \N__43034\,
            I => pin_out_11
        );

    \I__10004\ : CascadeMux
    port map (
            O => \N__43029\,
            I => \n7_adj_827_cascade_\
        );

    \I__10003\ : IoInMux
    port map (
            O => \N__43026\,
            I => \N__43023\
        );

    \I__10002\ : LocalMux
    port map (
            O => \N__43023\,
            I => \N__43020\
        );

    \I__10001\ : Span4Mux_s3_v
    port map (
            O => \N__43020\,
            I => \N__43017\
        );

    \I__10000\ : Sp12to4
    port map (
            O => \N__43017\,
            I => \N__43014\
        );

    \I__9999\ : Span12Mux_h
    port map (
            O => \N__43014\,
            I => \N__43011\
        );

    \I__9998\ : Span12Mux_v
    port map (
            O => \N__43011\,
            I => \N__43006\
        );

    \I__9997\ : InMux
    port map (
            O => \N__43010\,
            I => \N__43001\
        );

    \I__9996\ : InMux
    port map (
            O => \N__43009\,
            I => \N__43001\
        );

    \I__9995\ : Odrv12
    port map (
            O => \N__43006\,
            I => pin_out_10
        );

    \I__9994\ : LocalMux
    port map (
            O => \N__43001\,
            I => pin_out_10
        );

    \I__9993\ : CascadeMux
    port map (
            O => \N__42996\,
            I => \n9675_cascade_\
        );

    \I__9992\ : CascadeMux
    port map (
            O => \N__42993\,
            I => \n7_adj_823_cascade_\
        );

    \I__9991\ : IoInMux
    port map (
            O => \N__42990\,
            I => \N__42987\
        );

    \I__9990\ : LocalMux
    port map (
            O => \N__42987\,
            I => \N__42984\
        );

    \I__9989\ : IoSpan4Mux
    port map (
            O => \N__42984\,
            I => \N__42981\
        );

    \I__9988\ : Sp12to4
    port map (
            O => \N__42981\,
            I => \N__42978\
        );

    \I__9987\ : Span12Mux_v
    port map (
            O => \N__42978\,
            I => \N__42974\
        );

    \I__9986\ : InMux
    port map (
            O => \N__42977\,
            I => \N__42971\
        );

    \I__9985\ : Odrv12
    port map (
            O => \N__42974\,
            I => pin_oe_19
        );

    \I__9984\ : LocalMux
    port map (
            O => \N__42971\,
            I => pin_oe_19
        );

    \I__9983\ : IoInMux
    port map (
            O => \N__42966\,
            I => \N__42963\
        );

    \I__9982\ : LocalMux
    port map (
            O => \N__42963\,
            I => \N__42960\
        );

    \I__9981\ : IoSpan4Mux
    port map (
            O => \N__42960\,
            I => \N__42957\
        );

    \I__9980\ : Span4Mux_s3_h
    port map (
            O => \N__42957\,
            I => \N__42954\
        );

    \I__9979\ : Sp12to4
    port map (
            O => \N__42954\,
            I => \N__42951\
        );

    \I__9978\ : Span12Mux_v
    port map (
            O => \N__42951\,
            I => \N__42947\
        );

    \I__9977\ : InMux
    port map (
            O => \N__42950\,
            I => \N__42943\
        );

    \I__9976\ : Span12Mux_h
    port map (
            O => \N__42947\,
            I => \N__42940\
        );

    \I__9975\ : InMux
    port map (
            O => \N__42946\,
            I => \N__42937\
        );

    \I__9974\ : LocalMux
    port map (
            O => \N__42943\,
            I => \N__42934\
        );

    \I__9973\ : Odrv12
    port map (
            O => \N__42940\,
            I => pin_out_7
        );

    \I__9972\ : LocalMux
    port map (
            O => \N__42937\,
            I => pin_out_7
        );

    \I__9971\ : Odrv4
    port map (
            O => \N__42934\,
            I => pin_out_7
        );

    \I__9970\ : IoInMux
    port map (
            O => \N__42927\,
            I => \N__42924\
        );

    \I__9969\ : LocalMux
    port map (
            O => \N__42924\,
            I => \N__42921\
        );

    \I__9968\ : Span4Mux_s3_h
    port map (
            O => \N__42921\,
            I => \N__42918\
        );

    \I__9967\ : Span4Mux_v
    port map (
            O => \N__42918\,
            I => \N__42915\
        );

    \I__9966\ : Span4Mux_v
    port map (
            O => \N__42915\,
            I => \N__42912\
        );

    \I__9965\ : Sp12to4
    port map (
            O => \N__42912\,
            I => \N__42909\
        );

    \I__9964\ : Span12Mux_h
    port map (
            O => \N__42909\,
            I => \N__42904\
        );

    \I__9963\ : InMux
    port map (
            O => \N__42908\,
            I => \N__42899\
        );

    \I__9962\ : InMux
    port map (
            O => \N__42907\,
            I => \N__42899\
        );

    \I__9961\ : Odrv12
    port map (
            O => \N__42904\,
            I => pin_out_6
        );

    \I__9960\ : LocalMux
    port map (
            O => \N__42899\,
            I => pin_out_6
        );

    \I__9959\ : InMux
    port map (
            O => \N__42894\,
            I => \N__42891\
        );

    \I__9958\ : LocalMux
    port map (
            O => \N__42891\,
            I => n13358
        );

    \I__9957\ : InMux
    port map (
            O => \N__42888\,
            I => \N__42884\
        );

    \I__9956\ : InMux
    port map (
            O => \N__42887\,
            I => \N__42881\
        );

    \I__9955\ : LocalMux
    port map (
            O => \N__42884\,
            I => \N__42869\
        );

    \I__9954\ : LocalMux
    port map (
            O => \N__42881\,
            I => \N__42869\
        );

    \I__9953\ : InMux
    port map (
            O => \N__42880\,
            I => \N__42862\
        );

    \I__9952\ : InMux
    port map (
            O => \N__42879\,
            I => \N__42862\
        );

    \I__9951\ : InMux
    port map (
            O => \N__42878\,
            I => \N__42862\
        );

    \I__9950\ : InMux
    port map (
            O => \N__42877\,
            I => \N__42853\
        );

    \I__9949\ : InMux
    port map (
            O => \N__42876\,
            I => \N__42853\
        );

    \I__9948\ : InMux
    port map (
            O => \N__42875\,
            I => \N__42853\
        );

    \I__9947\ : InMux
    port map (
            O => \N__42874\,
            I => \N__42853\
        );

    \I__9946\ : Span4Mux_v
    port map (
            O => \N__42869\,
            I => \N__42850\
        );

    \I__9945\ : LocalMux
    port map (
            O => \N__42862\,
            I => n3762
        );

    \I__9944\ : LocalMux
    port map (
            O => \N__42853\,
            I => n3762
        );

    \I__9943\ : Odrv4
    port map (
            O => \N__42850\,
            I => n3762
        );

    \I__9942\ : InMux
    port map (
            O => \N__42843\,
            I => \N__42840\
        );

    \I__9941\ : LocalMux
    port map (
            O => \N__42840\,
            I => \N__42837\
        );

    \I__9940\ : Odrv4
    port map (
            O => \N__42837\,
            I => n11964
        );

    \I__9939\ : IoInMux
    port map (
            O => \N__42834\,
            I => \N__42831\
        );

    \I__9938\ : LocalMux
    port map (
            O => \N__42831\,
            I => \N__42828\
        );

    \I__9937\ : IoSpan4Mux
    port map (
            O => \N__42828\,
            I => \N__42825\
        );

    \I__9936\ : Span4Mux_s0_h
    port map (
            O => \N__42825\,
            I => \N__42822\
        );

    \I__9935\ : Sp12to4
    port map (
            O => \N__42822\,
            I => \N__42819\
        );

    \I__9934\ : Span12Mux_h
    port map (
            O => \N__42819\,
            I => \N__42815\
        );

    \I__9933\ : InMux
    port map (
            O => \N__42818\,
            I => \N__42812\
        );

    \I__9932\ : Odrv12
    port map (
            O => \N__42815\,
            I => pin_oe_16
        );

    \I__9931\ : LocalMux
    port map (
            O => \N__42812\,
            I => pin_oe_16
        );

    \I__9930\ : InMux
    port map (
            O => \N__42807\,
            I => \N__42804\
        );

    \I__9929\ : LocalMux
    port map (
            O => \N__42804\,
            I => n11820
        );

    \I__9928\ : CascadeMux
    port map (
            O => \N__42801\,
            I => \N__42798\
        );

    \I__9927\ : InMux
    port map (
            O => \N__42798\,
            I => \N__42794\
        );

    \I__9926\ : InMux
    port map (
            O => \N__42797\,
            I => \N__42791\
        );

    \I__9925\ : LocalMux
    port map (
            O => \N__42794\,
            I => counter_7
        );

    \I__9924\ : LocalMux
    port map (
            O => \N__42791\,
            I => counter_7
        );

    \I__9923\ : InMux
    port map (
            O => \N__42786\,
            I => \N__42782\
        );

    \I__9922\ : InMux
    port map (
            O => \N__42785\,
            I => \N__42779\
        );

    \I__9921\ : LocalMux
    port map (
            O => \N__42782\,
            I => \N__42776\
        );

    \I__9920\ : LocalMux
    port map (
            O => \N__42779\,
            I => counter_0
        );

    \I__9919\ : Odrv4
    port map (
            O => \N__42776\,
            I => counter_0
        );

    \I__9918\ : CascadeMux
    port map (
            O => \N__42771\,
            I => \N__42768\
        );

    \I__9917\ : InMux
    port map (
            O => \N__42768\,
            I => \N__42764\
        );

    \I__9916\ : InMux
    port map (
            O => \N__42767\,
            I => \N__42761\
        );

    \I__9915\ : LocalMux
    port map (
            O => \N__42764\,
            I => counter_6
        );

    \I__9914\ : LocalMux
    port map (
            O => \N__42761\,
            I => counter_6
        );

    \I__9913\ : InMux
    port map (
            O => \N__42756\,
            I => \N__42752\
        );

    \I__9912\ : InMux
    port map (
            O => \N__42755\,
            I => \N__42749\
        );

    \I__9911\ : LocalMux
    port map (
            O => \N__42752\,
            I => counter_1
        );

    \I__9910\ : LocalMux
    port map (
            O => \N__42749\,
            I => counter_1
        );

    \I__9909\ : CascadeMux
    port map (
            O => \N__42744\,
            I => \n10_cascade_\
        );

    \I__9908\ : CascadeMux
    port map (
            O => \N__42741\,
            I => \n9_adj_824_cascade_\
        );

    \I__9907\ : CascadeMux
    port map (
            O => \N__42738\,
            I => \n8_adj_822_cascade_\
        );

    \I__9906\ : IoInMux
    port map (
            O => \N__42735\,
            I => \N__42732\
        );

    \I__9905\ : LocalMux
    port map (
            O => \N__42732\,
            I => \N__42729\
        );

    \I__9904\ : Span12Mux_s5_h
    port map (
            O => \N__42729\,
            I => \N__42725\
        );

    \I__9903\ : InMux
    port map (
            O => \N__42728\,
            I => \N__42721\
        );

    \I__9902\ : Span12Mux_v
    port map (
            O => \N__42725\,
            I => \N__42718\
        );

    \I__9901\ : InMux
    port map (
            O => \N__42724\,
            I => \N__42715\
        );

    \I__9900\ : LocalMux
    port map (
            O => \N__42721\,
            I => \N__42712\
        );

    \I__9899\ : Odrv12
    port map (
            O => \N__42718\,
            I => pin_out_5
        );

    \I__9898\ : LocalMux
    port map (
            O => \N__42715\,
            I => pin_out_5
        );

    \I__9897\ : Odrv4
    port map (
            O => \N__42712\,
            I => pin_out_5
        );

    \I__9896\ : IoInMux
    port map (
            O => \N__42705\,
            I => \N__42702\
        );

    \I__9895\ : LocalMux
    port map (
            O => \N__42702\,
            I => \N__42699\
        );

    \I__9894\ : Span12Mux_s4_h
    port map (
            O => \N__42699\,
            I => \N__42695\
        );

    \I__9893\ : InMux
    port map (
            O => \N__42698\,
            I => \N__42691\
        );

    \I__9892\ : Span12Mux_v
    port map (
            O => \N__42695\,
            I => \N__42688\
        );

    \I__9891\ : InMux
    port map (
            O => \N__42694\,
            I => \N__42685\
        );

    \I__9890\ : LocalMux
    port map (
            O => \N__42691\,
            I => \N__42682\
        );

    \I__9889\ : Odrv12
    port map (
            O => \N__42688\,
            I => pin_out_4
        );

    \I__9888\ : LocalMux
    port map (
            O => \N__42685\,
            I => pin_out_4
        );

    \I__9887\ : Odrv4
    port map (
            O => \N__42682\,
            I => pin_out_4
        );

    \I__9886\ : CascadeMux
    port map (
            O => \N__42675\,
            I => \n13357_cascade_\
        );

    \I__9885\ : InMux
    port map (
            O => \N__42672\,
            I => \N__42669\
        );

    \I__9884\ : LocalMux
    port map (
            O => \N__42669\,
            I => n13625
        );

    \I__9883\ : CascadeMux
    port map (
            O => \N__42666\,
            I => \n6_adj_810_cascade_\
        );

    \I__9882\ : InMux
    port map (
            O => \N__42663\,
            I => \N__42660\
        );

    \I__9881\ : LocalMux
    port map (
            O => \N__42660\,
            I => \N__42657\
        );

    \I__9880\ : Span4Mux_h
    port map (
            O => \N__42657\,
            I => \N__42654\
        );

    \I__9879\ : Span4Mux_v
    port map (
            O => \N__42654\,
            I => \N__42651\
        );

    \I__9878\ : Odrv4
    port map (
            O => \N__42651\,
            I => n11874
        );

    \I__9877\ : CascadeMux
    port map (
            O => \N__42648\,
            I => \N__42645\
        );

    \I__9876\ : InMux
    port map (
            O => \N__42645\,
            I => \N__42642\
        );

    \I__9875\ : LocalMux
    port map (
            O => \N__42642\,
            I => n11823
        );

    \I__9874\ : InMux
    port map (
            O => \N__42639\,
            I => \N__42636\
        );

    \I__9873\ : LocalMux
    port map (
            O => \N__42636\,
            I => \N__42632\
        );

    \I__9872\ : InMux
    port map (
            O => \N__42635\,
            I => \N__42629\
        );

    \I__9871\ : Span4Mux_s3_h
    port map (
            O => \N__42632\,
            I => \N__42622\
        );

    \I__9870\ : LocalMux
    port map (
            O => \N__42629\,
            I => \N__42622\
        );

    \I__9869\ : InMux
    port map (
            O => \N__42628\,
            I => \N__42619\
        );

    \I__9868\ : InMux
    port map (
            O => \N__42627\,
            I => \N__42616\
        );

    \I__9867\ : Span4Mux_v
    port map (
            O => \N__42622\,
            I => \N__42610\
        );

    \I__9866\ : LocalMux
    port map (
            O => \N__42619\,
            I => \N__42605\
        );

    \I__9865\ : LocalMux
    port map (
            O => \N__42616\,
            I => \N__42605\
        );

    \I__9864\ : InMux
    port map (
            O => \N__42615\,
            I => \N__42600\
        );

    \I__9863\ : InMux
    port map (
            O => \N__42614\,
            I => \N__42595\
        );

    \I__9862\ : InMux
    port map (
            O => \N__42613\,
            I => \N__42595\
        );

    \I__9861\ : Span4Mux_h
    port map (
            O => \N__42610\,
            I => \N__42592\
        );

    \I__9860\ : Span4Mux_v
    port map (
            O => \N__42605\,
            I => \N__42589\
        );

    \I__9859\ : InMux
    port map (
            O => \N__42604\,
            I => \N__42584\
        );

    \I__9858\ : InMux
    port map (
            O => \N__42603\,
            I => \N__42579\
        );

    \I__9857\ : LocalMux
    port map (
            O => \N__42600\,
            I => \N__42575\
        );

    \I__9856\ : LocalMux
    port map (
            O => \N__42595\,
            I => \N__42572\
        );

    \I__9855\ : Span4Mux_h
    port map (
            O => \N__42592\,
            I => \N__42569\
        );

    \I__9854\ : Span4Mux_h
    port map (
            O => \N__42589\,
            I => \N__42566\
        );

    \I__9853\ : InMux
    port map (
            O => \N__42588\,
            I => \N__42561\
        );

    \I__9852\ : InMux
    port map (
            O => \N__42587\,
            I => \N__42561\
        );

    \I__9851\ : LocalMux
    port map (
            O => \N__42584\,
            I => \N__42558\
        );

    \I__9850\ : InMux
    port map (
            O => \N__42583\,
            I => \N__42553\
        );

    \I__9849\ : InMux
    port map (
            O => \N__42582\,
            I => \N__42553\
        );

    \I__9848\ : LocalMux
    port map (
            O => \N__42579\,
            I => \N__42550\
        );

    \I__9847\ : InMux
    port map (
            O => \N__42578\,
            I => \N__42547\
        );

    \I__9846\ : Span4Mux_v
    port map (
            O => \N__42575\,
            I => \N__42542\
        );

    \I__9845\ : Span4Mux_v
    port map (
            O => \N__42572\,
            I => \N__42542\
        );

    \I__9844\ : Span4Mux_h
    port map (
            O => \N__42569\,
            I => \N__42539\
        );

    \I__9843\ : Span4Mux_h
    port map (
            O => \N__42566\,
            I => \N__42536\
        );

    \I__9842\ : LocalMux
    port map (
            O => \N__42561\,
            I => n7
        );

    \I__9841\ : Odrv12
    port map (
            O => \N__42558\,
            I => n7
        );

    \I__9840\ : LocalMux
    port map (
            O => \N__42553\,
            I => n7
        );

    \I__9839\ : Odrv4
    port map (
            O => \N__42550\,
            I => n7
        );

    \I__9838\ : LocalMux
    port map (
            O => \N__42547\,
            I => n7
        );

    \I__9837\ : Odrv4
    port map (
            O => \N__42542\,
            I => n7
        );

    \I__9836\ : Odrv4
    port map (
            O => \N__42539\,
            I => n7
        );

    \I__9835\ : Odrv4
    port map (
            O => \N__42536\,
            I => n7
        );

    \I__9834\ : InMux
    port map (
            O => \N__42519\,
            I => n10576
        );

    \I__9833\ : InMux
    port map (
            O => \N__42516\,
            I => n10577
        );

    \I__9832\ : InMux
    port map (
            O => \N__42513\,
            I => n10578
        );

    \I__9831\ : InMux
    port map (
            O => \N__42510\,
            I => \N__42506\
        );

    \I__9830\ : InMux
    port map (
            O => \N__42509\,
            I => \N__42503\
        );

    \I__9829\ : LocalMux
    port map (
            O => \N__42506\,
            I => current_pin_5
        );

    \I__9828\ : LocalMux
    port map (
            O => \N__42503\,
            I => current_pin_5
        );

    \I__9827\ : InMux
    port map (
            O => \N__42498\,
            I => n10579
        );

    \I__9826\ : InMux
    port map (
            O => \N__42495\,
            I => \N__42491\
        );

    \I__9825\ : InMux
    port map (
            O => \N__42494\,
            I => \N__42488\
        );

    \I__9824\ : LocalMux
    port map (
            O => \N__42491\,
            I => current_pin_6
        );

    \I__9823\ : LocalMux
    port map (
            O => \N__42488\,
            I => current_pin_6
        );

    \I__9822\ : InMux
    port map (
            O => \N__42483\,
            I => n10580
        );

    \I__9821\ : InMux
    port map (
            O => \N__42480\,
            I => n10581
        );

    \I__9820\ : InMux
    port map (
            O => \N__42477\,
            I => \N__42473\
        );

    \I__9819\ : InMux
    port map (
            O => \N__42476\,
            I => \N__42470\
        );

    \I__9818\ : LocalMux
    port map (
            O => \N__42473\,
            I => current_pin_7
        );

    \I__9817\ : LocalMux
    port map (
            O => \N__42470\,
            I => current_pin_7
        );

    \I__9816\ : SRMux
    port map (
            O => \N__42465\,
            I => \N__42462\
        );

    \I__9815\ : LocalMux
    port map (
            O => \N__42462\,
            I => \N__42459\
        );

    \I__9814\ : Odrv4
    port map (
            O => \N__42459\,
            I => n7985
        );

    \I__9813\ : CEMux
    port map (
            O => \N__42456\,
            I => \N__42452\
        );

    \I__9812\ : InMux
    port map (
            O => \N__42455\,
            I => \N__42449\
        );

    \I__9811\ : LocalMux
    port map (
            O => \N__42452\,
            I => n7635
        );

    \I__9810\ : LocalMux
    port map (
            O => \N__42449\,
            I => n7635
        );

    \I__9809\ : InMux
    port map (
            O => \N__42444\,
            I => n10703
        );

    \I__9808\ : InMux
    port map (
            O => \N__42441\,
            I => n10704
        );

    \I__9807\ : InMux
    port map (
            O => \N__42438\,
            I => n10705
        );

    \I__9806\ : CascadeMux
    port map (
            O => \N__42435\,
            I => \N__42428\
        );

    \I__9805\ : CascadeMux
    port map (
            O => \N__42434\,
            I => \N__42424\
        );

    \I__9804\ : CascadeMux
    port map (
            O => \N__42433\,
            I => \N__42420\
        );

    \I__9803\ : InMux
    port map (
            O => \N__42432\,
            I => \N__42405\
        );

    \I__9802\ : InMux
    port map (
            O => \N__42431\,
            I => \N__42405\
        );

    \I__9801\ : InMux
    port map (
            O => \N__42428\,
            I => \N__42405\
        );

    \I__9800\ : InMux
    port map (
            O => \N__42427\,
            I => \N__42405\
        );

    \I__9799\ : InMux
    port map (
            O => \N__42424\,
            I => \N__42405\
        );

    \I__9798\ : InMux
    port map (
            O => \N__42423\,
            I => \N__42405\
        );

    \I__9797\ : InMux
    port map (
            O => \N__42420\,
            I => \N__42405\
        );

    \I__9796\ : LocalMux
    port map (
            O => \N__42405\,
            I => n13603
        );

    \I__9795\ : InMux
    port map (
            O => \N__42402\,
            I => n10706
        );

    \I__9794\ : CEMux
    port map (
            O => \N__42399\,
            I => \N__42395\
        );

    \I__9793\ : CEMux
    port map (
            O => \N__42398\,
            I => \N__42392\
        );

    \I__9792\ : LocalMux
    port map (
            O => \N__42395\,
            I => \N__42387\
        );

    \I__9791\ : LocalMux
    port map (
            O => \N__42392\,
            I => \N__42387\
        );

    \I__9790\ : Span4Mux_v
    port map (
            O => \N__42387\,
            I => \N__42384\
        );

    \I__9789\ : Odrv4
    port map (
            O => \N__42384\,
            I => n7681
        );

    \I__9788\ : InMux
    port map (
            O => \N__42381\,
            I => \N__42378\
        );

    \I__9787\ : LocalMux
    port map (
            O => \N__42378\,
            I => \N__42375\
        );

    \I__9786\ : Span4Mux_h
    port map (
            O => \N__42375\,
            I => \N__42372\
        );

    \I__9785\ : Odrv4
    port map (
            O => \N__42372\,
            I => n11824
        );

    \I__9784\ : InMux
    port map (
            O => \N__42369\,
            I => \bfn_17_17_0_\
        );

    \I__9783\ : InMux
    port map (
            O => \N__42366\,
            I => n10575
        );

    \I__9782\ : CascadeMux
    port map (
            O => \N__42363\,
            I => \N__42359\
        );

    \I__9781\ : CascadeMux
    port map (
            O => \N__42362\,
            I => \N__42356\
        );

    \I__9780\ : InMux
    port map (
            O => \N__42359\,
            I => \N__42353\
        );

    \I__9779\ : InMux
    port map (
            O => \N__42356\,
            I => \N__42350\
        );

    \I__9778\ : LocalMux
    port map (
            O => \N__42353\,
            I => \nx.n2491\
        );

    \I__9777\ : LocalMux
    port map (
            O => \N__42350\,
            I => \nx.n2491\
        );

    \I__9776\ : InMux
    port map (
            O => \N__42345\,
            I => \N__42342\
        );

    \I__9775\ : LocalMux
    port map (
            O => \N__42342\,
            I => \nx.n2558\
        );

    \I__9774\ : InMux
    port map (
            O => \N__42339\,
            I => \nx.n10956\
        );

    \I__9773\ : CascadeMux
    port map (
            O => \N__42336\,
            I => \N__42333\
        );

    \I__9772\ : InMux
    port map (
            O => \N__42333\,
            I => \N__42329\
        );

    \I__9771\ : CascadeMux
    port map (
            O => \N__42332\,
            I => \N__42326\
        );

    \I__9770\ : LocalMux
    port map (
            O => \N__42329\,
            I => \N__42323\
        );

    \I__9769\ : InMux
    port map (
            O => \N__42326\,
            I => \N__42320\
        );

    \I__9768\ : Span4Mux_v
    port map (
            O => \N__42323\,
            I => \N__42317\
        );

    \I__9767\ : LocalMux
    port map (
            O => \N__42320\,
            I => \nx.n2490\
        );

    \I__9766\ : Odrv4
    port map (
            O => \N__42317\,
            I => \nx.n2490\
        );

    \I__9765\ : InMux
    port map (
            O => \N__42312\,
            I => \N__42309\
        );

    \I__9764\ : LocalMux
    port map (
            O => \N__42309\,
            I => \N__42306\
        );

    \I__9763\ : Odrv4
    port map (
            O => \N__42306\,
            I => \nx.n2557\
        );

    \I__9762\ : InMux
    port map (
            O => \N__42303\,
            I => \nx.n10957\
        );

    \I__9761\ : CascadeMux
    port map (
            O => \N__42300\,
            I => \N__42290\
        );

    \I__9760\ : CascadeMux
    port map (
            O => \N__42299\,
            I => \N__42284\
        );

    \I__9759\ : CascadeMux
    port map (
            O => \N__42298\,
            I => \N__42276\
        );

    \I__9758\ : CascadeMux
    port map (
            O => \N__42297\,
            I => \N__42271\
        );

    \I__9757\ : CascadeMux
    port map (
            O => \N__42296\,
            I => \N__42264\
        );

    \I__9756\ : CascadeMux
    port map (
            O => \N__42295\,
            I => \N__42259\
        );

    \I__9755\ : InMux
    port map (
            O => \N__42294\,
            I => \N__42244\
        );

    \I__9754\ : InMux
    port map (
            O => \N__42293\,
            I => \N__42244\
        );

    \I__9753\ : InMux
    port map (
            O => \N__42290\,
            I => \N__42244\
        );

    \I__9752\ : InMux
    port map (
            O => \N__42289\,
            I => \N__42239\
        );

    \I__9751\ : InMux
    port map (
            O => \N__42288\,
            I => \N__42239\
        );

    \I__9750\ : InMux
    port map (
            O => \N__42287\,
            I => \N__42230\
        );

    \I__9749\ : InMux
    port map (
            O => \N__42284\,
            I => \N__42230\
        );

    \I__9748\ : InMux
    port map (
            O => \N__42283\,
            I => \N__42230\
        );

    \I__9747\ : InMux
    port map (
            O => \N__42282\,
            I => \N__42230\
        );

    \I__9746\ : CascadeMux
    port map (
            O => \N__42281\,
            I => \N__42226\
        );

    \I__9745\ : InMux
    port map (
            O => \N__42280\,
            I => \N__42188\
        );

    \I__9744\ : InMux
    port map (
            O => \N__42279\,
            I => \N__42188\
        );

    \I__9743\ : InMux
    port map (
            O => \N__42276\,
            I => \N__42176\
        );

    \I__9742\ : InMux
    port map (
            O => \N__42275\,
            I => \N__42176\
        );

    \I__9741\ : InMux
    port map (
            O => \N__42274\,
            I => \N__42176\
        );

    \I__9740\ : InMux
    port map (
            O => \N__42271\,
            I => \N__42176\
        );

    \I__9739\ : InMux
    port map (
            O => \N__42270\,
            I => \N__42176\
        );

    \I__9738\ : InMux
    port map (
            O => \N__42269\,
            I => \N__42163\
        );

    \I__9737\ : InMux
    port map (
            O => \N__42268\,
            I => \N__42163\
        );

    \I__9736\ : InMux
    port map (
            O => \N__42267\,
            I => \N__42154\
        );

    \I__9735\ : InMux
    port map (
            O => \N__42264\,
            I => \N__42154\
        );

    \I__9734\ : InMux
    port map (
            O => \N__42263\,
            I => \N__42154\
        );

    \I__9733\ : InMux
    port map (
            O => \N__42262\,
            I => \N__42154\
        );

    \I__9732\ : InMux
    port map (
            O => \N__42259\,
            I => \N__42145\
        );

    \I__9731\ : InMux
    port map (
            O => \N__42258\,
            I => \N__42145\
        );

    \I__9730\ : InMux
    port map (
            O => \N__42257\,
            I => \N__42145\
        );

    \I__9729\ : InMux
    port map (
            O => \N__42256\,
            I => \N__42145\
        );

    \I__9728\ : InMux
    port map (
            O => \N__42255\,
            I => \N__42142\
        );

    \I__9727\ : InMux
    port map (
            O => \N__42254\,
            I => \N__42129\
        );

    \I__9726\ : InMux
    port map (
            O => \N__42253\,
            I => \N__42129\
        );

    \I__9725\ : InMux
    port map (
            O => \N__42252\,
            I => \N__42129\
        );

    \I__9724\ : InMux
    port map (
            O => \N__42251\,
            I => \N__42129\
        );

    \I__9723\ : LocalMux
    port map (
            O => \N__42244\,
            I => \N__42113\
        );

    \I__9722\ : LocalMux
    port map (
            O => \N__42239\,
            I => \N__42113\
        );

    \I__9721\ : LocalMux
    port map (
            O => \N__42230\,
            I => \N__42113\
        );

    \I__9720\ : InMux
    port map (
            O => \N__42229\,
            I => \N__42110\
        );

    \I__9719\ : InMux
    port map (
            O => \N__42226\,
            I => \N__42105\
        );

    \I__9718\ : InMux
    port map (
            O => \N__42225\,
            I => \N__42105\
        );

    \I__9717\ : InMux
    port map (
            O => \N__42224\,
            I => \N__42102\
        );

    \I__9716\ : InMux
    port map (
            O => \N__42223\,
            I => \N__42099\
        );

    \I__9715\ : InMux
    port map (
            O => \N__42222\,
            I => \N__42077\
        );

    \I__9714\ : InMux
    port map (
            O => \N__42221\,
            I => \N__42077\
        );

    \I__9713\ : InMux
    port map (
            O => \N__42220\,
            I => \N__42077\
        );

    \I__9712\ : InMux
    port map (
            O => \N__42219\,
            I => \N__42077\
        );

    \I__9711\ : InMux
    port map (
            O => \N__42218\,
            I => \N__42072\
        );

    \I__9710\ : InMux
    port map (
            O => \N__42217\,
            I => \N__42072\
        );

    \I__9709\ : InMux
    port map (
            O => \N__42216\,
            I => \N__42068\
        );

    \I__9708\ : InMux
    port map (
            O => \N__42215\,
            I => \N__42044\
        );

    \I__9707\ : InMux
    port map (
            O => \N__42214\,
            I => \N__42034\
        );

    \I__9706\ : InMux
    port map (
            O => \N__42213\,
            I => \N__42034\
        );

    \I__9705\ : InMux
    port map (
            O => \N__42212\,
            I => \N__42034\
        );

    \I__9704\ : CascadeMux
    port map (
            O => \N__42211\,
            I => \N__42027\
        );

    \I__9703\ : CascadeMux
    port map (
            O => \N__42210\,
            I => \N__42016\
        );

    \I__9702\ : CascadeMux
    port map (
            O => \N__42209\,
            I => \N__42006\
        );

    \I__9701\ : InMux
    port map (
            O => \N__42208\,
            I => \N__41988\
        );

    \I__9700\ : InMux
    port map (
            O => \N__42207\,
            I => \N__41988\
        );

    \I__9699\ : InMux
    port map (
            O => \N__42206\,
            I => \N__41988\
        );

    \I__9698\ : InMux
    port map (
            O => \N__42205\,
            I => \N__41988\
        );

    \I__9697\ : InMux
    port map (
            O => \N__42204\,
            I => \N__41979\
        );

    \I__9696\ : InMux
    port map (
            O => \N__42203\,
            I => \N__41979\
        );

    \I__9695\ : InMux
    port map (
            O => \N__42202\,
            I => \N__41979\
        );

    \I__9694\ : InMux
    port map (
            O => \N__42201\,
            I => \N__41979\
        );

    \I__9693\ : InMux
    port map (
            O => \N__42200\,
            I => \N__41969\
        );

    \I__9692\ : InMux
    port map (
            O => \N__42199\,
            I => \N__41969\
        );

    \I__9691\ : InMux
    port map (
            O => \N__42198\,
            I => \N__41960\
        );

    \I__9690\ : InMux
    port map (
            O => \N__42197\,
            I => \N__41953\
        );

    \I__9689\ : InMux
    port map (
            O => \N__42196\,
            I => \N__41953\
        );

    \I__9688\ : InMux
    port map (
            O => \N__42195\,
            I => \N__41953\
        );

    \I__9687\ : InMux
    port map (
            O => \N__42194\,
            I => \N__41948\
        );

    \I__9686\ : InMux
    port map (
            O => \N__42193\,
            I => \N__41948\
        );

    \I__9685\ : LocalMux
    port map (
            O => \N__42188\,
            I => \N__41945\
        );

    \I__9684\ : CascadeMux
    port map (
            O => \N__42187\,
            I => \N__41940\
        );

    \I__9683\ : LocalMux
    port map (
            O => \N__42176\,
            I => \N__41932\
        );

    \I__9682\ : InMux
    port map (
            O => \N__42175\,
            I => \N__41923\
        );

    \I__9681\ : InMux
    port map (
            O => \N__42174\,
            I => \N__41923\
        );

    \I__9680\ : InMux
    port map (
            O => \N__42173\,
            I => \N__41923\
        );

    \I__9679\ : InMux
    port map (
            O => \N__42172\,
            I => \N__41923\
        );

    \I__9678\ : InMux
    port map (
            O => \N__42171\,
            I => \N__41914\
        );

    \I__9677\ : InMux
    port map (
            O => \N__42170\,
            I => \N__41914\
        );

    \I__9676\ : InMux
    port map (
            O => \N__42169\,
            I => \N__41914\
        );

    \I__9675\ : InMux
    port map (
            O => \N__42168\,
            I => \N__41914\
        );

    \I__9674\ : LocalMux
    port map (
            O => \N__42163\,
            I => \N__41905\
        );

    \I__9673\ : LocalMux
    port map (
            O => \N__42154\,
            I => \N__41905\
        );

    \I__9672\ : LocalMux
    port map (
            O => \N__42145\,
            I => \N__41905\
        );

    \I__9671\ : LocalMux
    port map (
            O => \N__42142\,
            I => \N__41905\
        );

    \I__9670\ : InMux
    port map (
            O => \N__42141\,
            I => \N__41896\
        );

    \I__9669\ : InMux
    port map (
            O => \N__42140\,
            I => \N__41896\
        );

    \I__9668\ : InMux
    port map (
            O => \N__42139\,
            I => \N__41896\
        );

    \I__9667\ : InMux
    port map (
            O => \N__42138\,
            I => \N__41896\
        );

    \I__9666\ : LocalMux
    port map (
            O => \N__42129\,
            I => \N__41893\
        );

    \I__9665\ : InMux
    port map (
            O => \N__42128\,
            I => \N__41886\
        );

    \I__9664\ : InMux
    port map (
            O => \N__42127\,
            I => \N__41886\
        );

    \I__9663\ : InMux
    port map (
            O => \N__42126\,
            I => \N__41886\
        );

    \I__9662\ : InMux
    port map (
            O => \N__42125\,
            I => \N__41879\
        );

    \I__9661\ : InMux
    port map (
            O => \N__42124\,
            I => \N__41879\
        );

    \I__9660\ : InMux
    port map (
            O => \N__42123\,
            I => \N__41879\
        );

    \I__9659\ : CascadeMux
    port map (
            O => \N__42122\,
            I => \N__41876\
        );

    \I__9658\ : CascadeMux
    port map (
            O => \N__42121\,
            I => \N__41872\
        );

    \I__9657\ : CascadeMux
    port map (
            O => \N__42120\,
            I => \N__41869\
        );

    \I__9656\ : Span4Mux_v
    port map (
            O => \N__42113\,
            I => \N__41855\
        );

    \I__9655\ : LocalMux
    port map (
            O => \N__42110\,
            I => \N__41855\
        );

    \I__9654\ : LocalMux
    port map (
            O => \N__42105\,
            I => \N__41855\
        );

    \I__9653\ : LocalMux
    port map (
            O => \N__42102\,
            I => \N__41850\
        );

    \I__9652\ : LocalMux
    port map (
            O => \N__42099\,
            I => \N__41850\
        );

    \I__9651\ : InMux
    port map (
            O => \N__42098\,
            I => \N__41843\
        );

    \I__9650\ : InMux
    port map (
            O => \N__42097\,
            I => \N__41843\
        );

    \I__9649\ : InMux
    port map (
            O => \N__42096\,
            I => \N__41843\
        );

    \I__9648\ : InMux
    port map (
            O => \N__42095\,
            I => \N__41836\
        );

    \I__9647\ : InMux
    port map (
            O => \N__42094\,
            I => \N__41836\
        );

    \I__9646\ : InMux
    port map (
            O => \N__42093\,
            I => \N__41836\
        );

    \I__9645\ : InMux
    port map (
            O => \N__42092\,
            I => \N__41827\
        );

    \I__9644\ : InMux
    port map (
            O => \N__42091\,
            I => \N__41827\
        );

    \I__9643\ : InMux
    port map (
            O => \N__42090\,
            I => \N__41827\
        );

    \I__9642\ : InMux
    port map (
            O => \N__42089\,
            I => \N__41827\
        );

    \I__9641\ : InMux
    port map (
            O => \N__42088\,
            I => \N__41820\
        );

    \I__9640\ : InMux
    port map (
            O => \N__42087\,
            I => \N__41820\
        );

    \I__9639\ : InMux
    port map (
            O => \N__42086\,
            I => \N__41820\
        );

    \I__9638\ : LocalMux
    port map (
            O => \N__42077\,
            I => \N__41815\
        );

    \I__9637\ : LocalMux
    port map (
            O => \N__42072\,
            I => \N__41815\
        );

    \I__9636\ : CascadeMux
    port map (
            O => \N__42071\,
            I => \N__41807\
        );

    \I__9635\ : LocalMux
    port map (
            O => \N__42068\,
            I => \N__41802\
        );

    \I__9634\ : InMux
    port map (
            O => \N__42067\,
            I => \N__41793\
        );

    \I__9633\ : InMux
    port map (
            O => \N__42066\,
            I => \N__41793\
        );

    \I__9632\ : InMux
    port map (
            O => \N__42065\,
            I => \N__41793\
        );

    \I__9631\ : InMux
    port map (
            O => \N__42064\,
            I => \N__41793\
        );

    \I__9630\ : InMux
    port map (
            O => \N__42063\,
            I => \N__41786\
        );

    \I__9629\ : InMux
    port map (
            O => \N__42062\,
            I => \N__41786\
        );

    \I__9628\ : InMux
    port map (
            O => \N__42061\,
            I => \N__41786\
        );

    \I__9627\ : InMux
    port map (
            O => \N__42060\,
            I => \N__41783\
        );

    \I__9626\ : InMux
    port map (
            O => \N__42059\,
            I => \N__41772\
        );

    \I__9625\ : InMux
    port map (
            O => \N__42058\,
            I => \N__41772\
        );

    \I__9624\ : InMux
    port map (
            O => \N__42057\,
            I => \N__41772\
        );

    \I__9623\ : InMux
    port map (
            O => \N__42056\,
            I => \N__41772\
        );

    \I__9622\ : InMux
    port map (
            O => \N__42055\,
            I => \N__41772\
        );

    \I__9621\ : InMux
    port map (
            O => \N__42054\,
            I => \N__41763\
        );

    \I__9620\ : InMux
    port map (
            O => \N__42053\,
            I => \N__41763\
        );

    \I__9619\ : InMux
    port map (
            O => \N__42052\,
            I => \N__41763\
        );

    \I__9618\ : InMux
    port map (
            O => \N__42051\,
            I => \N__41763\
        );

    \I__9617\ : InMux
    port map (
            O => \N__42050\,
            I => \N__41754\
        );

    \I__9616\ : InMux
    port map (
            O => \N__42049\,
            I => \N__41754\
        );

    \I__9615\ : InMux
    port map (
            O => \N__42048\,
            I => \N__41754\
        );

    \I__9614\ : InMux
    port map (
            O => \N__42047\,
            I => \N__41754\
        );

    \I__9613\ : LocalMux
    port map (
            O => \N__42044\,
            I => \N__41739\
        );

    \I__9612\ : InMux
    port map (
            O => \N__42043\,
            I => \N__41732\
        );

    \I__9611\ : InMux
    port map (
            O => \N__42042\,
            I => \N__41732\
        );

    \I__9610\ : InMux
    port map (
            O => \N__42041\,
            I => \N__41732\
        );

    \I__9609\ : LocalMux
    port map (
            O => \N__42034\,
            I => \N__41729\
        );

    \I__9608\ : InMux
    port map (
            O => \N__42033\,
            I => \N__41724\
        );

    \I__9607\ : InMux
    port map (
            O => \N__42032\,
            I => \N__41724\
        );

    \I__9606\ : InMux
    port map (
            O => \N__42031\,
            I => \N__41713\
        );

    \I__9605\ : InMux
    port map (
            O => \N__42030\,
            I => \N__41713\
        );

    \I__9604\ : InMux
    port map (
            O => \N__42027\,
            I => \N__41713\
        );

    \I__9603\ : InMux
    port map (
            O => \N__42026\,
            I => \N__41713\
        );

    \I__9602\ : InMux
    port map (
            O => \N__42025\,
            I => \N__41713\
        );

    \I__9601\ : InMux
    port map (
            O => \N__42024\,
            I => \N__41704\
        );

    \I__9600\ : InMux
    port map (
            O => \N__42023\,
            I => \N__41704\
        );

    \I__9599\ : InMux
    port map (
            O => \N__42022\,
            I => \N__41704\
        );

    \I__9598\ : InMux
    port map (
            O => \N__42021\,
            I => \N__41704\
        );

    \I__9597\ : InMux
    port map (
            O => \N__42020\,
            I => \N__41695\
        );

    \I__9596\ : InMux
    port map (
            O => \N__42019\,
            I => \N__41695\
        );

    \I__9595\ : InMux
    port map (
            O => \N__42016\,
            I => \N__41695\
        );

    \I__9594\ : InMux
    port map (
            O => \N__42015\,
            I => \N__41695\
        );

    \I__9593\ : InMux
    port map (
            O => \N__42014\,
            I => \N__41688\
        );

    \I__9592\ : InMux
    port map (
            O => \N__42013\,
            I => \N__41688\
        );

    \I__9591\ : InMux
    port map (
            O => \N__42012\,
            I => \N__41688\
        );

    \I__9590\ : InMux
    port map (
            O => \N__42011\,
            I => \N__41681\
        );

    \I__9589\ : InMux
    port map (
            O => \N__42010\,
            I => \N__41681\
        );

    \I__9588\ : InMux
    port map (
            O => \N__42009\,
            I => \N__41681\
        );

    \I__9587\ : InMux
    port map (
            O => \N__42006\,
            I => \N__41672\
        );

    \I__9586\ : InMux
    port map (
            O => \N__42005\,
            I => \N__41672\
        );

    \I__9585\ : InMux
    port map (
            O => \N__42004\,
            I => \N__41672\
        );

    \I__9584\ : InMux
    port map (
            O => \N__42003\,
            I => \N__41663\
        );

    \I__9583\ : InMux
    port map (
            O => \N__42002\,
            I => \N__41663\
        );

    \I__9582\ : InMux
    port map (
            O => \N__42001\,
            I => \N__41663\
        );

    \I__9581\ : InMux
    port map (
            O => \N__42000\,
            I => \N__41663\
        );

    \I__9580\ : InMux
    port map (
            O => \N__41999\,
            I => \N__41658\
        );

    \I__9579\ : InMux
    port map (
            O => \N__41998\,
            I => \N__41658\
        );

    \I__9578\ : CascadeMux
    port map (
            O => \N__41997\,
            I => \N__41649\
        );

    \I__9577\ : LocalMux
    port map (
            O => \N__41988\,
            I => \N__41633\
        );

    \I__9576\ : LocalMux
    port map (
            O => \N__41979\,
            I => \N__41633\
        );

    \I__9575\ : InMux
    port map (
            O => \N__41978\,
            I => \N__41620\
        );

    \I__9574\ : InMux
    port map (
            O => \N__41977\,
            I => \N__41620\
        );

    \I__9573\ : InMux
    port map (
            O => \N__41976\,
            I => \N__41620\
        );

    \I__9572\ : CascadeMux
    port map (
            O => \N__41975\,
            I => \N__41601\
        );

    \I__9571\ : CascadeMux
    port map (
            O => \N__41974\,
            I => \N__41593\
        );

    \I__9570\ : LocalMux
    port map (
            O => \N__41969\,
            I => \N__41586\
        );

    \I__9569\ : InMux
    port map (
            O => \N__41968\,
            I => \N__41579\
        );

    \I__9568\ : InMux
    port map (
            O => \N__41967\,
            I => \N__41579\
        );

    \I__9567\ : InMux
    port map (
            O => \N__41966\,
            I => \N__41579\
        );

    \I__9566\ : CascadeMux
    port map (
            O => \N__41965\,
            I => \N__41574\
        );

    \I__9565\ : CascadeMux
    port map (
            O => \N__41964\,
            I => \N__41569\
        );

    \I__9564\ : CascadeMux
    port map (
            O => \N__41963\,
            I => \N__41562\
        );

    \I__9563\ : LocalMux
    port map (
            O => \N__41960\,
            I => \N__41552\
        );

    \I__9562\ : LocalMux
    port map (
            O => \N__41953\,
            I => \N__41552\
        );

    \I__9561\ : LocalMux
    port map (
            O => \N__41948\,
            I => \N__41552\
        );

    \I__9560\ : Span4Mux_v
    port map (
            O => \N__41945\,
            I => \N__41549\
        );

    \I__9559\ : InMux
    port map (
            O => \N__41944\,
            I => \N__41540\
        );

    \I__9558\ : InMux
    port map (
            O => \N__41943\,
            I => \N__41540\
        );

    \I__9557\ : InMux
    port map (
            O => \N__41940\,
            I => \N__41540\
        );

    \I__9556\ : InMux
    port map (
            O => \N__41939\,
            I => \N__41540\
        );

    \I__9555\ : InMux
    port map (
            O => \N__41938\,
            I => \N__41531\
        );

    \I__9554\ : InMux
    port map (
            O => \N__41937\,
            I => \N__41531\
        );

    \I__9553\ : InMux
    port map (
            O => \N__41936\,
            I => \N__41531\
        );

    \I__9552\ : InMux
    port map (
            O => \N__41935\,
            I => \N__41531\
        );

    \I__9551\ : Span4Mux_v
    port map (
            O => \N__41932\,
            I => \N__41524\
        );

    \I__9550\ : LocalMux
    port map (
            O => \N__41923\,
            I => \N__41524\
        );

    \I__9549\ : LocalMux
    port map (
            O => \N__41914\,
            I => \N__41524\
        );

    \I__9548\ : Span4Mux_v
    port map (
            O => \N__41905\,
            I => \N__41519\
        );

    \I__9547\ : LocalMux
    port map (
            O => \N__41896\,
            I => \N__41519\
        );

    \I__9546\ : Span4Mux_v
    port map (
            O => \N__41893\,
            I => \N__41512\
        );

    \I__9545\ : LocalMux
    port map (
            O => \N__41886\,
            I => \N__41512\
        );

    \I__9544\ : LocalMux
    port map (
            O => \N__41879\,
            I => \N__41512\
        );

    \I__9543\ : InMux
    port map (
            O => \N__41876\,
            I => \N__41509\
        );

    \I__9542\ : InMux
    port map (
            O => \N__41875\,
            I => \N__41502\
        );

    \I__9541\ : InMux
    port map (
            O => \N__41872\,
            I => \N__41502\
        );

    \I__9540\ : InMux
    port map (
            O => \N__41869\,
            I => \N__41502\
        );

    \I__9539\ : CascadeMux
    port map (
            O => \N__41868\,
            I => \N__41499\
        );

    \I__9538\ : CascadeMux
    port map (
            O => \N__41867\,
            I => \N__41496\
        );

    \I__9537\ : CascadeMux
    port map (
            O => \N__41866\,
            I => \N__41493\
        );

    \I__9536\ : CascadeMux
    port map (
            O => \N__41865\,
            I => \N__41490\
        );

    \I__9535\ : CascadeMux
    port map (
            O => \N__41864\,
            I => \N__41487\
        );

    \I__9534\ : CascadeMux
    port map (
            O => \N__41863\,
            I => \N__41484\
        );

    \I__9533\ : CascadeMux
    port map (
            O => \N__41862\,
            I => \N__41480\
        );

    \I__9532\ : Span4Mux_v
    port map (
            O => \N__41855\,
            I => \N__41467\
        );

    \I__9531\ : Span4Mux_v
    port map (
            O => \N__41850\,
            I => \N__41467\
        );

    \I__9530\ : LocalMux
    port map (
            O => \N__41843\,
            I => \N__41462\
        );

    \I__9529\ : LocalMux
    port map (
            O => \N__41836\,
            I => \N__41462\
        );

    \I__9528\ : LocalMux
    port map (
            O => \N__41827\,
            I => \N__41457\
        );

    \I__9527\ : LocalMux
    port map (
            O => \N__41820\,
            I => \N__41457\
        );

    \I__9526\ : Span4Mux_v
    port map (
            O => \N__41815\,
            I => \N__41454\
        );

    \I__9525\ : InMux
    port map (
            O => \N__41814\,
            I => \N__41445\
        );

    \I__9524\ : InMux
    port map (
            O => \N__41813\,
            I => \N__41445\
        );

    \I__9523\ : InMux
    port map (
            O => \N__41812\,
            I => \N__41445\
        );

    \I__9522\ : InMux
    port map (
            O => \N__41811\,
            I => \N__41445\
        );

    \I__9521\ : InMux
    port map (
            O => \N__41810\,
            I => \N__41436\
        );

    \I__9520\ : InMux
    port map (
            O => \N__41807\,
            I => \N__41436\
        );

    \I__9519\ : InMux
    port map (
            O => \N__41806\,
            I => \N__41436\
        );

    \I__9518\ : InMux
    port map (
            O => \N__41805\,
            I => \N__41436\
        );

    \I__9517\ : Span4Mux_v
    port map (
            O => \N__41802\,
            I => \N__41421\
        );

    \I__9516\ : LocalMux
    port map (
            O => \N__41793\,
            I => \N__41421\
        );

    \I__9515\ : LocalMux
    port map (
            O => \N__41786\,
            I => \N__41421\
        );

    \I__9514\ : LocalMux
    port map (
            O => \N__41783\,
            I => \N__41421\
        );

    \I__9513\ : LocalMux
    port map (
            O => \N__41772\,
            I => \N__41421\
        );

    \I__9512\ : LocalMux
    port map (
            O => \N__41763\,
            I => \N__41421\
        );

    \I__9511\ : LocalMux
    port map (
            O => \N__41754\,
            I => \N__41421\
        );

    \I__9510\ : InMux
    port map (
            O => \N__41753\,
            I => \N__41414\
        );

    \I__9509\ : InMux
    port map (
            O => \N__41752\,
            I => \N__41414\
        );

    \I__9508\ : InMux
    port map (
            O => \N__41751\,
            I => \N__41414\
        );

    \I__9507\ : InMux
    port map (
            O => \N__41750\,
            I => \N__41407\
        );

    \I__9506\ : InMux
    port map (
            O => \N__41749\,
            I => \N__41407\
        );

    \I__9505\ : InMux
    port map (
            O => \N__41748\,
            I => \N__41407\
        );

    \I__9504\ : InMux
    port map (
            O => \N__41747\,
            I => \N__41400\
        );

    \I__9503\ : InMux
    port map (
            O => \N__41746\,
            I => \N__41400\
        );

    \I__9502\ : InMux
    port map (
            O => \N__41745\,
            I => \N__41400\
        );

    \I__9501\ : InMux
    port map (
            O => \N__41744\,
            I => \N__41393\
        );

    \I__9500\ : InMux
    port map (
            O => \N__41743\,
            I => \N__41393\
        );

    \I__9499\ : InMux
    port map (
            O => \N__41742\,
            I => \N__41393\
        );

    \I__9498\ : Span4Mux_v
    port map (
            O => \N__41739\,
            I => \N__41390\
        );

    \I__9497\ : LocalMux
    port map (
            O => \N__41732\,
            I => \N__41387\
        );

    \I__9496\ : Span4Mux_v
    port map (
            O => \N__41729\,
            I => \N__41372\
        );

    \I__9495\ : LocalMux
    port map (
            O => \N__41724\,
            I => \N__41372\
        );

    \I__9494\ : LocalMux
    port map (
            O => \N__41713\,
            I => \N__41372\
        );

    \I__9493\ : LocalMux
    port map (
            O => \N__41704\,
            I => \N__41372\
        );

    \I__9492\ : LocalMux
    port map (
            O => \N__41695\,
            I => \N__41372\
        );

    \I__9491\ : LocalMux
    port map (
            O => \N__41688\,
            I => \N__41372\
        );

    \I__9490\ : LocalMux
    port map (
            O => \N__41681\,
            I => \N__41372\
        );

    \I__9489\ : InMux
    port map (
            O => \N__41680\,
            I => \N__41367\
        );

    \I__9488\ : InMux
    port map (
            O => \N__41679\,
            I => \N__41367\
        );

    \I__9487\ : LocalMux
    port map (
            O => \N__41672\,
            I => \N__41360\
        );

    \I__9486\ : LocalMux
    port map (
            O => \N__41663\,
            I => \N__41360\
        );

    \I__9485\ : LocalMux
    port map (
            O => \N__41658\,
            I => \N__41360\
        );

    \I__9484\ : InMux
    port map (
            O => \N__41657\,
            I => \N__41353\
        );

    \I__9483\ : InMux
    port map (
            O => \N__41656\,
            I => \N__41353\
        );

    \I__9482\ : InMux
    port map (
            O => \N__41655\,
            I => \N__41353\
        );

    \I__9481\ : InMux
    port map (
            O => \N__41654\,
            I => \N__41342\
        );

    \I__9480\ : InMux
    port map (
            O => \N__41653\,
            I => \N__41342\
        );

    \I__9479\ : InMux
    port map (
            O => \N__41652\,
            I => \N__41342\
        );

    \I__9478\ : InMux
    port map (
            O => \N__41649\,
            I => \N__41342\
        );

    \I__9477\ : InMux
    port map (
            O => \N__41648\,
            I => \N__41342\
        );

    \I__9476\ : InMux
    port map (
            O => \N__41647\,
            I => \N__41333\
        );

    \I__9475\ : InMux
    port map (
            O => \N__41646\,
            I => \N__41333\
        );

    \I__9474\ : InMux
    port map (
            O => \N__41645\,
            I => \N__41333\
        );

    \I__9473\ : InMux
    port map (
            O => \N__41644\,
            I => \N__41333\
        );

    \I__9472\ : InMux
    port map (
            O => \N__41643\,
            I => \N__41324\
        );

    \I__9471\ : InMux
    port map (
            O => \N__41642\,
            I => \N__41324\
        );

    \I__9470\ : InMux
    port map (
            O => \N__41641\,
            I => \N__41324\
        );

    \I__9469\ : InMux
    port map (
            O => \N__41640\,
            I => \N__41324\
        );

    \I__9468\ : CascadeMux
    port map (
            O => \N__41639\,
            I => \N__41318\
        );

    \I__9467\ : CascadeMux
    port map (
            O => \N__41638\,
            I => \N__41311\
        );

    \I__9466\ : Span4Mux_v
    port map (
            O => \N__41633\,
            I => \N__41305\
        );

    \I__9465\ : InMux
    port map (
            O => \N__41632\,
            I => \N__41298\
        );

    \I__9464\ : InMux
    port map (
            O => \N__41631\,
            I => \N__41298\
        );

    \I__9463\ : InMux
    port map (
            O => \N__41630\,
            I => \N__41298\
        );

    \I__9462\ : InMux
    port map (
            O => \N__41629\,
            I => \N__41291\
        );

    \I__9461\ : InMux
    port map (
            O => \N__41628\,
            I => \N__41291\
        );

    \I__9460\ : InMux
    port map (
            O => \N__41627\,
            I => \N__41291\
        );

    \I__9459\ : LocalMux
    port map (
            O => \N__41620\,
            I => \N__41288\
        );

    \I__9458\ : InMux
    port map (
            O => \N__41619\,
            I => \N__41285\
        );

    \I__9457\ : InMux
    port map (
            O => \N__41618\,
            I => \N__41278\
        );

    \I__9456\ : InMux
    port map (
            O => \N__41617\,
            I => \N__41278\
        );

    \I__9455\ : InMux
    port map (
            O => \N__41616\,
            I => \N__41278\
        );

    \I__9454\ : InMux
    port map (
            O => \N__41615\,
            I => \N__41271\
        );

    \I__9453\ : InMux
    port map (
            O => \N__41614\,
            I => \N__41271\
        );

    \I__9452\ : InMux
    port map (
            O => \N__41613\,
            I => \N__41271\
        );

    \I__9451\ : InMux
    port map (
            O => \N__41612\,
            I => \N__41264\
        );

    \I__9450\ : InMux
    port map (
            O => \N__41611\,
            I => \N__41264\
        );

    \I__9449\ : InMux
    port map (
            O => \N__41610\,
            I => \N__41264\
        );

    \I__9448\ : InMux
    port map (
            O => \N__41609\,
            I => \N__41259\
        );

    \I__9447\ : InMux
    port map (
            O => \N__41608\,
            I => \N__41259\
        );

    \I__9446\ : InMux
    port map (
            O => \N__41607\,
            I => \N__41252\
        );

    \I__9445\ : InMux
    port map (
            O => \N__41606\,
            I => \N__41252\
        );

    \I__9444\ : InMux
    port map (
            O => \N__41605\,
            I => \N__41252\
        );

    \I__9443\ : InMux
    port map (
            O => \N__41604\,
            I => \N__41241\
        );

    \I__9442\ : InMux
    port map (
            O => \N__41601\,
            I => \N__41241\
        );

    \I__9441\ : InMux
    port map (
            O => \N__41600\,
            I => \N__41241\
        );

    \I__9440\ : InMux
    port map (
            O => \N__41599\,
            I => \N__41241\
        );

    \I__9439\ : InMux
    port map (
            O => \N__41598\,
            I => \N__41241\
        );

    \I__9438\ : InMux
    port map (
            O => \N__41597\,
            I => \N__41232\
        );

    \I__9437\ : InMux
    port map (
            O => \N__41596\,
            I => \N__41232\
        );

    \I__9436\ : InMux
    port map (
            O => \N__41593\,
            I => \N__41232\
        );

    \I__9435\ : InMux
    port map (
            O => \N__41592\,
            I => \N__41232\
        );

    \I__9434\ : InMux
    port map (
            O => \N__41591\,
            I => \N__41227\
        );

    \I__9433\ : InMux
    port map (
            O => \N__41590\,
            I => \N__41227\
        );

    \I__9432\ : InMux
    port map (
            O => \N__41589\,
            I => \N__41224\
        );

    \I__9431\ : Span4Mux_v
    port map (
            O => \N__41586\,
            I => \N__41219\
        );

    \I__9430\ : LocalMux
    port map (
            O => \N__41579\,
            I => \N__41219\
        );

    \I__9429\ : InMux
    port map (
            O => \N__41578\,
            I => \N__41210\
        );

    \I__9428\ : InMux
    port map (
            O => \N__41577\,
            I => \N__41210\
        );

    \I__9427\ : InMux
    port map (
            O => \N__41574\,
            I => \N__41210\
        );

    \I__9426\ : InMux
    port map (
            O => \N__41573\,
            I => \N__41210\
        );

    \I__9425\ : InMux
    port map (
            O => \N__41572\,
            I => \N__41201\
        );

    \I__9424\ : InMux
    port map (
            O => \N__41569\,
            I => \N__41201\
        );

    \I__9423\ : InMux
    port map (
            O => \N__41568\,
            I => \N__41201\
        );

    \I__9422\ : InMux
    port map (
            O => \N__41567\,
            I => \N__41201\
        );

    \I__9421\ : InMux
    port map (
            O => \N__41566\,
            I => \N__41192\
        );

    \I__9420\ : InMux
    port map (
            O => \N__41565\,
            I => \N__41192\
        );

    \I__9419\ : InMux
    port map (
            O => \N__41562\,
            I => \N__41192\
        );

    \I__9418\ : InMux
    port map (
            O => \N__41561\,
            I => \N__41192\
        );

    \I__9417\ : InMux
    port map (
            O => \N__41560\,
            I => \N__41187\
        );

    \I__9416\ : InMux
    port map (
            O => \N__41559\,
            I => \N__41187\
        );

    \I__9415\ : Span4Mux_v
    port map (
            O => \N__41552\,
            I => \N__41184\
        );

    \I__9414\ : Span4Mux_h
    port map (
            O => \N__41549\,
            I => \N__41177\
        );

    \I__9413\ : LocalMux
    port map (
            O => \N__41540\,
            I => \N__41177\
        );

    \I__9412\ : LocalMux
    port map (
            O => \N__41531\,
            I => \N__41177\
        );

    \I__9411\ : Span4Mux_v
    port map (
            O => \N__41524\,
            I => \N__41174\
        );

    \I__9410\ : Span4Mux_v
    port map (
            O => \N__41519\,
            I => \N__41169\
        );

    \I__9409\ : Span4Mux_v
    port map (
            O => \N__41512\,
            I => \N__41169\
        );

    \I__9408\ : LocalMux
    port map (
            O => \N__41509\,
            I => \N__41164\
        );

    \I__9407\ : LocalMux
    port map (
            O => \N__41502\,
            I => \N__41164\
        );

    \I__9406\ : InMux
    port map (
            O => \N__41499\,
            I => \N__41157\
        );

    \I__9405\ : InMux
    port map (
            O => \N__41496\,
            I => \N__41157\
        );

    \I__9404\ : InMux
    port map (
            O => \N__41493\,
            I => \N__41157\
        );

    \I__9403\ : InMux
    port map (
            O => \N__41490\,
            I => \N__41146\
        );

    \I__9402\ : InMux
    port map (
            O => \N__41487\,
            I => \N__41146\
        );

    \I__9401\ : InMux
    port map (
            O => \N__41484\,
            I => \N__41146\
        );

    \I__9400\ : InMux
    port map (
            O => \N__41483\,
            I => \N__41146\
        );

    \I__9399\ : InMux
    port map (
            O => \N__41480\,
            I => \N__41146\
        );

    \I__9398\ : InMux
    port map (
            O => \N__41479\,
            I => \N__41137\
        );

    \I__9397\ : InMux
    port map (
            O => \N__41478\,
            I => \N__41137\
        );

    \I__9396\ : InMux
    port map (
            O => \N__41477\,
            I => \N__41137\
        );

    \I__9395\ : InMux
    port map (
            O => \N__41476\,
            I => \N__41137\
        );

    \I__9394\ : InMux
    port map (
            O => \N__41475\,
            I => \N__41128\
        );

    \I__9393\ : InMux
    port map (
            O => \N__41474\,
            I => \N__41128\
        );

    \I__9392\ : InMux
    port map (
            O => \N__41473\,
            I => \N__41128\
        );

    \I__9391\ : InMux
    port map (
            O => \N__41472\,
            I => \N__41128\
        );

    \I__9390\ : Span4Mux_h
    port map (
            O => \N__41467\,
            I => \N__41123\
        );

    \I__9389\ : Span4Mux_v
    port map (
            O => \N__41462\,
            I => \N__41123\
        );

    \I__9388\ : Span4Mux_v
    port map (
            O => \N__41457\,
            I => \N__41116\
        );

    \I__9387\ : Span4Mux_h
    port map (
            O => \N__41454\,
            I => \N__41116\
        );

    \I__9386\ : LocalMux
    port map (
            O => \N__41445\,
            I => \N__41116\
        );

    \I__9385\ : LocalMux
    port map (
            O => \N__41436\,
            I => \N__41103\
        );

    \I__9384\ : Span4Mux_v
    port map (
            O => \N__41421\,
            I => \N__41103\
        );

    \I__9383\ : LocalMux
    port map (
            O => \N__41414\,
            I => \N__41103\
        );

    \I__9382\ : LocalMux
    port map (
            O => \N__41407\,
            I => \N__41103\
        );

    \I__9381\ : LocalMux
    port map (
            O => \N__41400\,
            I => \N__41103\
        );

    \I__9380\ : LocalMux
    port map (
            O => \N__41393\,
            I => \N__41103\
        );

    \I__9379\ : Span4Mux_v
    port map (
            O => \N__41390\,
            I => \N__41094\
        );

    \I__9378\ : Span4Mux_h
    port map (
            O => \N__41387\,
            I => \N__41094\
        );

    \I__9377\ : Span4Mux_v
    port map (
            O => \N__41372\,
            I => \N__41094\
        );

    \I__9376\ : LocalMux
    port map (
            O => \N__41367\,
            I => \N__41094\
        );

    \I__9375\ : Span4Mux_v
    port map (
            O => \N__41360\,
            I => \N__41083\
        );

    \I__9374\ : LocalMux
    port map (
            O => \N__41353\,
            I => \N__41083\
        );

    \I__9373\ : LocalMux
    port map (
            O => \N__41342\,
            I => \N__41083\
        );

    \I__9372\ : LocalMux
    port map (
            O => \N__41333\,
            I => \N__41083\
        );

    \I__9371\ : LocalMux
    port map (
            O => \N__41324\,
            I => \N__41083\
        );

    \I__9370\ : InMux
    port map (
            O => \N__41323\,
            I => \N__41078\
        );

    \I__9369\ : InMux
    port map (
            O => \N__41322\,
            I => \N__41078\
        );

    \I__9368\ : InMux
    port map (
            O => \N__41321\,
            I => \N__41069\
        );

    \I__9367\ : InMux
    port map (
            O => \N__41318\,
            I => \N__41069\
        );

    \I__9366\ : InMux
    port map (
            O => \N__41317\,
            I => \N__41069\
        );

    \I__9365\ : InMux
    port map (
            O => \N__41316\,
            I => \N__41069\
        );

    \I__9364\ : InMux
    port map (
            O => \N__41315\,
            I => \N__41064\
        );

    \I__9363\ : InMux
    port map (
            O => \N__41314\,
            I => \N__41064\
        );

    \I__9362\ : InMux
    port map (
            O => \N__41311\,
            I => \N__41055\
        );

    \I__9361\ : InMux
    port map (
            O => \N__41310\,
            I => \N__41055\
        );

    \I__9360\ : InMux
    port map (
            O => \N__41309\,
            I => \N__41055\
        );

    \I__9359\ : InMux
    port map (
            O => \N__41308\,
            I => \N__41055\
        );

    \I__9358\ : Sp12to4
    port map (
            O => \N__41305\,
            I => \N__41042\
        );

    \I__9357\ : LocalMux
    port map (
            O => \N__41298\,
            I => \N__41042\
        );

    \I__9356\ : LocalMux
    port map (
            O => \N__41291\,
            I => \N__41042\
        );

    \I__9355\ : Span12Mux_h
    port map (
            O => \N__41288\,
            I => \N__41042\
        );

    \I__9354\ : LocalMux
    port map (
            O => \N__41285\,
            I => \N__41042\
        );

    \I__9353\ : LocalMux
    port map (
            O => \N__41278\,
            I => \N__41042\
        );

    \I__9352\ : LocalMux
    port map (
            O => \N__41271\,
            I => \N__41037\
        );

    \I__9351\ : LocalMux
    port map (
            O => \N__41264\,
            I => \N__41037\
        );

    \I__9350\ : LocalMux
    port map (
            O => \N__41259\,
            I => \N__41014\
        );

    \I__9349\ : LocalMux
    port map (
            O => \N__41252\,
            I => \N__41014\
        );

    \I__9348\ : LocalMux
    port map (
            O => \N__41241\,
            I => \N__41014\
        );

    \I__9347\ : LocalMux
    port map (
            O => \N__41232\,
            I => \N__41014\
        );

    \I__9346\ : LocalMux
    port map (
            O => \N__41227\,
            I => \N__41014\
        );

    \I__9345\ : LocalMux
    port map (
            O => \N__41224\,
            I => \N__41014\
        );

    \I__9344\ : Sp12to4
    port map (
            O => \N__41219\,
            I => \N__41014\
        );

    \I__9343\ : LocalMux
    port map (
            O => \N__41210\,
            I => \N__41014\
        );

    \I__9342\ : LocalMux
    port map (
            O => \N__41201\,
            I => \N__41014\
        );

    \I__9341\ : LocalMux
    port map (
            O => \N__41192\,
            I => \N__41014\
        );

    \I__9340\ : LocalMux
    port map (
            O => \N__41187\,
            I => \N__41014\
        );

    \I__9339\ : Span4Mux_h
    port map (
            O => \N__41184\,
            I => \N__41009\
        );

    \I__9338\ : Span4Mux_v
    port map (
            O => \N__41177\,
            I => \N__41009\
        );

    \I__9337\ : Span4Mux_h
    port map (
            O => \N__41174\,
            I => \N__40994\
        );

    \I__9336\ : Span4Mux_h
    port map (
            O => \N__41169\,
            I => \N__40994\
        );

    \I__9335\ : Span4Mux_v
    port map (
            O => \N__41164\,
            I => \N__40994\
        );

    \I__9334\ : LocalMux
    port map (
            O => \N__41157\,
            I => \N__40994\
        );

    \I__9333\ : LocalMux
    port map (
            O => \N__41146\,
            I => \N__40994\
        );

    \I__9332\ : LocalMux
    port map (
            O => \N__41137\,
            I => \N__40994\
        );

    \I__9331\ : LocalMux
    port map (
            O => \N__41128\,
            I => \N__40994\
        );

    \I__9330\ : Span4Mux_h
    port map (
            O => \N__41123\,
            I => \N__40987\
        );

    \I__9329\ : Span4Mux_v
    port map (
            O => \N__41116\,
            I => \N__40987\
        );

    \I__9328\ : Span4Mux_v
    port map (
            O => \N__41103\,
            I => \N__40987\
        );

    \I__9327\ : Span4Mux_v
    port map (
            O => \N__41094\,
            I => \N__40974\
        );

    \I__9326\ : Span4Mux_v
    port map (
            O => \N__41083\,
            I => \N__40974\
        );

    \I__9325\ : LocalMux
    port map (
            O => \N__41078\,
            I => \N__40974\
        );

    \I__9324\ : LocalMux
    port map (
            O => \N__41069\,
            I => \N__40974\
        );

    \I__9323\ : LocalMux
    port map (
            O => \N__41064\,
            I => \N__40974\
        );

    \I__9322\ : LocalMux
    port map (
            O => \N__41055\,
            I => \N__40974\
        );

    \I__9321\ : Span12Mux_v
    port map (
            O => \N__41042\,
            I => \N__40971\
        );

    \I__9320\ : Span12Mux_s10_h
    port map (
            O => \N__41037\,
            I => \N__40966\
        );

    \I__9319\ : Span12Mux_s9_v
    port map (
            O => \N__41014\,
            I => \N__40966\
        );

    \I__9318\ : Span4Mux_v
    port map (
            O => \N__41009\,
            I => \N__40961\
        );

    \I__9317\ : Span4Mux_v
    port map (
            O => \N__40994\,
            I => \N__40961\
        );

    \I__9316\ : Span4Mux_v
    port map (
            O => \N__40987\,
            I => \N__40956\
        );

    \I__9315\ : Span4Mux_v
    port map (
            O => \N__40974\,
            I => \N__40956\
        );

    \I__9314\ : Odrv12
    port map (
            O => \N__40971\,
            I => \CONSTANT_ONE_NET\
        );

    \I__9313\ : Odrv12
    port map (
            O => \N__40966\,
            I => \CONSTANT_ONE_NET\
        );

    \I__9312\ : Odrv4
    port map (
            O => \N__40961\,
            I => \CONSTANT_ONE_NET\
        );

    \I__9311\ : Odrv4
    port map (
            O => \N__40956\,
            I => \CONSTANT_ONE_NET\
        );

    \I__9310\ : InMux
    port map (
            O => \N__40947\,
            I => \N__40943\
        );

    \I__9309\ : InMux
    port map (
            O => \N__40946\,
            I => \N__40940\
        );

    \I__9308\ : LocalMux
    port map (
            O => \N__40943\,
            I => \N__40937\
        );

    \I__9307\ : LocalMux
    port map (
            O => \N__40940\,
            I => \N__40934\
        );

    \I__9306\ : Odrv4
    port map (
            O => \N__40937\,
            I => \nx.n2489\
        );

    \I__9305\ : Odrv4
    port map (
            O => \N__40934\,
            I => \nx.n2489\
        );

    \I__9304\ : CascadeMux
    port map (
            O => \N__40929\,
            I => \N__40923\
        );

    \I__9303\ : InMux
    port map (
            O => \N__40928\,
            I => \N__40918\
        );

    \I__9302\ : CascadeMux
    port map (
            O => \N__40927\,
            I => \N__40915\
        );

    \I__9301\ : InMux
    port map (
            O => \N__40926\,
            I => \N__40911\
        );

    \I__9300\ : InMux
    port map (
            O => \N__40923\,
            I => \N__40908\
        );

    \I__9299\ : CascadeMux
    port map (
            O => \N__40922\,
            I => \N__40904\
        );

    \I__9298\ : CascadeMux
    port map (
            O => \N__40921\,
            I => \N__40895\
        );

    \I__9297\ : LocalMux
    port map (
            O => \N__40918\,
            I => \N__40891\
        );

    \I__9296\ : InMux
    port map (
            O => \N__40915\,
            I => \N__40886\
        );

    \I__9295\ : InMux
    port map (
            O => \N__40914\,
            I => \N__40886\
        );

    \I__9294\ : LocalMux
    port map (
            O => \N__40911\,
            I => \N__40881\
        );

    \I__9293\ : LocalMux
    port map (
            O => \N__40908\,
            I => \N__40881\
        );

    \I__9292\ : InMux
    port map (
            O => \N__40907\,
            I => \N__40874\
        );

    \I__9291\ : InMux
    port map (
            O => \N__40904\,
            I => \N__40874\
        );

    \I__9290\ : InMux
    port map (
            O => \N__40903\,
            I => \N__40874\
        );

    \I__9289\ : InMux
    port map (
            O => \N__40902\,
            I => \N__40871\
        );

    \I__9288\ : InMux
    port map (
            O => \N__40901\,
            I => \N__40868\
        );

    \I__9287\ : CascadeMux
    port map (
            O => \N__40900\,
            I => \N__40865\
        );

    \I__9286\ : InMux
    port map (
            O => \N__40899\,
            I => \N__40856\
        );

    \I__9285\ : InMux
    port map (
            O => \N__40898\,
            I => \N__40849\
        );

    \I__9284\ : InMux
    port map (
            O => \N__40895\,
            I => \N__40849\
        );

    \I__9283\ : InMux
    port map (
            O => \N__40894\,
            I => \N__40849\
        );

    \I__9282\ : Span4Mux_v
    port map (
            O => \N__40891\,
            I => \N__40840\
        );

    \I__9281\ : LocalMux
    port map (
            O => \N__40886\,
            I => \N__40840\
        );

    \I__9280\ : Span4Mux_v
    port map (
            O => \N__40881\,
            I => \N__40840\
        );

    \I__9279\ : LocalMux
    port map (
            O => \N__40874\,
            I => \N__40840\
        );

    \I__9278\ : LocalMux
    port map (
            O => \N__40871\,
            I => \N__40835\
        );

    \I__9277\ : LocalMux
    port map (
            O => \N__40868\,
            I => \N__40835\
        );

    \I__9276\ : InMux
    port map (
            O => \N__40865\,
            I => \N__40828\
        );

    \I__9275\ : InMux
    port map (
            O => \N__40864\,
            I => \N__40828\
        );

    \I__9274\ : InMux
    port map (
            O => \N__40863\,
            I => \N__40828\
        );

    \I__9273\ : InMux
    port map (
            O => \N__40862\,
            I => \N__40819\
        );

    \I__9272\ : InMux
    port map (
            O => \N__40861\,
            I => \N__40819\
        );

    \I__9271\ : InMux
    port map (
            O => \N__40860\,
            I => \N__40819\
        );

    \I__9270\ : InMux
    port map (
            O => \N__40859\,
            I => \N__40819\
        );

    \I__9269\ : LocalMux
    port map (
            O => \N__40856\,
            I => \nx.n2522\
        );

    \I__9268\ : LocalMux
    port map (
            O => \N__40849\,
            I => \nx.n2522\
        );

    \I__9267\ : Odrv4
    port map (
            O => \N__40840\,
            I => \nx.n2522\
        );

    \I__9266\ : Odrv4
    port map (
            O => \N__40835\,
            I => \nx.n2522\
        );

    \I__9265\ : LocalMux
    port map (
            O => \N__40828\,
            I => \nx.n2522\
        );

    \I__9264\ : LocalMux
    port map (
            O => \N__40819\,
            I => \nx.n2522\
        );

    \I__9263\ : InMux
    port map (
            O => \N__40806\,
            I => \nx.n10958\
        );

    \I__9262\ : CascadeMux
    port map (
            O => \N__40803\,
            I => \N__40799\
        );

    \I__9261\ : InMux
    port map (
            O => \N__40802\,
            I => \N__40796\
        );

    \I__9260\ : InMux
    port map (
            O => \N__40799\,
            I => \N__40793\
        );

    \I__9259\ : LocalMux
    port map (
            O => \N__40796\,
            I => \N__40790\
        );

    \I__9258\ : LocalMux
    port map (
            O => \N__40793\,
            I => \N__40787\
        );

    \I__9257\ : Span4Mux_v
    port map (
            O => \N__40790\,
            I => \N__40784\
        );

    \I__9256\ : Odrv4
    port map (
            O => \N__40787\,
            I => \nx.n2588\
        );

    \I__9255\ : Odrv4
    port map (
            O => \N__40784\,
            I => \nx.n2588\
        );

    \I__9254\ : IoInMux
    port map (
            O => \N__40779\,
            I => \N__40776\
        );

    \I__9253\ : LocalMux
    port map (
            O => \N__40776\,
            I => \N__40773\
        );

    \I__9252\ : Span12Mux_s11_h
    port map (
            O => \N__40773\,
            I => \N__40770\
        );

    \I__9251\ : Span12Mux_v
    port map (
            O => \N__40770\,
            I => \N__40766\
        );

    \I__9250\ : InMux
    port map (
            O => \N__40769\,
            I => \N__40763\
        );

    \I__9249\ : Odrv12
    port map (
            O => \N__40766\,
            I => pin_oe_12
        );

    \I__9248\ : LocalMux
    port map (
            O => \N__40763\,
            I => pin_oe_12
        );

    \I__9247\ : InMux
    port map (
            O => \N__40758\,
            I => \N__40755\
        );

    \I__9246\ : LocalMux
    port map (
            O => \N__40755\,
            I => n45
        );

    \I__9245\ : InMux
    port map (
            O => \N__40752\,
            I => \bfn_17_15_0_\
        );

    \I__9244\ : InMux
    port map (
            O => \N__40749\,
            I => n10700
        );

    \I__9243\ : InMux
    port map (
            O => \N__40746\,
            I => n10701
        );

    \I__9242\ : InMux
    port map (
            O => \N__40743\,
            I => n10702
        );

    \I__9241\ : CascadeMux
    port map (
            O => \N__40740\,
            I => \N__40737\
        );

    \I__9240\ : InMux
    port map (
            O => \N__40737\,
            I => \N__40733\
        );

    \I__9239\ : InMux
    port map (
            O => \N__40736\,
            I => \N__40730\
        );

    \I__9238\ : LocalMux
    port map (
            O => \N__40733\,
            I => \N__40726\
        );

    \I__9237\ : LocalMux
    port map (
            O => \N__40730\,
            I => \N__40723\
        );

    \I__9236\ : InMux
    port map (
            O => \N__40729\,
            I => \N__40720\
        );

    \I__9235\ : Span4Mux_h
    port map (
            O => \N__40726\,
            I => \N__40717\
        );

    \I__9234\ : Span4Mux_h
    port map (
            O => \N__40723\,
            I => \N__40714\
        );

    \I__9233\ : LocalMux
    port map (
            O => \N__40720\,
            I => \nx.n2498\
        );

    \I__9232\ : Odrv4
    port map (
            O => \N__40717\,
            I => \nx.n2498\
        );

    \I__9231\ : Odrv4
    port map (
            O => \N__40714\,
            I => \nx.n2498\
        );

    \I__9230\ : InMux
    port map (
            O => \N__40707\,
            I => \N__40704\
        );

    \I__9229\ : LocalMux
    port map (
            O => \N__40704\,
            I => \N__40701\
        );

    \I__9228\ : Span4Mux_v
    port map (
            O => \N__40701\,
            I => \N__40698\
        );

    \I__9227\ : Odrv4
    port map (
            O => \N__40698\,
            I => \nx.n2565\
        );

    \I__9226\ : InMux
    port map (
            O => \N__40695\,
            I => \nx.n10949\
        );

    \I__9225\ : InMux
    port map (
            O => \N__40692\,
            I => \N__40687\
        );

    \I__9224\ : InMux
    port map (
            O => \N__40691\,
            I => \N__40684\
        );

    \I__9223\ : InMux
    port map (
            O => \N__40690\,
            I => \N__40681\
        );

    \I__9222\ : LocalMux
    port map (
            O => \N__40687\,
            I => \nx.n2497\
        );

    \I__9221\ : LocalMux
    port map (
            O => \N__40684\,
            I => \nx.n2497\
        );

    \I__9220\ : LocalMux
    port map (
            O => \N__40681\,
            I => \nx.n2497\
        );

    \I__9219\ : CascadeMux
    port map (
            O => \N__40674\,
            I => \N__40671\
        );

    \I__9218\ : InMux
    port map (
            O => \N__40671\,
            I => \N__40668\
        );

    \I__9217\ : LocalMux
    port map (
            O => \N__40668\,
            I => \N__40665\
        );

    \I__9216\ : Odrv4
    port map (
            O => \N__40665\,
            I => \nx.n2564\
        );

    \I__9215\ : InMux
    port map (
            O => \N__40662\,
            I => \nx.n10950\
        );

    \I__9214\ : InMux
    port map (
            O => \N__40659\,
            I => \N__40655\
        );

    \I__9213\ : InMux
    port map (
            O => \N__40658\,
            I => \N__40652\
        );

    \I__9212\ : LocalMux
    port map (
            O => \N__40655\,
            I => \nx.n2496\
        );

    \I__9211\ : LocalMux
    port map (
            O => \N__40652\,
            I => \nx.n2496\
        );

    \I__9210\ : InMux
    port map (
            O => \N__40647\,
            I => \N__40644\
        );

    \I__9209\ : LocalMux
    port map (
            O => \N__40644\,
            I => \nx.n2563\
        );

    \I__9208\ : InMux
    port map (
            O => \N__40641\,
            I => \nx.n10951\
        );

    \I__9207\ : CascadeMux
    port map (
            O => \N__40638\,
            I => \N__40634\
        );

    \I__9206\ : InMux
    port map (
            O => \N__40637\,
            I => \N__40631\
        );

    \I__9205\ : InMux
    port map (
            O => \N__40634\,
            I => \N__40628\
        );

    \I__9204\ : LocalMux
    port map (
            O => \N__40631\,
            I => \nx.n2495\
        );

    \I__9203\ : LocalMux
    port map (
            O => \N__40628\,
            I => \nx.n2495\
        );

    \I__9202\ : CascadeMux
    port map (
            O => \N__40623\,
            I => \N__40620\
        );

    \I__9201\ : InMux
    port map (
            O => \N__40620\,
            I => \N__40617\
        );

    \I__9200\ : LocalMux
    port map (
            O => \N__40617\,
            I => \N__40614\
        );

    \I__9199\ : Odrv4
    port map (
            O => \N__40614\,
            I => \nx.n2562\
        );

    \I__9198\ : InMux
    port map (
            O => \N__40611\,
            I => \nx.n10952\
        );

    \I__9197\ : CascadeMux
    port map (
            O => \N__40608\,
            I => \N__40605\
        );

    \I__9196\ : InMux
    port map (
            O => \N__40605\,
            I => \N__40601\
        );

    \I__9195\ : InMux
    port map (
            O => \N__40604\,
            I => \N__40597\
        );

    \I__9194\ : LocalMux
    port map (
            O => \N__40601\,
            I => \N__40594\
        );

    \I__9193\ : InMux
    port map (
            O => \N__40600\,
            I => \N__40591\
        );

    \I__9192\ : LocalMux
    port map (
            O => \N__40597\,
            I => \nx.n2494\
        );

    \I__9191\ : Odrv4
    port map (
            O => \N__40594\,
            I => \nx.n2494\
        );

    \I__9190\ : LocalMux
    port map (
            O => \N__40591\,
            I => \nx.n2494\
        );

    \I__9189\ : CascadeMux
    port map (
            O => \N__40584\,
            I => \N__40581\
        );

    \I__9188\ : InMux
    port map (
            O => \N__40581\,
            I => \N__40578\
        );

    \I__9187\ : LocalMux
    port map (
            O => \N__40578\,
            I => \N__40575\
        );

    \I__9186\ : Odrv4
    port map (
            O => \N__40575\,
            I => \nx.n2561\
        );

    \I__9185\ : InMux
    port map (
            O => \N__40572\,
            I => \bfn_16_26_0_\
        );

    \I__9184\ : CascadeMux
    port map (
            O => \N__40569\,
            I => \N__40566\
        );

    \I__9183\ : InMux
    port map (
            O => \N__40566\,
            I => \N__40562\
        );

    \I__9182\ : CascadeMux
    port map (
            O => \N__40565\,
            I => \N__40559\
        );

    \I__9181\ : LocalMux
    port map (
            O => \N__40562\,
            I => \N__40555\
        );

    \I__9180\ : InMux
    port map (
            O => \N__40559\,
            I => \N__40552\
        );

    \I__9179\ : InMux
    port map (
            O => \N__40558\,
            I => \N__40549\
        );

    \I__9178\ : Odrv4
    port map (
            O => \N__40555\,
            I => \nx.n2493\
        );

    \I__9177\ : LocalMux
    port map (
            O => \N__40552\,
            I => \nx.n2493\
        );

    \I__9176\ : LocalMux
    port map (
            O => \N__40549\,
            I => \nx.n2493\
        );

    \I__9175\ : InMux
    port map (
            O => \N__40542\,
            I => \N__40539\
        );

    \I__9174\ : LocalMux
    port map (
            O => \N__40539\,
            I => \N__40536\
        );

    \I__9173\ : Span4Mux_h
    port map (
            O => \N__40536\,
            I => \N__40533\
        );

    \I__9172\ : Odrv4
    port map (
            O => \N__40533\,
            I => \nx.n2560\
        );

    \I__9171\ : InMux
    port map (
            O => \N__40530\,
            I => \nx.n10954\
        );

    \I__9170\ : InMux
    port map (
            O => \N__40527\,
            I => \N__40524\
        );

    \I__9169\ : LocalMux
    port map (
            O => \N__40524\,
            I => \N__40520\
        );

    \I__9168\ : CascadeMux
    port map (
            O => \N__40523\,
            I => \N__40517\
        );

    \I__9167\ : Span4Mux_v
    port map (
            O => \N__40520\,
            I => \N__40513\
        );

    \I__9166\ : InMux
    port map (
            O => \N__40517\,
            I => \N__40510\
        );

    \I__9165\ : InMux
    port map (
            O => \N__40516\,
            I => \N__40507\
        );

    \I__9164\ : Odrv4
    port map (
            O => \N__40513\,
            I => \nx.n2492\
        );

    \I__9163\ : LocalMux
    port map (
            O => \N__40510\,
            I => \nx.n2492\
        );

    \I__9162\ : LocalMux
    port map (
            O => \N__40507\,
            I => \nx.n2492\
        );

    \I__9161\ : CascadeMux
    port map (
            O => \N__40500\,
            I => \N__40497\
        );

    \I__9160\ : InMux
    port map (
            O => \N__40497\,
            I => \N__40494\
        );

    \I__9159\ : LocalMux
    port map (
            O => \N__40494\,
            I => \N__40491\
        );

    \I__9158\ : Span4Mux_v
    port map (
            O => \N__40491\,
            I => \N__40488\
        );

    \I__9157\ : Odrv4
    port map (
            O => \N__40488\,
            I => \nx.n2559\
        );

    \I__9156\ : InMux
    port map (
            O => \N__40485\,
            I => \nx.n10955\
        );

    \I__9155\ : CascadeMux
    port map (
            O => \N__40482\,
            I => \N__40479\
        );

    \I__9154\ : InMux
    port map (
            O => \N__40479\,
            I => \N__40476\
        );

    \I__9153\ : LocalMux
    port map (
            O => \N__40476\,
            I => \N__40471\
        );

    \I__9152\ : InMux
    port map (
            O => \N__40475\,
            I => \N__40466\
        );

    \I__9151\ : InMux
    port map (
            O => \N__40474\,
            I => \N__40466\
        );

    \I__9150\ : Span4Mux_h
    port map (
            O => \N__40471\,
            I => \N__40463\
        );

    \I__9149\ : LocalMux
    port map (
            O => \N__40466\,
            I => \nx.n2506\
        );

    \I__9148\ : Odrv4
    port map (
            O => \N__40463\,
            I => \nx.n2506\
        );

    \I__9147\ : InMux
    port map (
            O => \N__40458\,
            I => \N__40455\
        );

    \I__9146\ : LocalMux
    port map (
            O => \N__40455\,
            I => \N__40452\
        );

    \I__9145\ : Odrv4
    port map (
            O => \N__40452\,
            I => \nx.n2573\
        );

    \I__9144\ : InMux
    port map (
            O => \N__40449\,
            I => \nx.n10941\
        );

    \I__9143\ : CascadeMux
    port map (
            O => \N__40446\,
            I => \N__40442\
        );

    \I__9142\ : CascadeMux
    port map (
            O => \N__40445\,
            I => \N__40439\
        );

    \I__9141\ : InMux
    port map (
            O => \N__40442\,
            I => \N__40436\
        );

    \I__9140\ : InMux
    port map (
            O => \N__40439\,
            I => \N__40433\
        );

    \I__9139\ : LocalMux
    port map (
            O => \N__40436\,
            I => \nx.n2505\
        );

    \I__9138\ : LocalMux
    port map (
            O => \N__40433\,
            I => \nx.n2505\
        );

    \I__9137\ : InMux
    port map (
            O => \N__40428\,
            I => \N__40425\
        );

    \I__9136\ : LocalMux
    port map (
            O => \N__40425\,
            I => \nx.n2572\
        );

    \I__9135\ : InMux
    port map (
            O => \N__40422\,
            I => \nx.n10942\
        );

    \I__9134\ : CascadeMux
    port map (
            O => \N__40419\,
            I => \N__40416\
        );

    \I__9133\ : InMux
    port map (
            O => \N__40416\,
            I => \N__40412\
        );

    \I__9132\ : CascadeMux
    port map (
            O => \N__40415\,
            I => \N__40409\
        );

    \I__9131\ : LocalMux
    port map (
            O => \N__40412\,
            I => \N__40405\
        );

    \I__9130\ : InMux
    port map (
            O => \N__40409\,
            I => \N__40402\
        );

    \I__9129\ : InMux
    port map (
            O => \N__40408\,
            I => \N__40399\
        );

    \I__9128\ : Span4Mux_h
    port map (
            O => \N__40405\,
            I => \N__40396\
        );

    \I__9127\ : LocalMux
    port map (
            O => \N__40402\,
            I => \nx.n2504\
        );

    \I__9126\ : LocalMux
    port map (
            O => \N__40399\,
            I => \nx.n2504\
        );

    \I__9125\ : Odrv4
    port map (
            O => \N__40396\,
            I => \nx.n2504\
        );

    \I__9124\ : InMux
    port map (
            O => \N__40389\,
            I => \N__40386\
        );

    \I__9123\ : LocalMux
    port map (
            O => \N__40386\,
            I => \N__40383\
        );

    \I__9122\ : Span4Mux_h
    port map (
            O => \N__40383\,
            I => \N__40380\
        );

    \I__9121\ : Odrv4
    port map (
            O => \N__40380\,
            I => \nx.n2571\
        );

    \I__9120\ : InMux
    port map (
            O => \N__40377\,
            I => \nx.n10943\
        );

    \I__9119\ : InMux
    port map (
            O => \N__40374\,
            I => \N__40369\
        );

    \I__9118\ : InMux
    port map (
            O => \N__40373\,
            I => \N__40366\
        );

    \I__9117\ : InMux
    port map (
            O => \N__40372\,
            I => \N__40363\
        );

    \I__9116\ : LocalMux
    port map (
            O => \N__40369\,
            I => \N__40360\
        );

    \I__9115\ : LocalMux
    port map (
            O => \N__40366\,
            I => \N__40357\
        );

    \I__9114\ : LocalMux
    port map (
            O => \N__40363\,
            I => \N__40354\
        );

    \I__9113\ : Odrv4
    port map (
            O => \N__40360\,
            I => \nx.n2503\
        );

    \I__9112\ : Odrv4
    port map (
            O => \N__40357\,
            I => \nx.n2503\
        );

    \I__9111\ : Odrv4
    port map (
            O => \N__40354\,
            I => \nx.n2503\
        );

    \I__9110\ : CascadeMux
    port map (
            O => \N__40347\,
            I => \N__40344\
        );

    \I__9109\ : InMux
    port map (
            O => \N__40344\,
            I => \N__40341\
        );

    \I__9108\ : LocalMux
    port map (
            O => \N__40341\,
            I => \N__40338\
        );

    \I__9107\ : Span4Mux_h
    port map (
            O => \N__40338\,
            I => \N__40335\
        );

    \I__9106\ : Odrv4
    port map (
            O => \N__40335\,
            I => \nx.n2570\
        );

    \I__9105\ : InMux
    port map (
            O => \N__40332\,
            I => \nx.n10944\
        );

    \I__9104\ : CascadeMux
    port map (
            O => \N__40329\,
            I => \N__40326\
        );

    \I__9103\ : InMux
    port map (
            O => \N__40326\,
            I => \N__40323\
        );

    \I__9102\ : LocalMux
    port map (
            O => \N__40323\,
            I => \N__40318\
        );

    \I__9101\ : InMux
    port map (
            O => \N__40322\,
            I => \N__40315\
        );

    \I__9100\ : InMux
    port map (
            O => \N__40321\,
            I => \N__40312\
        );

    \I__9099\ : Span4Mux_h
    port map (
            O => \N__40318\,
            I => \N__40309\
        );

    \I__9098\ : LocalMux
    port map (
            O => \N__40315\,
            I => \nx.n2502\
        );

    \I__9097\ : LocalMux
    port map (
            O => \N__40312\,
            I => \nx.n2502\
        );

    \I__9096\ : Odrv4
    port map (
            O => \N__40309\,
            I => \nx.n2502\
        );

    \I__9095\ : InMux
    port map (
            O => \N__40302\,
            I => \N__40299\
        );

    \I__9094\ : LocalMux
    port map (
            O => \N__40299\,
            I => \N__40296\
        );

    \I__9093\ : Span4Mux_h
    port map (
            O => \N__40296\,
            I => \N__40293\
        );

    \I__9092\ : Odrv4
    port map (
            O => \N__40293\,
            I => \nx.n2569\
        );

    \I__9091\ : InMux
    port map (
            O => \N__40290\,
            I => \bfn_16_25_0_\
        );

    \I__9090\ : CascadeMux
    port map (
            O => \N__40287\,
            I => \N__40284\
        );

    \I__9089\ : InMux
    port map (
            O => \N__40284\,
            I => \N__40280\
        );

    \I__9088\ : CascadeMux
    port map (
            O => \N__40283\,
            I => \N__40277\
        );

    \I__9087\ : LocalMux
    port map (
            O => \N__40280\,
            I => \N__40274\
        );

    \I__9086\ : InMux
    port map (
            O => \N__40277\,
            I => \N__40271\
        );

    \I__9085\ : Span4Mux_h
    port map (
            O => \N__40274\,
            I => \N__40268\
        );

    \I__9084\ : LocalMux
    port map (
            O => \N__40271\,
            I => \nx.n2501\
        );

    \I__9083\ : Odrv4
    port map (
            O => \N__40268\,
            I => \nx.n2501\
        );

    \I__9082\ : InMux
    port map (
            O => \N__40263\,
            I => \N__40260\
        );

    \I__9081\ : LocalMux
    port map (
            O => \N__40260\,
            I => \N__40257\
        );

    \I__9080\ : Span4Mux_h
    port map (
            O => \N__40257\,
            I => \N__40254\
        );

    \I__9079\ : Odrv4
    port map (
            O => \N__40254\,
            I => \nx.n2568\
        );

    \I__9078\ : InMux
    port map (
            O => \N__40251\,
            I => \nx.n10946\
        );

    \I__9077\ : CascadeMux
    port map (
            O => \N__40248\,
            I => \N__40245\
        );

    \I__9076\ : InMux
    port map (
            O => \N__40245\,
            I => \N__40242\
        );

    \I__9075\ : LocalMux
    port map (
            O => \N__40242\,
            I => \N__40238\
        );

    \I__9074\ : InMux
    port map (
            O => \N__40241\,
            I => \N__40234\
        );

    \I__9073\ : Span4Mux_h
    port map (
            O => \N__40238\,
            I => \N__40231\
        );

    \I__9072\ : InMux
    port map (
            O => \N__40237\,
            I => \N__40228\
        );

    \I__9071\ : LocalMux
    port map (
            O => \N__40234\,
            I => \nx.n2500\
        );

    \I__9070\ : Odrv4
    port map (
            O => \N__40231\,
            I => \nx.n2500\
        );

    \I__9069\ : LocalMux
    port map (
            O => \N__40228\,
            I => \nx.n2500\
        );

    \I__9068\ : CascadeMux
    port map (
            O => \N__40221\,
            I => \N__40218\
        );

    \I__9067\ : InMux
    port map (
            O => \N__40218\,
            I => \N__40215\
        );

    \I__9066\ : LocalMux
    port map (
            O => \N__40215\,
            I => \N__40212\
        );

    \I__9065\ : Span4Mux_v
    port map (
            O => \N__40212\,
            I => \N__40209\
        );

    \I__9064\ : Odrv4
    port map (
            O => \N__40209\,
            I => \nx.n2567\
        );

    \I__9063\ : InMux
    port map (
            O => \N__40206\,
            I => \nx.n10947\
        );

    \I__9062\ : CascadeMux
    port map (
            O => \N__40203\,
            I => \N__40198\
        );

    \I__9061\ : CascadeMux
    port map (
            O => \N__40202\,
            I => \N__40195\
        );

    \I__9060\ : InMux
    port map (
            O => \N__40201\,
            I => \N__40192\
        );

    \I__9059\ : InMux
    port map (
            O => \N__40198\,
            I => \N__40189\
        );

    \I__9058\ : InMux
    port map (
            O => \N__40195\,
            I => \N__40186\
        );

    \I__9057\ : LocalMux
    port map (
            O => \N__40192\,
            I => \N__40181\
        );

    \I__9056\ : LocalMux
    port map (
            O => \N__40189\,
            I => \N__40181\
        );

    \I__9055\ : LocalMux
    port map (
            O => \N__40186\,
            I => \nx.n2499\
        );

    \I__9054\ : Odrv4
    port map (
            O => \N__40181\,
            I => \nx.n2499\
        );

    \I__9053\ : InMux
    port map (
            O => \N__40176\,
            I => \N__40173\
        );

    \I__9052\ : LocalMux
    port map (
            O => \N__40173\,
            I => \N__40170\
        );

    \I__9051\ : Odrv4
    port map (
            O => \N__40170\,
            I => \nx.n2566\
        );

    \I__9050\ : InMux
    port map (
            O => \N__40167\,
            I => \nx.n10948\
        );

    \I__9049\ : CascadeMux
    port map (
            O => \N__40164\,
            I => \N__40160\
        );

    \I__9048\ : CascadeMux
    port map (
            O => \N__40163\,
            I => \N__40156\
        );

    \I__9047\ : InMux
    port map (
            O => \N__40160\,
            I => \N__40153\
        );

    \I__9046\ : InMux
    port map (
            O => \N__40159\,
            I => \N__40148\
        );

    \I__9045\ : InMux
    port map (
            O => \N__40156\,
            I => \N__40148\
        );

    \I__9044\ : LocalMux
    port map (
            O => \N__40153\,
            I => \N__40145\
        );

    \I__9043\ : LocalMux
    port map (
            O => \N__40148\,
            I => \N__40142\
        );

    \I__9042\ : Span4Mux_h
    port map (
            O => \N__40145\,
            I => \N__40137\
        );

    \I__9041\ : Span4Mux_h
    port map (
            O => \N__40142\,
            I => \N__40137\
        );

    \I__9040\ : Odrv4
    port map (
            O => \N__40137\,
            I => \nx.n2590\
        );

    \I__9039\ : CascadeMux
    port map (
            O => \N__40134\,
            I => \N__40131\
        );

    \I__9038\ : InMux
    port map (
            O => \N__40131\,
            I => \N__40128\
        );

    \I__9037\ : LocalMux
    port map (
            O => \N__40128\,
            I => \N__40125\
        );

    \I__9036\ : Odrv12
    port map (
            O => \N__40125\,
            I => \nx.n2657\
        );

    \I__9035\ : InMux
    port map (
            O => \N__40122\,
            I => \nx.n10978\
        );

    \I__9034\ : InMux
    port map (
            O => \N__40119\,
            I => \N__40116\
        );

    \I__9033\ : LocalMux
    port map (
            O => \N__40116\,
            I => \N__40113\
        );

    \I__9032\ : Odrv12
    port map (
            O => \N__40113\,
            I => \nx.n2656\
        );

    \I__9031\ : InMux
    port map (
            O => \N__40110\,
            I => \nx.n10979\
        );

    \I__9030\ : CascadeMux
    port map (
            O => \N__40107\,
            I => \N__40102\
        );

    \I__9029\ : InMux
    port map (
            O => \N__40106\,
            I => \N__40088\
        );

    \I__9028\ : InMux
    port map (
            O => \N__40105\,
            I => \N__40085\
        );

    \I__9027\ : InMux
    port map (
            O => \N__40102\,
            I => \N__40080\
        );

    \I__9026\ : InMux
    port map (
            O => \N__40101\,
            I => \N__40080\
        );

    \I__9025\ : InMux
    port map (
            O => \N__40100\,
            I => \N__40065\
        );

    \I__9024\ : InMux
    port map (
            O => \N__40099\,
            I => \N__40065\
        );

    \I__9023\ : InMux
    port map (
            O => \N__40098\,
            I => \N__40065\
        );

    \I__9022\ : InMux
    port map (
            O => \N__40097\,
            I => \N__40065\
        );

    \I__9021\ : InMux
    port map (
            O => \N__40096\,
            I => \N__40065\
        );

    \I__9020\ : InMux
    port map (
            O => \N__40095\,
            I => \N__40062\
        );

    \I__9019\ : CascadeMux
    port map (
            O => \N__40094\,
            I => \N__40059\
        );

    \I__9018\ : CascadeMux
    port map (
            O => \N__40093\,
            I => \N__40055\
        );

    \I__9017\ : CascadeMux
    port map (
            O => \N__40092\,
            I => \N__40052\
        );

    \I__9016\ : CascadeMux
    port map (
            O => \N__40091\,
            I => \N__40048\
        );

    \I__9015\ : LocalMux
    port map (
            O => \N__40088\,
            I => \N__40039\
        );

    \I__9014\ : LocalMux
    port map (
            O => \N__40085\,
            I => \N__40039\
        );

    \I__9013\ : LocalMux
    port map (
            O => \N__40080\,
            I => \N__40039\
        );

    \I__9012\ : InMux
    port map (
            O => \N__40079\,
            I => \N__40034\
        );

    \I__9011\ : InMux
    port map (
            O => \N__40078\,
            I => \N__40034\
        );

    \I__9010\ : InMux
    port map (
            O => \N__40077\,
            I => \N__40031\
        );

    \I__9009\ : InMux
    port map (
            O => \N__40076\,
            I => \N__40028\
        );

    \I__9008\ : LocalMux
    port map (
            O => \N__40065\,
            I => \N__40023\
        );

    \I__9007\ : LocalMux
    port map (
            O => \N__40062\,
            I => \N__40023\
        );

    \I__9006\ : InMux
    port map (
            O => \N__40059\,
            I => \N__40012\
        );

    \I__9005\ : InMux
    port map (
            O => \N__40058\,
            I => \N__40012\
        );

    \I__9004\ : InMux
    port map (
            O => \N__40055\,
            I => \N__40012\
        );

    \I__9003\ : InMux
    port map (
            O => \N__40052\,
            I => \N__40012\
        );

    \I__9002\ : InMux
    port map (
            O => \N__40051\,
            I => \N__40012\
        );

    \I__9001\ : InMux
    port map (
            O => \N__40048\,
            I => \N__40005\
        );

    \I__9000\ : InMux
    port map (
            O => \N__40047\,
            I => \N__40005\
        );

    \I__8999\ : InMux
    port map (
            O => \N__40046\,
            I => \N__40005\
        );

    \I__8998\ : Span4Mux_h
    port map (
            O => \N__40039\,
            I => \N__40002\
        );

    \I__8997\ : LocalMux
    port map (
            O => \N__40034\,
            I => \nx.n2621\
        );

    \I__8996\ : LocalMux
    port map (
            O => \N__40031\,
            I => \nx.n2621\
        );

    \I__8995\ : LocalMux
    port map (
            O => \N__40028\,
            I => \nx.n2621\
        );

    \I__8994\ : Odrv12
    port map (
            O => \N__40023\,
            I => \nx.n2621\
        );

    \I__8993\ : LocalMux
    port map (
            O => \N__40012\,
            I => \nx.n2621\
        );

    \I__8992\ : LocalMux
    port map (
            O => \N__40005\,
            I => \nx.n2621\
        );

    \I__8991\ : Odrv4
    port map (
            O => \N__40002\,
            I => \nx.n2621\
        );

    \I__8990\ : InMux
    port map (
            O => \N__39987\,
            I => \nx.n10980\
        );

    \I__8989\ : CascadeMux
    port map (
            O => \N__39984\,
            I => \N__39980\
        );

    \I__8988\ : InMux
    port map (
            O => \N__39983\,
            I => \N__39977\
        );

    \I__8987\ : InMux
    port map (
            O => \N__39980\,
            I => \N__39974\
        );

    \I__8986\ : LocalMux
    port map (
            O => \N__39977\,
            I => \N__39971\
        );

    \I__8985\ : LocalMux
    port map (
            O => \N__39974\,
            I => \N__39968\
        );

    \I__8984\ : Span4Mux_h
    port map (
            O => \N__39971\,
            I => \N__39965\
        );

    \I__8983\ : Span4Mux_h
    port map (
            O => \N__39968\,
            I => \N__39962\
        );

    \I__8982\ : Span4Mux_h
    port map (
            O => \N__39965\,
            I => \N__39959\
        );

    \I__8981\ : Span4Mux_h
    port map (
            O => \N__39962\,
            I => \N__39956\
        );

    \I__8980\ : Odrv4
    port map (
            O => \N__39959\,
            I => \nx.n2687\
        );

    \I__8979\ : Odrv4
    port map (
            O => \N__39956\,
            I => \nx.n2687\
        );

    \I__8978\ : InMux
    port map (
            O => \N__39951\,
            I => \N__39944\
        );

    \I__8977\ : InMux
    port map (
            O => \N__39950\,
            I => \N__39944\
        );

    \I__8976\ : CascadeMux
    port map (
            O => \N__39949\,
            I => \N__39941\
        );

    \I__8975\ : LocalMux
    port map (
            O => \N__39944\,
            I => \N__39938\
        );

    \I__8974\ : InMux
    port map (
            O => \N__39941\,
            I => \N__39935\
        );

    \I__8973\ : Span4Mux_h
    port map (
            O => \N__39938\,
            I => \N__39932\
        );

    \I__8972\ : LocalMux
    port map (
            O => \N__39935\,
            I => \nx.n2589\
        );

    \I__8971\ : Odrv4
    port map (
            O => \N__39932\,
            I => \nx.n2589\
        );

    \I__8970\ : InMux
    port map (
            O => \N__39927\,
            I => \N__39924\
        );

    \I__8969\ : LocalMux
    port map (
            O => \N__39924\,
            I => \N__39918\
        );

    \I__8968\ : InMux
    port map (
            O => \N__39923\,
            I => \N__39915\
        );

    \I__8967\ : InMux
    port map (
            O => \N__39922\,
            I => \N__39912\
        );

    \I__8966\ : InMux
    port map (
            O => \N__39921\,
            I => \N__39909\
        );

    \I__8965\ : Span4Mux_h
    port map (
            O => \N__39918\,
            I => \N__39906\
        );

    \I__8964\ : LocalMux
    port map (
            O => \N__39915\,
            I => \N__39903\
        );

    \I__8963\ : LocalMux
    port map (
            O => \N__39912\,
            I => \N__39900\
        );

    \I__8962\ : LocalMux
    port map (
            O => \N__39909\,
            I => \N__39896\
        );

    \I__8961\ : Span4Mux_h
    port map (
            O => \N__39906\,
            I => \N__39893\
        );

    \I__8960\ : Span4Mux_v
    port map (
            O => \N__39903\,
            I => \N__39890\
        );

    \I__8959\ : Span4Mux_h
    port map (
            O => \N__39900\,
            I => \N__39887\
        );

    \I__8958\ : InMux
    port map (
            O => \N__39899\,
            I => \N__39884\
        );

    \I__8957\ : Sp12to4
    port map (
            O => \N__39896\,
            I => \N__39881\
        );

    \I__8956\ : Span4Mux_h
    port map (
            O => \N__39893\,
            I => \N__39878\
        );

    \I__8955\ : Span4Mux_h
    port map (
            O => \N__39890\,
            I => \N__39873\
        );

    \I__8954\ : Span4Mux_h
    port map (
            O => \N__39887\,
            I => \N__39873\
        );

    \I__8953\ : LocalMux
    port map (
            O => \N__39884\,
            I => \nx.bit_ctr_10\
        );

    \I__8952\ : Odrv12
    port map (
            O => \N__39881\,
            I => \nx.bit_ctr_10\
        );

    \I__8951\ : Odrv4
    port map (
            O => \N__39878\,
            I => \nx.bit_ctr_10\
        );

    \I__8950\ : Odrv4
    port map (
            O => \N__39873\,
            I => \nx.bit_ctr_10\
        );

    \I__8949\ : InMux
    port map (
            O => \N__39864\,
            I => \N__39861\
        );

    \I__8948\ : LocalMux
    port map (
            O => \N__39861\,
            I => \N__39858\
        );

    \I__8947\ : Span4Mux_v
    port map (
            O => \N__39858\,
            I => \N__39855\
        );

    \I__8946\ : Odrv4
    port map (
            O => \N__39855\,
            I => \nx.n2577\
        );

    \I__8945\ : InMux
    port map (
            O => \N__39852\,
            I => \bfn_16_24_0_\
        );

    \I__8944\ : CascadeMux
    port map (
            O => \N__39849\,
            I => \N__39845\
        );

    \I__8943\ : InMux
    port map (
            O => \N__39848\,
            I => \N__39842\
        );

    \I__8942\ : InMux
    port map (
            O => \N__39845\,
            I => \N__39839\
        );

    \I__8941\ : LocalMux
    port map (
            O => \N__39842\,
            I => \N__39835\
        );

    \I__8940\ : LocalMux
    port map (
            O => \N__39839\,
            I => \N__39832\
        );

    \I__8939\ : InMux
    port map (
            O => \N__39838\,
            I => \N__39829\
        );

    \I__8938\ : Span4Mux_v
    port map (
            O => \N__39835\,
            I => \N__39824\
        );

    \I__8937\ : Span4Mux_v
    port map (
            O => \N__39832\,
            I => \N__39824\
        );

    \I__8936\ : LocalMux
    port map (
            O => \N__39829\,
            I => \nx.n2509\
        );

    \I__8935\ : Odrv4
    port map (
            O => \N__39824\,
            I => \nx.n2509\
        );

    \I__8934\ : InMux
    port map (
            O => \N__39819\,
            I => \N__39816\
        );

    \I__8933\ : LocalMux
    port map (
            O => \N__39816\,
            I => \N__39813\
        );

    \I__8932\ : Odrv4
    port map (
            O => \N__39813\,
            I => \nx.n2576\
        );

    \I__8931\ : InMux
    port map (
            O => \N__39810\,
            I => \nx.n10938\
        );

    \I__8930\ : CascadeMux
    port map (
            O => \N__39807\,
            I => \N__39802\
        );

    \I__8929\ : InMux
    port map (
            O => \N__39806\,
            I => \N__39797\
        );

    \I__8928\ : InMux
    port map (
            O => \N__39805\,
            I => \N__39797\
        );

    \I__8927\ : InMux
    port map (
            O => \N__39802\,
            I => \N__39794\
        );

    \I__8926\ : LocalMux
    port map (
            O => \N__39797\,
            I => \nx.n2508\
        );

    \I__8925\ : LocalMux
    port map (
            O => \N__39794\,
            I => \nx.n2508\
        );

    \I__8924\ : CascadeMux
    port map (
            O => \N__39789\,
            I => \N__39786\
        );

    \I__8923\ : InMux
    port map (
            O => \N__39786\,
            I => \N__39783\
        );

    \I__8922\ : LocalMux
    port map (
            O => \N__39783\,
            I => \N__39780\
        );

    \I__8921\ : Odrv4
    port map (
            O => \N__39780\,
            I => \nx.n2575\
        );

    \I__8920\ : InMux
    port map (
            O => \N__39777\,
            I => \nx.n10939\
        );

    \I__8919\ : CascadeMux
    port map (
            O => \N__39774\,
            I => \N__39771\
        );

    \I__8918\ : InMux
    port map (
            O => \N__39771\,
            I => \N__39767\
        );

    \I__8917\ : InMux
    port map (
            O => \N__39770\,
            I => \N__39764\
        );

    \I__8916\ : LocalMux
    port map (
            O => \N__39767\,
            I => \N__39761\
        );

    \I__8915\ : LocalMux
    port map (
            O => \N__39764\,
            I => \N__39758\
        );

    \I__8914\ : Span4Mux_h
    port map (
            O => \N__39761\,
            I => \N__39755\
        );

    \I__8913\ : Span4Mux_v
    port map (
            O => \N__39758\,
            I => \N__39752\
        );

    \I__8912\ : Odrv4
    port map (
            O => \N__39755\,
            I => \nx.n2507\
        );

    \I__8911\ : Odrv4
    port map (
            O => \N__39752\,
            I => \nx.n2507\
        );

    \I__8910\ : InMux
    port map (
            O => \N__39747\,
            I => \N__39744\
        );

    \I__8909\ : LocalMux
    port map (
            O => \N__39744\,
            I => \N__39741\
        );

    \I__8908\ : Odrv4
    port map (
            O => \N__39741\,
            I => \nx.n2574\
        );

    \I__8907\ : InMux
    port map (
            O => \N__39738\,
            I => \nx.n10940\
        );

    \I__8906\ : CascadeMux
    port map (
            O => \N__39735\,
            I => \N__39732\
        );

    \I__8905\ : InMux
    port map (
            O => \N__39732\,
            I => \N__39728\
        );

    \I__8904\ : CascadeMux
    port map (
            O => \N__39731\,
            I => \N__39724\
        );

    \I__8903\ : LocalMux
    port map (
            O => \N__39728\,
            I => \N__39721\
        );

    \I__8902\ : InMux
    port map (
            O => \N__39727\,
            I => \N__39718\
        );

    \I__8901\ : InMux
    port map (
            O => \N__39724\,
            I => \N__39715\
        );

    \I__8900\ : Span4Mux_v
    port map (
            O => \N__39721\,
            I => \N__39710\
        );

    \I__8899\ : LocalMux
    port map (
            O => \N__39718\,
            I => \N__39710\
        );

    \I__8898\ : LocalMux
    port map (
            O => \N__39715\,
            I => \nx.n2598\
        );

    \I__8897\ : Odrv4
    port map (
            O => \N__39710\,
            I => \nx.n2598\
        );

    \I__8896\ : InMux
    port map (
            O => \N__39705\,
            I => \N__39702\
        );

    \I__8895\ : LocalMux
    port map (
            O => \N__39702\,
            I => \N__39699\
        );

    \I__8894\ : Span4Mux_v
    port map (
            O => \N__39699\,
            I => \N__39696\
        );

    \I__8893\ : Span4Mux_h
    port map (
            O => \N__39696\,
            I => \N__39693\
        );

    \I__8892\ : Odrv4
    port map (
            O => \N__39693\,
            I => \nx.n2665\
        );

    \I__8891\ : InMux
    port map (
            O => \N__39690\,
            I => \nx.n10970\
        );

    \I__8890\ : CascadeMux
    port map (
            O => \N__39687\,
            I => \N__39684\
        );

    \I__8889\ : InMux
    port map (
            O => \N__39684\,
            I => \N__39680\
        );

    \I__8888\ : InMux
    port map (
            O => \N__39683\,
            I => \N__39677\
        );

    \I__8887\ : LocalMux
    port map (
            O => \N__39680\,
            I => \N__39674\
        );

    \I__8886\ : LocalMux
    port map (
            O => \N__39677\,
            I => \nx.n2597\
        );

    \I__8885\ : Odrv12
    port map (
            O => \N__39674\,
            I => \nx.n2597\
        );

    \I__8884\ : CascadeMux
    port map (
            O => \N__39669\,
            I => \N__39666\
        );

    \I__8883\ : InMux
    port map (
            O => \N__39666\,
            I => \N__39663\
        );

    \I__8882\ : LocalMux
    port map (
            O => \N__39663\,
            I => \N__39660\
        );

    \I__8881\ : Span4Mux_v
    port map (
            O => \N__39660\,
            I => \N__39657\
        );

    \I__8880\ : Span4Mux_h
    port map (
            O => \N__39657\,
            I => \N__39654\
        );

    \I__8879\ : Odrv4
    port map (
            O => \N__39654\,
            I => \nx.n2664\
        );

    \I__8878\ : InMux
    port map (
            O => \N__39651\,
            I => \nx.n10971\
        );

    \I__8877\ : InMux
    port map (
            O => \N__39648\,
            I => \N__39645\
        );

    \I__8876\ : LocalMux
    port map (
            O => \N__39645\,
            I => \N__39640\
        );

    \I__8875\ : CascadeMux
    port map (
            O => \N__39644\,
            I => \N__39637\
        );

    \I__8874\ : InMux
    port map (
            O => \N__39643\,
            I => \N__39634\
        );

    \I__8873\ : Span4Mux_v
    port map (
            O => \N__39640\,
            I => \N__39631\
        );

    \I__8872\ : InMux
    port map (
            O => \N__39637\,
            I => \N__39628\
        );

    \I__8871\ : LocalMux
    port map (
            O => \N__39634\,
            I => \N__39625\
        );

    \I__8870\ : Odrv4
    port map (
            O => \N__39631\,
            I => \nx.n2596\
        );

    \I__8869\ : LocalMux
    port map (
            O => \N__39628\,
            I => \nx.n2596\
        );

    \I__8868\ : Odrv4
    port map (
            O => \N__39625\,
            I => \nx.n2596\
        );

    \I__8867\ : CascadeMux
    port map (
            O => \N__39618\,
            I => \N__39615\
        );

    \I__8866\ : InMux
    port map (
            O => \N__39615\,
            I => \N__39612\
        );

    \I__8865\ : LocalMux
    port map (
            O => \N__39612\,
            I => \N__39609\
        );

    \I__8864\ : Span4Mux_v
    port map (
            O => \N__39609\,
            I => \N__39606\
        );

    \I__8863\ : Odrv4
    port map (
            O => \N__39606\,
            I => \nx.n2663\
        );

    \I__8862\ : InMux
    port map (
            O => \N__39603\,
            I => \nx.n10972\
        );

    \I__8861\ : InMux
    port map (
            O => \N__39600\,
            I => \N__39596\
        );

    \I__8860\ : CascadeMux
    port map (
            O => \N__39599\,
            I => \N__39593\
        );

    \I__8859\ : LocalMux
    port map (
            O => \N__39596\,
            I => \N__39589\
        );

    \I__8858\ : InMux
    port map (
            O => \N__39593\,
            I => \N__39586\
        );

    \I__8857\ : InMux
    port map (
            O => \N__39592\,
            I => \N__39583\
        );

    \I__8856\ : Span4Mux_h
    port map (
            O => \N__39589\,
            I => \N__39580\
        );

    \I__8855\ : LocalMux
    port map (
            O => \N__39586\,
            I => \N__39577\
        );

    \I__8854\ : LocalMux
    port map (
            O => \N__39583\,
            I => \N__39574\
        );

    \I__8853\ : Odrv4
    port map (
            O => \N__39580\,
            I => \nx.n2595\
        );

    \I__8852\ : Odrv4
    port map (
            O => \N__39577\,
            I => \nx.n2595\
        );

    \I__8851\ : Odrv12
    port map (
            O => \N__39574\,
            I => \nx.n2595\
        );

    \I__8850\ : InMux
    port map (
            O => \N__39567\,
            I => \N__39564\
        );

    \I__8849\ : LocalMux
    port map (
            O => \N__39564\,
            I => \N__39561\
        );

    \I__8848\ : Span4Mux_h
    port map (
            O => \N__39561\,
            I => \N__39558\
        );

    \I__8847\ : Span4Mux_h
    port map (
            O => \N__39558\,
            I => \N__39555\
        );

    \I__8846\ : Odrv4
    port map (
            O => \N__39555\,
            I => \nx.n2662\
        );

    \I__8845\ : InMux
    port map (
            O => \N__39552\,
            I => \nx.n10973\
        );

    \I__8844\ : InMux
    port map (
            O => \N__39549\,
            I => \N__39546\
        );

    \I__8843\ : LocalMux
    port map (
            O => \N__39546\,
            I => \N__39542\
        );

    \I__8842\ : CascadeMux
    port map (
            O => \N__39545\,
            I => \N__39539\
        );

    \I__8841\ : Span4Mux_h
    port map (
            O => \N__39542\,
            I => \N__39535\
        );

    \I__8840\ : InMux
    port map (
            O => \N__39539\,
            I => \N__39532\
        );

    \I__8839\ : InMux
    port map (
            O => \N__39538\,
            I => \N__39529\
        );

    \I__8838\ : Odrv4
    port map (
            O => \N__39535\,
            I => \nx.n2594\
        );

    \I__8837\ : LocalMux
    port map (
            O => \N__39532\,
            I => \nx.n2594\
        );

    \I__8836\ : LocalMux
    port map (
            O => \N__39529\,
            I => \nx.n2594\
        );

    \I__8835\ : CascadeMux
    port map (
            O => \N__39522\,
            I => \N__39519\
        );

    \I__8834\ : InMux
    port map (
            O => \N__39519\,
            I => \N__39516\
        );

    \I__8833\ : LocalMux
    port map (
            O => \N__39516\,
            I => \N__39513\
        );

    \I__8832\ : Span4Mux_h
    port map (
            O => \N__39513\,
            I => \N__39510\
        );

    \I__8831\ : Span4Mux_h
    port map (
            O => \N__39510\,
            I => \N__39507\
        );

    \I__8830\ : Odrv4
    port map (
            O => \N__39507\,
            I => \nx.n2661\
        );

    \I__8829\ : InMux
    port map (
            O => \N__39504\,
            I => \bfn_16_23_0_\
        );

    \I__8828\ : CascadeMux
    port map (
            O => \N__39501\,
            I => \N__39498\
        );

    \I__8827\ : InMux
    port map (
            O => \N__39498\,
            I => \N__39495\
        );

    \I__8826\ : LocalMux
    port map (
            O => \N__39495\,
            I => \N__39491\
        );

    \I__8825\ : CascadeMux
    port map (
            O => \N__39494\,
            I => \N__39488\
        );

    \I__8824\ : Span4Mux_v
    port map (
            O => \N__39491\,
            I => \N__39484\
        );

    \I__8823\ : InMux
    port map (
            O => \N__39488\,
            I => \N__39481\
        );

    \I__8822\ : InMux
    port map (
            O => \N__39487\,
            I => \N__39478\
        );

    \I__8821\ : Odrv4
    port map (
            O => \N__39484\,
            I => \nx.n2593\
        );

    \I__8820\ : LocalMux
    port map (
            O => \N__39481\,
            I => \nx.n2593\
        );

    \I__8819\ : LocalMux
    port map (
            O => \N__39478\,
            I => \nx.n2593\
        );

    \I__8818\ : InMux
    port map (
            O => \N__39471\,
            I => \N__39468\
        );

    \I__8817\ : LocalMux
    port map (
            O => \N__39468\,
            I => \N__39465\
        );

    \I__8816\ : Span4Mux_h
    port map (
            O => \N__39465\,
            I => \N__39462\
        );

    \I__8815\ : Span4Mux_h
    port map (
            O => \N__39462\,
            I => \N__39459\
        );

    \I__8814\ : Odrv4
    port map (
            O => \N__39459\,
            I => \nx.n2660\
        );

    \I__8813\ : InMux
    port map (
            O => \N__39456\,
            I => \nx.n10975\
        );

    \I__8812\ : InMux
    port map (
            O => \N__39453\,
            I => \N__39449\
        );

    \I__8811\ : CascadeMux
    port map (
            O => \N__39452\,
            I => \N__39446\
        );

    \I__8810\ : LocalMux
    port map (
            O => \N__39449\,
            I => \N__39443\
        );

    \I__8809\ : InMux
    port map (
            O => \N__39446\,
            I => \N__39440\
        );

    \I__8808\ : Odrv12
    port map (
            O => \N__39443\,
            I => \nx.n2592\
        );

    \I__8807\ : LocalMux
    port map (
            O => \N__39440\,
            I => \nx.n2592\
        );

    \I__8806\ : CascadeMux
    port map (
            O => \N__39435\,
            I => \N__39432\
        );

    \I__8805\ : InMux
    port map (
            O => \N__39432\,
            I => \N__39429\
        );

    \I__8804\ : LocalMux
    port map (
            O => \N__39429\,
            I => \N__39426\
        );

    \I__8803\ : Span4Mux_v
    port map (
            O => \N__39426\,
            I => \N__39423\
        );

    \I__8802\ : Span4Mux_h
    port map (
            O => \N__39423\,
            I => \N__39420\
        );

    \I__8801\ : Odrv4
    port map (
            O => \N__39420\,
            I => \nx.n2659\
        );

    \I__8800\ : InMux
    port map (
            O => \N__39417\,
            I => \nx.n10976\
        );

    \I__8799\ : CascadeMux
    port map (
            O => \N__39414\,
            I => \N__39411\
        );

    \I__8798\ : InMux
    port map (
            O => \N__39411\,
            I => \N__39407\
        );

    \I__8797\ : CascadeMux
    port map (
            O => \N__39410\,
            I => \N__39404\
        );

    \I__8796\ : LocalMux
    port map (
            O => \N__39407\,
            I => \N__39401\
        );

    \I__8795\ : InMux
    port map (
            O => \N__39404\,
            I => \N__39397\
        );

    \I__8794\ : Span4Mux_h
    port map (
            O => \N__39401\,
            I => \N__39394\
        );

    \I__8793\ : InMux
    port map (
            O => \N__39400\,
            I => \N__39391\
        );

    \I__8792\ : LocalMux
    port map (
            O => \N__39397\,
            I => \nx.n2591\
        );

    \I__8791\ : Odrv4
    port map (
            O => \N__39394\,
            I => \nx.n2591\
        );

    \I__8790\ : LocalMux
    port map (
            O => \N__39391\,
            I => \nx.n2591\
        );

    \I__8789\ : InMux
    port map (
            O => \N__39384\,
            I => \N__39381\
        );

    \I__8788\ : LocalMux
    port map (
            O => \N__39381\,
            I => \N__39378\
        );

    \I__8787\ : Odrv12
    port map (
            O => \N__39378\,
            I => \nx.n2658\
        );

    \I__8786\ : InMux
    port map (
            O => \N__39375\,
            I => \nx.n10977\
        );

    \I__8785\ : InMux
    port map (
            O => \N__39372\,
            I => \N__39369\
        );

    \I__8784\ : LocalMux
    port map (
            O => \N__39369\,
            I => \N__39365\
        );

    \I__8783\ : CascadeMux
    port map (
            O => \N__39368\,
            I => \N__39362\
        );

    \I__8782\ : Span4Mux_v
    port map (
            O => \N__39365\,
            I => \N__39359\
        );

    \I__8781\ : InMux
    port map (
            O => \N__39362\,
            I => \N__39356\
        );

    \I__8780\ : Odrv4
    port map (
            O => \N__39359\,
            I => \nx.n2606\
        );

    \I__8779\ : LocalMux
    port map (
            O => \N__39356\,
            I => \nx.n2606\
        );

    \I__8778\ : InMux
    port map (
            O => \N__39351\,
            I => \N__39348\
        );

    \I__8777\ : LocalMux
    port map (
            O => \N__39348\,
            I => \nx.n2673\
        );

    \I__8776\ : InMux
    port map (
            O => \N__39345\,
            I => \nx.n10962\
        );

    \I__8775\ : InMux
    port map (
            O => \N__39342\,
            I => \N__39339\
        );

    \I__8774\ : LocalMux
    port map (
            O => \N__39339\,
            I => \N__39334\
        );

    \I__8773\ : CascadeMux
    port map (
            O => \N__39338\,
            I => \N__39331\
        );

    \I__8772\ : InMux
    port map (
            O => \N__39337\,
            I => \N__39328\
        );

    \I__8771\ : Span4Mux_v
    port map (
            O => \N__39334\,
            I => \N__39325\
        );

    \I__8770\ : InMux
    port map (
            O => \N__39331\,
            I => \N__39322\
        );

    \I__8769\ : LocalMux
    port map (
            O => \N__39328\,
            I => \nx.n2605\
        );

    \I__8768\ : Odrv4
    port map (
            O => \N__39325\,
            I => \nx.n2605\
        );

    \I__8767\ : LocalMux
    port map (
            O => \N__39322\,
            I => \nx.n2605\
        );

    \I__8766\ : InMux
    port map (
            O => \N__39315\,
            I => \N__39312\
        );

    \I__8765\ : LocalMux
    port map (
            O => \N__39312\,
            I => \nx.n2672\
        );

    \I__8764\ : InMux
    port map (
            O => \N__39309\,
            I => \nx.n10963\
        );

    \I__8763\ : CascadeMux
    port map (
            O => \N__39306\,
            I => \N__39301\
        );

    \I__8762\ : CascadeMux
    port map (
            O => \N__39305\,
            I => \N__39298\
        );

    \I__8761\ : InMux
    port map (
            O => \N__39304\,
            I => \N__39295\
        );

    \I__8760\ : InMux
    port map (
            O => \N__39301\,
            I => \N__39292\
        );

    \I__8759\ : InMux
    port map (
            O => \N__39298\,
            I => \N__39289\
        );

    \I__8758\ : LocalMux
    port map (
            O => \N__39295\,
            I => \N__39284\
        );

    \I__8757\ : LocalMux
    port map (
            O => \N__39292\,
            I => \N__39284\
        );

    \I__8756\ : LocalMux
    port map (
            O => \N__39289\,
            I => \N__39281\
        );

    \I__8755\ : Span4Mux_h
    port map (
            O => \N__39284\,
            I => \N__39278\
        );

    \I__8754\ : Odrv4
    port map (
            O => \N__39281\,
            I => \nx.n2604\
        );

    \I__8753\ : Odrv4
    port map (
            O => \N__39278\,
            I => \nx.n2604\
        );

    \I__8752\ : CascadeMux
    port map (
            O => \N__39273\,
            I => \N__39270\
        );

    \I__8751\ : InMux
    port map (
            O => \N__39270\,
            I => \N__39267\
        );

    \I__8750\ : LocalMux
    port map (
            O => \N__39267\,
            I => \N__39264\
        );

    \I__8749\ : Odrv4
    port map (
            O => \N__39264\,
            I => \nx.n2671\
        );

    \I__8748\ : InMux
    port map (
            O => \N__39261\,
            I => \nx.n10964\
        );

    \I__8747\ : CascadeMux
    port map (
            O => \N__39258\,
            I => \N__39255\
        );

    \I__8746\ : InMux
    port map (
            O => \N__39255\,
            I => \N__39252\
        );

    \I__8745\ : LocalMux
    port map (
            O => \N__39252\,
            I => \N__39248\
        );

    \I__8744\ : InMux
    port map (
            O => \N__39251\,
            I => \N__39245\
        );

    \I__8743\ : Span4Mux_v
    port map (
            O => \N__39248\,
            I => \N__39242\
        );

    \I__8742\ : LocalMux
    port map (
            O => \N__39245\,
            I => \nx.n2603\
        );

    \I__8741\ : Odrv4
    port map (
            O => \N__39242\,
            I => \nx.n2603\
        );

    \I__8740\ : InMux
    port map (
            O => \N__39237\,
            I => \N__39234\
        );

    \I__8739\ : LocalMux
    port map (
            O => \N__39234\,
            I => \N__39231\
        );

    \I__8738\ : Span4Mux_h
    port map (
            O => \N__39231\,
            I => \N__39228\
        );

    \I__8737\ : Odrv4
    port map (
            O => \N__39228\,
            I => \nx.n2670\
        );

    \I__8736\ : InMux
    port map (
            O => \N__39225\,
            I => \nx.n10965\
        );

    \I__8735\ : CascadeMux
    port map (
            O => \N__39222\,
            I => \N__39218\
        );

    \I__8734\ : InMux
    port map (
            O => \N__39221\,
            I => \N__39215\
        );

    \I__8733\ : InMux
    port map (
            O => \N__39218\,
            I => \N__39211\
        );

    \I__8732\ : LocalMux
    port map (
            O => \N__39215\,
            I => \N__39208\
        );

    \I__8731\ : InMux
    port map (
            O => \N__39214\,
            I => \N__39205\
        );

    \I__8730\ : LocalMux
    port map (
            O => \N__39211\,
            I => \N__39202\
        );

    \I__8729\ : Odrv4
    port map (
            O => \N__39208\,
            I => \nx.n2602\
        );

    \I__8728\ : LocalMux
    port map (
            O => \N__39205\,
            I => \nx.n2602\
        );

    \I__8727\ : Odrv12
    port map (
            O => \N__39202\,
            I => \nx.n2602\
        );

    \I__8726\ : InMux
    port map (
            O => \N__39195\,
            I => \N__39192\
        );

    \I__8725\ : LocalMux
    port map (
            O => \N__39192\,
            I => \N__39189\
        );

    \I__8724\ : Span4Mux_v
    port map (
            O => \N__39189\,
            I => \N__39186\
        );

    \I__8723\ : Span4Mux_h
    port map (
            O => \N__39186\,
            I => \N__39183\
        );

    \I__8722\ : Odrv4
    port map (
            O => \N__39183\,
            I => \nx.n2669\
        );

    \I__8721\ : InMux
    port map (
            O => \N__39180\,
            I => \bfn_16_22_0_\
        );

    \I__8720\ : CascadeMux
    port map (
            O => \N__39177\,
            I => \N__39174\
        );

    \I__8719\ : InMux
    port map (
            O => \N__39174\,
            I => \N__39170\
        );

    \I__8718\ : InMux
    port map (
            O => \N__39173\,
            I => \N__39166\
        );

    \I__8717\ : LocalMux
    port map (
            O => \N__39170\,
            I => \N__39163\
        );

    \I__8716\ : InMux
    port map (
            O => \N__39169\,
            I => \N__39160\
        );

    \I__8715\ : LocalMux
    port map (
            O => \N__39166\,
            I => \nx.n2601\
        );

    \I__8714\ : Odrv4
    port map (
            O => \N__39163\,
            I => \nx.n2601\
        );

    \I__8713\ : LocalMux
    port map (
            O => \N__39160\,
            I => \nx.n2601\
        );

    \I__8712\ : CascadeMux
    port map (
            O => \N__39153\,
            I => \N__39150\
        );

    \I__8711\ : InMux
    port map (
            O => \N__39150\,
            I => \N__39147\
        );

    \I__8710\ : LocalMux
    port map (
            O => \N__39147\,
            I => \N__39144\
        );

    \I__8709\ : Odrv12
    port map (
            O => \N__39144\,
            I => \nx.n2668\
        );

    \I__8708\ : InMux
    port map (
            O => \N__39141\,
            I => \nx.n10967\
        );

    \I__8707\ : InMux
    port map (
            O => \N__39138\,
            I => \N__39134\
        );

    \I__8706\ : CascadeMux
    port map (
            O => \N__39137\,
            I => \N__39131\
        );

    \I__8705\ : LocalMux
    port map (
            O => \N__39134\,
            I => \N__39128\
        );

    \I__8704\ : InMux
    port map (
            O => \N__39131\,
            I => \N__39125\
        );

    \I__8703\ : Span4Mux_h
    port map (
            O => \N__39128\,
            I => \N__39121\
        );

    \I__8702\ : LocalMux
    port map (
            O => \N__39125\,
            I => \N__39118\
        );

    \I__8701\ : InMux
    port map (
            O => \N__39124\,
            I => \N__39115\
        );

    \I__8700\ : Odrv4
    port map (
            O => \N__39121\,
            I => \nx.n2600\
        );

    \I__8699\ : Odrv4
    port map (
            O => \N__39118\,
            I => \nx.n2600\
        );

    \I__8698\ : LocalMux
    port map (
            O => \N__39115\,
            I => \nx.n2600\
        );

    \I__8697\ : CascadeMux
    port map (
            O => \N__39108\,
            I => \N__39105\
        );

    \I__8696\ : InMux
    port map (
            O => \N__39105\,
            I => \N__39102\
        );

    \I__8695\ : LocalMux
    port map (
            O => \N__39102\,
            I => \N__39099\
        );

    \I__8694\ : Span4Mux_v
    port map (
            O => \N__39099\,
            I => \N__39096\
        );

    \I__8693\ : Span4Mux_h
    port map (
            O => \N__39096\,
            I => \N__39093\
        );

    \I__8692\ : Odrv4
    port map (
            O => \N__39093\,
            I => \nx.n2667\
        );

    \I__8691\ : InMux
    port map (
            O => \N__39090\,
            I => \nx.n10968\
        );

    \I__8690\ : CascadeMux
    port map (
            O => \N__39087\,
            I => \N__39083\
        );

    \I__8689\ : InMux
    port map (
            O => \N__39086\,
            I => \N__39080\
        );

    \I__8688\ : InMux
    port map (
            O => \N__39083\,
            I => \N__39076\
        );

    \I__8687\ : LocalMux
    port map (
            O => \N__39080\,
            I => \N__39073\
        );

    \I__8686\ : InMux
    port map (
            O => \N__39079\,
            I => \N__39070\
        );

    \I__8685\ : LocalMux
    port map (
            O => \N__39076\,
            I => \N__39067\
        );

    \I__8684\ : Span4Mux_v
    port map (
            O => \N__39073\,
            I => \N__39062\
        );

    \I__8683\ : LocalMux
    port map (
            O => \N__39070\,
            I => \N__39062\
        );

    \I__8682\ : Odrv4
    port map (
            O => \N__39067\,
            I => \nx.n2599\
        );

    \I__8681\ : Odrv4
    port map (
            O => \N__39062\,
            I => \nx.n2599\
        );

    \I__8680\ : InMux
    port map (
            O => \N__39057\,
            I => \N__39054\
        );

    \I__8679\ : LocalMux
    port map (
            O => \N__39054\,
            I => \N__39051\
        );

    \I__8678\ : Span4Mux_v
    port map (
            O => \N__39051\,
            I => \N__39048\
        );

    \I__8677\ : Span4Mux_h
    port map (
            O => \N__39048\,
            I => \N__39045\
        );

    \I__8676\ : Odrv4
    port map (
            O => \N__39045\,
            I => \nx.n2666\
        );

    \I__8675\ : InMux
    port map (
            O => \N__39042\,
            I => \nx.n10969\
        );

    \I__8674\ : CascadeMux
    port map (
            O => \N__39039\,
            I => \n7_adj_840_cascade_\
        );

    \I__8673\ : IoInMux
    port map (
            O => \N__39036\,
            I => \N__39033\
        );

    \I__8672\ : LocalMux
    port map (
            O => \N__39033\,
            I => \N__39030\
        );

    \I__8671\ : IoSpan4Mux
    port map (
            O => \N__39030\,
            I => \N__39027\
        );

    \I__8670\ : Span4Mux_s2_v
    port map (
            O => \N__39027\,
            I => \N__39024\
        );

    \I__8669\ : Sp12to4
    port map (
            O => \N__39024\,
            I => \N__39021\
        );

    \I__8668\ : Span12Mux_h
    port map (
            O => \N__39021\,
            I => \N__39016\
        );

    \I__8667\ : InMux
    port map (
            O => \N__39020\,
            I => \N__39013\
        );

    \I__8666\ : InMux
    port map (
            O => \N__39019\,
            I => \N__39010\
        );

    \I__8665\ : Odrv12
    port map (
            O => \N__39016\,
            I => pin_out_0
        );

    \I__8664\ : LocalMux
    port map (
            O => \N__39013\,
            I => pin_out_0
        );

    \I__8663\ : LocalMux
    port map (
            O => \N__39010\,
            I => pin_out_0
        );

    \I__8662\ : InMux
    port map (
            O => \N__39003\,
            I => \N__39000\
        );

    \I__8661\ : LocalMux
    port map (
            O => \N__39000\,
            I => n8_adj_817
        );

    \I__8660\ : IoInMux
    port map (
            O => \N__38997\,
            I => \N__38994\
        );

    \I__8659\ : LocalMux
    port map (
            O => \N__38994\,
            I => \N__38991\
        );

    \I__8658\ : IoSpan4Mux
    port map (
            O => \N__38991\,
            I => \N__38988\
        );

    \I__8657\ : Span4Mux_s2_v
    port map (
            O => \N__38988\,
            I => \N__38985\
        );

    \I__8656\ : Sp12to4
    port map (
            O => \N__38985\,
            I => \N__38982\
        );

    \I__8655\ : Span12Mux_s8_v
    port map (
            O => \N__38982\,
            I => \N__38979\
        );

    \I__8654\ : Span12Mux_h
    port map (
            O => \N__38979\,
            I => \N__38974\
        );

    \I__8653\ : InMux
    port map (
            O => \N__38978\,
            I => \N__38969\
        );

    \I__8652\ : InMux
    port map (
            O => \N__38977\,
            I => \N__38969\
        );

    \I__8651\ : Odrv12
    port map (
            O => \N__38974\,
            I => pin_out_1
        );

    \I__8650\ : LocalMux
    port map (
            O => \N__38969\,
            I => pin_out_1
        );

    \I__8649\ : InMux
    port map (
            O => \N__38964\,
            I => \N__38961\
        );

    \I__8648\ : LocalMux
    port map (
            O => \N__38961\,
            I => \N__38958\
        );

    \I__8647\ : Span12Mux_v
    port map (
            O => \N__38958\,
            I => \N__38955\
        );

    \I__8646\ : Odrv12
    port map (
            O => \N__38955\,
            I => n11952
        );

    \I__8645\ : IoInMux
    port map (
            O => \N__38952\,
            I => \N__38949\
        );

    \I__8644\ : LocalMux
    port map (
            O => \N__38949\,
            I => \N__38946\
        );

    \I__8643\ : Span12Mux_s5_v
    port map (
            O => \N__38946\,
            I => \N__38943\
        );

    \I__8642\ : Span12Mux_h
    port map (
            O => \N__38943\,
            I => \N__38939\
        );

    \I__8641\ : InMux
    port map (
            O => \N__38942\,
            I => \N__38936\
        );

    \I__8640\ : Odrv12
    port map (
            O => \N__38939\,
            I => pin_oe_8
        );

    \I__8639\ : LocalMux
    port map (
            O => \N__38936\,
            I => pin_oe_8
        );

    \I__8638\ : InMux
    port map (
            O => \N__38931\,
            I => \N__38928\
        );

    \I__8637\ : LocalMux
    port map (
            O => \N__38928\,
            I => \N__38924\
        );

    \I__8636\ : InMux
    port map (
            O => \N__38927\,
            I => \N__38921\
        );

    \I__8635\ : Span4Mux_v
    port map (
            O => \N__38924\,
            I => \N__38917\
        );

    \I__8634\ : LocalMux
    port map (
            O => \N__38921\,
            I => \N__38914\
        );

    \I__8633\ : InMux
    port map (
            O => \N__38920\,
            I => \N__38909\
        );

    \I__8632\ : Span4Mux_h
    port map (
            O => \N__38917\,
            I => \N__38906\
        );

    \I__8631\ : Span4Mux_v
    port map (
            O => \N__38914\,
            I => \N__38903\
        );

    \I__8630\ : InMux
    port map (
            O => \N__38913\,
            I => \N__38900\
        );

    \I__8629\ : InMux
    port map (
            O => \N__38912\,
            I => \N__38897\
        );

    \I__8628\ : LocalMux
    port map (
            O => \N__38909\,
            I => \N__38890\
        );

    \I__8627\ : Sp12to4
    port map (
            O => \N__38906\,
            I => \N__38890\
        );

    \I__8626\ : Sp12to4
    port map (
            O => \N__38903\,
            I => \N__38890\
        );

    \I__8625\ : LocalMux
    port map (
            O => \N__38900\,
            I => \nx.bit_ctr_9\
        );

    \I__8624\ : LocalMux
    port map (
            O => \N__38897\,
            I => \nx.bit_ctr_9\
        );

    \I__8623\ : Odrv12
    port map (
            O => \N__38890\,
            I => \nx.bit_ctr_9\
        );

    \I__8622\ : InMux
    port map (
            O => \N__38883\,
            I => \N__38880\
        );

    \I__8621\ : LocalMux
    port map (
            O => \N__38880\,
            I => \N__38877\
        );

    \I__8620\ : Span4Mux_v
    port map (
            O => \N__38877\,
            I => \N__38874\
        );

    \I__8619\ : Span4Mux_h
    port map (
            O => \N__38874\,
            I => \N__38871\
        );

    \I__8618\ : Odrv4
    port map (
            O => \N__38871\,
            I => \nx.n2677\
        );

    \I__8617\ : InMux
    port map (
            O => \N__38868\,
            I => \bfn_16_21_0_\
        );

    \I__8616\ : InMux
    port map (
            O => \N__38865\,
            I => \N__38862\
        );

    \I__8615\ : LocalMux
    port map (
            O => \N__38862\,
            I => \N__38858\
        );

    \I__8614\ : CascadeMux
    port map (
            O => \N__38861\,
            I => \N__38855\
        );

    \I__8613\ : Span4Mux_h
    port map (
            O => \N__38858\,
            I => \N__38852\
        );

    \I__8612\ : InMux
    port map (
            O => \N__38855\,
            I => \N__38849\
        );

    \I__8611\ : Odrv4
    port map (
            O => \N__38852\,
            I => \nx.n2609\
        );

    \I__8610\ : LocalMux
    port map (
            O => \N__38849\,
            I => \nx.n2609\
        );

    \I__8609\ : InMux
    port map (
            O => \N__38844\,
            I => \N__38841\
        );

    \I__8608\ : LocalMux
    port map (
            O => \N__38841\,
            I => \N__38838\
        );

    \I__8607\ : Span4Mux_h
    port map (
            O => \N__38838\,
            I => \N__38835\
        );

    \I__8606\ : Odrv4
    port map (
            O => \N__38835\,
            I => \nx.n2676\
        );

    \I__8605\ : InMux
    port map (
            O => \N__38832\,
            I => \nx.n10959\
        );

    \I__8604\ : InMux
    port map (
            O => \N__38829\,
            I => \N__38826\
        );

    \I__8603\ : LocalMux
    port map (
            O => \N__38826\,
            I => \N__38822\
        );

    \I__8602\ : CascadeMux
    port map (
            O => \N__38825\,
            I => \N__38818\
        );

    \I__8601\ : Span4Mux_h
    port map (
            O => \N__38822\,
            I => \N__38815\
        );

    \I__8600\ : InMux
    port map (
            O => \N__38821\,
            I => \N__38812\
        );

    \I__8599\ : InMux
    port map (
            O => \N__38818\,
            I => \N__38809\
        );

    \I__8598\ : Odrv4
    port map (
            O => \N__38815\,
            I => \nx.n2608\
        );

    \I__8597\ : LocalMux
    port map (
            O => \N__38812\,
            I => \nx.n2608\
        );

    \I__8596\ : LocalMux
    port map (
            O => \N__38809\,
            I => \nx.n2608\
        );

    \I__8595\ : CascadeMux
    port map (
            O => \N__38802\,
            I => \N__38799\
        );

    \I__8594\ : InMux
    port map (
            O => \N__38799\,
            I => \N__38796\
        );

    \I__8593\ : LocalMux
    port map (
            O => \N__38796\,
            I => \N__38793\
        );

    \I__8592\ : Span4Mux_v
    port map (
            O => \N__38793\,
            I => \N__38790\
        );

    \I__8591\ : Odrv4
    port map (
            O => \N__38790\,
            I => \nx.n2675\
        );

    \I__8590\ : InMux
    port map (
            O => \N__38787\,
            I => \nx.n10960\
        );

    \I__8589\ : InMux
    port map (
            O => \N__38784\,
            I => \N__38781\
        );

    \I__8588\ : LocalMux
    port map (
            O => \N__38781\,
            I => \N__38777\
        );

    \I__8587\ : CascadeMux
    port map (
            O => \N__38780\,
            I => \N__38774\
        );

    \I__8586\ : Span4Mux_h
    port map (
            O => \N__38777\,
            I => \N__38770\
        );

    \I__8585\ : InMux
    port map (
            O => \N__38774\,
            I => \N__38767\
        );

    \I__8584\ : InMux
    port map (
            O => \N__38773\,
            I => \N__38764\
        );

    \I__8583\ : Odrv4
    port map (
            O => \N__38770\,
            I => \nx.n2607\
        );

    \I__8582\ : LocalMux
    port map (
            O => \N__38767\,
            I => \nx.n2607\
        );

    \I__8581\ : LocalMux
    port map (
            O => \N__38764\,
            I => \nx.n2607\
        );

    \I__8580\ : CascadeMux
    port map (
            O => \N__38757\,
            I => \N__38754\
        );

    \I__8579\ : InMux
    port map (
            O => \N__38754\,
            I => \N__38751\
        );

    \I__8578\ : LocalMux
    port map (
            O => \N__38751\,
            I => \N__38748\
        );

    \I__8577\ : Span4Mux_v
    port map (
            O => \N__38748\,
            I => \N__38745\
        );

    \I__8576\ : Span4Mux_h
    port map (
            O => \N__38745\,
            I => \N__38742\
        );

    \I__8575\ : Odrv4
    port map (
            O => \N__38742\,
            I => \nx.n2674\
        );

    \I__8574\ : InMux
    port map (
            O => \N__38739\,
            I => \nx.n10961\
        );

    \I__8573\ : CascadeMux
    port map (
            O => \N__38736\,
            I => \n9488_cascade_\
        );

    \I__8572\ : CascadeMux
    port map (
            O => \N__38733\,
            I => \n7_adj_818_cascade_\
        );

    \I__8571\ : CascadeMux
    port map (
            O => \N__38730\,
            I => \N__38727\
        );

    \I__8570\ : InMux
    port map (
            O => \N__38727\,
            I => \N__38724\
        );

    \I__8569\ : LocalMux
    port map (
            O => \N__38724\,
            I => n7_adj_821
        );

    \I__8568\ : IoInMux
    port map (
            O => \N__38721\,
            I => \N__38718\
        );

    \I__8567\ : LocalMux
    port map (
            O => \N__38718\,
            I => \N__38715\
        );

    \I__8566\ : Span12Mux_s3_h
    port map (
            O => \N__38715\,
            I => \N__38712\
        );

    \I__8565\ : Span12Mux_v
    port map (
            O => \N__38712\,
            I => \N__38708\
        );

    \I__8564\ : InMux
    port map (
            O => \N__38711\,
            I => \N__38704\
        );

    \I__8563\ : Span12Mux_h
    port map (
            O => \N__38708\,
            I => \N__38701\
        );

    \I__8562\ : InMux
    port map (
            O => \N__38707\,
            I => \N__38698\
        );

    \I__8561\ : LocalMux
    port map (
            O => \N__38704\,
            I => \N__38695\
        );

    \I__8560\ : Odrv12
    port map (
            O => \N__38701\,
            I => pin_out_3
        );

    \I__8559\ : LocalMux
    port map (
            O => \N__38698\,
            I => pin_out_3
        );

    \I__8558\ : Odrv4
    port map (
            O => \N__38695\,
            I => pin_out_3
        );

    \I__8557\ : IoInMux
    port map (
            O => \N__38688\,
            I => \N__38685\
        );

    \I__8556\ : LocalMux
    port map (
            O => \N__38685\,
            I => \N__38682\
        );

    \I__8555\ : Span4Mux_s3_h
    port map (
            O => \N__38682\,
            I => \N__38679\
        );

    \I__8554\ : Span4Mux_h
    port map (
            O => \N__38679\,
            I => \N__38676\
        );

    \I__8553\ : Span4Mux_h
    port map (
            O => \N__38676\,
            I => \N__38673\
        );

    \I__8552\ : Span4Mux_h
    port map (
            O => \N__38673\,
            I => \N__38668\
        );

    \I__8551\ : InMux
    port map (
            O => \N__38672\,
            I => \N__38665\
        );

    \I__8550\ : InMux
    port map (
            O => \N__38671\,
            I => \N__38662\
        );

    \I__8549\ : Odrv4
    port map (
            O => \N__38668\,
            I => pin_out_2
        );

    \I__8548\ : LocalMux
    port map (
            O => \N__38665\,
            I => pin_out_2
        );

    \I__8547\ : LocalMux
    port map (
            O => \N__38662\,
            I => pin_out_2
        );

    \I__8546\ : CascadeMux
    port map (
            O => \N__38655\,
            I => \n13355_cascade_\
        );

    \I__8545\ : InMux
    port map (
            O => \N__38652\,
            I => \N__38649\
        );

    \I__8544\ : LocalMux
    port map (
            O => \N__38649\,
            I => n13354
        );

    \I__8543\ : InMux
    port map (
            O => \N__38646\,
            I => \N__38643\
        );

    \I__8542\ : LocalMux
    port map (
            O => \N__38643\,
            I => n9
        );

    \I__8541\ : CascadeMux
    port map (
            O => \N__38640\,
            I => \n9_cascade_\
        );

    \I__8540\ : CascadeMux
    port map (
            O => \N__38637\,
            I => \n8_adj_820_cascade_\
        );

    \I__8539\ : CascadeMux
    port map (
            O => \N__38634\,
            I => \n6_adj_805_cascade_\
        );

    \I__8538\ : InMux
    port map (
            O => \N__38631\,
            I => \N__38628\
        );

    \I__8537\ : LocalMux
    port map (
            O => \N__38628\,
            I => \N__38624\
        );

    \I__8536\ : InMux
    port map (
            O => \N__38627\,
            I => \N__38621\
        );

    \I__8535\ : Odrv12
    port map (
            O => \N__38624\,
            I => n1788
        );

    \I__8534\ : LocalMux
    port map (
            O => \N__38621\,
            I => n1788
        );

    \I__8533\ : IoInMux
    port map (
            O => \N__38616\,
            I => \N__38613\
        );

    \I__8532\ : LocalMux
    port map (
            O => \N__38613\,
            I => \N__38610\
        );

    \I__8531\ : Span4Mux_s3_v
    port map (
            O => \N__38610\,
            I => \N__38607\
        );

    \I__8530\ : Span4Mux_h
    port map (
            O => \N__38607\,
            I => \N__38604\
        );

    \I__8529\ : Span4Mux_v
    port map (
            O => \N__38604\,
            I => \N__38600\
        );

    \I__8528\ : InMux
    port map (
            O => \N__38603\,
            I => \N__38597\
        );

    \I__8527\ : Odrv4
    port map (
            O => \N__38600\,
            I => pin_oe_22
        );

    \I__8526\ : LocalMux
    port map (
            O => \N__38597\,
            I => pin_oe_22
        );

    \I__8525\ : InMux
    port map (
            O => \N__38592\,
            I => \N__38588\
        );

    \I__8524\ : CascadeMux
    port map (
            O => \N__38591\,
            I => \N__38585\
        );

    \I__8523\ : LocalMux
    port map (
            O => \N__38588\,
            I => \N__38582\
        );

    \I__8522\ : InMux
    port map (
            O => \N__38585\,
            I => \N__38579\
        );

    \I__8521\ : Span4Mux_v
    port map (
            O => \N__38582\,
            I => \N__38574\
        );

    \I__8520\ : LocalMux
    port map (
            O => \N__38579\,
            I => \N__38574\
        );

    \I__8519\ : Span4Mux_h
    port map (
            O => \N__38574\,
            I => \N__38570\
        );

    \I__8518\ : InMux
    port map (
            O => \N__38573\,
            I => \N__38567\
        );

    \I__8517\ : Odrv4
    port map (
            O => \N__38570\,
            I => \nx.n2392\
        );

    \I__8516\ : LocalMux
    port map (
            O => \N__38567\,
            I => \nx.n2392\
        );

    \I__8515\ : CascadeMux
    port map (
            O => \N__38562\,
            I => \N__38559\
        );

    \I__8514\ : InMux
    port map (
            O => \N__38559\,
            I => \N__38556\
        );

    \I__8513\ : LocalMux
    port map (
            O => \N__38556\,
            I => \nx.n2459\
        );

    \I__8512\ : CascadeMux
    port map (
            O => \N__38553\,
            I => \nx.n2491_cascade_\
        );

    \I__8511\ : InMux
    port map (
            O => \N__38550\,
            I => \N__38547\
        );

    \I__8510\ : LocalMux
    port map (
            O => \N__38547\,
            I => \N__38544\
        );

    \I__8509\ : Odrv12
    port map (
            O => \N__38544\,
            I => \nx.n33_adj_767\
        );

    \I__8508\ : InMux
    port map (
            O => \N__38541\,
            I => \N__38538\
        );

    \I__8507\ : LocalMux
    port map (
            O => \N__38538\,
            I => \nx.n2460\
        );

    \I__8506\ : CascadeMux
    port map (
            O => \N__38535\,
            I => \N__38532\
        );

    \I__8505\ : InMux
    port map (
            O => \N__38532\,
            I => \N__38528\
        );

    \I__8504\ : CascadeMux
    port map (
            O => \N__38531\,
            I => \N__38525\
        );

    \I__8503\ : LocalMux
    port map (
            O => \N__38528\,
            I => \N__38522\
        );

    \I__8502\ : InMux
    port map (
            O => \N__38525\,
            I => \N__38519\
        );

    \I__8501\ : Span4Mux_h
    port map (
            O => \N__38522\,
            I => \N__38513\
        );

    \I__8500\ : LocalMux
    port map (
            O => \N__38519\,
            I => \N__38513\
        );

    \I__8499\ : InMux
    port map (
            O => \N__38518\,
            I => \N__38510\
        );

    \I__8498\ : Odrv4
    port map (
            O => \N__38513\,
            I => \nx.n2393\
        );

    \I__8497\ : LocalMux
    port map (
            O => \N__38510\,
            I => \nx.n2393\
        );

    \I__8496\ : CascadeMux
    port map (
            O => \N__38505\,
            I => \N__38493\
        );

    \I__8495\ : CascadeMux
    port map (
            O => \N__38504\,
            I => \N__38489\
        );

    \I__8494\ : InMux
    port map (
            O => \N__38503\,
            I => \N__38482\
        );

    \I__8493\ : InMux
    port map (
            O => \N__38502\,
            I => \N__38482\
        );

    \I__8492\ : InMux
    port map (
            O => \N__38501\,
            I => \N__38479\
        );

    \I__8491\ : InMux
    port map (
            O => \N__38500\,
            I => \N__38475\
        );

    \I__8490\ : CascadeMux
    port map (
            O => \N__38499\,
            I => \N__38471\
        );

    \I__8489\ : CascadeMux
    port map (
            O => \N__38498\,
            I => \N__38466\
        );

    \I__8488\ : CascadeMux
    port map (
            O => \N__38497\,
            I => \N__38462\
        );

    \I__8487\ : CascadeMux
    port map (
            O => \N__38496\,
            I => \N__38457\
        );

    \I__8486\ : InMux
    port map (
            O => \N__38493\,
            I => \N__38445\
        );

    \I__8485\ : InMux
    port map (
            O => \N__38492\,
            I => \N__38445\
        );

    \I__8484\ : InMux
    port map (
            O => \N__38489\,
            I => \N__38445\
        );

    \I__8483\ : InMux
    port map (
            O => \N__38488\,
            I => \N__38445\
        );

    \I__8482\ : InMux
    port map (
            O => \N__38487\,
            I => \N__38445\
        );

    \I__8481\ : LocalMux
    port map (
            O => \N__38482\,
            I => \N__38440\
        );

    \I__8480\ : LocalMux
    port map (
            O => \N__38479\,
            I => \N__38440\
        );

    \I__8479\ : InMux
    port map (
            O => \N__38478\,
            I => \N__38437\
        );

    \I__8478\ : LocalMux
    port map (
            O => \N__38475\,
            I => \N__38434\
        );

    \I__8477\ : InMux
    port map (
            O => \N__38474\,
            I => \N__38431\
        );

    \I__8476\ : InMux
    port map (
            O => \N__38471\,
            I => \N__38424\
        );

    \I__8475\ : InMux
    port map (
            O => \N__38470\,
            I => \N__38424\
        );

    \I__8474\ : InMux
    port map (
            O => \N__38469\,
            I => \N__38424\
        );

    \I__8473\ : InMux
    port map (
            O => \N__38466\,
            I => \N__38419\
        );

    \I__8472\ : InMux
    port map (
            O => \N__38465\,
            I => \N__38419\
        );

    \I__8471\ : InMux
    port map (
            O => \N__38462\,
            I => \N__38408\
        );

    \I__8470\ : InMux
    port map (
            O => \N__38461\,
            I => \N__38408\
        );

    \I__8469\ : InMux
    port map (
            O => \N__38460\,
            I => \N__38408\
        );

    \I__8468\ : InMux
    port map (
            O => \N__38457\,
            I => \N__38408\
        );

    \I__8467\ : InMux
    port map (
            O => \N__38456\,
            I => \N__38408\
        );

    \I__8466\ : LocalMux
    port map (
            O => \N__38445\,
            I => \nx.n2423\
        );

    \I__8465\ : Odrv4
    port map (
            O => \N__38440\,
            I => \nx.n2423\
        );

    \I__8464\ : LocalMux
    port map (
            O => \N__38437\,
            I => \nx.n2423\
        );

    \I__8463\ : Odrv4
    port map (
            O => \N__38434\,
            I => \nx.n2423\
        );

    \I__8462\ : LocalMux
    port map (
            O => \N__38431\,
            I => \nx.n2423\
        );

    \I__8461\ : LocalMux
    port map (
            O => \N__38424\,
            I => \nx.n2423\
        );

    \I__8460\ : LocalMux
    port map (
            O => \N__38419\,
            I => \nx.n2423\
        );

    \I__8459\ : LocalMux
    port map (
            O => \N__38408\,
            I => \nx.n2423\
        );

    \I__8458\ : SRMux
    port map (
            O => \N__38391\,
            I => \N__38387\
        );

    \I__8457\ : SRMux
    port map (
            O => \N__38390\,
            I => \N__38384\
        );

    \I__8456\ : LocalMux
    port map (
            O => \N__38387\,
            I => \N__38379\
        );

    \I__8455\ : LocalMux
    port map (
            O => \N__38384\,
            I => \N__38379\
        );

    \I__8454\ : Span4Mux_v
    port map (
            O => \N__38379\,
            I => \N__38376\
        );

    \I__8453\ : Span4Mux_h
    port map (
            O => \N__38376\,
            I => \N__38373\
        );

    \I__8452\ : Odrv4
    port map (
            O => \N__38373\,
            I => n7992
        );

    \I__8451\ : InMux
    port map (
            O => \N__38370\,
            I => \N__38367\
        );

    \I__8450\ : LocalMux
    port map (
            O => \N__38367\,
            I => n7602
        );

    \I__8449\ : IoInMux
    port map (
            O => \N__38364\,
            I => \N__38361\
        );

    \I__8448\ : LocalMux
    port map (
            O => \N__38361\,
            I => \N__38358\
        );

    \I__8447\ : IoSpan4Mux
    port map (
            O => \N__38358\,
            I => \N__38355\
        );

    \I__8446\ : Span4Mux_s0_h
    port map (
            O => \N__38355\,
            I => \N__38352\
        );

    \I__8445\ : Sp12to4
    port map (
            O => \N__38352\,
            I => \N__38349\
        );

    \I__8444\ : Span12Mux_s11_h
    port map (
            O => \N__38349\,
            I => \N__38346\
        );

    \I__8443\ : Span12Mux_v
    port map (
            O => \N__38346\,
            I => \N__38342\
        );

    \I__8442\ : InMux
    port map (
            O => \N__38345\,
            I => \N__38339\
        );

    \I__8441\ : Odrv12
    port map (
            O => \N__38342\,
            I => pin_oe_11
        );

    \I__8440\ : LocalMux
    port map (
            O => \N__38339\,
            I => pin_oe_11
        );

    \I__8439\ : InMux
    port map (
            O => \N__38334\,
            I => \N__38331\
        );

    \I__8438\ : LocalMux
    port map (
            O => \N__38331\,
            I => \nx.n2476\
        );

    \I__8437\ : CascadeMux
    port map (
            O => \N__38328\,
            I => \N__38325\
        );

    \I__8436\ : InMux
    port map (
            O => \N__38325\,
            I => \N__38322\
        );

    \I__8435\ : LocalMux
    port map (
            O => \N__38322\,
            I => \N__38318\
        );

    \I__8434\ : CascadeMux
    port map (
            O => \N__38321\,
            I => \N__38314\
        );

    \I__8433\ : Span4Mux_h
    port map (
            O => \N__38318\,
            I => \N__38311\
        );

    \I__8432\ : InMux
    port map (
            O => \N__38317\,
            I => \N__38308\
        );

    \I__8431\ : InMux
    port map (
            O => \N__38314\,
            I => \N__38305\
        );

    \I__8430\ : Odrv4
    port map (
            O => \N__38311\,
            I => \nx.n2409\
        );

    \I__8429\ : LocalMux
    port map (
            O => \N__38308\,
            I => \nx.n2409\
        );

    \I__8428\ : LocalMux
    port map (
            O => \N__38305\,
            I => \nx.n2409\
        );

    \I__8427\ : InMux
    port map (
            O => \N__38298\,
            I => \N__38294\
        );

    \I__8426\ : CascadeMux
    port map (
            O => \N__38297\,
            I => \N__38291\
        );

    \I__8425\ : LocalMux
    port map (
            O => \N__38294\,
            I => \N__38287\
        );

    \I__8424\ : InMux
    port map (
            O => \N__38291\,
            I => \N__38284\
        );

    \I__8423\ : InMux
    port map (
            O => \N__38290\,
            I => \N__38281\
        );

    \I__8422\ : Span4Mux_h
    port map (
            O => \N__38287\,
            I => \N__38278\
        );

    \I__8421\ : LocalMux
    port map (
            O => \N__38284\,
            I => \N__38273\
        );

    \I__8420\ : LocalMux
    port map (
            O => \N__38281\,
            I => \N__38273\
        );

    \I__8419\ : Odrv4
    port map (
            O => \N__38278\,
            I => \nx.n2400\
        );

    \I__8418\ : Odrv12
    port map (
            O => \N__38273\,
            I => \nx.n2400\
        );

    \I__8417\ : CascadeMux
    port map (
            O => \N__38268\,
            I => \N__38265\
        );

    \I__8416\ : InMux
    port map (
            O => \N__38265\,
            I => \N__38262\
        );

    \I__8415\ : LocalMux
    port map (
            O => \N__38262\,
            I => \nx.n2467\
        );

    \I__8414\ : CascadeMux
    port map (
            O => \N__38259\,
            I => \N__38255\
        );

    \I__8413\ : InMux
    port map (
            O => \N__38258\,
            I => \N__38251\
        );

    \I__8412\ : InMux
    port map (
            O => \N__38255\,
            I => \N__38248\
        );

    \I__8411\ : InMux
    port map (
            O => \N__38254\,
            I => \N__38245\
        );

    \I__8410\ : LocalMux
    port map (
            O => \N__38251\,
            I => \N__38242\
        );

    \I__8409\ : LocalMux
    port map (
            O => \N__38248\,
            I => \N__38239\
        );

    \I__8408\ : LocalMux
    port map (
            O => \N__38245\,
            I => \N__38236\
        );

    \I__8407\ : Odrv4
    port map (
            O => \N__38242\,
            I => \nx.n2396\
        );

    \I__8406\ : Odrv4
    port map (
            O => \N__38239\,
            I => \nx.n2396\
        );

    \I__8405\ : Odrv12
    port map (
            O => \N__38236\,
            I => \nx.n2396\
        );

    \I__8404\ : InMux
    port map (
            O => \N__38229\,
            I => \N__38226\
        );

    \I__8403\ : LocalMux
    port map (
            O => \N__38226\,
            I => \N__38223\
        );

    \I__8402\ : Odrv4
    port map (
            O => \N__38223\,
            I => \nx.n2463\
        );

    \I__8401\ : CascadeMux
    port map (
            O => \N__38220\,
            I => \nx.n2495_cascade_\
        );

    \I__8400\ : InMux
    port map (
            O => \N__38217\,
            I => \N__38214\
        );

    \I__8399\ : LocalMux
    port map (
            O => \N__38214\,
            I => \N__38211\
        );

    \I__8398\ : Odrv4
    port map (
            O => \N__38211\,
            I => \nx.n34_adj_758\
        );

    \I__8397\ : InMux
    port map (
            O => \N__38208\,
            I => \N__38205\
        );

    \I__8396\ : LocalMux
    port map (
            O => \N__38205\,
            I => \N__38201\
        );

    \I__8395\ : CascadeMux
    port map (
            O => \N__38204\,
            I => \N__38198\
        );

    \I__8394\ : Span4Mux_h
    port map (
            O => \N__38201\,
            I => \N__38195\
        );

    \I__8393\ : InMux
    port map (
            O => \N__38198\,
            I => \N__38192\
        );

    \I__8392\ : Odrv4
    port map (
            O => \N__38195\,
            I => \nx.n2398\
        );

    \I__8391\ : LocalMux
    port map (
            O => \N__38192\,
            I => \nx.n2398\
        );

    \I__8390\ : InMux
    port map (
            O => \N__38187\,
            I => \N__38184\
        );

    \I__8389\ : LocalMux
    port map (
            O => \N__38184\,
            I => \nx.n2465\
        );

    \I__8388\ : InMux
    port map (
            O => \N__38181\,
            I => \N__38177\
        );

    \I__8387\ : CascadeMux
    port map (
            O => \N__38180\,
            I => \N__38174\
        );

    \I__8386\ : LocalMux
    port map (
            O => \N__38177\,
            I => \N__38170\
        );

    \I__8385\ : InMux
    port map (
            O => \N__38174\,
            I => \N__38167\
        );

    \I__8384\ : InMux
    port map (
            O => \N__38173\,
            I => \N__38164\
        );

    \I__8383\ : Odrv4
    port map (
            O => \N__38170\,
            I => \nx.n2395\
        );

    \I__8382\ : LocalMux
    port map (
            O => \N__38167\,
            I => \nx.n2395\
        );

    \I__8381\ : LocalMux
    port map (
            O => \N__38164\,
            I => \nx.n2395\
        );

    \I__8380\ : CascadeMux
    port map (
            O => \N__38157\,
            I => \N__38154\
        );

    \I__8379\ : InMux
    port map (
            O => \N__38154\,
            I => \N__38151\
        );

    \I__8378\ : LocalMux
    port map (
            O => \N__38151\,
            I => \nx.n2462\
        );

    \I__8377\ : CascadeMux
    port map (
            O => \N__38148\,
            I => \N__38144\
        );

    \I__8376\ : InMux
    port map (
            O => \N__38147\,
            I => \N__38140\
        );

    \I__8375\ : InMux
    port map (
            O => \N__38144\,
            I => \N__38137\
        );

    \I__8374\ : InMux
    port map (
            O => \N__38143\,
            I => \N__38134\
        );

    \I__8373\ : LocalMux
    port map (
            O => \N__38140\,
            I => \N__38131\
        );

    \I__8372\ : LocalMux
    port map (
            O => \N__38137\,
            I => \N__38128\
        );

    \I__8371\ : LocalMux
    port map (
            O => \N__38134\,
            I => \N__38125\
        );

    \I__8370\ : Odrv4
    port map (
            O => \N__38131\,
            I => \nx.n2397\
        );

    \I__8369\ : Odrv4
    port map (
            O => \N__38128\,
            I => \nx.n2397\
        );

    \I__8368\ : Odrv12
    port map (
            O => \N__38125\,
            I => \nx.n2397\
        );

    \I__8367\ : CascadeMux
    port map (
            O => \N__38118\,
            I => \N__38115\
        );

    \I__8366\ : InMux
    port map (
            O => \N__38115\,
            I => \N__38112\
        );

    \I__8365\ : LocalMux
    port map (
            O => \N__38112\,
            I => \nx.n2464\
        );

    \I__8364\ : CascadeMux
    port map (
            O => \N__38109\,
            I => \nx.n2496_cascade_\
        );

    \I__8363\ : InMux
    port map (
            O => \N__38106\,
            I => \N__38101\
        );

    \I__8362\ : CascadeMux
    port map (
            O => \N__38105\,
            I => \N__38098\
        );

    \I__8361\ : InMux
    port map (
            O => \N__38104\,
            I => \N__38095\
        );

    \I__8360\ : LocalMux
    port map (
            O => \N__38101\,
            I => \N__38092\
        );

    \I__8359\ : InMux
    port map (
            O => \N__38098\,
            I => \N__38089\
        );

    \I__8358\ : LocalMux
    port map (
            O => \N__38095\,
            I => \N__38086\
        );

    \I__8357\ : Odrv4
    port map (
            O => \N__38092\,
            I => \nx.n2394\
        );

    \I__8356\ : LocalMux
    port map (
            O => \N__38089\,
            I => \nx.n2394\
        );

    \I__8355\ : Odrv12
    port map (
            O => \N__38086\,
            I => \nx.n2394\
        );

    \I__8354\ : CascadeMux
    port map (
            O => \N__38079\,
            I => \N__38076\
        );

    \I__8353\ : InMux
    port map (
            O => \N__38076\,
            I => \N__38073\
        );

    \I__8352\ : LocalMux
    port map (
            O => \N__38073\,
            I => \nx.n2461\
        );

    \I__8351\ : CascadeMux
    port map (
            O => \N__38070\,
            I => \nx.n2592_cascade_\
        );

    \I__8350\ : InMux
    port map (
            O => \N__38067\,
            I => \N__38064\
        );

    \I__8349\ : LocalMux
    port map (
            O => \N__38064\,
            I => \nx.n35\
        );

    \I__8348\ : InMux
    port map (
            O => \N__38061\,
            I => \N__38058\
        );

    \I__8347\ : LocalMux
    port map (
            O => \N__38058\,
            I => \N__38055\
        );

    \I__8346\ : Span4Mux_v
    port map (
            O => \N__38055\,
            I => \N__38051\
        );

    \I__8345\ : InMux
    port map (
            O => \N__38054\,
            I => \N__38048\
        );

    \I__8344\ : Span4Mux_h
    port map (
            O => \N__38051\,
            I => \N__38043\
        );

    \I__8343\ : LocalMux
    port map (
            O => \N__38048\,
            I => \N__38043\
        );

    \I__8342\ : Odrv4
    port map (
            O => \N__38043\,
            I => \nx.n2391\
        );

    \I__8341\ : InMux
    port map (
            O => \N__38040\,
            I => \N__38037\
        );

    \I__8340\ : LocalMux
    port map (
            O => \N__38037\,
            I => \N__38034\
        );

    \I__8339\ : Odrv4
    port map (
            O => \N__38034\,
            I => \nx.n2458\
        );

    \I__8338\ : CascadeMux
    port map (
            O => \N__38031\,
            I => \nx.n2490_cascade_\
        );

    \I__8337\ : InMux
    port map (
            O => \N__38028\,
            I => \N__38025\
        );

    \I__8336\ : LocalMux
    port map (
            O => \N__38025\,
            I => \nx.n22_adj_755\
        );

    \I__8335\ : InMux
    port map (
            O => \N__38022\,
            I => \N__38018\
        );

    \I__8334\ : CascadeMux
    port map (
            O => \N__38021\,
            I => \N__38005\
        );

    \I__8333\ : LocalMux
    port map (
            O => \N__38018\,
            I => \N__38001\
        );

    \I__8332\ : CascadeMux
    port map (
            O => \N__38017\,
            I => \N__37996\
        );

    \I__8331\ : CascadeMux
    port map (
            O => \N__38016\,
            I => \N__37992\
        );

    \I__8330\ : CascadeMux
    port map (
            O => \N__38015\,
            I => \N__37989\
        );

    \I__8329\ : InMux
    port map (
            O => \N__38014\,
            I => \N__37978\
        );

    \I__8328\ : InMux
    port map (
            O => \N__38013\,
            I => \N__37978\
        );

    \I__8327\ : InMux
    port map (
            O => \N__38012\,
            I => \N__37978\
        );

    \I__8326\ : InMux
    port map (
            O => \N__38011\,
            I => \N__37978\
        );

    \I__8325\ : CascadeMux
    port map (
            O => \N__38010\,
            I => \N__37975\
        );

    \I__8324\ : CascadeMux
    port map (
            O => \N__38009\,
            I => \N__37972\
        );

    \I__8323\ : CascadeMux
    port map (
            O => \N__38008\,
            I => \N__37969\
        );

    \I__8322\ : InMux
    port map (
            O => \N__38005\,
            I => \N__37964\
        );

    \I__8321\ : InMux
    port map (
            O => \N__38004\,
            I => \N__37961\
        );

    \I__8320\ : Span4Mux_h
    port map (
            O => \N__38001\,
            I => \N__37958\
        );

    \I__8319\ : InMux
    port map (
            O => \N__38000\,
            I => \N__37949\
        );

    \I__8318\ : InMux
    port map (
            O => \N__37999\,
            I => \N__37949\
        );

    \I__8317\ : InMux
    port map (
            O => \N__37996\,
            I => \N__37949\
        );

    \I__8316\ : InMux
    port map (
            O => \N__37995\,
            I => \N__37949\
        );

    \I__8315\ : InMux
    port map (
            O => \N__37992\,
            I => \N__37944\
        );

    \I__8314\ : InMux
    port map (
            O => \N__37989\,
            I => \N__37944\
        );

    \I__8313\ : InMux
    port map (
            O => \N__37988\,
            I => \N__37939\
        );

    \I__8312\ : InMux
    port map (
            O => \N__37987\,
            I => \N__37939\
        );

    \I__8311\ : LocalMux
    port map (
            O => \N__37978\,
            I => \N__37936\
        );

    \I__8310\ : InMux
    port map (
            O => \N__37975\,
            I => \N__37925\
        );

    \I__8309\ : InMux
    port map (
            O => \N__37972\,
            I => \N__37925\
        );

    \I__8308\ : InMux
    port map (
            O => \N__37969\,
            I => \N__37925\
        );

    \I__8307\ : InMux
    port map (
            O => \N__37968\,
            I => \N__37925\
        );

    \I__8306\ : InMux
    port map (
            O => \N__37967\,
            I => \N__37925\
        );

    \I__8305\ : LocalMux
    port map (
            O => \N__37964\,
            I => \N__37920\
        );

    \I__8304\ : LocalMux
    port map (
            O => \N__37961\,
            I => \N__37920\
        );

    \I__8303\ : Odrv4
    port map (
            O => \N__37958\,
            I => \nx.n2324\
        );

    \I__8302\ : LocalMux
    port map (
            O => \N__37949\,
            I => \nx.n2324\
        );

    \I__8301\ : LocalMux
    port map (
            O => \N__37944\,
            I => \nx.n2324\
        );

    \I__8300\ : LocalMux
    port map (
            O => \N__37939\,
            I => \nx.n2324\
        );

    \I__8299\ : Odrv4
    port map (
            O => \N__37936\,
            I => \nx.n2324\
        );

    \I__8298\ : LocalMux
    port map (
            O => \N__37925\,
            I => \nx.n2324\
        );

    \I__8297\ : Odrv4
    port map (
            O => \N__37920\,
            I => \nx.n2324\
        );

    \I__8296\ : CascadeMux
    port map (
            O => \N__37905\,
            I => \N__37902\
        );

    \I__8295\ : InMux
    port map (
            O => \N__37902\,
            I => \N__37899\
        );

    \I__8294\ : LocalMux
    port map (
            O => \N__37899\,
            I => \N__37893\
        );

    \I__8293\ : InMux
    port map (
            O => \N__37898\,
            I => \N__37890\
        );

    \I__8292\ : CascadeMux
    port map (
            O => \N__37897\,
            I => \N__37887\
        );

    \I__8291\ : InMux
    port map (
            O => \N__37896\,
            I => \N__37884\
        );

    \I__8290\ : Span4Mux_h
    port map (
            O => \N__37893\,
            I => \N__37879\
        );

    \I__8289\ : LocalMux
    port map (
            O => \N__37890\,
            I => \N__37879\
        );

    \I__8288\ : InMux
    port map (
            O => \N__37887\,
            I => \N__37876\
        );

    \I__8287\ : LocalMux
    port map (
            O => \N__37884\,
            I => \nx.n2307\
        );

    \I__8286\ : Odrv4
    port map (
            O => \N__37879\,
            I => \nx.n2307\
        );

    \I__8285\ : LocalMux
    port map (
            O => \N__37876\,
            I => \nx.n2307\
        );

    \I__8284\ : InMux
    port map (
            O => \N__37869\,
            I => \N__37866\
        );

    \I__8283\ : LocalMux
    port map (
            O => \N__37866\,
            I => \nx.n13321\
        );

    \I__8282\ : CascadeMux
    port map (
            O => \N__37863\,
            I => \nx.n2505_cascade_\
        );

    \I__8281\ : CascadeMux
    port map (
            O => \N__37860\,
            I => \nx.n2606_cascade_\
        );

    \I__8280\ : CascadeMux
    port map (
            O => \N__37857\,
            I => \N__37853\
        );

    \I__8279\ : InMux
    port map (
            O => \N__37856\,
            I => \N__37850\
        );

    \I__8278\ : InMux
    port map (
            O => \N__37853\,
            I => \N__37847\
        );

    \I__8277\ : LocalMux
    port map (
            O => \N__37850\,
            I => \N__37843\
        );

    \I__8276\ : LocalMux
    port map (
            O => \N__37847\,
            I => \N__37840\
        );

    \I__8275\ : CascadeMux
    port map (
            O => \N__37846\,
            I => \N__37837\
        );

    \I__8274\ : Span4Mux_v
    port map (
            O => \N__37843\,
            I => \N__37832\
        );

    \I__8273\ : Span4Mux_h
    port map (
            O => \N__37840\,
            I => \N__37832\
        );

    \I__8272\ : InMux
    port map (
            O => \N__37837\,
            I => \N__37829\
        );

    \I__8271\ : Span4Mux_h
    port map (
            O => \N__37832\,
            I => \N__37826\
        );

    \I__8270\ : LocalMux
    port map (
            O => \N__37829\,
            I => \nx.n2705\
        );

    \I__8269\ : Odrv4
    port map (
            O => \N__37826\,
            I => \nx.n2705\
        );

    \I__8268\ : CascadeMux
    port map (
            O => \N__37821\,
            I => \N__37818\
        );

    \I__8267\ : InMux
    port map (
            O => \N__37818\,
            I => \N__37814\
        );

    \I__8266\ : InMux
    port map (
            O => \N__37817\,
            I => \N__37811\
        );

    \I__8265\ : LocalMux
    port map (
            O => \N__37814\,
            I => \N__37808\
        );

    \I__8264\ : LocalMux
    port map (
            O => \N__37811\,
            I => \N__37805\
        );

    \I__8263\ : Span4Mux_h
    port map (
            O => \N__37808\,
            I => \N__37801\
        );

    \I__8262\ : Span4Mux_h
    port map (
            O => \N__37805\,
            I => \N__37798\
        );

    \I__8261\ : InMux
    port map (
            O => \N__37804\,
            I => \N__37795\
        );

    \I__8260\ : Span4Mux_h
    port map (
            O => \N__37801\,
            I => \N__37792\
        );

    \I__8259\ : Odrv4
    port map (
            O => \N__37798\,
            I => \nx.n2704\
        );

    \I__8258\ : LocalMux
    port map (
            O => \N__37795\,
            I => \nx.n2704\
        );

    \I__8257\ : Odrv4
    port map (
            O => \N__37792\,
            I => \nx.n2704\
        );

    \I__8256\ : CascadeMux
    port map (
            O => \N__37785\,
            I => \nx.n37_adj_772_cascade_\
        );

    \I__8255\ : InMux
    port map (
            O => \N__37782\,
            I => \N__37779\
        );

    \I__8254\ : LocalMux
    port map (
            O => \N__37779\,
            I => \nx.n39_adj_773\
        );

    \I__8253\ : CascadeMux
    port map (
            O => \N__37776\,
            I => \nx.n2522_cascade_\
        );

    \I__8252\ : InMux
    port map (
            O => \N__37773\,
            I => \N__37770\
        );

    \I__8251\ : LocalMux
    port map (
            O => \N__37770\,
            I => \N__37767\
        );

    \I__8250\ : Span4Mux_h
    port map (
            O => \N__37767\,
            I => \N__37763\
        );

    \I__8249\ : InMux
    port map (
            O => \N__37766\,
            I => \N__37759\
        );

    \I__8248\ : Span4Mux_v
    port map (
            O => \N__37763\,
            I => \N__37756\
        );

    \I__8247\ : InMux
    port map (
            O => \N__37762\,
            I => \N__37753\
        );

    \I__8246\ : LocalMux
    port map (
            O => \N__37759\,
            I => \N__37750\
        );

    \I__8245\ : Odrv4
    port map (
            O => \N__37756\,
            I => \nx.n2793\
        );

    \I__8244\ : LocalMux
    port map (
            O => \N__37753\,
            I => \nx.n2793\
        );

    \I__8243\ : Odrv12
    port map (
            O => \N__37750\,
            I => \nx.n2793\
        );

    \I__8242\ : CascadeMux
    port map (
            O => \N__37743\,
            I => \N__37740\
        );

    \I__8241\ : InMux
    port map (
            O => \N__37740\,
            I => \N__37737\
        );

    \I__8240\ : LocalMux
    port map (
            O => \N__37737\,
            I => \N__37734\
        );

    \I__8239\ : Span4Mux_h
    port map (
            O => \N__37734\,
            I => \N__37731\
        );

    \I__8238\ : Span4Mux_h
    port map (
            O => \N__37731\,
            I => \N__37728\
        );

    \I__8237\ : Odrv4
    port map (
            O => \N__37728\,
            I => \nx.n2860\
        );

    \I__8236\ : CascadeMux
    port map (
            O => \N__37725\,
            I => \N__37722\
        );

    \I__8235\ : InMux
    port map (
            O => \N__37722\,
            I => \N__37719\
        );

    \I__8234\ : LocalMux
    port map (
            O => \N__37719\,
            I => \N__37715\
        );

    \I__8233\ : CascadeMux
    port map (
            O => \N__37718\,
            I => \N__37711\
        );

    \I__8232\ : Span4Mux_h
    port map (
            O => \N__37715\,
            I => \N__37708\
        );

    \I__8231\ : InMux
    port map (
            O => \N__37714\,
            I => \N__37705\
        );

    \I__8230\ : InMux
    port map (
            O => \N__37711\,
            I => \N__37702\
        );

    \I__8229\ : Odrv4
    port map (
            O => \N__37708\,
            I => \nx.n2892\
        );

    \I__8228\ : LocalMux
    port map (
            O => \N__37705\,
            I => \nx.n2892\
        );

    \I__8227\ : LocalMux
    port map (
            O => \N__37702\,
            I => \nx.n2892\
        );

    \I__8226\ : CascadeMux
    port map (
            O => \N__37695\,
            I => \N__37692\
        );

    \I__8225\ : InMux
    port map (
            O => \N__37692\,
            I => \N__37689\
        );

    \I__8224\ : LocalMux
    port map (
            O => \N__37689\,
            I => \nx.n2960\
        );

    \I__8223\ : InMux
    port map (
            O => \N__37686\,
            I => \N__37682\
        );

    \I__8222\ : InMux
    port map (
            O => \N__37685\,
            I => \N__37679\
        );

    \I__8221\ : LocalMux
    port map (
            O => \N__37682\,
            I => \N__37674\
        );

    \I__8220\ : LocalMux
    port map (
            O => \N__37679\,
            I => \N__37674\
        );

    \I__8219\ : Span4Mux_h
    port map (
            O => \N__37674\,
            I => \N__37670\
        );

    \I__8218\ : InMux
    port map (
            O => \N__37673\,
            I => \N__37667\
        );

    \I__8217\ : Odrv4
    port map (
            O => \N__37670\,
            I => \nx.n2992\
        );

    \I__8216\ : LocalMux
    port map (
            O => \N__37667\,
            I => \nx.n2992\
        );

    \I__8215\ : InMux
    port map (
            O => \N__37662\,
            I => \N__37659\
        );

    \I__8214\ : LocalMux
    port map (
            O => \N__37659\,
            I => \N__37655\
        );

    \I__8213\ : InMux
    port map (
            O => \N__37658\,
            I => \N__37651\
        );

    \I__8212\ : Span4Mux_h
    port map (
            O => \N__37655\,
            I => \N__37648\
        );

    \I__8211\ : CascadeMux
    port map (
            O => \N__37654\,
            I => \N__37645\
        );

    \I__8210\ : LocalMux
    port map (
            O => \N__37651\,
            I => \N__37642\
        );

    \I__8209\ : Span4Mux_v
    port map (
            O => \N__37648\,
            I => \N__37639\
        );

    \I__8208\ : InMux
    port map (
            O => \N__37645\,
            I => \N__37636\
        );

    \I__8207\ : Span4Mux_v
    port map (
            O => \N__37642\,
            I => \N__37633\
        );

    \I__8206\ : Odrv4
    port map (
            O => \N__37639\,
            I => \nx.n2794\
        );

    \I__8205\ : LocalMux
    port map (
            O => \N__37636\,
            I => \nx.n2794\
        );

    \I__8204\ : Odrv4
    port map (
            O => \N__37633\,
            I => \nx.n2794\
        );

    \I__8203\ : CascadeMux
    port map (
            O => \N__37626\,
            I => \N__37623\
        );

    \I__8202\ : InMux
    port map (
            O => \N__37623\,
            I => \N__37620\
        );

    \I__8201\ : LocalMux
    port map (
            O => \N__37620\,
            I => \N__37617\
        );

    \I__8200\ : Span4Mux_h
    port map (
            O => \N__37617\,
            I => \N__37614\
        );

    \I__8199\ : Span4Mux_h
    port map (
            O => \N__37614\,
            I => \N__37611\
        );

    \I__8198\ : Odrv4
    port map (
            O => \N__37611\,
            I => \nx.n2861\
        );

    \I__8197\ : CascadeMux
    port map (
            O => \N__37608\,
            I => \N__37599\
        );

    \I__8196\ : InMux
    port map (
            O => \N__37607\,
            I => \N__37592\
        );

    \I__8195\ : CascadeMux
    port map (
            O => \N__37606\,
            I => \N__37589\
        );

    \I__8194\ : InMux
    port map (
            O => \N__37605\,
            I => \N__37581\
        );

    \I__8193\ : InMux
    port map (
            O => \N__37604\,
            I => \N__37581\
        );

    \I__8192\ : InMux
    port map (
            O => \N__37603\,
            I => \N__37581\
        );

    \I__8191\ : CascadeMux
    port map (
            O => \N__37602\,
            I => \N__37576\
        );

    \I__8190\ : InMux
    port map (
            O => \N__37599\,
            I => \N__37570\
        );

    \I__8189\ : InMux
    port map (
            O => \N__37598\,
            I => \N__37570\
        );

    \I__8188\ : InMux
    port map (
            O => \N__37597\,
            I => \N__37567\
        );

    \I__8187\ : InMux
    port map (
            O => \N__37596\,
            I => \N__37561\
        );

    \I__8186\ : CascadeMux
    port map (
            O => \N__37595\,
            I => \N__37557\
        );

    \I__8185\ : LocalMux
    port map (
            O => \N__37592\,
            I => \N__37552\
        );

    \I__8184\ : InMux
    port map (
            O => \N__37589\,
            I => \N__37547\
        );

    \I__8183\ : InMux
    port map (
            O => \N__37588\,
            I => \N__37547\
        );

    \I__8182\ : LocalMux
    port map (
            O => \N__37581\,
            I => \N__37544\
        );

    \I__8181\ : InMux
    port map (
            O => \N__37580\,
            I => \N__37539\
        );

    \I__8180\ : InMux
    port map (
            O => \N__37579\,
            I => \N__37539\
        );

    \I__8179\ : InMux
    port map (
            O => \N__37576\,
            I => \N__37534\
        );

    \I__8178\ : InMux
    port map (
            O => \N__37575\,
            I => \N__37534\
        );

    \I__8177\ : LocalMux
    port map (
            O => \N__37570\,
            I => \N__37531\
        );

    \I__8176\ : LocalMux
    port map (
            O => \N__37567\,
            I => \N__37528\
        );

    \I__8175\ : CascadeMux
    port map (
            O => \N__37566\,
            I => \N__37525\
        );

    \I__8174\ : CascadeMux
    port map (
            O => \N__37565\,
            I => \N__37522\
        );

    \I__8173\ : CascadeMux
    port map (
            O => \N__37564\,
            I => \N__37518\
        );

    \I__8172\ : LocalMux
    port map (
            O => \N__37561\,
            I => \N__37514\
        );

    \I__8171\ : InMux
    port map (
            O => \N__37560\,
            I => \N__37506\
        );

    \I__8170\ : InMux
    port map (
            O => \N__37557\,
            I => \N__37506\
        );

    \I__8169\ : InMux
    port map (
            O => \N__37556\,
            I => \N__37506\
        );

    \I__8168\ : InMux
    port map (
            O => \N__37555\,
            I => \N__37503\
        );

    \I__8167\ : Span4Mux_v
    port map (
            O => \N__37552\,
            I => \N__37500\
        );

    \I__8166\ : LocalMux
    port map (
            O => \N__37547\,
            I => \N__37493\
        );

    \I__8165\ : Span4Mux_h
    port map (
            O => \N__37544\,
            I => \N__37493\
        );

    \I__8164\ : LocalMux
    port map (
            O => \N__37539\,
            I => \N__37493\
        );

    \I__8163\ : LocalMux
    port map (
            O => \N__37534\,
            I => \N__37486\
        );

    \I__8162\ : Span4Mux_h
    port map (
            O => \N__37531\,
            I => \N__37486\
        );

    \I__8161\ : Span4Mux_h
    port map (
            O => \N__37528\,
            I => \N__37486\
        );

    \I__8160\ : InMux
    port map (
            O => \N__37525\,
            I => \N__37479\
        );

    \I__8159\ : InMux
    port map (
            O => \N__37522\,
            I => \N__37479\
        );

    \I__8158\ : InMux
    port map (
            O => \N__37521\,
            I => \N__37479\
        );

    \I__8157\ : InMux
    port map (
            O => \N__37518\,
            I => \N__37474\
        );

    \I__8156\ : InMux
    port map (
            O => \N__37517\,
            I => \N__37474\
        );

    \I__8155\ : Span4Mux_v
    port map (
            O => \N__37514\,
            I => \N__37471\
        );

    \I__8154\ : InMux
    port map (
            O => \N__37513\,
            I => \N__37468\
        );

    \I__8153\ : LocalMux
    port map (
            O => \N__37506\,
            I => \nx.n2819\
        );

    \I__8152\ : LocalMux
    port map (
            O => \N__37503\,
            I => \nx.n2819\
        );

    \I__8151\ : Odrv4
    port map (
            O => \N__37500\,
            I => \nx.n2819\
        );

    \I__8150\ : Odrv4
    port map (
            O => \N__37493\,
            I => \nx.n2819\
        );

    \I__8149\ : Odrv4
    port map (
            O => \N__37486\,
            I => \nx.n2819\
        );

    \I__8148\ : LocalMux
    port map (
            O => \N__37479\,
            I => \nx.n2819\
        );

    \I__8147\ : LocalMux
    port map (
            O => \N__37474\,
            I => \nx.n2819\
        );

    \I__8146\ : Odrv4
    port map (
            O => \N__37471\,
            I => \nx.n2819\
        );

    \I__8145\ : LocalMux
    port map (
            O => \N__37468\,
            I => \nx.n2819\
        );

    \I__8144\ : InMux
    port map (
            O => \N__37449\,
            I => \N__37445\
        );

    \I__8143\ : InMux
    port map (
            O => \N__37448\,
            I => \N__37442\
        );

    \I__8142\ : LocalMux
    port map (
            O => \N__37445\,
            I => \nx.n2893\
        );

    \I__8141\ : LocalMux
    port map (
            O => \N__37442\,
            I => \nx.n2893\
        );

    \I__8140\ : CascadeMux
    port map (
            O => \N__37437\,
            I => \N__37433\
        );

    \I__8139\ : InMux
    port map (
            O => \N__37436\,
            I => \N__37430\
        );

    \I__8138\ : InMux
    port map (
            O => \N__37433\,
            I => \N__37427\
        );

    \I__8137\ : LocalMux
    port map (
            O => \N__37430\,
            I => \N__37422\
        );

    \I__8136\ : LocalMux
    port map (
            O => \N__37427\,
            I => \N__37422\
        );

    \I__8135\ : Odrv4
    port map (
            O => \N__37422\,
            I => \nx.n2898\
        );

    \I__8134\ : InMux
    port map (
            O => \N__37419\,
            I => \N__37414\
        );

    \I__8133\ : CascadeMux
    port map (
            O => \N__37418\,
            I => \N__37411\
        );

    \I__8132\ : InMux
    port map (
            O => \N__37417\,
            I => \N__37408\
        );

    \I__8131\ : LocalMux
    port map (
            O => \N__37414\,
            I => \N__37405\
        );

    \I__8130\ : InMux
    port map (
            O => \N__37411\,
            I => \N__37402\
        );

    \I__8129\ : LocalMux
    port map (
            O => \N__37408\,
            I => \nx.n2904\
        );

    \I__8128\ : Odrv4
    port map (
            O => \N__37405\,
            I => \nx.n2904\
        );

    \I__8127\ : LocalMux
    port map (
            O => \N__37402\,
            I => \nx.n2904\
        );

    \I__8126\ : CascadeMux
    port map (
            O => \N__37395\,
            I => \nx.n2893_cascade_\
        );

    \I__8125\ : CascadeMux
    port map (
            O => \N__37392\,
            I => \N__37389\
        );

    \I__8124\ : InMux
    port map (
            O => \N__37389\,
            I => \N__37386\
        );

    \I__8123\ : LocalMux
    port map (
            O => \N__37386\,
            I => \N__37383\
        );

    \I__8122\ : Span4Mux_v
    port map (
            O => \N__37383\,
            I => \N__37378\
        );

    \I__8121\ : InMux
    port map (
            O => \N__37382\,
            I => \N__37375\
        );

    \I__8120\ : CascadeMux
    port map (
            O => \N__37381\,
            I => \N__37372\
        );

    \I__8119\ : Span4Mux_h
    port map (
            O => \N__37378\,
            I => \N__37367\
        );

    \I__8118\ : LocalMux
    port map (
            O => \N__37375\,
            I => \N__37367\
        );

    \I__8117\ : InMux
    port map (
            O => \N__37372\,
            I => \N__37364\
        );

    \I__8116\ : Odrv4
    port map (
            O => \N__37367\,
            I => \nx.n2897\
        );

    \I__8115\ : LocalMux
    port map (
            O => \N__37364\,
            I => \nx.n2897\
        );

    \I__8114\ : InMux
    port map (
            O => \N__37359\,
            I => \N__37356\
        );

    \I__8113\ : LocalMux
    port map (
            O => \N__37356\,
            I => \nx.n41_adj_768\
        );

    \I__8112\ : CascadeMux
    port map (
            O => \N__37353\,
            I => \N__37350\
        );

    \I__8111\ : InMux
    port map (
            O => \N__37350\,
            I => \N__37346\
        );

    \I__8110\ : InMux
    port map (
            O => \N__37349\,
            I => \N__37343\
        );

    \I__8109\ : LocalMux
    port map (
            O => \N__37346\,
            I => \N__37340\
        );

    \I__8108\ : LocalMux
    port map (
            O => \N__37343\,
            I => \N__37336\
        );

    \I__8107\ : Span4Mux_h
    port map (
            O => \N__37340\,
            I => \N__37333\
        );

    \I__8106\ : InMux
    port map (
            O => \N__37339\,
            I => \N__37330\
        );

    \I__8105\ : Odrv12
    port map (
            O => \N__37336\,
            I => \nx.n2894\
        );

    \I__8104\ : Odrv4
    port map (
            O => \N__37333\,
            I => \nx.n2894\
        );

    \I__8103\ : LocalMux
    port map (
            O => \N__37330\,
            I => \nx.n2894\
        );

    \I__8102\ : CascadeMux
    port map (
            O => \N__37323\,
            I => \N__37314\
        );

    \I__8101\ : CascadeMux
    port map (
            O => \N__37322\,
            I => \N__37308\
        );

    \I__8100\ : InMux
    port map (
            O => \N__37321\,
            I => \N__37300\
        );

    \I__8099\ : CascadeMux
    port map (
            O => \N__37320\,
            I => \N__37295\
        );

    \I__8098\ : InMux
    port map (
            O => \N__37319\,
            I => \N__37288\
        );

    \I__8097\ : InMux
    port map (
            O => \N__37318\,
            I => \N__37288\
        );

    \I__8096\ : InMux
    port map (
            O => \N__37317\,
            I => \N__37285\
        );

    \I__8095\ : InMux
    port map (
            O => \N__37314\,
            I => \N__37280\
        );

    \I__8094\ : InMux
    port map (
            O => \N__37313\,
            I => \N__37280\
        );

    \I__8093\ : InMux
    port map (
            O => \N__37312\,
            I => \N__37277\
        );

    \I__8092\ : InMux
    port map (
            O => \N__37311\,
            I => \N__37269\
        );

    \I__8091\ : InMux
    port map (
            O => \N__37308\,
            I => \N__37269\
        );

    \I__8090\ : InMux
    port map (
            O => \N__37307\,
            I => \N__37269\
        );

    \I__8089\ : InMux
    port map (
            O => \N__37306\,
            I => \N__37264\
        );

    \I__8088\ : InMux
    port map (
            O => \N__37305\,
            I => \N__37264\
        );

    \I__8087\ : CascadeMux
    port map (
            O => \N__37304\,
            I => \N__37259\
        );

    \I__8086\ : CascadeMux
    port map (
            O => \N__37303\,
            I => \N__37256\
        );

    \I__8085\ : LocalMux
    port map (
            O => \N__37300\,
            I => \N__37252\
        );

    \I__8084\ : InMux
    port map (
            O => \N__37299\,
            I => \N__37241\
        );

    \I__8083\ : InMux
    port map (
            O => \N__37298\,
            I => \N__37241\
        );

    \I__8082\ : InMux
    port map (
            O => \N__37295\,
            I => \N__37241\
        );

    \I__8081\ : InMux
    port map (
            O => \N__37294\,
            I => \N__37241\
        );

    \I__8080\ : InMux
    port map (
            O => \N__37293\,
            I => \N__37241\
        );

    \I__8079\ : LocalMux
    port map (
            O => \N__37288\,
            I => \N__37232\
        );

    \I__8078\ : LocalMux
    port map (
            O => \N__37285\,
            I => \N__37232\
        );

    \I__8077\ : LocalMux
    port map (
            O => \N__37280\,
            I => \N__37232\
        );

    \I__8076\ : LocalMux
    port map (
            O => \N__37277\,
            I => \N__37232\
        );

    \I__8075\ : CascadeMux
    port map (
            O => \N__37276\,
            I => \N__37228\
        );

    \I__8074\ : LocalMux
    port map (
            O => \N__37269\,
            I => \N__37224\
        );

    \I__8073\ : LocalMux
    port map (
            O => \N__37264\,
            I => \N__37221\
        );

    \I__8072\ : InMux
    port map (
            O => \N__37263\,
            I => \N__37218\
        );

    \I__8071\ : InMux
    port map (
            O => \N__37262\,
            I => \N__37215\
        );

    \I__8070\ : InMux
    port map (
            O => \N__37259\,
            I => \N__37208\
        );

    \I__8069\ : InMux
    port map (
            O => \N__37256\,
            I => \N__37208\
        );

    \I__8068\ : InMux
    port map (
            O => \N__37255\,
            I => \N__37208\
        );

    \I__8067\ : Span4Mux_h
    port map (
            O => \N__37252\,
            I => \N__37201\
        );

    \I__8066\ : LocalMux
    port map (
            O => \N__37241\,
            I => \N__37201\
        );

    \I__8065\ : Span4Mux_v
    port map (
            O => \N__37232\,
            I => \N__37201\
        );

    \I__8064\ : InMux
    port map (
            O => \N__37231\,
            I => \N__37194\
        );

    \I__8063\ : InMux
    port map (
            O => \N__37228\,
            I => \N__37194\
        );

    \I__8062\ : InMux
    port map (
            O => \N__37227\,
            I => \N__37194\
        );

    \I__8061\ : Span4Mux_h
    port map (
            O => \N__37224\,
            I => \N__37189\
        );

    \I__8060\ : Span4Mux_v
    port map (
            O => \N__37221\,
            I => \N__37189\
        );

    \I__8059\ : LocalMux
    port map (
            O => \N__37218\,
            I => \N__37186\
        );

    \I__8058\ : LocalMux
    port map (
            O => \N__37215\,
            I => \nx.n2918\
        );

    \I__8057\ : LocalMux
    port map (
            O => \N__37208\,
            I => \nx.n2918\
        );

    \I__8056\ : Odrv4
    port map (
            O => \N__37201\,
            I => \nx.n2918\
        );

    \I__8055\ : LocalMux
    port map (
            O => \N__37194\,
            I => \nx.n2918\
        );

    \I__8054\ : Odrv4
    port map (
            O => \N__37189\,
            I => \nx.n2918\
        );

    \I__8053\ : Odrv4
    port map (
            O => \N__37186\,
            I => \nx.n2918\
        );

    \I__8052\ : InMux
    port map (
            O => \N__37173\,
            I => \N__37170\
        );

    \I__8051\ : LocalMux
    port map (
            O => \N__37170\,
            I => \nx.n2961\
        );

    \I__8050\ : InMux
    port map (
            O => \N__37167\,
            I => \N__37163\
        );

    \I__8049\ : InMux
    port map (
            O => \N__37166\,
            I => \N__37160\
        );

    \I__8048\ : LocalMux
    port map (
            O => \N__37163\,
            I => \N__37154\
        );

    \I__8047\ : LocalMux
    port map (
            O => \N__37160\,
            I => \N__37154\
        );

    \I__8046\ : InMux
    port map (
            O => \N__37159\,
            I => \N__37151\
        );

    \I__8045\ : Odrv12
    port map (
            O => \N__37154\,
            I => \nx.n2993\
        );

    \I__8044\ : LocalMux
    port map (
            O => \N__37151\,
            I => \nx.n2993\
        );

    \I__8043\ : InMux
    port map (
            O => \N__37146\,
            I => \N__37143\
        );

    \I__8042\ : LocalMux
    port map (
            O => \N__37143\,
            I => \N__37140\
        );

    \I__8041\ : Span4Mux_h
    port map (
            O => \N__37140\,
            I => \N__37137\
        );

    \I__8040\ : Odrv4
    port map (
            O => \N__37137\,
            I => \nx.n40\
        );

    \I__8039\ : CascadeMux
    port map (
            O => \N__37134\,
            I => \nx.n2609_cascade_\
        );

    \I__8038\ : CascadeMux
    port map (
            O => \N__37131\,
            I => \N__37128\
        );

    \I__8037\ : InMux
    port map (
            O => \N__37128\,
            I => \N__37125\
        );

    \I__8036\ : LocalMux
    port map (
            O => \N__37125\,
            I => \nx.n28\
        );

    \I__8035\ : CascadeMux
    port map (
            O => \N__37122\,
            I => \n6_adj_813_cascade_\
        );

    \I__8034\ : InMux
    port map (
            O => \N__37119\,
            I => \N__37116\
        );

    \I__8033\ : LocalMux
    port map (
            O => \N__37116\,
            I => \N__37113\
        );

    \I__8032\ : Span4Mux_v
    port map (
            O => \N__37113\,
            I => \N__37110\
        );

    \I__8031\ : Odrv4
    port map (
            O => \N__37110\,
            I => n11974
        );

    \I__8030\ : CascadeMux
    port map (
            O => \N__37107\,
            I => \N__37104\
        );

    \I__8029\ : InMux
    port map (
            O => \N__37104\,
            I => \N__37099\
        );

    \I__8028\ : CascadeMux
    port map (
            O => \N__37103\,
            I => \N__37096\
        );

    \I__8027\ : InMux
    port map (
            O => \N__37102\,
            I => \N__37093\
        );

    \I__8026\ : LocalMux
    port map (
            O => \N__37099\,
            I => \N__37090\
        );

    \I__8025\ : InMux
    port map (
            O => \N__37096\,
            I => \N__37087\
        );

    \I__8024\ : LocalMux
    port map (
            O => \N__37093\,
            I => \N__37084\
        );

    \I__8023\ : Span4Mux_h
    port map (
            O => \N__37090\,
            I => \N__37081\
        );

    \I__8022\ : LocalMux
    port map (
            O => \N__37087\,
            I => \N__37076\
        );

    \I__8021\ : Span4Mux_h
    port map (
            O => \N__37084\,
            I => \N__37076\
        );

    \I__8020\ : Span4Mux_h
    port map (
            O => \N__37081\,
            I => \N__37073\
        );

    \I__8019\ : Span4Mux_h
    port map (
            O => \N__37076\,
            I => \N__37070\
        );

    \I__8018\ : Odrv4
    port map (
            O => \N__37073\,
            I => \nx.n2890\
        );

    \I__8017\ : Odrv4
    port map (
            O => \N__37070\,
            I => \nx.n2890\
        );

    \I__8016\ : CascadeMux
    port map (
            O => \N__37065\,
            I => \N__37062\
        );

    \I__8015\ : InMux
    port map (
            O => \N__37062\,
            I => \N__37059\
        );

    \I__8014\ : LocalMux
    port map (
            O => \N__37059\,
            I => \N__37056\
        );

    \I__8013\ : Span4Mux_v
    port map (
            O => \N__37056\,
            I => \N__37053\
        );

    \I__8012\ : Span4Mux_h
    port map (
            O => \N__37053\,
            I => \N__37050\
        );

    \I__8011\ : Odrv4
    port map (
            O => \N__37050\,
            I => \nx.n30_adj_759\
        );

    \I__8010\ : InMux
    port map (
            O => \N__37047\,
            I => \N__37044\
        );

    \I__8009\ : LocalMux
    port map (
            O => \N__37044\,
            I => \N__37041\
        );

    \I__8008\ : Span4Mux_v
    port map (
            O => \N__37041\,
            I => \N__37038\
        );

    \I__8007\ : Odrv4
    port map (
            O => \N__37038\,
            I => \nx.n39_adj_761\
        );

    \I__8006\ : InMux
    port map (
            O => \N__37035\,
            I => \N__37032\
        );

    \I__8005\ : LocalMux
    port map (
            O => \N__37032\,
            I => \N__37029\
        );

    \I__8004\ : Span4Mux_v
    port map (
            O => \N__37029\,
            I => \N__37026\
        );

    \I__8003\ : Span4Mux_h
    port map (
            O => \N__37026\,
            I => \N__37023\
        );

    \I__8002\ : Odrv4
    port map (
            O => \N__37023\,
            I => \nx.n42_adj_765\
        );

    \I__8001\ : CascadeMux
    port map (
            O => \N__37020\,
            I => \nx.n45_adj_769_cascade_\
        );

    \I__8000\ : InMux
    port map (
            O => \N__37017\,
            I => \N__37014\
        );

    \I__7999\ : LocalMux
    port map (
            O => \N__37014\,
            I => \nx.n47_adj_770\
        );

    \I__7998\ : CascadeMux
    port map (
            O => \N__37011\,
            I => \N__37008\
        );

    \I__7997\ : InMux
    port map (
            O => \N__37008\,
            I => \N__37004\
        );

    \I__7996\ : InMux
    port map (
            O => \N__37007\,
            I => \N__37001\
        );

    \I__7995\ : LocalMux
    port map (
            O => \N__37004\,
            I => \N__36998\
        );

    \I__7994\ : LocalMux
    port map (
            O => \N__37001\,
            I => \nx.n2896\
        );

    \I__7993\ : Odrv4
    port map (
            O => \N__36998\,
            I => \nx.n2896\
        );

    \I__7992\ : CascadeMux
    port map (
            O => \N__36993\,
            I => \nx.n2918_cascade_\
        );

    \I__7991\ : InMux
    port map (
            O => \N__36990\,
            I => \N__36987\
        );

    \I__7990\ : LocalMux
    port map (
            O => \N__36987\,
            I => \nx.n2963\
        );

    \I__7989\ : InMux
    port map (
            O => \N__36984\,
            I => \N__36981\
        );

    \I__7988\ : LocalMux
    port map (
            O => \N__36981\,
            I => \nx.n2970\
        );

    \I__7987\ : InMux
    port map (
            O => \N__36978\,
            I => \N__36974\
        );

    \I__7986\ : InMux
    port map (
            O => \N__36977\,
            I => \N__36971\
        );

    \I__7985\ : LocalMux
    port map (
            O => \N__36974\,
            I => \N__36966\
        );

    \I__7984\ : LocalMux
    port map (
            O => \N__36971\,
            I => \N__36966\
        );

    \I__7983\ : Span4Mux_h
    port map (
            O => \N__36966\,
            I => \N__36963\
        );

    \I__7982\ : Odrv4
    port map (
            O => \N__36963\,
            I => \nx.n3002\
        );

    \I__7981\ : InMux
    port map (
            O => \N__36960\,
            I => \N__36956\
        );

    \I__7980\ : InMux
    port map (
            O => \N__36959\,
            I => \N__36953\
        );

    \I__7979\ : LocalMux
    port map (
            O => \N__36956\,
            I => \N__36948\
        );

    \I__7978\ : LocalMux
    port map (
            O => \N__36953\,
            I => \N__36948\
        );

    \I__7977\ : Span4Mux_h
    port map (
            O => \N__36948\,
            I => \N__36944\
        );

    \I__7976\ : InMux
    port map (
            O => \N__36947\,
            I => \N__36941\
        );

    \I__7975\ : Odrv4
    port map (
            O => \N__36944\,
            I => \nx.n2995\
        );

    \I__7974\ : LocalMux
    port map (
            O => \N__36941\,
            I => \nx.n2995\
        );

    \I__7973\ : CascadeMux
    port map (
            O => \N__36936\,
            I => \nx.n3002_cascade_\
        );

    \I__7972\ : InMux
    port map (
            O => \N__36933\,
            I => \N__36930\
        );

    \I__7971\ : LocalMux
    port map (
            O => \N__36930\,
            I => \N__36927\
        );

    \I__7970\ : Span4Mux_h
    port map (
            O => \N__36927\,
            I => \N__36924\
        );

    \I__7969\ : Odrv4
    port map (
            O => \N__36924\,
            I => \nx.n42\
        );

    \I__7968\ : InMux
    port map (
            O => \N__36921\,
            I => \N__36918\
        );

    \I__7967\ : LocalMux
    port map (
            O => \N__36918\,
            I => \nx.n2958\
        );

    \I__7966\ : CascadeMux
    port map (
            O => \N__36915\,
            I => \N__36912\
        );

    \I__7965\ : InMux
    port map (
            O => \N__36912\,
            I => \N__36908\
        );

    \I__7964\ : CascadeMux
    port map (
            O => \N__36911\,
            I => \N__36905\
        );

    \I__7963\ : LocalMux
    port map (
            O => \N__36908\,
            I => \N__36901\
        );

    \I__7962\ : InMux
    port map (
            O => \N__36905\,
            I => \N__36898\
        );

    \I__7961\ : CascadeMux
    port map (
            O => \N__36904\,
            I => \N__36895\
        );

    \I__7960\ : Span4Mux_h
    port map (
            O => \N__36901\,
            I => \N__36892\
        );

    \I__7959\ : LocalMux
    port map (
            O => \N__36898\,
            I => \N__36889\
        );

    \I__7958\ : InMux
    port map (
            O => \N__36895\,
            I => \N__36886\
        );

    \I__7957\ : Span4Mux_h
    port map (
            O => \N__36892\,
            I => \N__36883\
        );

    \I__7956\ : Span4Mux_h
    port map (
            O => \N__36889\,
            I => \N__36878\
        );

    \I__7955\ : LocalMux
    port map (
            O => \N__36886\,
            I => \N__36878\
        );

    \I__7954\ : Odrv4
    port map (
            O => \N__36883\,
            I => \nx.n2891\
        );

    \I__7953\ : Odrv4
    port map (
            O => \N__36878\,
            I => \nx.n2891\
        );

    \I__7952\ : InMux
    port map (
            O => \N__36873\,
            I => \N__36868\
        );

    \I__7951\ : InMux
    port map (
            O => \N__36872\,
            I => \N__36865\
        );

    \I__7950\ : InMux
    port map (
            O => \N__36871\,
            I => \N__36862\
        );

    \I__7949\ : LocalMux
    port map (
            O => \N__36868\,
            I => \N__36857\
        );

    \I__7948\ : LocalMux
    port map (
            O => \N__36865\,
            I => \N__36857\
        );

    \I__7947\ : LocalMux
    port map (
            O => \N__36862\,
            I => \N__36854\
        );

    \I__7946\ : Odrv12
    port map (
            O => \N__36857\,
            I => \nx.n2990\
        );

    \I__7945\ : Odrv4
    port map (
            O => \N__36854\,
            I => \nx.n2990\
        );

    \I__7944\ : InMux
    port map (
            O => \N__36849\,
            I => \N__36846\
        );

    \I__7943\ : LocalMux
    port map (
            O => \N__36846\,
            I => \N__36842\
        );

    \I__7942\ : CascadeMux
    port map (
            O => \N__36845\,
            I => \N__36838\
        );

    \I__7941\ : Span12Mux_h
    port map (
            O => \N__36842\,
            I => \N__36835\
        );

    \I__7940\ : InMux
    port map (
            O => \N__36841\,
            I => \N__36832\
        );

    \I__7939\ : InMux
    port map (
            O => \N__36838\,
            I => \N__36829\
        );

    \I__7938\ : Odrv12
    port map (
            O => \N__36835\,
            I => \nx.n2804\
        );

    \I__7937\ : LocalMux
    port map (
            O => \N__36832\,
            I => \nx.n2804\
        );

    \I__7936\ : LocalMux
    port map (
            O => \N__36829\,
            I => \nx.n2804\
        );

    \I__7935\ : CascadeMux
    port map (
            O => \N__36822\,
            I => \N__36819\
        );

    \I__7934\ : InMux
    port map (
            O => \N__36819\,
            I => \N__36816\
        );

    \I__7933\ : LocalMux
    port map (
            O => \N__36816\,
            I => \N__36813\
        );

    \I__7932\ : Span4Mux_h
    port map (
            O => \N__36813\,
            I => \N__36810\
        );

    \I__7931\ : Span4Mux_h
    port map (
            O => \N__36810\,
            I => \N__36807\
        );

    \I__7930\ : Odrv4
    port map (
            O => \N__36807\,
            I => \nx.n2871\
        );

    \I__7929\ : CascadeMux
    port map (
            O => \N__36804\,
            I => \N__36799\
        );

    \I__7928\ : InMux
    port map (
            O => \N__36803\,
            I => \N__36796\
        );

    \I__7927\ : CascadeMux
    port map (
            O => \N__36802\,
            I => \N__36793\
        );

    \I__7926\ : InMux
    port map (
            O => \N__36799\,
            I => \N__36790\
        );

    \I__7925\ : LocalMux
    port map (
            O => \N__36796\,
            I => \N__36787\
        );

    \I__7924\ : InMux
    port map (
            O => \N__36793\,
            I => \N__36784\
        );

    \I__7923\ : LocalMux
    port map (
            O => \N__36790\,
            I => \nx.n2903\
        );

    \I__7922\ : Odrv4
    port map (
            O => \N__36787\,
            I => \nx.n2903\
        );

    \I__7921\ : LocalMux
    port map (
            O => \N__36784\,
            I => \nx.n2903\
        );

    \I__7920\ : IoInMux
    port map (
            O => \N__36777\,
            I => \N__36774\
        );

    \I__7919\ : LocalMux
    port map (
            O => \N__36774\,
            I => \N__36771\
        );

    \I__7918\ : Span12Mux_s4_v
    port map (
            O => \N__36771\,
            I => \N__36768\
        );

    \I__7917\ : Span12Mux_h
    port map (
            O => \N__36768\,
            I => \N__36764\
        );

    \I__7916\ : InMux
    port map (
            O => \N__36767\,
            I => \N__36761\
        );

    \I__7915\ : Odrv12
    port map (
            O => \N__36764\,
            I => pin_oe_9
        );

    \I__7914\ : LocalMux
    port map (
            O => \N__36761\,
            I => pin_oe_9
        );

    \I__7913\ : IoInMux
    port map (
            O => \N__36756\,
            I => \N__36753\
        );

    \I__7912\ : LocalMux
    port map (
            O => \N__36753\,
            I => \N__36750\
        );

    \I__7911\ : Span12Mux_s6_v
    port map (
            O => \N__36750\,
            I => \N__36747\
        );

    \I__7910\ : Span12Mux_h
    port map (
            O => \N__36747\,
            I => \N__36743\
        );

    \I__7909\ : InMux
    port map (
            O => \N__36746\,
            I => \N__36740\
        );

    \I__7908\ : Odrv12
    port map (
            O => \N__36743\,
            I => pin_oe_10
        );

    \I__7907\ : LocalMux
    port map (
            O => \N__36740\,
            I => pin_oe_10
        );

    \I__7906\ : InMux
    port map (
            O => \N__36735\,
            I => \N__36732\
        );

    \I__7905\ : LocalMux
    port map (
            O => \N__36732\,
            I => n11960
        );

    \I__7904\ : InMux
    port map (
            O => \N__36729\,
            I => \N__36726\
        );

    \I__7903\ : LocalMux
    port map (
            O => \N__36726\,
            I => n2618
        );

    \I__7902\ : IoInMux
    port map (
            O => \N__36723\,
            I => \N__36720\
        );

    \I__7901\ : LocalMux
    port map (
            O => \N__36720\,
            I => \N__36717\
        );

    \I__7900\ : Span12Mux_s2_h
    port map (
            O => \N__36717\,
            I => \N__36714\
        );

    \I__7899\ : Span12Mux_h
    port map (
            O => \N__36714\,
            I => \N__36710\
        );

    \I__7898\ : InMux
    port map (
            O => \N__36713\,
            I => \N__36707\
        );

    \I__7897\ : Odrv12
    port map (
            O => \N__36710\,
            I => pin_oe_3
        );

    \I__7896\ : LocalMux
    port map (
            O => \N__36707\,
            I => pin_oe_3
        );

    \I__7895\ : CascadeMux
    port map (
            O => \N__36702\,
            I => \n8_adj_825_cascade_\
        );

    \I__7894\ : IoInMux
    port map (
            O => \N__36699\,
            I => \N__36696\
        );

    \I__7893\ : LocalMux
    port map (
            O => \N__36696\,
            I => \N__36693\
        );

    \I__7892\ : Span12Mux_s7_v
    port map (
            O => \N__36693\,
            I => \N__36690\
        );

    \I__7891\ : Span12Mux_h
    port map (
            O => \N__36690\,
            I => \N__36685\
        );

    \I__7890\ : InMux
    port map (
            O => \N__36689\,
            I => \N__36682\
        );

    \I__7889\ : InMux
    port map (
            O => \N__36688\,
            I => \N__36679\
        );

    \I__7888\ : Odrv12
    port map (
            O => \N__36685\,
            I => pin_out_9
        );

    \I__7887\ : LocalMux
    port map (
            O => \N__36682\,
            I => pin_out_9
        );

    \I__7886\ : LocalMux
    port map (
            O => \N__36679\,
            I => pin_out_9
        );

    \I__7885\ : InMux
    port map (
            O => \N__36672\,
            I => \N__36668\
        );

    \I__7884\ : CascadeMux
    port map (
            O => \N__36671\,
            I => \N__36665\
        );

    \I__7883\ : LocalMux
    port map (
            O => \N__36668\,
            I => \N__36661\
        );

    \I__7882\ : InMux
    port map (
            O => \N__36665\,
            I => \N__36658\
        );

    \I__7881\ : InMux
    port map (
            O => \N__36664\,
            I => \N__36655\
        );

    \I__7880\ : Odrv4
    port map (
            O => \N__36661\,
            I => \nx.n2297\
        );

    \I__7879\ : LocalMux
    port map (
            O => \N__36658\,
            I => \nx.n2297\
        );

    \I__7878\ : LocalMux
    port map (
            O => \N__36655\,
            I => \nx.n2297\
        );

    \I__7877\ : CascadeMux
    port map (
            O => \N__36648\,
            I => \N__36645\
        );

    \I__7876\ : InMux
    port map (
            O => \N__36645\,
            I => \N__36642\
        );

    \I__7875\ : LocalMux
    port map (
            O => \N__36642\,
            I => \nx.n2364\
        );

    \I__7874\ : InMux
    port map (
            O => \N__36639\,
            I => \N__36635\
        );

    \I__7873\ : CascadeMux
    port map (
            O => \N__36638\,
            I => \N__36632\
        );

    \I__7872\ : LocalMux
    port map (
            O => \N__36635\,
            I => \N__36628\
        );

    \I__7871\ : InMux
    port map (
            O => \N__36632\,
            I => \N__36625\
        );

    \I__7870\ : InMux
    port map (
            O => \N__36631\,
            I => \N__36622\
        );

    \I__7869\ : Odrv4
    port map (
            O => \N__36628\,
            I => \nx.n2298\
        );

    \I__7868\ : LocalMux
    port map (
            O => \N__36625\,
            I => \nx.n2298\
        );

    \I__7867\ : LocalMux
    port map (
            O => \N__36622\,
            I => \nx.n2298\
        );

    \I__7866\ : CascadeMux
    port map (
            O => \N__36615\,
            I => \N__36612\
        );

    \I__7865\ : InMux
    port map (
            O => \N__36612\,
            I => \N__36609\
        );

    \I__7864\ : LocalMux
    port map (
            O => \N__36609\,
            I => \nx.n2365\
        );

    \I__7863\ : InMux
    port map (
            O => \N__36606\,
            I => \N__36603\
        );

    \I__7862\ : LocalMux
    port map (
            O => \N__36603\,
            I => \N__36600\
        );

    \I__7861\ : Span4Mux_h
    port map (
            O => \N__36600\,
            I => \N__36597\
        );

    \I__7860\ : Odrv4
    port map (
            O => \N__36597\,
            I => \nx.n2168\
        );

    \I__7859\ : CascadeMux
    port map (
            O => \N__36594\,
            I => \N__36590\
        );

    \I__7858\ : CascadeMux
    port map (
            O => \N__36593\,
            I => \N__36587\
        );

    \I__7857\ : InMux
    port map (
            O => \N__36590\,
            I => \N__36584\
        );

    \I__7856\ : InMux
    port map (
            O => \N__36587\,
            I => \N__36581\
        );

    \I__7855\ : LocalMux
    port map (
            O => \N__36584\,
            I => \N__36577\
        );

    \I__7854\ : LocalMux
    port map (
            O => \N__36581\,
            I => \N__36574\
        );

    \I__7853\ : InMux
    port map (
            O => \N__36580\,
            I => \N__36571\
        );

    \I__7852\ : Odrv12
    port map (
            O => \N__36577\,
            I => \nx.n2101\
        );

    \I__7851\ : Odrv4
    port map (
            O => \N__36574\,
            I => \nx.n2101\
        );

    \I__7850\ : LocalMux
    port map (
            O => \N__36571\,
            I => \nx.n2101\
        );

    \I__7849\ : CascadeMux
    port map (
            O => \N__36564\,
            I => \N__36554\
        );

    \I__7848\ : CascadeMux
    port map (
            O => \N__36563\,
            I => \N__36549\
        );

    \I__7847\ : InMux
    port map (
            O => \N__36562\,
            I => \N__36545\
        );

    \I__7846\ : CascadeMux
    port map (
            O => \N__36561\,
            I => \N__36542\
        );

    \I__7845\ : CascadeMux
    port map (
            O => \N__36560\,
            I => \N__36539\
        );

    \I__7844\ : CascadeMux
    port map (
            O => \N__36559\,
            I => \N__36535\
        );

    \I__7843\ : CascadeMux
    port map (
            O => \N__36558\,
            I => \N__36529\
        );

    \I__7842\ : CascadeMux
    port map (
            O => \N__36557\,
            I => \N__36526\
        );

    \I__7841\ : InMux
    port map (
            O => \N__36554\,
            I => \N__36519\
        );

    \I__7840\ : InMux
    port map (
            O => \N__36553\,
            I => \N__36519\
        );

    \I__7839\ : InMux
    port map (
            O => \N__36552\,
            I => \N__36512\
        );

    \I__7838\ : InMux
    port map (
            O => \N__36549\,
            I => \N__36512\
        );

    \I__7837\ : InMux
    port map (
            O => \N__36548\,
            I => \N__36512\
        );

    \I__7836\ : LocalMux
    port map (
            O => \N__36545\,
            I => \N__36509\
        );

    \I__7835\ : InMux
    port map (
            O => \N__36542\,
            I => \N__36506\
        );

    \I__7834\ : InMux
    port map (
            O => \N__36539\,
            I => \N__36501\
        );

    \I__7833\ : InMux
    port map (
            O => \N__36538\,
            I => \N__36501\
        );

    \I__7832\ : InMux
    port map (
            O => \N__36535\,
            I => \N__36496\
        );

    \I__7831\ : InMux
    port map (
            O => \N__36534\,
            I => \N__36496\
        );

    \I__7830\ : InMux
    port map (
            O => \N__36533\,
            I => \N__36491\
        );

    \I__7829\ : InMux
    port map (
            O => \N__36532\,
            I => \N__36491\
        );

    \I__7828\ : InMux
    port map (
            O => \N__36529\,
            I => \N__36482\
        );

    \I__7827\ : InMux
    port map (
            O => \N__36526\,
            I => \N__36482\
        );

    \I__7826\ : InMux
    port map (
            O => \N__36525\,
            I => \N__36482\
        );

    \I__7825\ : InMux
    port map (
            O => \N__36524\,
            I => \N__36482\
        );

    \I__7824\ : LocalMux
    port map (
            O => \N__36519\,
            I => \N__36475\
        );

    \I__7823\ : LocalMux
    port map (
            O => \N__36512\,
            I => \N__36475\
        );

    \I__7822\ : Span4Mux_v
    port map (
            O => \N__36509\,
            I => \N__36475\
        );

    \I__7821\ : LocalMux
    port map (
            O => \N__36506\,
            I => \N__36472\
        );

    \I__7820\ : LocalMux
    port map (
            O => \N__36501\,
            I => \nx.n2126\
        );

    \I__7819\ : LocalMux
    port map (
            O => \N__36496\,
            I => \nx.n2126\
        );

    \I__7818\ : LocalMux
    port map (
            O => \N__36491\,
            I => \nx.n2126\
        );

    \I__7817\ : LocalMux
    port map (
            O => \N__36482\,
            I => \nx.n2126\
        );

    \I__7816\ : Odrv4
    port map (
            O => \N__36475\,
            I => \nx.n2126\
        );

    \I__7815\ : Odrv12
    port map (
            O => \N__36472\,
            I => \nx.n2126\
        );

    \I__7814\ : CascadeMux
    port map (
            O => \N__36459\,
            I => \N__36456\
        );

    \I__7813\ : InMux
    port map (
            O => \N__36456\,
            I => \N__36451\
        );

    \I__7812\ : InMux
    port map (
            O => \N__36455\,
            I => \N__36448\
        );

    \I__7811\ : InMux
    port map (
            O => \N__36454\,
            I => \N__36445\
        );

    \I__7810\ : LocalMux
    port map (
            O => \N__36451\,
            I => \N__36442\
        );

    \I__7809\ : LocalMux
    port map (
            O => \N__36448\,
            I => \N__36439\
        );

    \I__7808\ : LocalMux
    port map (
            O => \N__36445\,
            I => \N__36436\
        );

    \I__7807\ : Span4Mux_h
    port map (
            O => \N__36442\,
            I => \N__36433\
        );

    \I__7806\ : Span4Mux_h
    port map (
            O => \N__36439\,
            I => \N__36430\
        );

    \I__7805\ : Odrv4
    port map (
            O => \N__36436\,
            I => \nx.n2200\
        );

    \I__7804\ : Odrv4
    port map (
            O => \N__36433\,
            I => \nx.n2200\
        );

    \I__7803\ : Odrv4
    port map (
            O => \N__36430\,
            I => \nx.n2200\
        );

    \I__7802\ : InMux
    port map (
            O => \N__36423\,
            I => \N__36419\
        );

    \I__7801\ : CascadeMux
    port map (
            O => \N__36422\,
            I => \N__36416\
        );

    \I__7800\ : LocalMux
    port map (
            O => \N__36419\,
            I => \N__36412\
        );

    \I__7799\ : InMux
    port map (
            O => \N__36416\,
            I => \N__36409\
        );

    \I__7798\ : InMux
    port map (
            O => \N__36415\,
            I => \N__36406\
        );

    \I__7797\ : Span4Mux_h
    port map (
            O => \N__36412\,
            I => \N__36401\
        );

    \I__7796\ : LocalMux
    port map (
            O => \N__36409\,
            I => \N__36401\
        );

    \I__7795\ : LocalMux
    port map (
            O => \N__36406\,
            I => \nx.n2301\
        );

    \I__7794\ : Odrv4
    port map (
            O => \N__36401\,
            I => \nx.n2301\
        );

    \I__7793\ : CascadeMux
    port map (
            O => \N__36396\,
            I => \N__36393\
        );

    \I__7792\ : InMux
    port map (
            O => \N__36393\,
            I => \N__36390\
        );

    \I__7791\ : LocalMux
    port map (
            O => \N__36390\,
            I => \nx.n2368\
        );

    \I__7790\ : CascadeMux
    port map (
            O => \N__36387\,
            I => \n7602_cascade_\
        );

    \I__7789\ : CascadeMux
    port map (
            O => \N__36384\,
            I => \n7730_cascade_\
        );

    \I__7788\ : InMux
    port map (
            O => \N__36381\,
            I => \nx.n10931\
        );

    \I__7787\ : InMux
    port map (
            O => \N__36378\,
            I => \nx.n10932\
        );

    \I__7786\ : InMux
    port map (
            O => \N__36375\,
            I => \bfn_14_26_0_\
        );

    \I__7785\ : InMux
    port map (
            O => \N__36372\,
            I => \nx.n10934\
        );

    \I__7784\ : InMux
    port map (
            O => \N__36369\,
            I => \nx.n10935\
        );

    \I__7783\ : InMux
    port map (
            O => \N__36366\,
            I => \nx.n10936\
        );

    \I__7782\ : CascadeMux
    port map (
            O => \N__36363\,
            I => \N__36360\
        );

    \I__7781\ : InMux
    port map (
            O => \N__36360\,
            I => \N__36356\
        );

    \I__7780\ : InMux
    port map (
            O => \N__36359\,
            I => \N__36353\
        );

    \I__7779\ : LocalMux
    port map (
            O => \N__36356\,
            I => \N__36350\
        );

    \I__7778\ : LocalMux
    port map (
            O => \N__36353\,
            I => \N__36347\
        );

    \I__7777\ : Odrv4
    port map (
            O => \N__36350\,
            I => \nx.n2390\
        );

    \I__7776\ : Odrv4
    port map (
            O => \N__36347\,
            I => \nx.n2390\
        );

    \I__7775\ : InMux
    port map (
            O => \N__36342\,
            I => \nx.n10937\
        );

    \I__7774\ : IoInMux
    port map (
            O => \N__36339\,
            I => \N__36336\
        );

    \I__7773\ : LocalMux
    port map (
            O => \N__36336\,
            I => \N__36333\
        );

    \I__7772\ : Span12Mux_s6_v
    port map (
            O => \N__36333\,
            I => \N__36330\
        );

    \I__7771\ : Span12Mux_h
    port map (
            O => \N__36330\,
            I => \N__36326\
        );

    \I__7770\ : InMux
    port map (
            O => \N__36329\,
            I => \N__36323\
        );

    \I__7769\ : Odrv12
    port map (
            O => \N__36326\,
            I => pin_oe_18
        );

    \I__7768\ : LocalMux
    port map (
            O => \N__36323\,
            I => pin_oe_18
        );

    \I__7767\ : CascadeMux
    port map (
            O => \N__36318\,
            I => \N__36314\
        );

    \I__7766\ : InMux
    port map (
            O => \N__36317\,
            I => \N__36311\
        );

    \I__7765\ : InMux
    port map (
            O => \N__36314\,
            I => \N__36308\
        );

    \I__7764\ : LocalMux
    port map (
            O => \N__36311\,
            I => \N__36302\
        );

    \I__7763\ : LocalMux
    port map (
            O => \N__36308\,
            I => \N__36302\
        );

    \I__7762\ : InMux
    port map (
            O => \N__36307\,
            I => \N__36299\
        );

    \I__7761\ : Odrv4
    port map (
            O => \N__36302\,
            I => \nx.n2295\
        );

    \I__7760\ : LocalMux
    port map (
            O => \N__36299\,
            I => \nx.n2295\
        );

    \I__7759\ : CascadeMux
    port map (
            O => \N__36294\,
            I => \N__36291\
        );

    \I__7758\ : InMux
    port map (
            O => \N__36291\,
            I => \N__36288\
        );

    \I__7757\ : LocalMux
    port map (
            O => \N__36288\,
            I => \nx.n2362\
        );

    \I__7756\ : InMux
    port map (
            O => \N__36285\,
            I => \nx.n10922\
        );

    \I__7755\ : CascadeMux
    port map (
            O => \N__36282\,
            I => \N__36278\
        );

    \I__7754\ : CascadeMux
    port map (
            O => \N__36281\,
            I => \N__36275\
        );

    \I__7753\ : InMux
    port map (
            O => \N__36278\,
            I => \N__36271\
        );

    \I__7752\ : InMux
    port map (
            O => \N__36275\,
            I => \N__36268\
        );

    \I__7751\ : InMux
    port map (
            O => \N__36274\,
            I => \N__36265\
        );

    \I__7750\ : LocalMux
    port map (
            O => \N__36271\,
            I => \nx.n2404\
        );

    \I__7749\ : LocalMux
    port map (
            O => \N__36268\,
            I => \nx.n2404\
        );

    \I__7748\ : LocalMux
    port map (
            O => \N__36265\,
            I => \nx.n2404\
        );

    \I__7747\ : InMux
    port map (
            O => \N__36258\,
            I => \N__36255\
        );

    \I__7746\ : LocalMux
    port map (
            O => \N__36255\,
            I => \nx.n2471\
        );

    \I__7745\ : InMux
    port map (
            O => \N__36252\,
            I => \nx.n10923\
        );

    \I__7744\ : CascadeMux
    port map (
            O => \N__36249\,
            I => \N__36246\
        );

    \I__7743\ : InMux
    port map (
            O => \N__36246\,
            I => \N__36242\
        );

    \I__7742\ : CascadeMux
    port map (
            O => \N__36245\,
            I => \N__36239\
        );

    \I__7741\ : LocalMux
    port map (
            O => \N__36242\,
            I => \N__36235\
        );

    \I__7740\ : InMux
    port map (
            O => \N__36239\,
            I => \N__36232\
        );

    \I__7739\ : InMux
    port map (
            O => \N__36238\,
            I => \N__36229\
        );

    \I__7738\ : Odrv4
    port map (
            O => \N__36235\,
            I => \nx.n2403\
        );

    \I__7737\ : LocalMux
    port map (
            O => \N__36232\,
            I => \nx.n2403\
        );

    \I__7736\ : LocalMux
    port map (
            O => \N__36229\,
            I => \nx.n2403\
        );

    \I__7735\ : InMux
    port map (
            O => \N__36222\,
            I => \N__36219\
        );

    \I__7734\ : LocalMux
    port map (
            O => \N__36219\,
            I => \nx.n2470\
        );

    \I__7733\ : InMux
    port map (
            O => \N__36216\,
            I => \nx.n10924\
        );

    \I__7732\ : CascadeMux
    port map (
            O => \N__36213\,
            I => \N__36209\
        );

    \I__7731\ : InMux
    port map (
            O => \N__36212\,
            I => \N__36206\
        );

    \I__7730\ : InMux
    port map (
            O => \N__36209\,
            I => \N__36203\
        );

    \I__7729\ : LocalMux
    port map (
            O => \N__36206\,
            I => \N__36199\
        );

    \I__7728\ : LocalMux
    port map (
            O => \N__36203\,
            I => \N__36196\
        );

    \I__7727\ : InMux
    port map (
            O => \N__36202\,
            I => \N__36193\
        );

    \I__7726\ : Odrv4
    port map (
            O => \N__36199\,
            I => \nx.n2402\
        );

    \I__7725\ : Odrv4
    port map (
            O => \N__36196\,
            I => \nx.n2402\
        );

    \I__7724\ : LocalMux
    port map (
            O => \N__36193\,
            I => \nx.n2402\
        );

    \I__7723\ : InMux
    port map (
            O => \N__36186\,
            I => \N__36183\
        );

    \I__7722\ : LocalMux
    port map (
            O => \N__36183\,
            I => \N__36180\
        );

    \I__7721\ : Odrv4
    port map (
            O => \N__36180\,
            I => \nx.n2469\
        );

    \I__7720\ : InMux
    port map (
            O => \N__36177\,
            I => \bfn_14_25_0_\
        );

    \I__7719\ : CascadeMux
    port map (
            O => \N__36174\,
            I => \N__36171\
        );

    \I__7718\ : InMux
    port map (
            O => \N__36171\,
            I => \N__36167\
        );

    \I__7717\ : CascadeMux
    port map (
            O => \N__36170\,
            I => \N__36164\
        );

    \I__7716\ : LocalMux
    port map (
            O => \N__36167\,
            I => \N__36161\
        );

    \I__7715\ : InMux
    port map (
            O => \N__36164\,
            I => \N__36158\
        );

    \I__7714\ : Span4Mux_h
    port map (
            O => \N__36161\,
            I => \N__36155\
        );

    \I__7713\ : LocalMux
    port map (
            O => \N__36158\,
            I => \N__36152\
        );

    \I__7712\ : Odrv4
    port map (
            O => \N__36155\,
            I => \nx.n2401\
        );

    \I__7711\ : Odrv4
    port map (
            O => \N__36152\,
            I => \nx.n2401\
        );

    \I__7710\ : InMux
    port map (
            O => \N__36147\,
            I => \N__36144\
        );

    \I__7709\ : LocalMux
    port map (
            O => \N__36144\,
            I => \N__36141\
        );

    \I__7708\ : Odrv4
    port map (
            O => \N__36141\,
            I => \nx.n2468\
        );

    \I__7707\ : InMux
    port map (
            O => \N__36138\,
            I => \nx.n10926\
        );

    \I__7706\ : InMux
    port map (
            O => \N__36135\,
            I => \nx.n10927\
        );

    \I__7705\ : CascadeMux
    port map (
            O => \N__36132\,
            I => \N__36128\
        );

    \I__7704\ : CascadeMux
    port map (
            O => \N__36131\,
            I => \N__36124\
        );

    \I__7703\ : InMux
    port map (
            O => \N__36128\,
            I => \N__36121\
        );

    \I__7702\ : CascadeMux
    port map (
            O => \N__36127\,
            I => \N__36118\
        );

    \I__7701\ : InMux
    port map (
            O => \N__36124\,
            I => \N__36115\
        );

    \I__7700\ : LocalMux
    port map (
            O => \N__36121\,
            I => \N__36112\
        );

    \I__7699\ : InMux
    port map (
            O => \N__36118\,
            I => \N__36109\
        );

    \I__7698\ : LocalMux
    port map (
            O => \N__36115\,
            I => \N__36106\
        );

    \I__7697\ : Odrv4
    port map (
            O => \N__36112\,
            I => \nx.n2399\
        );

    \I__7696\ : LocalMux
    port map (
            O => \N__36109\,
            I => \nx.n2399\
        );

    \I__7695\ : Odrv4
    port map (
            O => \N__36106\,
            I => \nx.n2399\
        );

    \I__7694\ : InMux
    port map (
            O => \N__36099\,
            I => \N__36096\
        );

    \I__7693\ : LocalMux
    port map (
            O => \N__36096\,
            I => \N__36093\
        );

    \I__7692\ : Span4Mux_h
    port map (
            O => \N__36093\,
            I => \N__36090\
        );

    \I__7691\ : Odrv4
    port map (
            O => \N__36090\,
            I => \nx.n2466\
        );

    \I__7690\ : InMux
    port map (
            O => \N__36087\,
            I => \nx.n10928\
        );

    \I__7689\ : InMux
    port map (
            O => \N__36084\,
            I => \nx.n10929\
        );

    \I__7688\ : InMux
    port map (
            O => \N__36081\,
            I => \nx.n10930\
        );

    \I__7687\ : CascadeMux
    port map (
            O => \N__36078\,
            I => \nx.n2423_cascade_\
        );

    \I__7686\ : InMux
    port map (
            O => \N__36075\,
            I => \N__36072\
        );

    \I__7685\ : LocalMux
    port map (
            O => \N__36072\,
            I => \N__36068\
        );

    \I__7684\ : InMux
    port map (
            O => \N__36071\,
            I => \N__36065\
        );

    \I__7683\ : Odrv4
    port map (
            O => \N__36068\,
            I => \nx.n2374\
        );

    \I__7682\ : LocalMux
    port map (
            O => \N__36065\,
            I => \nx.n2374\
        );

    \I__7681\ : InMux
    port map (
            O => \N__36060\,
            I => \N__36054\
        );

    \I__7680\ : InMux
    port map (
            O => \N__36059\,
            I => \N__36049\
        );

    \I__7679\ : InMux
    port map (
            O => \N__36058\,
            I => \N__36049\
        );

    \I__7678\ : InMux
    port map (
            O => \N__36057\,
            I => \N__36046\
        );

    \I__7677\ : LocalMux
    port map (
            O => \N__36054\,
            I => \N__36042\
        );

    \I__7676\ : LocalMux
    port map (
            O => \N__36049\,
            I => \N__36039\
        );

    \I__7675\ : LocalMux
    port map (
            O => \N__36046\,
            I => \N__36036\
        );

    \I__7674\ : InMux
    port map (
            O => \N__36045\,
            I => \N__36033\
        );

    \I__7673\ : Span4Mux_v
    port map (
            O => \N__36042\,
            I => \N__36030\
        );

    \I__7672\ : Span12Mux_h
    port map (
            O => \N__36039\,
            I => \N__36027\
        );

    \I__7671\ : Span12Mux_h
    port map (
            O => \N__36036\,
            I => \N__36024\
        );

    \I__7670\ : LocalMux
    port map (
            O => \N__36033\,
            I => \nx.bit_ctr_11\
        );

    \I__7669\ : Odrv4
    port map (
            O => \N__36030\,
            I => \nx.bit_ctr_11\
        );

    \I__7668\ : Odrv12
    port map (
            O => \N__36027\,
            I => \nx.bit_ctr_11\
        );

    \I__7667\ : Odrv12
    port map (
            O => \N__36024\,
            I => \nx.bit_ctr_11\
        );

    \I__7666\ : InMux
    port map (
            O => \N__36015\,
            I => \N__36012\
        );

    \I__7665\ : LocalMux
    port map (
            O => \N__36012\,
            I => \nx.n2477\
        );

    \I__7664\ : InMux
    port map (
            O => \N__36009\,
            I => \bfn_14_24_0_\
        );

    \I__7663\ : InMux
    port map (
            O => \N__36006\,
            I => \nx.n10918\
        );

    \I__7662\ : CascadeMux
    port map (
            O => \N__36003\,
            I => \N__35999\
        );

    \I__7661\ : CascadeMux
    port map (
            O => \N__36002\,
            I => \N__35996\
        );

    \I__7660\ : InMux
    port map (
            O => \N__35999\,
            I => \N__35992\
        );

    \I__7659\ : InMux
    port map (
            O => \N__35996\,
            I => \N__35989\
        );

    \I__7658\ : InMux
    port map (
            O => \N__35995\,
            I => \N__35986\
        );

    \I__7657\ : LocalMux
    port map (
            O => \N__35992\,
            I => \nx.n2408\
        );

    \I__7656\ : LocalMux
    port map (
            O => \N__35989\,
            I => \nx.n2408\
        );

    \I__7655\ : LocalMux
    port map (
            O => \N__35986\,
            I => \nx.n2408\
        );

    \I__7654\ : InMux
    port map (
            O => \N__35979\,
            I => \N__35976\
        );

    \I__7653\ : LocalMux
    port map (
            O => \N__35976\,
            I => \nx.n2475\
        );

    \I__7652\ : InMux
    port map (
            O => \N__35973\,
            I => \nx.n10919\
        );

    \I__7651\ : CascadeMux
    port map (
            O => \N__35970\,
            I => \N__35965\
        );

    \I__7650\ : CascadeMux
    port map (
            O => \N__35969\,
            I => \N__35962\
        );

    \I__7649\ : InMux
    port map (
            O => \N__35968\,
            I => \N__35957\
        );

    \I__7648\ : InMux
    port map (
            O => \N__35965\,
            I => \N__35957\
        );

    \I__7647\ : InMux
    port map (
            O => \N__35962\,
            I => \N__35954\
        );

    \I__7646\ : LocalMux
    port map (
            O => \N__35957\,
            I => \nx.n2407\
        );

    \I__7645\ : LocalMux
    port map (
            O => \N__35954\,
            I => \nx.n2407\
        );

    \I__7644\ : InMux
    port map (
            O => \N__35949\,
            I => \N__35946\
        );

    \I__7643\ : LocalMux
    port map (
            O => \N__35946\,
            I => \nx.n2474\
        );

    \I__7642\ : InMux
    port map (
            O => \N__35943\,
            I => \nx.n10920\
        );

    \I__7641\ : CascadeMux
    port map (
            O => \N__35940\,
            I => \N__35937\
        );

    \I__7640\ : InMux
    port map (
            O => \N__35937\,
            I => \N__35933\
        );

    \I__7639\ : InMux
    port map (
            O => \N__35936\,
            I => \N__35930\
        );

    \I__7638\ : LocalMux
    port map (
            O => \N__35933\,
            I => \nx.n2406\
        );

    \I__7637\ : LocalMux
    port map (
            O => \N__35930\,
            I => \nx.n2406\
        );

    \I__7636\ : CascadeMux
    port map (
            O => \N__35925\,
            I => \N__35922\
        );

    \I__7635\ : InMux
    port map (
            O => \N__35922\,
            I => \N__35919\
        );

    \I__7634\ : LocalMux
    port map (
            O => \N__35919\,
            I => \nx.n2473\
        );

    \I__7633\ : InMux
    port map (
            O => \N__35916\,
            I => \nx.n10921\
        );

    \I__7632\ : InMux
    port map (
            O => \N__35913\,
            I => \N__35909\
        );

    \I__7631\ : CascadeMux
    port map (
            O => \N__35912\,
            I => \N__35906\
        );

    \I__7630\ : LocalMux
    port map (
            O => \N__35909\,
            I => \N__35902\
        );

    \I__7629\ : InMux
    port map (
            O => \N__35906\,
            I => \N__35899\
        );

    \I__7628\ : InMux
    port map (
            O => \N__35905\,
            I => \N__35896\
        );

    \I__7627\ : Odrv4
    port map (
            O => \N__35902\,
            I => \nx.n2405\
        );

    \I__7626\ : LocalMux
    port map (
            O => \N__35899\,
            I => \nx.n2405\
        );

    \I__7625\ : LocalMux
    port map (
            O => \N__35896\,
            I => \nx.n2405\
        );

    \I__7624\ : InMux
    port map (
            O => \N__35889\,
            I => \N__35886\
        );

    \I__7623\ : LocalMux
    port map (
            O => \N__35886\,
            I => \nx.n2472\
        );

    \I__7622\ : InMux
    port map (
            O => \N__35883\,
            I => \N__35880\
        );

    \I__7621\ : LocalMux
    port map (
            O => \N__35880\,
            I => \N__35877\
        );

    \I__7620\ : Odrv12
    port map (
            O => \N__35877\,
            I => \nx.n2953\
        );

    \I__7619\ : InMux
    port map (
            O => \N__35874\,
            I => \bfn_14_22_0_\
        );

    \I__7618\ : CascadeMux
    port map (
            O => \N__35871\,
            I => \N__35868\
        );

    \I__7617\ : InMux
    port map (
            O => \N__35868\,
            I => \N__35865\
        );

    \I__7616\ : LocalMux
    port map (
            O => \N__35865\,
            I => \N__35862\
        );

    \I__7615\ : Span4Mux_v
    port map (
            O => \N__35862\,
            I => \N__35858\
        );

    \I__7614\ : InMux
    port map (
            O => \N__35861\,
            I => \N__35855\
        );

    \I__7613\ : Span4Mux_h
    port map (
            O => \N__35858\,
            I => \N__35850\
        );

    \I__7612\ : LocalMux
    port map (
            O => \N__35855\,
            I => \N__35850\
        );

    \I__7611\ : Odrv4
    port map (
            O => \N__35850\,
            I => \nx.n2885\
        );

    \I__7610\ : InMux
    port map (
            O => \N__35847\,
            I => \nx.n11052\
        );

    \I__7609\ : InMux
    port map (
            O => \N__35844\,
            I => \N__35840\
        );

    \I__7608\ : InMux
    port map (
            O => \N__35843\,
            I => \N__35837\
        );

    \I__7607\ : LocalMux
    port map (
            O => \N__35840\,
            I => \N__35831\
        );

    \I__7606\ : LocalMux
    port map (
            O => \N__35837\,
            I => \N__35831\
        );

    \I__7605\ : InMux
    port map (
            O => \N__35836\,
            I => \N__35828\
        );

    \I__7604\ : Span4Mux_v
    port map (
            O => \N__35831\,
            I => \N__35823\
        );

    \I__7603\ : LocalMux
    port map (
            O => \N__35828\,
            I => \N__35823\
        );

    \I__7602\ : Span4Mux_h
    port map (
            O => \N__35823\,
            I => \N__35820\
        );

    \I__7601\ : Odrv4
    port map (
            O => \N__35820\,
            I => \nx.n2984\
        );

    \I__7600\ : InMux
    port map (
            O => \N__35817\,
            I => \N__35814\
        );

    \I__7599\ : LocalMux
    port map (
            O => \N__35814\,
            I => \nx.n27_adj_757\
        );

    \I__7598\ : InMux
    port map (
            O => \N__35811\,
            I => \N__35808\
        );

    \I__7597\ : LocalMux
    port map (
            O => \N__35808\,
            I => \nx.n36_adj_756\
        );

    \I__7596\ : InMux
    port map (
            O => \N__35805\,
            I => \N__35800\
        );

    \I__7595\ : InMux
    port map (
            O => \N__35804\,
            I => \N__35797\
        );

    \I__7594\ : CascadeMux
    port map (
            O => \N__35803\,
            I => \N__35794\
        );

    \I__7593\ : LocalMux
    port map (
            O => \N__35800\,
            I => \N__35791\
        );

    \I__7592\ : LocalMux
    port map (
            O => \N__35797\,
            I => \N__35788\
        );

    \I__7591\ : InMux
    port map (
            O => \N__35794\,
            I => \N__35785\
        );

    \I__7590\ : Span4Mux_v
    port map (
            O => \N__35791\,
            I => \N__35778\
        );

    \I__7589\ : Span4Mux_v
    port map (
            O => \N__35788\,
            I => \N__35778\
        );

    \I__7588\ : LocalMux
    port map (
            O => \N__35785\,
            I => \N__35778\
        );

    \I__7587\ : Odrv4
    port map (
            O => \N__35778\,
            I => \nx.n2708\
        );

    \I__7586\ : CascadeMux
    port map (
            O => \N__35775\,
            I => \N__35772\
        );

    \I__7585\ : InMux
    port map (
            O => \N__35772\,
            I => \N__35768\
        );

    \I__7584\ : InMux
    port map (
            O => \N__35771\,
            I => \N__35765\
        );

    \I__7583\ : LocalMux
    port map (
            O => \N__35768\,
            I => \N__35761\
        );

    \I__7582\ : LocalMux
    port map (
            O => \N__35765\,
            I => \N__35758\
        );

    \I__7581\ : InMux
    port map (
            O => \N__35764\,
            I => \N__35755\
        );

    \I__7580\ : Span4Mux_h
    port map (
            O => \N__35761\,
            I => \N__35752\
        );

    \I__7579\ : Odrv12
    port map (
            O => \N__35758\,
            I => \nx.n2703\
        );

    \I__7578\ : LocalMux
    port map (
            O => \N__35755\,
            I => \nx.n2703\
        );

    \I__7577\ : Odrv4
    port map (
            O => \N__35752\,
            I => \nx.n2703\
        );

    \I__7576\ : InMux
    port map (
            O => \N__35745\,
            I => \N__35742\
        );

    \I__7575\ : LocalMux
    port map (
            O => \N__35742\,
            I => \N__35739\
        );

    \I__7574\ : Odrv12
    port map (
            O => \N__35739\,
            I => \nx.n39_adj_689\
        );

    \I__7573\ : CascadeMux
    port map (
            O => \N__35736\,
            I => \nx.n25_adj_702_cascade_\
        );

    \I__7572\ : InMux
    port map (
            O => \N__35733\,
            I => \N__35730\
        );

    \I__7571\ : LocalMux
    port map (
            O => \N__35730\,
            I => \N__35727\
        );

    \I__7570\ : Span4Mux_h
    port map (
            O => \N__35727\,
            I => \N__35724\
        );

    \I__7569\ : Odrv4
    port map (
            O => \N__35724\,
            I => \nx.n34_adj_701\
        );

    \I__7568\ : InMux
    port map (
            O => \N__35721\,
            I => \N__35718\
        );

    \I__7567\ : LocalMux
    port map (
            O => \N__35718\,
            I => \N__35715\
        );

    \I__7566\ : Odrv4
    port map (
            O => \N__35715\,
            I => \nx.n35_adj_708\
        );

    \I__7565\ : InMux
    port map (
            O => \N__35712\,
            I => \N__35709\
        );

    \I__7564\ : LocalMux
    port map (
            O => \N__35709\,
            I => \nx.n32_adj_703\
        );

    \I__7563\ : CascadeMux
    port map (
            O => \N__35706\,
            I => \nx.n37_adj_709_cascade_\
        );

    \I__7562\ : InMux
    port map (
            O => \N__35703\,
            I => \N__35700\
        );

    \I__7561\ : LocalMux
    port map (
            O => \N__35700\,
            I => \N__35697\
        );

    \I__7560\ : Span4Mux_v
    port map (
            O => \N__35697\,
            I => \N__35694\
        );

    \I__7559\ : Odrv4
    port map (
            O => \N__35694\,
            I => \nx.n31_adj_707\
        );

    \I__7558\ : InMux
    port map (
            O => \N__35691\,
            I => \bfn_14_21_0_\
        );

    \I__7557\ : InMux
    port map (
            O => \N__35688\,
            I => \nx.n11044\
        );

    \I__7556\ : InMux
    port map (
            O => \N__35685\,
            I => \N__35682\
        );

    \I__7555\ : LocalMux
    port map (
            O => \N__35682\,
            I => \nx.n2959\
        );

    \I__7554\ : InMux
    port map (
            O => \N__35679\,
            I => \nx.n11045\
        );

    \I__7553\ : InMux
    port map (
            O => \N__35676\,
            I => \nx.n11046\
        );

    \I__7552\ : InMux
    port map (
            O => \N__35673\,
            I => \N__35670\
        );

    \I__7551\ : LocalMux
    port map (
            O => \N__35670\,
            I => \N__35667\
        );

    \I__7550\ : Span4Mux_h
    port map (
            O => \N__35667\,
            I => \N__35664\
        );

    \I__7549\ : Odrv4
    port map (
            O => \N__35664\,
            I => \nx.n2957\
        );

    \I__7548\ : InMux
    port map (
            O => \N__35661\,
            I => \nx.n11047\
        );

    \I__7547\ : CascadeMux
    port map (
            O => \N__35658\,
            I => \N__35654\
        );

    \I__7546\ : InMux
    port map (
            O => \N__35657\,
            I => \N__35651\
        );

    \I__7545\ : InMux
    port map (
            O => \N__35654\,
            I => \N__35648\
        );

    \I__7544\ : LocalMux
    port map (
            O => \N__35651\,
            I => \N__35643\
        );

    \I__7543\ : LocalMux
    port map (
            O => \N__35648\,
            I => \N__35643\
        );

    \I__7542\ : Span4Mux_h
    port map (
            O => \N__35643\,
            I => \N__35640\
        );

    \I__7541\ : Odrv4
    port map (
            O => \N__35640\,
            I => \nx.n2889\
        );

    \I__7540\ : CascadeMux
    port map (
            O => \N__35637\,
            I => \N__35634\
        );

    \I__7539\ : InMux
    port map (
            O => \N__35634\,
            I => \N__35631\
        );

    \I__7538\ : LocalMux
    port map (
            O => \N__35631\,
            I => \N__35628\
        );

    \I__7537\ : Odrv4
    port map (
            O => \N__35628\,
            I => \nx.n2956\
        );

    \I__7536\ : InMux
    port map (
            O => \N__35625\,
            I => \nx.n11048\
        );

    \I__7535\ : CascadeMux
    port map (
            O => \N__35622\,
            I => \N__35619\
        );

    \I__7534\ : InMux
    port map (
            O => \N__35619\,
            I => \N__35616\
        );

    \I__7533\ : LocalMux
    port map (
            O => \N__35616\,
            I => \N__35613\
        );

    \I__7532\ : Span4Mux_v
    port map (
            O => \N__35613\,
            I => \N__35608\
        );

    \I__7531\ : InMux
    port map (
            O => \N__35612\,
            I => \N__35605\
        );

    \I__7530\ : InMux
    port map (
            O => \N__35611\,
            I => \N__35602\
        );

    \I__7529\ : Span4Mux_h
    port map (
            O => \N__35608\,
            I => \N__35599\
        );

    \I__7528\ : LocalMux
    port map (
            O => \N__35605\,
            I => \N__35596\
        );

    \I__7527\ : LocalMux
    port map (
            O => \N__35602\,
            I => \nx.n2888\
        );

    \I__7526\ : Odrv4
    port map (
            O => \N__35599\,
            I => \nx.n2888\
        );

    \I__7525\ : Odrv4
    port map (
            O => \N__35596\,
            I => \nx.n2888\
        );

    \I__7524\ : CascadeMux
    port map (
            O => \N__35589\,
            I => \N__35586\
        );

    \I__7523\ : InMux
    port map (
            O => \N__35586\,
            I => \N__35583\
        );

    \I__7522\ : LocalMux
    port map (
            O => \N__35583\,
            I => \N__35580\
        );

    \I__7521\ : Span4Mux_h
    port map (
            O => \N__35580\,
            I => \N__35577\
        );

    \I__7520\ : Odrv4
    port map (
            O => \N__35577\,
            I => \nx.n2955\
        );

    \I__7519\ : InMux
    port map (
            O => \N__35574\,
            I => \nx.n11049\
        );

    \I__7518\ : CascadeMux
    port map (
            O => \N__35571\,
            I => \N__35567\
        );

    \I__7517\ : InMux
    port map (
            O => \N__35570\,
            I => \N__35564\
        );

    \I__7516\ : InMux
    port map (
            O => \N__35567\,
            I => \N__35561\
        );

    \I__7515\ : LocalMux
    port map (
            O => \N__35564\,
            I => \N__35555\
        );

    \I__7514\ : LocalMux
    port map (
            O => \N__35561\,
            I => \N__35555\
        );

    \I__7513\ : InMux
    port map (
            O => \N__35560\,
            I => \N__35552\
        );

    \I__7512\ : Odrv4
    port map (
            O => \N__35555\,
            I => \nx.n2887\
        );

    \I__7511\ : LocalMux
    port map (
            O => \N__35552\,
            I => \nx.n2887\
        );

    \I__7510\ : CascadeMux
    port map (
            O => \N__35547\,
            I => \N__35544\
        );

    \I__7509\ : InMux
    port map (
            O => \N__35544\,
            I => \N__35541\
        );

    \I__7508\ : LocalMux
    port map (
            O => \N__35541\,
            I => \nx.n2954\
        );

    \I__7507\ : InMux
    port map (
            O => \N__35538\,
            I => \nx.n11050\
        );

    \I__7506\ : CascadeMux
    port map (
            O => \N__35535\,
            I => \N__35532\
        );

    \I__7505\ : InMux
    port map (
            O => \N__35532\,
            I => \N__35529\
        );

    \I__7504\ : LocalMux
    port map (
            O => \N__35529\,
            I => \N__35525\
        );

    \I__7503\ : InMux
    port map (
            O => \N__35528\,
            I => \N__35522\
        );

    \I__7502\ : Odrv4
    port map (
            O => \N__35525\,
            I => \nx.n2886\
        );

    \I__7501\ : LocalMux
    port map (
            O => \N__35522\,
            I => \nx.n2886\
        );

    \I__7500\ : CascadeMux
    port map (
            O => \N__35517\,
            I => \N__35512\
        );

    \I__7499\ : CascadeMux
    port map (
            O => \N__35516\,
            I => \N__35509\
        );

    \I__7498\ : InMux
    port map (
            O => \N__35515\,
            I => \N__35506\
        );

    \I__7497\ : InMux
    port map (
            O => \N__35512\,
            I => \N__35503\
        );

    \I__7496\ : InMux
    port map (
            O => \N__35509\,
            I => \N__35500\
        );

    \I__7495\ : LocalMux
    port map (
            O => \N__35506\,
            I => \N__35497\
        );

    \I__7494\ : LocalMux
    port map (
            O => \N__35503\,
            I => \N__35494\
        );

    \I__7493\ : LocalMux
    port map (
            O => \N__35500\,
            I => \N__35491\
        );

    \I__7492\ : Span4Mux_v
    port map (
            O => \N__35497\,
            I => \N__35486\
        );

    \I__7491\ : Span4Mux_h
    port map (
            O => \N__35494\,
            I => \N__35486\
        );

    \I__7490\ : Odrv4
    port map (
            O => \N__35491\,
            I => \nx.n2902\
        );

    \I__7489\ : Odrv4
    port map (
            O => \N__35486\,
            I => \nx.n2902\
        );

    \I__7488\ : CascadeMux
    port map (
            O => \N__35481\,
            I => \N__35478\
        );

    \I__7487\ : InMux
    port map (
            O => \N__35478\,
            I => \N__35475\
        );

    \I__7486\ : LocalMux
    port map (
            O => \N__35475\,
            I => \N__35472\
        );

    \I__7485\ : Span4Mux_v
    port map (
            O => \N__35472\,
            I => \N__35469\
        );

    \I__7484\ : Odrv4
    port map (
            O => \N__35469\,
            I => \nx.n2969\
        );

    \I__7483\ : InMux
    port map (
            O => \N__35466\,
            I => \bfn_14_20_0_\
        );

    \I__7482\ : CascadeMux
    port map (
            O => \N__35463\,
            I => \N__35459\
        );

    \I__7481\ : InMux
    port map (
            O => \N__35462\,
            I => \N__35456\
        );

    \I__7480\ : InMux
    port map (
            O => \N__35459\,
            I => \N__35453\
        );

    \I__7479\ : LocalMux
    port map (
            O => \N__35456\,
            I => \N__35450\
        );

    \I__7478\ : LocalMux
    port map (
            O => \N__35453\,
            I => \N__35446\
        );

    \I__7477\ : Span4Mux_v
    port map (
            O => \N__35450\,
            I => \N__35443\
        );

    \I__7476\ : InMux
    port map (
            O => \N__35449\,
            I => \N__35440\
        );

    \I__7475\ : Span4Mux_h
    port map (
            O => \N__35446\,
            I => \N__35437\
        );

    \I__7474\ : Odrv4
    port map (
            O => \N__35443\,
            I => \nx.n2901\
        );

    \I__7473\ : LocalMux
    port map (
            O => \N__35440\,
            I => \nx.n2901\
        );

    \I__7472\ : Odrv4
    port map (
            O => \N__35437\,
            I => \nx.n2901\
        );

    \I__7471\ : CascadeMux
    port map (
            O => \N__35430\,
            I => \N__35427\
        );

    \I__7470\ : InMux
    port map (
            O => \N__35427\,
            I => \N__35424\
        );

    \I__7469\ : LocalMux
    port map (
            O => \N__35424\,
            I => \N__35421\
        );

    \I__7468\ : Span4Mux_v
    port map (
            O => \N__35421\,
            I => \N__35418\
        );

    \I__7467\ : Odrv4
    port map (
            O => \N__35418\,
            I => \nx.n2968\
        );

    \I__7466\ : InMux
    port map (
            O => \N__35415\,
            I => \nx.n11036\
        );

    \I__7465\ : InMux
    port map (
            O => \N__35412\,
            I => \N__35408\
        );

    \I__7464\ : CascadeMux
    port map (
            O => \N__35411\,
            I => \N__35405\
        );

    \I__7463\ : LocalMux
    port map (
            O => \N__35408\,
            I => \N__35402\
        );

    \I__7462\ : InMux
    port map (
            O => \N__35405\,
            I => \N__35398\
        );

    \I__7461\ : Span4Mux_v
    port map (
            O => \N__35402\,
            I => \N__35395\
        );

    \I__7460\ : InMux
    port map (
            O => \N__35401\,
            I => \N__35392\
        );

    \I__7459\ : LocalMux
    port map (
            O => \N__35398\,
            I => \N__35389\
        );

    \I__7458\ : Odrv4
    port map (
            O => \N__35395\,
            I => \nx.n2900\
        );

    \I__7457\ : LocalMux
    port map (
            O => \N__35392\,
            I => \nx.n2900\
        );

    \I__7456\ : Odrv12
    port map (
            O => \N__35389\,
            I => \nx.n2900\
        );

    \I__7455\ : InMux
    port map (
            O => \N__35382\,
            I => \N__35379\
        );

    \I__7454\ : LocalMux
    port map (
            O => \N__35379\,
            I => \N__35376\
        );

    \I__7453\ : Odrv4
    port map (
            O => \N__35376\,
            I => \nx.n2967\
        );

    \I__7452\ : InMux
    port map (
            O => \N__35373\,
            I => \nx.n11037\
        );

    \I__7451\ : CascadeMux
    port map (
            O => \N__35370\,
            I => \N__35366\
        );

    \I__7450\ : InMux
    port map (
            O => \N__35369\,
            I => \N__35363\
        );

    \I__7449\ : InMux
    port map (
            O => \N__35366\,
            I => \N__35360\
        );

    \I__7448\ : LocalMux
    port map (
            O => \N__35363\,
            I => \N__35357\
        );

    \I__7447\ : LocalMux
    port map (
            O => \N__35360\,
            I => \N__35353\
        );

    \I__7446\ : Span4Mux_h
    port map (
            O => \N__35357\,
            I => \N__35350\
        );

    \I__7445\ : InMux
    port map (
            O => \N__35356\,
            I => \N__35347\
        );

    \I__7444\ : Span4Mux_h
    port map (
            O => \N__35353\,
            I => \N__35344\
        );

    \I__7443\ : Span4Mux_v
    port map (
            O => \N__35350\,
            I => \N__35341\
        );

    \I__7442\ : LocalMux
    port map (
            O => \N__35347\,
            I => \nx.n2899\
        );

    \I__7441\ : Odrv4
    port map (
            O => \N__35344\,
            I => \nx.n2899\
        );

    \I__7440\ : Odrv4
    port map (
            O => \N__35341\,
            I => \nx.n2899\
        );

    \I__7439\ : InMux
    port map (
            O => \N__35334\,
            I => \N__35331\
        );

    \I__7438\ : LocalMux
    port map (
            O => \N__35331\,
            I => \N__35328\
        );

    \I__7437\ : Span4Mux_h
    port map (
            O => \N__35328\,
            I => \N__35325\
        );

    \I__7436\ : Odrv4
    port map (
            O => \N__35325\,
            I => \nx.n2966\
        );

    \I__7435\ : InMux
    port map (
            O => \N__35322\,
            I => \nx.n11038\
        );

    \I__7434\ : InMux
    port map (
            O => \N__35319\,
            I => \N__35316\
        );

    \I__7433\ : LocalMux
    port map (
            O => \N__35316\,
            I => \N__35313\
        );

    \I__7432\ : Odrv12
    port map (
            O => \N__35313\,
            I => \nx.n2965\
        );

    \I__7431\ : InMux
    port map (
            O => \N__35310\,
            I => \nx.n11039\
        );

    \I__7430\ : InMux
    port map (
            O => \N__35307\,
            I => \N__35304\
        );

    \I__7429\ : LocalMux
    port map (
            O => \N__35304\,
            I => \N__35301\
        );

    \I__7428\ : Span4Mux_v
    port map (
            O => \N__35301\,
            I => \N__35298\
        );

    \I__7427\ : Odrv4
    port map (
            O => \N__35298\,
            I => \nx.n2964\
        );

    \I__7426\ : InMux
    port map (
            O => \N__35295\,
            I => \nx.n11040\
        );

    \I__7425\ : InMux
    port map (
            O => \N__35292\,
            I => \nx.n11041\
        );

    \I__7424\ : CascadeMux
    port map (
            O => \N__35289\,
            I => \N__35286\
        );

    \I__7423\ : InMux
    port map (
            O => \N__35286\,
            I => \N__35283\
        );

    \I__7422\ : LocalMux
    port map (
            O => \N__35283\,
            I => \N__35279\
        );

    \I__7421\ : InMux
    port map (
            O => \N__35282\,
            I => \N__35276\
        );

    \I__7420\ : Odrv4
    port map (
            O => \N__35279\,
            I => \nx.n2895\
        );

    \I__7419\ : LocalMux
    port map (
            O => \N__35276\,
            I => \nx.n2895\
        );

    \I__7418\ : InMux
    port map (
            O => \N__35271\,
            I => \N__35268\
        );

    \I__7417\ : LocalMux
    port map (
            O => \N__35268\,
            I => \N__35265\
        );

    \I__7416\ : Odrv4
    port map (
            O => \N__35265\,
            I => \nx.n2962\
        );

    \I__7415\ : InMux
    port map (
            O => \N__35262\,
            I => \nx.n11042\
        );

    \I__7414\ : InMux
    port map (
            O => \N__35259\,
            I => \N__35254\
        );

    \I__7413\ : InMux
    port map (
            O => \N__35258\,
            I => \N__35251\
        );

    \I__7412\ : InMux
    port map (
            O => \N__35257\,
            I => \N__35248\
        );

    \I__7411\ : LocalMux
    port map (
            O => \N__35254\,
            I => \N__35245\
        );

    \I__7410\ : LocalMux
    port map (
            O => \N__35251\,
            I => \N__35242\
        );

    \I__7409\ : LocalMux
    port map (
            O => \N__35248\,
            I => \N__35239\
        );

    \I__7408\ : Span4Mux_h
    port map (
            O => \N__35245\,
            I => \N__35234\
        );

    \I__7407\ : Span4Mux_h
    port map (
            O => \N__35242\,
            I => \N__35234\
        );

    \I__7406\ : Span4Mux_h
    port map (
            O => \N__35239\,
            I => \N__35229\
        );

    \I__7405\ : Span4Mux_v
    port map (
            O => \N__35234\,
            I => \N__35226\
        );

    \I__7404\ : InMux
    port map (
            O => \N__35233\,
            I => \N__35223\
        );

    \I__7403\ : InMux
    port map (
            O => \N__35232\,
            I => \N__35220\
        );

    \I__7402\ : Span4Mux_h
    port map (
            O => \N__35229\,
            I => \N__35217\
        );

    \I__7401\ : Span4Mux_h
    port map (
            O => \N__35226\,
            I => \N__35214\
        );

    \I__7400\ : LocalMux
    port map (
            O => \N__35223\,
            I => \nx.bit_ctr_6\
        );

    \I__7399\ : LocalMux
    port map (
            O => \N__35220\,
            I => \nx.bit_ctr_6\
        );

    \I__7398\ : Odrv4
    port map (
            O => \N__35217\,
            I => \nx.bit_ctr_6\
        );

    \I__7397\ : Odrv4
    port map (
            O => \N__35214\,
            I => \nx.bit_ctr_6\
        );

    \I__7396\ : InMux
    port map (
            O => \N__35205\,
            I => \N__35202\
        );

    \I__7395\ : LocalMux
    port map (
            O => \N__35202\,
            I => \N__35199\
        );

    \I__7394\ : Span4Mux_h
    port map (
            O => \N__35199\,
            I => \N__35196\
        );

    \I__7393\ : Odrv4
    port map (
            O => \N__35196\,
            I => \nx.n2977\
        );

    \I__7392\ : InMux
    port map (
            O => \N__35193\,
            I => \bfn_14_19_0_\
        );

    \I__7391\ : CascadeMux
    port map (
            O => \N__35190\,
            I => \N__35187\
        );

    \I__7390\ : InMux
    port map (
            O => \N__35187\,
            I => \N__35182\
        );

    \I__7389\ : InMux
    port map (
            O => \N__35186\,
            I => \N__35179\
        );

    \I__7388\ : InMux
    port map (
            O => \N__35185\,
            I => \N__35176\
        );

    \I__7387\ : LocalMux
    port map (
            O => \N__35182\,
            I => \N__35173\
        );

    \I__7386\ : LocalMux
    port map (
            O => \N__35179\,
            I => \nx.n2909\
        );

    \I__7385\ : LocalMux
    port map (
            O => \N__35176\,
            I => \nx.n2909\
        );

    \I__7384\ : Odrv12
    port map (
            O => \N__35173\,
            I => \nx.n2909\
        );

    \I__7383\ : InMux
    port map (
            O => \N__35166\,
            I => \N__35163\
        );

    \I__7382\ : LocalMux
    port map (
            O => \N__35163\,
            I => \N__35160\
        );

    \I__7381\ : Span4Mux_h
    port map (
            O => \N__35160\,
            I => \N__35157\
        );

    \I__7380\ : Odrv4
    port map (
            O => \N__35157\,
            I => \nx.n2976\
        );

    \I__7379\ : InMux
    port map (
            O => \N__35154\,
            I => \nx.n11028\
        );

    \I__7378\ : InMux
    port map (
            O => \N__35151\,
            I => \N__35147\
        );

    \I__7377\ : CascadeMux
    port map (
            O => \N__35150\,
            I => \N__35143\
        );

    \I__7376\ : LocalMux
    port map (
            O => \N__35147\,
            I => \N__35140\
        );

    \I__7375\ : CascadeMux
    port map (
            O => \N__35146\,
            I => \N__35137\
        );

    \I__7374\ : InMux
    port map (
            O => \N__35143\,
            I => \N__35134\
        );

    \I__7373\ : Span4Mux_v
    port map (
            O => \N__35140\,
            I => \N__35131\
        );

    \I__7372\ : InMux
    port map (
            O => \N__35137\,
            I => \N__35128\
        );

    \I__7371\ : LocalMux
    port map (
            O => \N__35134\,
            I => \N__35121\
        );

    \I__7370\ : Sp12to4
    port map (
            O => \N__35131\,
            I => \N__35121\
        );

    \I__7369\ : LocalMux
    port map (
            O => \N__35128\,
            I => \N__35121\
        );

    \I__7368\ : Odrv12
    port map (
            O => \N__35121\,
            I => \nx.n2908\
        );

    \I__7367\ : InMux
    port map (
            O => \N__35118\,
            I => \N__35115\
        );

    \I__7366\ : LocalMux
    port map (
            O => \N__35115\,
            I => \N__35112\
        );

    \I__7365\ : Odrv12
    port map (
            O => \N__35112\,
            I => \nx.n2975\
        );

    \I__7364\ : InMux
    port map (
            O => \N__35109\,
            I => \nx.n11029\
        );

    \I__7363\ : InMux
    port map (
            O => \N__35106\,
            I => \N__35100\
        );

    \I__7362\ : InMux
    port map (
            O => \N__35105\,
            I => \N__35100\
        );

    \I__7361\ : LocalMux
    port map (
            O => \N__35100\,
            I => \N__35096\
        );

    \I__7360\ : CascadeMux
    port map (
            O => \N__35099\,
            I => \N__35093\
        );

    \I__7359\ : Span4Mux_v
    port map (
            O => \N__35096\,
            I => \N__35090\
        );

    \I__7358\ : InMux
    port map (
            O => \N__35093\,
            I => \N__35087\
        );

    \I__7357\ : Sp12to4
    port map (
            O => \N__35090\,
            I => \N__35082\
        );

    \I__7356\ : LocalMux
    port map (
            O => \N__35087\,
            I => \N__35082\
        );

    \I__7355\ : Odrv12
    port map (
            O => \N__35082\,
            I => \nx.n2907\
        );

    \I__7354\ : InMux
    port map (
            O => \N__35079\,
            I => \N__35076\
        );

    \I__7353\ : LocalMux
    port map (
            O => \N__35076\,
            I => \nx.n2974\
        );

    \I__7352\ : InMux
    port map (
            O => \N__35073\,
            I => \nx.n11030\
        );

    \I__7351\ : CascadeMux
    port map (
            O => \N__35070\,
            I => \N__35066\
        );

    \I__7350\ : InMux
    port map (
            O => \N__35069\,
            I => \N__35062\
        );

    \I__7349\ : InMux
    port map (
            O => \N__35066\,
            I => \N__35059\
        );

    \I__7348\ : CascadeMux
    port map (
            O => \N__35065\,
            I => \N__35056\
        );

    \I__7347\ : LocalMux
    port map (
            O => \N__35062\,
            I => \N__35051\
        );

    \I__7346\ : LocalMux
    port map (
            O => \N__35059\,
            I => \N__35051\
        );

    \I__7345\ : InMux
    port map (
            O => \N__35056\,
            I => \N__35048\
        );

    \I__7344\ : Span4Mux_h
    port map (
            O => \N__35051\,
            I => \N__35045\
        );

    \I__7343\ : LocalMux
    port map (
            O => \N__35048\,
            I => \nx.n2906\
        );

    \I__7342\ : Odrv4
    port map (
            O => \N__35045\,
            I => \nx.n2906\
        );

    \I__7341\ : InMux
    port map (
            O => \N__35040\,
            I => \N__35037\
        );

    \I__7340\ : LocalMux
    port map (
            O => \N__35037\,
            I => \N__35034\
        );

    \I__7339\ : Odrv4
    port map (
            O => \N__35034\,
            I => \nx.n2973\
        );

    \I__7338\ : InMux
    port map (
            O => \N__35031\,
            I => \nx.n11031\
        );

    \I__7337\ : InMux
    port map (
            O => \N__35028\,
            I => \N__35021\
        );

    \I__7336\ : InMux
    port map (
            O => \N__35027\,
            I => \N__35021\
        );

    \I__7335\ : InMux
    port map (
            O => \N__35026\,
            I => \N__35018\
        );

    \I__7334\ : LocalMux
    port map (
            O => \N__35021\,
            I => \nx.n2905\
        );

    \I__7333\ : LocalMux
    port map (
            O => \N__35018\,
            I => \nx.n2905\
        );

    \I__7332\ : CascadeMux
    port map (
            O => \N__35013\,
            I => \N__35010\
        );

    \I__7331\ : InMux
    port map (
            O => \N__35010\,
            I => \N__35007\
        );

    \I__7330\ : LocalMux
    port map (
            O => \N__35007\,
            I => \nx.n2972\
        );

    \I__7329\ : InMux
    port map (
            O => \N__35004\,
            I => \nx.n11032\
        );

    \I__7328\ : CascadeMux
    port map (
            O => \N__35001\,
            I => \N__34998\
        );

    \I__7327\ : InMux
    port map (
            O => \N__34998\,
            I => \N__34995\
        );

    \I__7326\ : LocalMux
    port map (
            O => \N__34995\,
            I => \N__34992\
        );

    \I__7325\ : Odrv4
    port map (
            O => \N__34992\,
            I => \nx.n2971\
        );

    \I__7324\ : InMux
    port map (
            O => \N__34989\,
            I => \nx.n11033\
        );

    \I__7323\ : InMux
    port map (
            O => \N__34986\,
            I => \nx.n11034\
        );

    \I__7322\ : CascadeMux
    port map (
            O => \N__34983\,
            I => \N__34980\
        );

    \I__7321\ : InMux
    port map (
            O => \N__34980\,
            I => \N__34977\
        );

    \I__7320\ : LocalMux
    port map (
            O => \N__34977\,
            I => \N__34974\
        );

    \I__7319\ : Span4Mux_h
    port map (
            O => \N__34974\,
            I => \N__34970\
        );

    \I__7318\ : InMux
    port map (
            O => \N__34973\,
            I => \N__34967\
        );

    \I__7317\ : Odrv4
    port map (
            O => \N__34970\,
            I => \nx.n2291\
        );

    \I__7316\ : LocalMux
    port map (
            O => \N__34967\,
            I => \nx.n2291\
        );

    \I__7315\ : InMux
    port map (
            O => \N__34962\,
            I => \nx.n10917\
        );

    \I__7314\ : InMux
    port map (
            O => \N__34959\,
            I => \N__34955\
        );

    \I__7313\ : InMux
    port map (
            O => \N__34958\,
            I => \N__34952\
        );

    \I__7312\ : LocalMux
    port map (
            O => \N__34955\,
            I => \N__34947\
        );

    \I__7311\ : LocalMux
    port map (
            O => \N__34952\,
            I => \N__34947\
        );

    \I__7310\ : Odrv12
    port map (
            O => \N__34947\,
            I => \nx.n3006\
        );

    \I__7309\ : InMux
    port map (
            O => \N__34944\,
            I => \N__34940\
        );

    \I__7308\ : InMux
    port map (
            O => \N__34943\,
            I => \N__34937\
        );

    \I__7307\ : LocalMux
    port map (
            O => \N__34940\,
            I => \N__34931\
        );

    \I__7306\ : LocalMux
    port map (
            O => \N__34937\,
            I => \N__34931\
        );

    \I__7305\ : InMux
    port map (
            O => \N__34936\,
            I => \N__34928\
        );

    \I__7304\ : Odrv12
    port map (
            O => \N__34931\,
            I => \nx.n3004\
        );

    \I__7303\ : LocalMux
    port map (
            O => \N__34928\,
            I => \nx.n3004\
        );

    \I__7302\ : CascadeMux
    port map (
            O => \N__34923\,
            I => \nx.n3006_cascade_\
        );

    \I__7301\ : InMux
    port map (
            O => \N__34920\,
            I => \N__34917\
        );

    \I__7300\ : LocalMux
    port map (
            O => \N__34917\,
            I => \N__34914\
        );

    \I__7299\ : Span4Mux_h
    port map (
            O => \N__34914\,
            I => \N__34911\
        );

    \I__7298\ : Odrv4
    port map (
            O => \N__34911\,
            I => \nx.n43\
        );

    \I__7297\ : InMux
    port map (
            O => \N__34908\,
            I => \N__34904\
        );

    \I__7296\ : InMux
    port map (
            O => \N__34907\,
            I => \N__34901\
        );

    \I__7295\ : LocalMux
    port map (
            O => \N__34904\,
            I => \N__34896\
        );

    \I__7294\ : LocalMux
    port map (
            O => \N__34901\,
            I => \N__34896\
        );

    \I__7293\ : Span4Mux_h
    port map (
            O => \N__34896\,
            I => \N__34892\
        );

    \I__7292\ : InMux
    port map (
            O => \N__34895\,
            I => \N__34889\
        );

    \I__7291\ : Odrv4
    port map (
            O => \N__34892\,
            I => \nx.n2999\
        );

    \I__7290\ : LocalMux
    port map (
            O => \N__34889\,
            I => \nx.n2999\
        );

    \I__7289\ : InMux
    port map (
            O => \N__34884\,
            I => \N__34879\
        );

    \I__7288\ : CascadeMux
    port map (
            O => \N__34883\,
            I => \N__34876\
        );

    \I__7287\ : CascadeMux
    port map (
            O => \N__34882\,
            I => \N__34873\
        );

    \I__7286\ : LocalMux
    port map (
            O => \N__34879\,
            I => \N__34870\
        );

    \I__7285\ : InMux
    port map (
            O => \N__34876\,
            I => \N__34867\
        );

    \I__7284\ : InMux
    port map (
            O => \N__34873\,
            I => \N__34864\
        );

    \I__7283\ : Span4Mux_h
    port map (
            O => \N__34870\,
            I => \N__34859\
        );

    \I__7282\ : LocalMux
    port map (
            O => \N__34867\,
            I => \N__34859\
        );

    \I__7281\ : LocalMux
    port map (
            O => \N__34864\,
            I => \N__34856\
        );

    \I__7280\ : Odrv4
    port map (
            O => \N__34859\,
            I => \nx.n2797\
        );

    \I__7279\ : Odrv4
    port map (
            O => \N__34856\,
            I => \nx.n2797\
        );

    \I__7278\ : InMux
    port map (
            O => \N__34851\,
            I => \N__34848\
        );

    \I__7277\ : LocalMux
    port map (
            O => \N__34848\,
            I => \N__34845\
        );

    \I__7276\ : Span4Mux_h
    port map (
            O => \N__34845\,
            I => \N__34842\
        );

    \I__7275\ : Span4Mux_h
    port map (
            O => \N__34842\,
            I => \N__34839\
        );

    \I__7274\ : Odrv4
    port map (
            O => \N__34839\,
            I => \nx.n2864\
        );

    \I__7273\ : CascadeMux
    port map (
            O => \N__34836\,
            I => \nx.n2896_cascade_\
        );

    \I__7272\ : CascadeMux
    port map (
            O => \N__34833\,
            I => \nx.n43_adj_763_cascade_\
        );

    \I__7271\ : InMux
    port map (
            O => \N__34830\,
            I => \N__34827\
        );

    \I__7270\ : LocalMux
    port map (
            O => \N__34827\,
            I => \N__34824\
        );

    \I__7269\ : Span4Mux_h
    port map (
            O => \N__34824\,
            I => \N__34821\
        );

    \I__7268\ : Odrv4
    port map (
            O => \N__34821\,
            I => \nx.n38_adj_762\
        );

    \I__7267\ : InMux
    port map (
            O => \N__34818\,
            I => \N__34814\
        );

    \I__7266\ : CascadeMux
    port map (
            O => \N__34817\,
            I => \N__34811\
        );

    \I__7265\ : LocalMux
    port map (
            O => \N__34814\,
            I => \N__34808\
        );

    \I__7264\ : InMux
    port map (
            O => \N__34811\,
            I => \N__34805\
        );

    \I__7263\ : Span4Mux_v
    port map (
            O => \N__34808\,
            I => \N__34801\
        );

    \I__7262\ : LocalMux
    port map (
            O => \N__34805\,
            I => \N__34798\
        );

    \I__7261\ : InMux
    port map (
            O => \N__34804\,
            I => \N__34795\
        );

    \I__7260\ : Span4Mux_h
    port map (
            O => \N__34801\,
            I => \N__34790\
        );

    \I__7259\ : Span4Mux_h
    port map (
            O => \N__34798\,
            I => \N__34790\
        );

    \I__7258\ : LocalMux
    port map (
            O => \N__34795\,
            I => \nx.n2806\
        );

    \I__7257\ : Odrv4
    port map (
            O => \N__34790\,
            I => \nx.n2806\
        );

    \I__7256\ : CascadeMux
    port map (
            O => \N__34785\,
            I => \N__34782\
        );

    \I__7255\ : InMux
    port map (
            O => \N__34782\,
            I => \N__34779\
        );

    \I__7254\ : LocalMux
    port map (
            O => \N__34779\,
            I => \N__34776\
        );

    \I__7253\ : Span4Mux_v
    port map (
            O => \N__34776\,
            I => \N__34773\
        );

    \I__7252\ : Span4Mux_h
    port map (
            O => \N__34773\,
            I => \N__34770\
        );

    \I__7251\ : Odrv4
    port map (
            O => \N__34770\,
            I => \nx.n2873\
        );

    \I__7250\ : InMux
    port map (
            O => \N__34767\,
            I => \N__34764\
        );

    \I__7249\ : LocalMux
    port map (
            O => \N__34764\,
            I => \N__34761\
        );

    \I__7248\ : Span4Mux_v
    port map (
            O => \N__34761\,
            I => \N__34757\
        );

    \I__7247\ : InMux
    port map (
            O => \N__34760\,
            I => \N__34754\
        );

    \I__7246\ : Odrv4
    port map (
            O => \N__34757\,
            I => \nx.n2299\
        );

    \I__7245\ : LocalMux
    port map (
            O => \N__34754\,
            I => \nx.n2299\
        );

    \I__7244\ : InMux
    port map (
            O => \N__34749\,
            I => \N__34746\
        );

    \I__7243\ : LocalMux
    port map (
            O => \N__34746\,
            I => \N__34743\
        );

    \I__7242\ : Odrv4
    port map (
            O => \N__34743\,
            I => \nx.n2366\
        );

    \I__7241\ : InMux
    port map (
            O => \N__34740\,
            I => \nx.n10909\
        );

    \I__7240\ : InMux
    port map (
            O => \N__34737\,
            I => \nx.n10910\
        );

    \I__7239\ : InMux
    port map (
            O => \N__34734\,
            I => \nx.n10911\
        );

    \I__7238\ : CascadeMux
    port map (
            O => \N__34731\,
            I => \N__34727\
        );

    \I__7237\ : CascadeMux
    port map (
            O => \N__34730\,
            I => \N__34724\
        );

    \I__7236\ : InMux
    port map (
            O => \N__34727\,
            I => \N__34721\
        );

    \I__7235\ : InMux
    port map (
            O => \N__34724\,
            I => \N__34718\
        );

    \I__7234\ : LocalMux
    port map (
            O => \N__34721\,
            I => \N__34714\
        );

    \I__7233\ : LocalMux
    port map (
            O => \N__34718\,
            I => \N__34711\
        );

    \I__7232\ : InMux
    port map (
            O => \N__34717\,
            I => \N__34708\
        );

    \I__7231\ : Span4Mux_v
    port map (
            O => \N__34714\,
            I => \N__34701\
        );

    \I__7230\ : Span4Mux_v
    port map (
            O => \N__34711\,
            I => \N__34701\
        );

    \I__7229\ : LocalMux
    port map (
            O => \N__34708\,
            I => \N__34701\
        );

    \I__7228\ : Span4Mux_h
    port map (
            O => \N__34701\,
            I => \N__34698\
        );

    \I__7227\ : Odrv4
    port map (
            O => \N__34698\,
            I => \nx.n2296\
        );

    \I__7226\ : InMux
    port map (
            O => \N__34695\,
            I => \N__34692\
        );

    \I__7225\ : LocalMux
    port map (
            O => \N__34692\,
            I => \N__34689\
        );

    \I__7224\ : Odrv12
    port map (
            O => \N__34689\,
            I => \nx.n2363\
        );

    \I__7223\ : InMux
    port map (
            O => \N__34686\,
            I => \nx.n10912\
        );

    \I__7222\ : InMux
    port map (
            O => \N__34683\,
            I => \nx.n10913\
        );

    \I__7221\ : CascadeMux
    port map (
            O => \N__34680\,
            I => \N__34675\
        );

    \I__7220\ : CascadeMux
    port map (
            O => \N__34679\,
            I => \N__34672\
        );

    \I__7219\ : InMux
    port map (
            O => \N__34678\,
            I => \N__34667\
        );

    \I__7218\ : InMux
    port map (
            O => \N__34675\,
            I => \N__34667\
        );

    \I__7217\ : InMux
    port map (
            O => \N__34672\,
            I => \N__34664\
        );

    \I__7216\ : LocalMux
    port map (
            O => \N__34667\,
            I => \N__34661\
        );

    \I__7215\ : LocalMux
    port map (
            O => \N__34664\,
            I => \nx.n2294\
        );

    \I__7214\ : Odrv4
    port map (
            O => \N__34661\,
            I => \nx.n2294\
        );

    \I__7213\ : InMux
    port map (
            O => \N__34656\,
            I => \N__34653\
        );

    \I__7212\ : LocalMux
    port map (
            O => \N__34653\,
            I => \N__34650\
        );

    \I__7211\ : Odrv4
    port map (
            O => \N__34650\,
            I => \nx.n2361\
        );

    \I__7210\ : InMux
    port map (
            O => \N__34647\,
            I => \bfn_13_28_0_\
        );

    \I__7209\ : CascadeMux
    port map (
            O => \N__34644\,
            I => \N__34639\
        );

    \I__7208\ : InMux
    port map (
            O => \N__34643\,
            I => \N__34636\
        );

    \I__7207\ : InMux
    port map (
            O => \N__34642\,
            I => \N__34633\
        );

    \I__7206\ : InMux
    port map (
            O => \N__34639\,
            I => \N__34630\
        );

    \I__7205\ : LocalMux
    port map (
            O => \N__34636\,
            I => \N__34627\
        );

    \I__7204\ : LocalMux
    port map (
            O => \N__34633\,
            I => \nx.n2293\
        );

    \I__7203\ : LocalMux
    port map (
            O => \N__34630\,
            I => \nx.n2293\
        );

    \I__7202\ : Odrv4
    port map (
            O => \N__34627\,
            I => \nx.n2293\
        );

    \I__7201\ : InMux
    port map (
            O => \N__34620\,
            I => \N__34617\
        );

    \I__7200\ : LocalMux
    port map (
            O => \N__34617\,
            I => \nx.n2360\
        );

    \I__7199\ : InMux
    port map (
            O => \N__34614\,
            I => \nx.n10915\
        );

    \I__7198\ : CascadeMux
    port map (
            O => \N__34611\,
            I => \N__34608\
        );

    \I__7197\ : InMux
    port map (
            O => \N__34608\,
            I => \N__34605\
        );

    \I__7196\ : LocalMux
    port map (
            O => \N__34605\,
            I => \N__34602\
        );

    \I__7195\ : Span4Mux_h
    port map (
            O => \N__34602\,
            I => \N__34597\
        );

    \I__7194\ : InMux
    port map (
            O => \N__34601\,
            I => \N__34592\
        );

    \I__7193\ : InMux
    port map (
            O => \N__34600\,
            I => \N__34592\
        );

    \I__7192\ : Odrv4
    port map (
            O => \N__34597\,
            I => \nx.n2292\
        );

    \I__7191\ : LocalMux
    port map (
            O => \N__34592\,
            I => \nx.n2292\
        );

    \I__7190\ : InMux
    port map (
            O => \N__34587\,
            I => \N__34584\
        );

    \I__7189\ : LocalMux
    port map (
            O => \N__34584\,
            I => \N__34581\
        );

    \I__7188\ : Odrv4
    port map (
            O => \N__34581\,
            I => \nx.n2359\
        );

    \I__7187\ : InMux
    port map (
            O => \N__34578\,
            I => \nx.n10916\
        );

    \I__7186\ : InMux
    port map (
            O => \N__34575\,
            I => \nx.n10901\
        );

    \I__7185\ : CascadeMux
    port map (
            O => \N__34572\,
            I => \N__34567\
        );

    \I__7184\ : InMux
    port map (
            O => \N__34571\,
            I => \N__34564\
        );

    \I__7183\ : InMux
    port map (
            O => \N__34570\,
            I => \N__34561\
        );

    \I__7182\ : InMux
    port map (
            O => \N__34567\,
            I => \N__34558\
        );

    \I__7181\ : LocalMux
    port map (
            O => \N__34564\,
            I => \N__34555\
        );

    \I__7180\ : LocalMux
    port map (
            O => \N__34561\,
            I => \nx.n2306\
        );

    \I__7179\ : LocalMux
    port map (
            O => \N__34558\,
            I => \nx.n2306\
        );

    \I__7178\ : Odrv4
    port map (
            O => \N__34555\,
            I => \nx.n2306\
        );

    \I__7177\ : CascadeMux
    port map (
            O => \N__34548\,
            I => \N__34545\
        );

    \I__7176\ : InMux
    port map (
            O => \N__34545\,
            I => \N__34542\
        );

    \I__7175\ : LocalMux
    port map (
            O => \N__34542\,
            I => \nx.n2373\
        );

    \I__7174\ : InMux
    port map (
            O => \N__34539\,
            I => \nx.n10902\
        );

    \I__7173\ : CascadeMux
    port map (
            O => \N__34536\,
            I => \N__34532\
        );

    \I__7172\ : CascadeMux
    port map (
            O => \N__34535\,
            I => \N__34529\
        );

    \I__7171\ : InMux
    port map (
            O => \N__34532\,
            I => \N__34525\
        );

    \I__7170\ : InMux
    port map (
            O => \N__34529\,
            I => \N__34522\
        );

    \I__7169\ : InMux
    port map (
            O => \N__34528\,
            I => \N__34519\
        );

    \I__7168\ : LocalMux
    port map (
            O => \N__34525\,
            I => \N__34516\
        );

    \I__7167\ : LocalMux
    port map (
            O => \N__34522\,
            I => \nx.n2305\
        );

    \I__7166\ : LocalMux
    port map (
            O => \N__34519\,
            I => \nx.n2305\
        );

    \I__7165\ : Odrv4
    port map (
            O => \N__34516\,
            I => \nx.n2305\
        );

    \I__7164\ : InMux
    port map (
            O => \N__34509\,
            I => \N__34506\
        );

    \I__7163\ : LocalMux
    port map (
            O => \N__34506\,
            I => \nx.n2372\
        );

    \I__7162\ : InMux
    port map (
            O => \N__34503\,
            I => \nx.n10903\
        );

    \I__7161\ : CascadeMux
    port map (
            O => \N__34500\,
            I => \N__34495\
        );

    \I__7160\ : InMux
    port map (
            O => \N__34499\,
            I => \N__34492\
        );

    \I__7159\ : InMux
    port map (
            O => \N__34498\,
            I => \N__34489\
        );

    \I__7158\ : InMux
    port map (
            O => \N__34495\,
            I => \N__34486\
        );

    \I__7157\ : LocalMux
    port map (
            O => \N__34492\,
            I => \nx.n2304\
        );

    \I__7156\ : LocalMux
    port map (
            O => \N__34489\,
            I => \nx.n2304\
        );

    \I__7155\ : LocalMux
    port map (
            O => \N__34486\,
            I => \nx.n2304\
        );

    \I__7154\ : InMux
    port map (
            O => \N__34479\,
            I => \N__34476\
        );

    \I__7153\ : LocalMux
    port map (
            O => \N__34476\,
            I => \nx.n2371\
        );

    \I__7152\ : InMux
    port map (
            O => \N__34473\,
            I => \nx.n10904\
        );

    \I__7151\ : CascadeMux
    port map (
            O => \N__34470\,
            I => \N__34466\
        );

    \I__7150\ : InMux
    port map (
            O => \N__34469\,
            I => \N__34463\
        );

    \I__7149\ : InMux
    port map (
            O => \N__34466\,
            I => \N__34460\
        );

    \I__7148\ : LocalMux
    port map (
            O => \N__34463\,
            I => \nx.n2303\
        );

    \I__7147\ : LocalMux
    port map (
            O => \N__34460\,
            I => \nx.n2303\
        );

    \I__7146\ : InMux
    port map (
            O => \N__34455\,
            I => \N__34452\
        );

    \I__7145\ : LocalMux
    port map (
            O => \N__34452\,
            I => \nx.n2370\
        );

    \I__7144\ : InMux
    port map (
            O => \N__34449\,
            I => \nx.n10905\
        );

    \I__7143\ : CascadeMux
    port map (
            O => \N__34446\,
            I => \N__34443\
        );

    \I__7142\ : InMux
    port map (
            O => \N__34443\,
            I => \N__34439\
        );

    \I__7141\ : InMux
    port map (
            O => \N__34442\,
            I => \N__34436\
        );

    \I__7140\ : LocalMux
    port map (
            O => \N__34439\,
            I => \N__34433\
        );

    \I__7139\ : LocalMux
    port map (
            O => \N__34436\,
            I => \nx.n2302\
        );

    \I__7138\ : Odrv4
    port map (
            O => \N__34433\,
            I => \nx.n2302\
        );

    \I__7137\ : InMux
    port map (
            O => \N__34428\,
            I => \N__34425\
        );

    \I__7136\ : LocalMux
    port map (
            O => \N__34425\,
            I => \N__34422\
        );

    \I__7135\ : Odrv4
    port map (
            O => \N__34422\,
            I => \nx.n2369\
        );

    \I__7134\ : InMux
    port map (
            O => \N__34419\,
            I => \bfn_13_27_0_\
        );

    \I__7133\ : InMux
    port map (
            O => \N__34416\,
            I => \nx.n10907\
        );

    \I__7132\ : InMux
    port map (
            O => \N__34413\,
            I => \N__34409\
        );

    \I__7131\ : CascadeMux
    port map (
            O => \N__34412\,
            I => \N__34406\
        );

    \I__7130\ : LocalMux
    port map (
            O => \N__34409\,
            I => \N__34402\
        );

    \I__7129\ : InMux
    port map (
            O => \N__34406\,
            I => \N__34399\
        );

    \I__7128\ : InMux
    port map (
            O => \N__34405\,
            I => \N__34396\
        );

    \I__7127\ : Odrv4
    port map (
            O => \N__34402\,
            I => \nx.n2300\
        );

    \I__7126\ : LocalMux
    port map (
            O => \N__34399\,
            I => \nx.n2300\
        );

    \I__7125\ : LocalMux
    port map (
            O => \N__34396\,
            I => \nx.n2300\
        );

    \I__7124\ : InMux
    port map (
            O => \N__34389\,
            I => \N__34386\
        );

    \I__7123\ : LocalMux
    port map (
            O => \N__34386\,
            I => \N__34383\
        );

    \I__7122\ : Odrv4
    port map (
            O => \N__34383\,
            I => \nx.n2367\
        );

    \I__7121\ : InMux
    port map (
            O => \N__34380\,
            I => \nx.n10908\
        );

    \I__7120\ : CascadeMux
    port map (
            O => \N__34377\,
            I => \nx.n2398_cascade_\
        );

    \I__7119\ : InMux
    port map (
            O => \N__34374\,
            I => \N__34371\
        );

    \I__7118\ : LocalMux
    port map (
            O => \N__34371\,
            I => \N__34368\
        );

    \I__7117\ : Odrv4
    port map (
            O => \N__34368\,
            I => \nx.n31_adj_700\
        );

    \I__7116\ : InMux
    port map (
            O => \N__34365\,
            I => \N__34362\
        );

    \I__7115\ : LocalMux
    port map (
            O => \N__34362\,
            I => \nx.n32_adj_698\
        );

    \I__7114\ : CascadeMux
    port map (
            O => \N__34359\,
            I => \N__34356\
        );

    \I__7113\ : InMux
    port map (
            O => \N__34356\,
            I => \N__34353\
        );

    \I__7112\ : LocalMux
    port map (
            O => \N__34353\,
            I => \nx.n33_adj_699\
        );

    \I__7111\ : InMux
    port map (
            O => \N__34350\,
            I => \N__34347\
        );

    \I__7110\ : LocalMux
    port map (
            O => \N__34347\,
            I => \nx.n34_adj_697\
        );

    \I__7109\ : CascadeMux
    port map (
            O => \N__34344\,
            I => \nx.n2324_cascade_\
        );

    \I__7108\ : InMux
    port map (
            O => \N__34341\,
            I => \N__34337\
        );

    \I__7107\ : InMux
    port map (
            O => \N__34340\,
            I => \N__34334\
        );

    \I__7106\ : LocalMux
    port map (
            O => \N__34337\,
            I => \N__34330\
        );

    \I__7105\ : LocalMux
    port map (
            O => \N__34334\,
            I => \N__34325\
        );

    \I__7104\ : InMux
    port map (
            O => \N__34333\,
            I => \N__34322\
        );

    \I__7103\ : Span4Mux_v
    port map (
            O => \N__34330\,
            I => \N__34319\
        );

    \I__7102\ : InMux
    port map (
            O => \N__34329\,
            I => \N__34316\
        );

    \I__7101\ : InMux
    port map (
            O => \N__34328\,
            I => \N__34313\
        );

    \I__7100\ : Span4Mux_h
    port map (
            O => \N__34325\,
            I => \N__34310\
        );

    \I__7099\ : LocalMux
    port map (
            O => \N__34322\,
            I => \N__34303\
        );

    \I__7098\ : Sp12to4
    port map (
            O => \N__34319\,
            I => \N__34303\
        );

    \I__7097\ : LocalMux
    port map (
            O => \N__34316\,
            I => \N__34303\
        );

    \I__7096\ : LocalMux
    port map (
            O => \N__34313\,
            I => \nx.bit_ctr_12\
        );

    \I__7095\ : Odrv4
    port map (
            O => \N__34310\,
            I => \nx.bit_ctr_12\
        );

    \I__7094\ : Odrv12
    port map (
            O => \N__34303\,
            I => \nx.bit_ctr_12\
        );

    \I__7093\ : InMux
    port map (
            O => \N__34296\,
            I => \N__34293\
        );

    \I__7092\ : LocalMux
    port map (
            O => \N__34293\,
            I => \N__34290\
        );

    \I__7091\ : Odrv4
    port map (
            O => \N__34290\,
            I => \nx.n2377\
        );

    \I__7090\ : InMux
    port map (
            O => \N__34287\,
            I => \bfn_13_26_0_\
        );

    \I__7089\ : CascadeMux
    port map (
            O => \N__34284\,
            I => \N__34281\
        );

    \I__7088\ : InMux
    port map (
            O => \N__34281\,
            I => \N__34277\
        );

    \I__7087\ : InMux
    port map (
            O => \N__34280\,
            I => \N__34274\
        );

    \I__7086\ : LocalMux
    port map (
            O => \N__34277\,
            I => \N__34271\
        );

    \I__7085\ : LocalMux
    port map (
            O => \N__34274\,
            I => \nx.n2309\
        );

    \I__7084\ : Odrv4
    port map (
            O => \N__34271\,
            I => \nx.n2309\
        );

    \I__7083\ : InMux
    port map (
            O => \N__34266\,
            I => \N__34263\
        );

    \I__7082\ : LocalMux
    port map (
            O => \N__34263\,
            I => \N__34260\
        );

    \I__7081\ : Odrv4
    port map (
            O => \N__34260\,
            I => \nx.n2376\
        );

    \I__7080\ : InMux
    port map (
            O => \N__34257\,
            I => \nx.n10899\
        );

    \I__7079\ : CascadeMux
    port map (
            O => \N__34254\,
            I => \N__34251\
        );

    \I__7078\ : InMux
    port map (
            O => \N__34251\,
            I => \N__34246\
        );

    \I__7077\ : InMux
    port map (
            O => \N__34250\,
            I => \N__34243\
        );

    \I__7076\ : InMux
    port map (
            O => \N__34249\,
            I => \N__34240\
        );

    \I__7075\ : LocalMux
    port map (
            O => \N__34246\,
            I => \N__34237\
        );

    \I__7074\ : LocalMux
    port map (
            O => \N__34243\,
            I => \nx.n2308\
        );

    \I__7073\ : LocalMux
    port map (
            O => \N__34240\,
            I => \nx.n2308\
        );

    \I__7072\ : Odrv4
    port map (
            O => \N__34237\,
            I => \nx.n2308\
        );

    \I__7071\ : CascadeMux
    port map (
            O => \N__34230\,
            I => \N__34227\
        );

    \I__7070\ : InMux
    port map (
            O => \N__34227\,
            I => \N__34224\
        );

    \I__7069\ : LocalMux
    port map (
            O => \N__34224\,
            I => \N__34221\
        );

    \I__7068\ : Odrv4
    port map (
            O => \N__34221\,
            I => \nx.n2375\
        );

    \I__7067\ : InMux
    port map (
            O => \N__34218\,
            I => \nx.n10900\
        );

    \I__7066\ : CascadeMux
    port map (
            O => \N__34215\,
            I => \nx.n2507_cascade_\
        );

    \I__7065\ : CascadeMux
    port map (
            O => \N__34212\,
            I => \nx.n2603_cascade_\
        );

    \I__7064\ : InMux
    port map (
            O => \N__34209\,
            I => \N__34205\
        );

    \I__7063\ : CascadeMux
    port map (
            O => \N__34208\,
            I => \N__34202\
        );

    \I__7062\ : LocalMux
    port map (
            O => \N__34205\,
            I => \N__34198\
        );

    \I__7061\ : InMux
    port map (
            O => \N__34202\,
            I => \N__34195\
        );

    \I__7060\ : InMux
    port map (
            O => \N__34201\,
            I => \N__34192\
        );

    \I__7059\ : Span4Mux_h
    port map (
            O => \N__34198\,
            I => \N__34187\
        );

    \I__7058\ : LocalMux
    port map (
            O => \N__34195\,
            I => \N__34187\
        );

    \I__7057\ : LocalMux
    port map (
            O => \N__34192\,
            I => \N__34184\
        );

    \I__7056\ : Span4Mux_h
    port map (
            O => \N__34187\,
            I => \N__34181\
        );

    \I__7055\ : Odrv4
    port map (
            O => \N__34184\,
            I => \nx.n2702\
        );

    \I__7054\ : Odrv4
    port map (
            O => \N__34181\,
            I => \nx.n2702\
        );

    \I__7053\ : InMux
    port map (
            O => \N__34176\,
            I => \N__34173\
        );

    \I__7052\ : LocalMux
    port map (
            O => \N__34173\,
            I => \N__34169\
        );

    \I__7051\ : CascadeMux
    port map (
            O => \N__34172\,
            I => \N__34165\
        );

    \I__7050\ : Span4Mux_h
    port map (
            O => \N__34169\,
            I => \N__34162\
        );

    \I__7049\ : InMux
    port map (
            O => \N__34168\,
            I => \N__34159\
        );

    \I__7048\ : InMux
    port map (
            O => \N__34165\,
            I => \N__34156\
        );

    \I__7047\ : Odrv4
    port map (
            O => \N__34162\,
            I => \nx.n2803\
        );

    \I__7046\ : LocalMux
    port map (
            O => \N__34159\,
            I => \nx.n2803\
        );

    \I__7045\ : LocalMux
    port map (
            O => \N__34156\,
            I => \nx.n2803\
        );

    \I__7044\ : CascadeMux
    port map (
            O => \N__34149\,
            I => \N__34146\
        );

    \I__7043\ : InMux
    port map (
            O => \N__34146\,
            I => \N__34143\
        );

    \I__7042\ : LocalMux
    port map (
            O => \N__34143\,
            I => \N__34140\
        );

    \I__7041\ : Span4Mux_h
    port map (
            O => \N__34140\,
            I => \N__34137\
        );

    \I__7040\ : Odrv4
    port map (
            O => \N__34137\,
            I => \nx.n2870\
        );

    \I__7039\ : CascadeMux
    port map (
            O => \N__34134\,
            I => \nx.n2501_cascade_\
        );

    \I__7038\ : InMux
    port map (
            O => \N__34131\,
            I => \N__34128\
        );

    \I__7037\ : LocalMux
    port map (
            O => \N__34128\,
            I => \N__34123\
        );

    \I__7036\ : InMux
    port map (
            O => \N__34127\,
            I => \N__34120\
        );

    \I__7035\ : InMux
    port map (
            O => \N__34126\,
            I => \N__34117\
        );

    \I__7034\ : Span4Mux_h
    port map (
            O => \N__34123\,
            I => \N__34112\
        );

    \I__7033\ : LocalMux
    port map (
            O => \N__34120\,
            I => \N__34112\
        );

    \I__7032\ : LocalMux
    port map (
            O => \N__34117\,
            I => \N__34109\
        );

    \I__7031\ : Span4Mux_v
    port map (
            O => \N__34112\,
            I => \N__34106\
        );

    \I__7030\ : Span4Mux_h
    port map (
            O => \N__34109\,
            I => \N__34103\
        );

    \I__7029\ : Odrv4
    port map (
            O => \N__34106\,
            I => \nx.n3085\
        );

    \I__7028\ : Odrv4
    port map (
            O => \N__34103\,
            I => \nx.n3085\
        );

    \I__7027\ : InMux
    port map (
            O => \N__34098\,
            I => \N__34095\
        );

    \I__7026\ : LocalMux
    port map (
            O => \N__34095\,
            I => \N__34092\
        );

    \I__7025\ : Span4Mux_h
    port map (
            O => \N__34092\,
            I => \N__34089\
        );

    \I__7024\ : Span4Mux_h
    port map (
            O => \N__34089\,
            I => \N__34086\
        );

    \I__7023\ : Odrv4
    port map (
            O => \N__34086\,
            I => \nx.n3152\
        );

    \I__7022\ : InMux
    port map (
            O => \N__34083\,
            I => \nx.n11103\
        );

    \I__7021\ : InMux
    port map (
            O => \N__34080\,
            I => \N__34075\
        );

    \I__7020\ : InMux
    port map (
            O => \N__34079\,
            I => \N__34072\
        );

    \I__7019\ : InMux
    port map (
            O => \N__34078\,
            I => \N__34069\
        );

    \I__7018\ : LocalMux
    port map (
            O => \N__34075\,
            I => \N__34066\
        );

    \I__7017\ : LocalMux
    port map (
            O => \N__34072\,
            I => \N__34063\
        );

    \I__7016\ : LocalMux
    port map (
            O => \N__34069\,
            I => \N__34060\
        );

    \I__7015\ : Span4Mux_v
    port map (
            O => \N__34066\,
            I => \N__34055\
        );

    \I__7014\ : Span4Mux_v
    port map (
            O => \N__34063\,
            I => \N__34055\
        );

    \I__7013\ : Span4Mux_h
    port map (
            O => \N__34060\,
            I => \N__34052\
        );

    \I__7012\ : Odrv4
    port map (
            O => \N__34055\,
            I => \nx.n3084\
        );

    \I__7011\ : Odrv4
    port map (
            O => \N__34052\,
            I => \nx.n3084\
        );

    \I__7010\ : InMux
    port map (
            O => \N__34047\,
            I => \N__34044\
        );

    \I__7009\ : LocalMux
    port map (
            O => \N__34044\,
            I => \N__34041\
        );

    \I__7008\ : Span12Mux_h
    port map (
            O => \N__34041\,
            I => \N__34038\
        );

    \I__7007\ : Odrv12
    port map (
            O => \N__34038\,
            I => \nx.n3151\
        );

    \I__7006\ : InMux
    port map (
            O => \N__34035\,
            I => \nx.n11104\
        );

    \I__7005\ : CascadeMux
    port map (
            O => \N__34032\,
            I => \N__34029\
        );

    \I__7004\ : InMux
    port map (
            O => \N__34029\,
            I => \N__34017\
        );

    \I__7003\ : InMux
    port map (
            O => \N__34028\,
            I => \N__34017\
        );

    \I__7002\ : InMux
    port map (
            O => \N__34027\,
            I => \N__34017\
        );

    \I__7001\ : InMux
    port map (
            O => \N__34026\,
            I => \N__34014\
        );

    \I__7000\ : CascadeMux
    port map (
            O => \N__34025\,
            I => \N__34011\
        );

    \I__6999\ : CascadeMux
    port map (
            O => \N__34024\,
            I => \N__34008\
        );

    \I__6998\ : LocalMux
    port map (
            O => \N__34017\,
            I => \N__33998\
        );

    \I__6997\ : LocalMux
    port map (
            O => \N__34014\,
            I => \N__33995\
        );

    \I__6996\ : InMux
    port map (
            O => \N__34011\,
            I => \N__33990\
        );

    \I__6995\ : InMux
    port map (
            O => \N__34008\,
            I => \N__33990\
        );

    \I__6994\ : CascadeMux
    port map (
            O => \N__34007\,
            I => \N__33981\
        );

    \I__6993\ : CascadeMux
    port map (
            O => \N__34006\,
            I => \N__33978\
        );

    \I__6992\ : CascadeMux
    port map (
            O => \N__34005\,
            I => \N__33974\
        );

    \I__6991\ : CascadeMux
    port map (
            O => \N__34004\,
            I => \N__33969\
        );

    \I__6990\ : CascadeMux
    port map (
            O => \N__34003\,
            I => \N__33963\
        );

    \I__6989\ : CascadeMux
    port map (
            O => \N__34002\,
            I => \N__33959\
        );

    \I__6988\ : CascadeMux
    port map (
            O => \N__34001\,
            I => \N__33956\
        );

    \I__6987\ : Span4Mux_v
    port map (
            O => \N__33998\,
            I => \N__33948\
        );

    \I__6986\ : Span4Mux_v
    port map (
            O => \N__33995\,
            I => \N__33948\
        );

    \I__6985\ : LocalMux
    port map (
            O => \N__33990\,
            I => \N__33948\
        );

    \I__6984\ : InMux
    port map (
            O => \N__33989\,
            I => \N__33943\
        );

    \I__6983\ : InMux
    port map (
            O => \N__33988\,
            I => \N__33943\
        );

    \I__6982\ : InMux
    port map (
            O => \N__33987\,
            I => \N__33930\
        );

    \I__6981\ : InMux
    port map (
            O => \N__33986\,
            I => \N__33930\
        );

    \I__6980\ : InMux
    port map (
            O => \N__33985\,
            I => \N__33930\
        );

    \I__6979\ : InMux
    port map (
            O => \N__33984\,
            I => \N__33930\
        );

    \I__6978\ : InMux
    port map (
            O => \N__33981\,
            I => \N__33930\
        );

    \I__6977\ : InMux
    port map (
            O => \N__33978\,
            I => \N__33930\
        );

    \I__6976\ : InMux
    port map (
            O => \N__33977\,
            I => \N__33915\
        );

    \I__6975\ : InMux
    port map (
            O => \N__33974\,
            I => \N__33915\
        );

    \I__6974\ : InMux
    port map (
            O => \N__33973\,
            I => \N__33915\
        );

    \I__6973\ : InMux
    port map (
            O => \N__33972\,
            I => \N__33915\
        );

    \I__6972\ : InMux
    port map (
            O => \N__33969\,
            I => \N__33915\
        );

    \I__6971\ : InMux
    port map (
            O => \N__33968\,
            I => \N__33915\
        );

    \I__6970\ : InMux
    port map (
            O => \N__33967\,
            I => \N__33915\
        );

    \I__6969\ : InMux
    port map (
            O => \N__33966\,
            I => \N__33902\
        );

    \I__6968\ : InMux
    port map (
            O => \N__33963\,
            I => \N__33902\
        );

    \I__6967\ : InMux
    port map (
            O => \N__33962\,
            I => \N__33902\
        );

    \I__6966\ : InMux
    port map (
            O => \N__33959\,
            I => \N__33902\
        );

    \I__6965\ : InMux
    port map (
            O => \N__33956\,
            I => \N__33902\
        );

    \I__6964\ : InMux
    port map (
            O => \N__33955\,
            I => \N__33902\
        );

    \I__6963\ : Odrv4
    port map (
            O => \N__33948\,
            I => \nx.n3116\
        );

    \I__6962\ : LocalMux
    port map (
            O => \N__33943\,
            I => \nx.n3116\
        );

    \I__6961\ : LocalMux
    port map (
            O => \N__33930\,
            I => \nx.n3116\
        );

    \I__6960\ : LocalMux
    port map (
            O => \N__33915\,
            I => \nx.n3116\
        );

    \I__6959\ : LocalMux
    port map (
            O => \N__33902\,
            I => \nx.n3116\
        );

    \I__6958\ : CascadeMux
    port map (
            O => \N__33891\,
            I => \N__33888\
        );

    \I__6957\ : InMux
    port map (
            O => \N__33888\,
            I => \N__33884\
        );

    \I__6956\ : InMux
    port map (
            O => \N__33887\,
            I => \N__33881\
        );

    \I__6955\ : LocalMux
    port map (
            O => \N__33884\,
            I => \N__33878\
        );

    \I__6954\ : LocalMux
    port map (
            O => \N__33881\,
            I => \N__33875\
        );

    \I__6953\ : Span4Mux_h
    port map (
            O => \N__33878\,
            I => \N__33872\
        );

    \I__6952\ : Span4Mux_h
    port map (
            O => \N__33875\,
            I => \N__33869\
        );

    \I__6951\ : Odrv4
    port map (
            O => \N__33872\,
            I => \nx.n3083\
        );

    \I__6950\ : Odrv4
    port map (
            O => \N__33869\,
            I => \nx.n3083\
        );

    \I__6949\ : InMux
    port map (
            O => \N__33864\,
            I => \nx.n11105\
        );

    \I__6948\ : InMux
    port map (
            O => \N__33861\,
            I => \N__33858\
        );

    \I__6947\ : LocalMux
    port map (
            O => \N__33858\,
            I => \N__33855\
        );

    \I__6946\ : Span4Mux_v
    port map (
            O => \N__33855\,
            I => \N__33852\
        );

    \I__6945\ : Odrv4
    port map (
            O => \N__33852\,
            I => \nx.n13280\
        );

    \I__6944\ : InMux
    port map (
            O => \N__33849\,
            I => \N__33846\
        );

    \I__6943\ : LocalMux
    port map (
            O => \N__33846\,
            I => \N__33841\
        );

    \I__6942\ : InMux
    port map (
            O => \N__33845\,
            I => \N__33838\
        );

    \I__6941\ : CascadeMux
    port map (
            O => \N__33844\,
            I => \N__33835\
        );

    \I__6940\ : Span4Mux_h
    port map (
            O => \N__33841\,
            I => \N__33832\
        );

    \I__6939\ : LocalMux
    port map (
            O => \N__33838\,
            I => \N__33829\
        );

    \I__6938\ : InMux
    port map (
            O => \N__33835\,
            I => \N__33826\
        );

    \I__6937\ : Odrv4
    port map (
            O => \N__33832\,
            I => \nx.n2805\
        );

    \I__6936\ : Odrv4
    port map (
            O => \N__33829\,
            I => \nx.n2805\
        );

    \I__6935\ : LocalMux
    port map (
            O => \N__33826\,
            I => \nx.n2805\
        );

    \I__6934\ : CascadeMux
    port map (
            O => \N__33819\,
            I => \N__33816\
        );

    \I__6933\ : InMux
    port map (
            O => \N__33816\,
            I => \N__33813\
        );

    \I__6932\ : LocalMux
    port map (
            O => \N__33813\,
            I => \N__33810\
        );

    \I__6931\ : Span4Mux_h
    port map (
            O => \N__33810\,
            I => \N__33807\
        );

    \I__6930\ : Odrv4
    port map (
            O => \N__33807\,
            I => \nx.n2872\
        );

    \I__6929\ : CascadeMux
    port map (
            O => \N__33804\,
            I => \N__33800\
        );

    \I__6928\ : InMux
    port map (
            O => \N__33803\,
            I => \N__33797\
        );

    \I__6927\ : InMux
    port map (
            O => \N__33800\,
            I => \N__33793\
        );

    \I__6926\ : LocalMux
    port map (
            O => \N__33797\,
            I => \N__33790\
        );

    \I__6925\ : InMux
    port map (
            O => \N__33796\,
            I => \N__33787\
        );

    \I__6924\ : LocalMux
    port map (
            O => \N__33793\,
            I => \N__33784\
        );

    \I__6923\ : Span4Mux_h
    port map (
            O => \N__33790\,
            I => \N__33779\
        );

    \I__6922\ : LocalMux
    port map (
            O => \N__33787\,
            I => \N__33779\
        );

    \I__6921\ : Span4Mux_h
    port map (
            O => \N__33784\,
            I => \N__33776\
        );

    \I__6920\ : Odrv4
    port map (
            O => \N__33779\,
            I => \nx.n2798\
        );

    \I__6919\ : Odrv4
    port map (
            O => \N__33776\,
            I => \nx.n2798\
        );

    \I__6918\ : CascadeMux
    port map (
            O => \N__33771\,
            I => \N__33768\
        );

    \I__6917\ : InMux
    port map (
            O => \N__33768\,
            I => \N__33765\
        );

    \I__6916\ : LocalMux
    port map (
            O => \N__33765\,
            I => \N__33762\
        );

    \I__6915\ : Span4Mux_v
    port map (
            O => \N__33762\,
            I => \N__33759\
        );

    \I__6914\ : Span4Mux_h
    port map (
            O => \N__33759\,
            I => \N__33756\
        );

    \I__6913\ : Odrv4
    port map (
            O => \N__33756\,
            I => \nx.n2865\
        );

    \I__6912\ : InMux
    port map (
            O => \N__33753\,
            I => \N__33749\
        );

    \I__6911\ : InMux
    port map (
            O => \N__33752\,
            I => \N__33746\
        );

    \I__6910\ : LocalMux
    port map (
            O => \N__33749\,
            I => \N__33740\
        );

    \I__6909\ : LocalMux
    port map (
            O => \N__33746\,
            I => \N__33740\
        );

    \I__6908\ : InMux
    port map (
            O => \N__33745\,
            I => \N__33737\
        );

    \I__6907\ : Odrv4
    port map (
            O => \N__33740\,
            I => \nx.n2986\
        );

    \I__6906\ : LocalMux
    port map (
            O => \N__33737\,
            I => \nx.n2986\
        );

    \I__6905\ : InMux
    port map (
            O => \N__33732\,
            I => \N__33728\
        );

    \I__6904\ : InMux
    port map (
            O => \N__33731\,
            I => \N__33725\
        );

    \I__6903\ : LocalMux
    port map (
            O => \N__33728\,
            I => \N__33720\
        );

    \I__6902\ : LocalMux
    port map (
            O => \N__33725\,
            I => \N__33720\
        );

    \I__6901\ : Span4Mux_h
    port map (
            O => \N__33720\,
            I => \N__33716\
        );

    \I__6900\ : InMux
    port map (
            O => \N__33719\,
            I => \N__33713\
        );

    \I__6899\ : Odrv4
    port map (
            O => \N__33716\,
            I => \nx.n2991\
        );

    \I__6898\ : LocalMux
    port map (
            O => \N__33713\,
            I => \nx.n2991\
        );

    \I__6897\ : InMux
    port map (
            O => \N__33708\,
            I => \N__33705\
        );

    \I__6896\ : LocalMux
    port map (
            O => \N__33705\,
            I => \N__33702\
        );

    \I__6895\ : Span4Mux_h
    port map (
            O => \N__33702\,
            I => \N__33699\
        );

    \I__6894\ : Odrv4
    port map (
            O => \N__33699\,
            I => \nx.n3160\
        );

    \I__6893\ : InMux
    port map (
            O => \N__33696\,
            I => \nx.n11095\
        );

    \I__6892\ : InMux
    port map (
            O => \N__33693\,
            I => \N__33689\
        );

    \I__6891\ : CascadeMux
    port map (
            O => \N__33692\,
            I => \N__33686\
        );

    \I__6890\ : LocalMux
    port map (
            O => \N__33689\,
            I => \N__33682\
        );

    \I__6889\ : InMux
    port map (
            O => \N__33686\,
            I => \N__33679\
        );

    \I__6888\ : InMux
    port map (
            O => \N__33685\,
            I => \N__33676\
        );

    \I__6887\ : Span4Mux_v
    port map (
            O => \N__33682\,
            I => \N__33673\
        );

    \I__6886\ : LocalMux
    port map (
            O => \N__33679\,
            I => \N__33668\
        );

    \I__6885\ : LocalMux
    port map (
            O => \N__33676\,
            I => \N__33668\
        );

    \I__6884\ : Odrv4
    port map (
            O => \N__33673\,
            I => \nx.n3092\
        );

    \I__6883\ : Odrv4
    port map (
            O => \N__33668\,
            I => \nx.n3092\
        );

    \I__6882\ : InMux
    port map (
            O => \N__33663\,
            I => \N__33660\
        );

    \I__6881\ : LocalMux
    port map (
            O => \N__33660\,
            I => \N__33657\
        );

    \I__6880\ : Span4Mux_v
    port map (
            O => \N__33657\,
            I => \N__33654\
        );

    \I__6879\ : Odrv4
    port map (
            O => \N__33654\,
            I => \nx.n3159\
        );

    \I__6878\ : InMux
    port map (
            O => \N__33651\,
            I => \nx.n11096\
        );

    \I__6877\ : InMux
    port map (
            O => \N__33648\,
            I => \N__33644\
        );

    \I__6876\ : InMux
    port map (
            O => \N__33647\,
            I => \N__33641\
        );

    \I__6875\ : LocalMux
    port map (
            O => \N__33644\,
            I => \N__33637\
        );

    \I__6874\ : LocalMux
    port map (
            O => \N__33641\,
            I => \N__33634\
        );

    \I__6873\ : InMux
    port map (
            O => \N__33640\,
            I => \N__33631\
        );

    \I__6872\ : Span4Mux_v
    port map (
            O => \N__33637\,
            I => \N__33626\
        );

    \I__6871\ : Span4Mux_h
    port map (
            O => \N__33634\,
            I => \N__33626\
        );

    \I__6870\ : LocalMux
    port map (
            O => \N__33631\,
            I => \N__33623\
        );

    \I__6869\ : Odrv4
    port map (
            O => \N__33626\,
            I => \nx.n3091\
        );

    \I__6868\ : Odrv4
    port map (
            O => \N__33623\,
            I => \nx.n3091\
        );

    \I__6867\ : InMux
    port map (
            O => \N__33618\,
            I => \N__33615\
        );

    \I__6866\ : LocalMux
    port map (
            O => \N__33615\,
            I => \N__33612\
        );

    \I__6865\ : Span4Mux_v
    port map (
            O => \N__33612\,
            I => \N__33609\
        );

    \I__6864\ : Odrv4
    port map (
            O => \N__33609\,
            I => \nx.n3158\
        );

    \I__6863\ : InMux
    port map (
            O => \N__33606\,
            I => \nx.n11097\
        );

    \I__6862\ : InMux
    port map (
            O => \N__33603\,
            I => \N__33599\
        );

    \I__6861\ : InMux
    port map (
            O => \N__33602\,
            I => \N__33596\
        );

    \I__6860\ : LocalMux
    port map (
            O => \N__33599\,
            I => \N__33592\
        );

    \I__6859\ : LocalMux
    port map (
            O => \N__33596\,
            I => \N__33589\
        );

    \I__6858\ : InMux
    port map (
            O => \N__33595\,
            I => \N__33586\
        );

    \I__6857\ : Span4Mux_v
    port map (
            O => \N__33592\,
            I => \N__33581\
        );

    \I__6856\ : Span4Mux_h
    port map (
            O => \N__33589\,
            I => \N__33581\
        );

    \I__6855\ : LocalMux
    port map (
            O => \N__33586\,
            I => \N__33578\
        );

    \I__6854\ : Odrv4
    port map (
            O => \N__33581\,
            I => \nx.n3090\
        );

    \I__6853\ : Odrv4
    port map (
            O => \N__33578\,
            I => \nx.n3090\
        );

    \I__6852\ : InMux
    port map (
            O => \N__33573\,
            I => \N__33570\
        );

    \I__6851\ : LocalMux
    port map (
            O => \N__33570\,
            I => \N__33567\
        );

    \I__6850\ : Span4Mux_h
    port map (
            O => \N__33567\,
            I => \N__33564\
        );

    \I__6849\ : Odrv4
    port map (
            O => \N__33564\,
            I => \nx.n3157\
        );

    \I__6848\ : InMux
    port map (
            O => \N__33561\,
            I => \nx.n11098\
        );

    \I__6847\ : InMux
    port map (
            O => \N__33558\,
            I => \N__33555\
        );

    \I__6846\ : LocalMux
    port map (
            O => \N__33555\,
            I => \N__33550\
        );

    \I__6845\ : InMux
    port map (
            O => \N__33554\,
            I => \N__33547\
        );

    \I__6844\ : InMux
    port map (
            O => \N__33553\,
            I => \N__33544\
        );

    \I__6843\ : Span4Mux_h
    port map (
            O => \N__33550\,
            I => \N__33541\
        );

    \I__6842\ : LocalMux
    port map (
            O => \N__33547\,
            I => \N__33536\
        );

    \I__6841\ : LocalMux
    port map (
            O => \N__33544\,
            I => \N__33536\
        );

    \I__6840\ : Odrv4
    port map (
            O => \N__33541\,
            I => \nx.n3089\
        );

    \I__6839\ : Odrv4
    port map (
            O => \N__33536\,
            I => \nx.n3089\
        );

    \I__6838\ : InMux
    port map (
            O => \N__33531\,
            I => \N__33528\
        );

    \I__6837\ : LocalMux
    port map (
            O => \N__33528\,
            I => \N__33525\
        );

    \I__6836\ : Span4Mux_h
    port map (
            O => \N__33525\,
            I => \N__33522\
        );

    \I__6835\ : Odrv4
    port map (
            O => \N__33522\,
            I => \nx.n3156\
        );

    \I__6834\ : InMux
    port map (
            O => \N__33519\,
            I => \nx.n11099\
        );

    \I__6833\ : InMux
    port map (
            O => \N__33516\,
            I => \N__33512\
        );

    \I__6832\ : InMux
    port map (
            O => \N__33515\,
            I => \N__33509\
        );

    \I__6831\ : LocalMux
    port map (
            O => \N__33512\,
            I => \N__33505\
        );

    \I__6830\ : LocalMux
    port map (
            O => \N__33509\,
            I => \N__33502\
        );

    \I__6829\ : InMux
    port map (
            O => \N__33508\,
            I => \N__33499\
        );

    \I__6828\ : Span4Mux_v
    port map (
            O => \N__33505\,
            I => \N__33496\
        );

    \I__6827\ : Span4Mux_h
    port map (
            O => \N__33502\,
            I => \N__33493\
        );

    \I__6826\ : LocalMux
    port map (
            O => \N__33499\,
            I => \N__33490\
        );

    \I__6825\ : Odrv4
    port map (
            O => \N__33496\,
            I => \nx.n3088\
        );

    \I__6824\ : Odrv4
    port map (
            O => \N__33493\,
            I => \nx.n3088\
        );

    \I__6823\ : Odrv4
    port map (
            O => \N__33490\,
            I => \nx.n3088\
        );

    \I__6822\ : InMux
    port map (
            O => \N__33483\,
            I => \N__33480\
        );

    \I__6821\ : LocalMux
    port map (
            O => \N__33480\,
            I => \N__33477\
        );

    \I__6820\ : Span4Mux_h
    port map (
            O => \N__33477\,
            I => \N__33474\
        );

    \I__6819\ : Odrv4
    port map (
            O => \N__33474\,
            I => \nx.n3155\
        );

    \I__6818\ : InMux
    port map (
            O => \N__33471\,
            I => \nx.n11100\
        );

    \I__6817\ : InMux
    port map (
            O => \N__33468\,
            I => \N__33463\
        );

    \I__6816\ : InMux
    port map (
            O => \N__33467\,
            I => \N__33460\
        );

    \I__6815\ : CascadeMux
    port map (
            O => \N__33466\,
            I => \N__33457\
        );

    \I__6814\ : LocalMux
    port map (
            O => \N__33463\,
            I => \N__33454\
        );

    \I__6813\ : LocalMux
    port map (
            O => \N__33460\,
            I => \N__33451\
        );

    \I__6812\ : InMux
    port map (
            O => \N__33457\,
            I => \N__33448\
        );

    \I__6811\ : Span4Mux_h
    port map (
            O => \N__33454\,
            I => \N__33445\
        );

    \I__6810\ : Span4Mux_h
    port map (
            O => \N__33451\,
            I => \N__33442\
        );

    \I__6809\ : LocalMux
    port map (
            O => \N__33448\,
            I => \N__33439\
        );

    \I__6808\ : Odrv4
    port map (
            O => \N__33445\,
            I => \nx.n3087\
        );

    \I__6807\ : Odrv4
    port map (
            O => \N__33442\,
            I => \nx.n3087\
        );

    \I__6806\ : Odrv12
    port map (
            O => \N__33439\,
            I => \nx.n3087\
        );

    \I__6805\ : InMux
    port map (
            O => \N__33432\,
            I => \N__33429\
        );

    \I__6804\ : LocalMux
    port map (
            O => \N__33429\,
            I => \N__33426\
        );

    \I__6803\ : Span4Mux_h
    port map (
            O => \N__33426\,
            I => \N__33423\
        );

    \I__6802\ : Odrv4
    port map (
            O => \N__33423\,
            I => \nx.n3154\
        );

    \I__6801\ : InMux
    port map (
            O => \N__33420\,
            I => \nx.n11101\
        );

    \I__6800\ : InMux
    port map (
            O => \N__33417\,
            I => \N__33414\
        );

    \I__6799\ : LocalMux
    port map (
            O => \N__33414\,
            I => \N__33409\
        );

    \I__6798\ : InMux
    port map (
            O => \N__33413\,
            I => \N__33406\
        );

    \I__6797\ : InMux
    port map (
            O => \N__33412\,
            I => \N__33403\
        );

    \I__6796\ : Span4Mux_h
    port map (
            O => \N__33409\,
            I => \N__33400\
        );

    \I__6795\ : LocalMux
    port map (
            O => \N__33406\,
            I => \N__33397\
        );

    \I__6794\ : LocalMux
    port map (
            O => \N__33403\,
            I => \N__33394\
        );

    \I__6793\ : Odrv4
    port map (
            O => \N__33400\,
            I => \nx.n3086\
        );

    \I__6792\ : Odrv12
    port map (
            O => \N__33397\,
            I => \nx.n3086\
        );

    \I__6791\ : Odrv12
    port map (
            O => \N__33394\,
            I => \nx.n3086\
        );

    \I__6790\ : InMux
    port map (
            O => \N__33387\,
            I => \N__33384\
        );

    \I__6789\ : LocalMux
    port map (
            O => \N__33384\,
            I => \N__33381\
        );

    \I__6788\ : Span4Mux_h
    port map (
            O => \N__33381\,
            I => \N__33378\
        );

    \I__6787\ : Odrv4
    port map (
            O => \N__33378\,
            I => \nx.n3153\
        );

    \I__6786\ : InMux
    port map (
            O => \N__33375\,
            I => \bfn_13_20_0_\
        );

    \I__6785\ : CascadeMux
    port map (
            O => \N__33372\,
            I => \N__33369\
        );

    \I__6784\ : InMux
    port map (
            O => \N__33369\,
            I => \N__33366\
        );

    \I__6783\ : LocalMux
    port map (
            O => \N__33366\,
            I => \N__33362\
        );

    \I__6782\ : InMux
    port map (
            O => \N__33365\,
            I => \N__33358\
        );

    \I__6781\ : Span4Mux_v
    port map (
            O => \N__33362\,
            I => \N__33355\
        );

    \I__6780\ : InMux
    port map (
            O => \N__33361\,
            I => \N__33352\
        );

    \I__6779\ : LocalMux
    port map (
            O => \N__33358\,
            I => \nx.n3100\
        );

    \I__6778\ : Odrv4
    port map (
            O => \N__33355\,
            I => \nx.n3100\
        );

    \I__6777\ : LocalMux
    port map (
            O => \N__33352\,
            I => \nx.n3100\
        );

    \I__6776\ : InMux
    port map (
            O => \N__33345\,
            I => \N__33342\
        );

    \I__6775\ : LocalMux
    port map (
            O => \N__33342\,
            I => \nx.n3167\
        );

    \I__6774\ : InMux
    port map (
            O => \N__33339\,
            I => \nx.n11088\
        );

    \I__6773\ : CascadeMux
    port map (
            O => \N__33336\,
            I => \N__33333\
        );

    \I__6772\ : InMux
    port map (
            O => \N__33333\,
            I => \N__33330\
        );

    \I__6771\ : LocalMux
    port map (
            O => \N__33330\,
            I => \N__33325\
        );

    \I__6770\ : InMux
    port map (
            O => \N__33329\,
            I => \N__33322\
        );

    \I__6769\ : InMux
    port map (
            O => \N__33328\,
            I => \N__33319\
        );

    \I__6768\ : Span4Mux_h
    port map (
            O => \N__33325\,
            I => \N__33316\
        );

    \I__6767\ : LocalMux
    port map (
            O => \N__33322\,
            I => \N__33311\
        );

    \I__6766\ : LocalMux
    port map (
            O => \N__33319\,
            I => \N__33311\
        );

    \I__6765\ : Odrv4
    port map (
            O => \N__33316\,
            I => \nx.n3099\
        );

    \I__6764\ : Odrv4
    port map (
            O => \N__33311\,
            I => \nx.n3099\
        );

    \I__6763\ : InMux
    port map (
            O => \N__33306\,
            I => \N__33303\
        );

    \I__6762\ : LocalMux
    port map (
            O => \N__33303\,
            I => \nx.n3166\
        );

    \I__6761\ : InMux
    port map (
            O => \N__33300\,
            I => \nx.n11089\
        );

    \I__6760\ : CascadeMux
    port map (
            O => \N__33297\,
            I => \N__33294\
        );

    \I__6759\ : InMux
    port map (
            O => \N__33294\,
            I => \N__33290\
        );

    \I__6758\ : InMux
    port map (
            O => \N__33293\,
            I => \N__33287\
        );

    \I__6757\ : LocalMux
    port map (
            O => \N__33290\,
            I => \N__33283\
        );

    \I__6756\ : LocalMux
    port map (
            O => \N__33287\,
            I => \N__33280\
        );

    \I__6755\ : InMux
    port map (
            O => \N__33286\,
            I => \N__33277\
        );

    \I__6754\ : Span4Mux_h
    port map (
            O => \N__33283\,
            I => \N__33274\
        );

    \I__6753\ : Span4Mux_v
    port map (
            O => \N__33280\,
            I => \N__33271\
        );

    \I__6752\ : LocalMux
    port map (
            O => \N__33277\,
            I => \nx.n3098\
        );

    \I__6751\ : Odrv4
    port map (
            O => \N__33274\,
            I => \nx.n3098\
        );

    \I__6750\ : Odrv4
    port map (
            O => \N__33271\,
            I => \nx.n3098\
        );

    \I__6749\ : InMux
    port map (
            O => \N__33264\,
            I => \N__33261\
        );

    \I__6748\ : LocalMux
    port map (
            O => \N__33261\,
            I => \N__33258\
        );

    \I__6747\ : Odrv12
    port map (
            O => \N__33258\,
            I => \nx.n3165\
        );

    \I__6746\ : InMux
    port map (
            O => \N__33255\,
            I => \nx.n11090\
        );

    \I__6745\ : CascadeMux
    port map (
            O => \N__33252\,
            I => \N__33249\
        );

    \I__6744\ : InMux
    port map (
            O => \N__33249\,
            I => \N__33245\
        );

    \I__6743\ : InMux
    port map (
            O => \N__33248\,
            I => \N__33242\
        );

    \I__6742\ : LocalMux
    port map (
            O => \N__33245\,
            I => \N__33239\
        );

    \I__6741\ : LocalMux
    port map (
            O => \N__33242\,
            I => \N__33235\
        );

    \I__6740\ : Span4Mux_h
    port map (
            O => \N__33239\,
            I => \N__33232\
        );

    \I__6739\ : InMux
    port map (
            O => \N__33238\,
            I => \N__33229\
        );

    \I__6738\ : Odrv4
    port map (
            O => \N__33235\,
            I => \nx.n3097\
        );

    \I__6737\ : Odrv4
    port map (
            O => \N__33232\,
            I => \nx.n3097\
        );

    \I__6736\ : LocalMux
    port map (
            O => \N__33229\,
            I => \nx.n3097\
        );

    \I__6735\ : InMux
    port map (
            O => \N__33222\,
            I => \N__33219\
        );

    \I__6734\ : LocalMux
    port map (
            O => \N__33219\,
            I => \nx.n3164\
        );

    \I__6733\ : InMux
    port map (
            O => \N__33216\,
            I => \nx.n11091\
        );

    \I__6732\ : CascadeMux
    port map (
            O => \N__33213\,
            I => \N__33210\
        );

    \I__6731\ : InMux
    port map (
            O => \N__33210\,
            I => \N__33206\
        );

    \I__6730\ : InMux
    port map (
            O => \N__33209\,
            I => \N__33202\
        );

    \I__6729\ : LocalMux
    port map (
            O => \N__33206\,
            I => \N__33199\
        );

    \I__6728\ : CascadeMux
    port map (
            O => \N__33205\,
            I => \N__33196\
        );

    \I__6727\ : LocalMux
    port map (
            O => \N__33202\,
            I => \N__33193\
        );

    \I__6726\ : Span4Mux_h
    port map (
            O => \N__33199\,
            I => \N__33190\
        );

    \I__6725\ : InMux
    port map (
            O => \N__33196\,
            I => \N__33187\
        );

    \I__6724\ : Odrv4
    port map (
            O => \N__33193\,
            I => \nx.n3096\
        );

    \I__6723\ : Odrv4
    port map (
            O => \N__33190\,
            I => \nx.n3096\
        );

    \I__6722\ : LocalMux
    port map (
            O => \N__33187\,
            I => \nx.n3096\
        );

    \I__6721\ : InMux
    port map (
            O => \N__33180\,
            I => \N__33177\
        );

    \I__6720\ : LocalMux
    port map (
            O => \N__33177\,
            I => \nx.n3163\
        );

    \I__6719\ : InMux
    port map (
            O => \N__33174\,
            I => \nx.n11092\
        );

    \I__6718\ : CascadeMux
    port map (
            O => \N__33171\,
            I => \N__33168\
        );

    \I__6717\ : InMux
    port map (
            O => \N__33168\,
            I => \N__33165\
        );

    \I__6716\ : LocalMux
    port map (
            O => \N__33165\,
            I => \N__33160\
        );

    \I__6715\ : InMux
    port map (
            O => \N__33164\,
            I => \N__33157\
        );

    \I__6714\ : InMux
    port map (
            O => \N__33163\,
            I => \N__33154\
        );

    \I__6713\ : Span4Mux_h
    port map (
            O => \N__33160\,
            I => \N__33151\
        );

    \I__6712\ : LocalMux
    port map (
            O => \N__33157\,
            I => \N__33148\
        );

    \I__6711\ : LocalMux
    port map (
            O => \N__33154\,
            I => \nx.n3095\
        );

    \I__6710\ : Odrv4
    port map (
            O => \N__33151\,
            I => \nx.n3095\
        );

    \I__6709\ : Odrv12
    port map (
            O => \N__33148\,
            I => \nx.n3095\
        );

    \I__6708\ : InMux
    port map (
            O => \N__33141\,
            I => \N__33138\
        );

    \I__6707\ : LocalMux
    port map (
            O => \N__33138\,
            I => \nx.n3162\
        );

    \I__6706\ : InMux
    port map (
            O => \N__33135\,
            I => \nx.n11093\
        );

    \I__6705\ : InMux
    port map (
            O => \N__33132\,
            I => \N__33128\
        );

    \I__6704\ : InMux
    port map (
            O => \N__33131\,
            I => \N__33125\
        );

    \I__6703\ : LocalMux
    port map (
            O => \N__33128\,
            I => \N__33121\
        );

    \I__6702\ : LocalMux
    port map (
            O => \N__33125\,
            I => \N__33118\
        );

    \I__6701\ : InMux
    port map (
            O => \N__33124\,
            I => \N__33115\
        );

    \I__6700\ : Span4Mux_h
    port map (
            O => \N__33121\,
            I => \N__33110\
        );

    \I__6699\ : Span4Mux_h
    port map (
            O => \N__33118\,
            I => \N__33110\
        );

    \I__6698\ : LocalMux
    port map (
            O => \N__33115\,
            I => \nx.n3094\
        );

    \I__6697\ : Odrv4
    port map (
            O => \N__33110\,
            I => \nx.n3094\
        );

    \I__6696\ : CascadeMux
    port map (
            O => \N__33105\,
            I => \N__33102\
        );

    \I__6695\ : InMux
    port map (
            O => \N__33102\,
            I => \N__33099\
        );

    \I__6694\ : LocalMux
    port map (
            O => \N__33099\,
            I => \nx.n3161\
        );

    \I__6693\ : InMux
    port map (
            O => \N__33096\,
            I => \bfn_13_19_0_\
        );

    \I__6692\ : CascadeMux
    port map (
            O => \N__33093\,
            I => \N__33089\
        );

    \I__6691\ : InMux
    port map (
            O => \N__33092\,
            I => \N__33086\
        );

    \I__6690\ : InMux
    port map (
            O => \N__33089\,
            I => \N__33082\
        );

    \I__6689\ : LocalMux
    port map (
            O => \N__33086\,
            I => \N__33079\
        );

    \I__6688\ : InMux
    port map (
            O => \N__33085\,
            I => \N__33076\
        );

    \I__6687\ : LocalMux
    port map (
            O => \N__33082\,
            I => \N__33073\
        );

    \I__6686\ : Span4Mux_v
    port map (
            O => \N__33079\,
            I => \N__33070\
        );

    \I__6685\ : LocalMux
    port map (
            O => \N__33076\,
            I => \N__33067\
        );

    \I__6684\ : Span4Mux_v
    port map (
            O => \N__33073\,
            I => \N__33064\
        );

    \I__6683\ : Span4Mux_h
    port map (
            O => \N__33070\,
            I => \N__33061\
        );

    \I__6682\ : Odrv4
    port map (
            O => \N__33067\,
            I => \nx.n3093\
        );

    \I__6681\ : Odrv4
    port map (
            O => \N__33064\,
            I => \nx.n3093\
        );

    \I__6680\ : Odrv4
    port map (
            O => \N__33061\,
            I => \nx.n3093\
        );

    \I__6679\ : CascadeMux
    port map (
            O => \N__33054\,
            I => \N__33051\
        );

    \I__6678\ : InMux
    port map (
            O => \N__33051\,
            I => \N__33047\
        );

    \I__6677\ : CascadeMux
    port map (
            O => \N__33050\,
            I => \N__33044\
        );

    \I__6676\ : LocalMux
    port map (
            O => \N__33047\,
            I => \N__33040\
        );

    \I__6675\ : InMux
    port map (
            O => \N__33044\,
            I => \N__33035\
        );

    \I__6674\ : InMux
    port map (
            O => \N__33043\,
            I => \N__33035\
        );

    \I__6673\ : Span4Mux_v
    port map (
            O => \N__33040\,
            I => \N__33032\
        );

    \I__6672\ : LocalMux
    port map (
            O => \N__33035\,
            I => \nx.n3108\
        );

    \I__6671\ : Odrv4
    port map (
            O => \N__33032\,
            I => \nx.n3108\
        );

    \I__6670\ : InMux
    port map (
            O => \N__33027\,
            I => \N__33024\
        );

    \I__6669\ : LocalMux
    port map (
            O => \N__33024\,
            I => \N__33021\
        );

    \I__6668\ : Span4Mux_h
    port map (
            O => \N__33021\,
            I => \N__33018\
        );

    \I__6667\ : Odrv4
    port map (
            O => \N__33018\,
            I => \nx.n3175\
        );

    \I__6666\ : InMux
    port map (
            O => \N__33015\,
            I => \nx.n11080\
        );

    \I__6665\ : CascadeMux
    port map (
            O => \N__33012\,
            I => \N__33009\
        );

    \I__6664\ : InMux
    port map (
            O => \N__33009\,
            I => \N__33006\
        );

    \I__6663\ : LocalMux
    port map (
            O => \N__33006\,
            I => \N__33001\
        );

    \I__6662\ : InMux
    port map (
            O => \N__33005\,
            I => \N__32998\
        );

    \I__6661\ : InMux
    port map (
            O => \N__33004\,
            I => \N__32995\
        );

    \I__6660\ : Span4Mux_h
    port map (
            O => \N__33001\,
            I => \N__32992\
        );

    \I__6659\ : LocalMux
    port map (
            O => \N__32998\,
            I => \nx.n3107\
        );

    \I__6658\ : LocalMux
    port map (
            O => \N__32995\,
            I => \nx.n3107\
        );

    \I__6657\ : Odrv4
    port map (
            O => \N__32992\,
            I => \nx.n3107\
        );

    \I__6656\ : InMux
    port map (
            O => \N__32985\,
            I => \N__32982\
        );

    \I__6655\ : LocalMux
    port map (
            O => \N__32982\,
            I => \nx.n3174\
        );

    \I__6654\ : InMux
    port map (
            O => \N__32979\,
            I => \nx.n11081\
        );

    \I__6653\ : CascadeMux
    port map (
            O => \N__32976\,
            I => \N__32972\
        );

    \I__6652\ : InMux
    port map (
            O => \N__32975\,
            I => \N__32969\
        );

    \I__6651\ : InMux
    port map (
            O => \N__32972\,
            I => \N__32966\
        );

    \I__6650\ : LocalMux
    port map (
            O => \N__32969\,
            I => \N__32963\
        );

    \I__6649\ : LocalMux
    port map (
            O => \N__32966\,
            I => \N__32959\
        );

    \I__6648\ : Span4Mux_v
    port map (
            O => \N__32963\,
            I => \N__32956\
        );

    \I__6647\ : InMux
    port map (
            O => \N__32962\,
            I => \N__32953\
        );

    \I__6646\ : Span4Mux_h
    port map (
            O => \N__32959\,
            I => \N__32948\
        );

    \I__6645\ : Span4Mux_h
    port map (
            O => \N__32956\,
            I => \N__32948\
        );

    \I__6644\ : LocalMux
    port map (
            O => \N__32953\,
            I => \nx.n3106\
        );

    \I__6643\ : Odrv4
    port map (
            O => \N__32948\,
            I => \nx.n3106\
        );

    \I__6642\ : InMux
    port map (
            O => \N__32943\,
            I => \N__32940\
        );

    \I__6641\ : LocalMux
    port map (
            O => \N__32940\,
            I => \N__32937\
        );

    \I__6640\ : Odrv4
    port map (
            O => \N__32937\,
            I => \nx.n3173\
        );

    \I__6639\ : InMux
    port map (
            O => \N__32934\,
            I => \nx.n11082\
        );

    \I__6638\ : CascadeMux
    port map (
            O => \N__32931\,
            I => \N__32928\
        );

    \I__6637\ : InMux
    port map (
            O => \N__32928\,
            I => \N__32925\
        );

    \I__6636\ : LocalMux
    port map (
            O => \N__32925\,
            I => \N__32920\
        );

    \I__6635\ : InMux
    port map (
            O => \N__32924\,
            I => \N__32917\
        );

    \I__6634\ : InMux
    port map (
            O => \N__32923\,
            I => \N__32914\
        );

    \I__6633\ : Span4Mux_h
    port map (
            O => \N__32920\,
            I => \N__32911\
        );

    \I__6632\ : LocalMux
    port map (
            O => \N__32917\,
            I => \nx.n3105\
        );

    \I__6631\ : LocalMux
    port map (
            O => \N__32914\,
            I => \nx.n3105\
        );

    \I__6630\ : Odrv4
    port map (
            O => \N__32911\,
            I => \nx.n3105\
        );

    \I__6629\ : InMux
    port map (
            O => \N__32904\,
            I => \N__32901\
        );

    \I__6628\ : LocalMux
    port map (
            O => \N__32901\,
            I => \N__32898\
        );

    \I__6627\ : Odrv4
    port map (
            O => \N__32898\,
            I => \nx.n3172\
        );

    \I__6626\ : InMux
    port map (
            O => \N__32895\,
            I => \nx.n11083\
        );

    \I__6625\ : CascadeMux
    port map (
            O => \N__32892\,
            I => \N__32888\
        );

    \I__6624\ : InMux
    port map (
            O => \N__32891\,
            I => \N__32885\
        );

    \I__6623\ : InMux
    port map (
            O => \N__32888\,
            I => \N__32881\
        );

    \I__6622\ : LocalMux
    port map (
            O => \N__32885\,
            I => \N__32878\
        );

    \I__6621\ : InMux
    port map (
            O => \N__32884\,
            I => \N__32875\
        );

    \I__6620\ : LocalMux
    port map (
            O => \N__32881\,
            I => \N__32872\
        );

    \I__6619\ : Span4Mux_v
    port map (
            O => \N__32878\,
            I => \N__32869\
        );

    \I__6618\ : LocalMux
    port map (
            O => \N__32875\,
            I => \N__32866\
        );

    \I__6617\ : Span4Mux_h
    port map (
            O => \N__32872\,
            I => \N__32861\
        );

    \I__6616\ : Span4Mux_h
    port map (
            O => \N__32869\,
            I => \N__32861\
        );

    \I__6615\ : Odrv4
    port map (
            O => \N__32866\,
            I => \nx.n3104\
        );

    \I__6614\ : Odrv4
    port map (
            O => \N__32861\,
            I => \nx.n3104\
        );

    \I__6613\ : InMux
    port map (
            O => \N__32856\,
            I => \N__32853\
        );

    \I__6612\ : LocalMux
    port map (
            O => \N__32853\,
            I => \nx.n3171\
        );

    \I__6611\ : InMux
    port map (
            O => \N__32850\,
            I => \nx.n11084\
        );

    \I__6610\ : CascadeMux
    port map (
            O => \N__32847\,
            I => \N__32844\
        );

    \I__6609\ : InMux
    port map (
            O => \N__32844\,
            I => \N__32840\
        );

    \I__6608\ : InMux
    port map (
            O => \N__32843\,
            I => \N__32837\
        );

    \I__6607\ : LocalMux
    port map (
            O => \N__32840\,
            I => \N__32834\
        );

    \I__6606\ : LocalMux
    port map (
            O => \N__32837\,
            I => \N__32830\
        );

    \I__6605\ : Span4Mux_v
    port map (
            O => \N__32834\,
            I => \N__32827\
        );

    \I__6604\ : InMux
    port map (
            O => \N__32833\,
            I => \N__32824\
        );

    \I__6603\ : Span4Mux_h
    port map (
            O => \N__32830\,
            I => \N__32821\
        );

    \I__6602\ : Span4Mux_h
    port map (
            O => \N__32827\,
            I => \N__32818\
        );

    \I__6601\ : LocalMux
    port map (
            O => \N__32824\,
            I => \nx.n3103\
        );

    \I__6600\ : Odrv4
    port map (
            O => \N__32821\,
            I => \nx.n3103\
        );

    \I__6599\ : Odrv4
    port map (
            O => \N__32818\,
            I => \nx.n3103\
        );

    \I__6598\ : InMux
    port map (
            O => \N__32811\,
            I => \N__32808\
        );

    \I__6597\ : LocalMux
    port map (
            O => \N__32808\,
            I => \nx.n3170\
        );

    \I__6596\ : InMux
    port map (
            O => \N__32805\,
            I => \nx.n11085\
        );

    \I__6595\ : CascadeMux
    port map (
            O => \N__32802\,
            I => \N__32799\
        );

    \I__6594\ : InMux
    port map (
            O => \N__32799\,
            I => \N__32795\
        );

    \I__6593\ : InMux
    port map (
            O => \N__32798\,
            I => \N__32791\
        );

    \I__6592\ : LocalMux
    port map (
            O => \N__32795\,
            I => \N__32788\
        );

    \I__6591\ : InMux
    port map (
            O => \N__32794\,
            I => \N__32785\
        );

    \I__6590\ : LocalMux
    port map (
            O => \N__32791\,
            I => \nx.n3102\
        );

    \I__6589\ : Odrv4
    port map (
            O => \N__32788\,
            I => \nx.n3102\
        );

    \I__6588\ : LocalMux
    port map (
            O => \N__32785\,
            I => \nx.n3102\
        );

    \I__6587\ : InMux
    port map (
            O => \N__32778\,
            I => \N__32775\
        );

    \I__6586\ : LocalMux
    port map (
            O => \N__32775\,
            I => \nx.n3169\
        );

    \I__6585\ : InMux
    port map (
            O => \N__32772\,
            I => \bfn_13_18_0_\
        );

    \I__6584\ : CascadeMux
    port map (
            O => \N__32769\,
            I => \N__32764\
        );

    \I__6583\ : CascadeMux
    port map (
            O => \N__32768\,
            I => \N__32761\
        );

    \I__6582\ : CascadeMux
    port map (
            O => \N__32767\,
            I => \N__32758\
        );

    \I__6581\ : InMux
    port map (
            O => \N__32764\,
            I => \N__32755\
        );

    \I__6580\ : InMux
    port map (
            O => \N__32761\,
            I => \N__32752\
        );

    \I__6579\ : InMux
    port map (
            O => \N__32758\,
            I => \N__32749\
        );

    \I__6578\ : LocalMux
    port map (
            O => \N__32755\,
            I => \N__32746\
        );

    \I__6577\ : LocalMux
    port map (
            O => \N__32752\,
            I => \N__32743\
        );

    \I__6576\ : LocalMux
    port map (
            O => \N__32749\,
            I => \N__32740\
        );

    \I__6575\ : Span4Mux_h
    port map (
            O => \N__32746\,
            I => \N__32737\
        );

    \I__6574\ : Span4Mux_v
    port map (
            O => \N__32743\,
            I => \N__32732\
        );

    \I__6573\ : Span4Mux_h
    port map (
            O => \N__32740\,
            I => \N__32732\
        );

    \I__6572\ : Odrv4
    port map (
            O => \N__32737\,
            I => \nx.n3101\
        );

    \I__6571\ : Odrv4
    port map (
            O => \N__32732\,
            I => \nx.n3101\
        );

    \I__6570\ : InMux
    port map (
            O => \N__32727\,
            I => \N__32724\
        );

    \I__6569\ : LocalMux
    port map (
            O => \N__32724\,
            I => \nx.n3168\
        );

    \I__6568\ : InMux
    port map (
            O => \N__32721\,
            I => \nx.n11087\
        );

    \I__6567\ : InMux
    port map (
            O => \N__32718\,
            I => \N__32715\
        );

    \I__6566\ : LocalMux
    port map (
            O => \N__32715\,
            I => \N__32712\
        );

    \I__6565\ : Odrv4
    port map (
            O => \N__32712\,
            I => \nx.n2169\
        );

    \I__6564\ : CascadeMux
    port map (
            O => \N__32709\,
            I => \N__32704\
        );

    \I__6563\ : CascadeMux
    port map (
            O => \N__32708\,
            I => \N__32701\
        );

    \I__6562\ : CascadeMux
    port map (
            O => \N__32707\,
            I => \N__32698\
        );

    \I__6561\ : InMux
    port map (
            O => \N__32704\,
            I => \N__32695\
        );

    \I__6560\ : InMux
    port map (
            O => \N__32701\,
            I => \N__32692\
        );

    \I__6559\ : InMux
    port map (
            O => \N__32698\,
            I => \N__32689\
        );

    \I__6558\ : LocalMux
    port map (
            O => \N__32695\,
            I => \N__32684\
        );

    \I__6557\ : LocalMux
    port map (
            O => \N__32692\,
            I => \N__32684\
        );

    \I__6556\ : LocalMux
    port map (
            O => \N__32689\,
            I => \N__32681\
        );

    \I__6555\ : Span4Mux_v
    port map (
            O => \N__32684\,
            I => \N__32678\
        );

    \I__6554\ : Odrv12
    port map (
            O => \N__32681\,
            I => \nx.n2102\
        );

    \I__6553\ : Odrv4
    port map (
            O => \N__32678\,
            I => \nx.n2102\
        );

    \I__6552\ : CascadeMux
    port map (
            O => \N__32673\,
            I => \N__32670\
        );

    \I__6551\ : InMux
    port map (
            O => \N__32670\,
            I => \N__32666\
        );

    \I__6550\ : InMux
    port map (
            O => \N__32669\,
            I => \N__32662\
        );

    \I__6549\ : LocalMux
    port map (
            O => \N__32666\,
            I => \N__32659\
        );

    \I__6548\ : InMux
    port map (
            O => \N__32665\,
            I => \N__32656\
        );

    \I__6547\ : LocalMux
    port map (
            O => \N__32662\,
            I => \nx.n2201\
        );

    \I__6546\ : Odrv4
    port map (
            O => \N__32659\,
            I => \nx.n2201\
        );

    \I__6545\ : LocalMux
    port map (
            O => \N__32656\,
            I => \nx.n2201\
        );

    \I__6544\ : InMux
    port map (
            O => \N__32649\,
            I => \N__32646\
        );

    \I__6543\ : LocalMux
    port map (
            O => \N__32646\,
            I => \nx.n2261\
        );

    \I__6542\ : CascadeMux
    port map (
            O => \N__32643\,
            I => \N__32639\
        );

    \I__6541\ : InMux
    port map (
            O => \N__32642\,
            I => \N__32635\
        );

    \I__6540\ : InMux
    port map (
            O => \N__32639\,
            I => \N__32632\
        );

    \I__6539\ : InMux
    port map (
            O => \N__32638\,
            I => \N__32629\
        );

    \I__6538\ : LocalMux
    port map (
            O => \N__32635\,
            I => \nx.n2194\
        );

    \I__6537\ : LocalMux
    port map (
            O => \N__32632\,
            I => \nx.n2194\
        );

    \I__6536\ : LocalMux
    port map (
            O => \N__32629\,
            I => \nx.n2194\
        );

    \I__6535\ : InMux
    port map (
            O => \N__32622\,
            I => \N__32619\
        );

    \I__6534\ : LocalMux
    port map (
            O => \N__32619\,
            I => \N__32616\
        );

    \I__6533\ : Odrv4
    port map (
            O => \N__32616\,
            I => \nx.n2262\
        );

    \I__6532\ : CascadeMux
    port map (
            O => \N__32613\,
            I => \N__32610\
        );

    \I__6531\ : InMux
    port map (
            O => \N__32610\,
            I => \N__32606\
        );

    \I__6530\ : CascadeMux
    port map (
            O => \N__32609\,
            I => \N__32603\
        );

    \I__6529\ : LocalMux
    port map (
            O => \N__32606\,
            I => \N__32600\
        );

    \I__6528\ : InMux
    port map (
            O => \N__32603\,
            I => \N__32597\
        );

    \I__6527\ : Span4Mux_v
    port map (
            O => \N__32600\,
            I => \N__32593\
        );

    \I__6526\ : LocalMux
    port map (
            O => \N__32597\,
            I => \N__32590\
        );

    \I__6525\ : InMux
    port map (
            O => \N__32596\,
            I => \N__32587\
        );

    \I__6524\ : Odrv4
    port map (
            O => \N__32593\,
            I => \nx.n2195\
        );

    \I__6523\ : Odrv4
    port map (
            O => \N__32590\,
            I => \nx.n2195\
        );

    \I__6522\ : LocalMux
    port map (
            O => \N__32587\,
            I => \nx.n2195\
        );

    \I__6521\ : CascadeMux
    port map (
            O => \N__32580\,
            I => \N__32573\
        );

    \I__6520\ : InMux
    port map (
            O => \N__32579\,
            I => \N__32566\
        );

    \I__6519\ : CascadeMux
    port map (
            O => \N__32578\,
            I => \N__32563\
        );

    \I__6518\ : CascadeMux
    port map (
            O => \N__32577\,
            I => \N__32555\
        );

    \I__6517\ : CascadeMux
    port map (
            O => \N__32576\,
            I => \N__32549\
        );

    \I__6516\ : InMux
    port map (
            O => \N__32573\,
            I => \N__32542\
        );

    \I__6515\ : InMux
    port map (
            O => \N__32572\,
            I => \N__32542\
        );

    \I__6514\ : InMux
    port map (
            O => \N__32571\,
            I => \N__32542\
        );

    \I__6513\ : CascadeMux
    port map (
            O => \N__32570\,
            I => \N__32539\
        );

    \I__6512\ : CascadeMux
    port map (
            O => \N__32569\,
            I => \N__32535\
        );

    \I__6511\ : LocalMux
    port map (
            O => \N__32566\,
            I => \N__32532\
        );

    \I__6510\ : InMux
    port map (
            O => \N__32563\,
            I => \N__32525\
        );

    \I__6509\ : InMux
    port map (
            O => \N__32562\,
            I => \N__32525\
        );

    \I__6508\ : InMux
    port map (
            O => \N__32561\,
            I => \N__32525\
        );

    \I__6507\ : InMux
    port map (
            O => \N__32560\,
            I => \N__32518\
        );

    \I__6506\ : InMux
    port map (
            O => \N__32559\,
            I => \N__32518\
        );

    \I__6505\ : InMux
    port map (
            O => \N__32558\,
            I => \N__32518\
        );

    \I__6504\ : InMux
    port map (
            O => \N__32555\,
            I => \N__32511\
        );

    \I__6503\ : InMux
    port map (
            O => \N__32554\,
            I => \N__32511\
        );

    \I__6502\ : InMux
    port map (
            O => \N__32553\,
            I => \N__32511\
        );

    \I__6501\ : InMux
    port map (
            O => \N__32552\,
            I => \N__32506\
        );

    \I__6500\ : InMux
    port map (
            O => \N__32549\,
            I => \N__32506\
        );

    \I__6499\ : LocalMux
    port map (
            O => \N__32542\,
            I => \N__32503\
        );

    \I__6498\ : InMux
    port map (
            O => \N__32539\,
            I => \N__32496\
        );

    \I__6497\ : InMux
    port map (
            O => \N__32538\,
            I => \N__32496\
        );

    \I__6496\ : InMux
    port map (
            O => \N__32535\,
            I => \N__32496\
        );

    \I__6495\ : Span4Mux_h
    port map (
            O => \N__32532\,
            I => \N__32493\
        );

    \I__6494\ : LocalMux
    port map (
            O => \N__32525\,
            I => \N__32490\
        );

    \I__6493\ : LocalMux
    port map (
            O => \N__32518\,
            I => \nx.n2225\
        );

    \I__6492\ : LocalMux
    port map (
            O => \N__32511\,
            I => \nx.n2225\
        );

    \I__6491\ : LocalMux
    port map (
            O => \N__32506\,
            I => \nx.n2225\
        );

    \I__6490\ : Odrv4
    port map (
            O => \N__32503\,
            I => \nx.n2225\
        );

    \I__6489\ : LocalMux
    port map (
            O => \N__32496\,
            I => \nx.n2225\
        );

    \I__6488\ : Odrv4
    port map (
            O => \N__32493\,
            I => \nx.n2225\
        );

    \I__6487\ : Odrv12
    port map (
            O => \N__32490\,
            I => \nx.n2225\
        );

    \I__6486\ : IoInMux
    port map (
            O => \N__32475\,
            I => \N__32472\
        );

    \I__6485\ : LocalMux
    port map (
            O => \N__32472\,
            I => \N__32469\
        );

    \I__6484\ : IoSpan4Mux
    port map (
            O => \N__32469\,
            I => \N__32466\
        );

    \I__6483\ : Sp12to4
    port map (
            O => \N__32466\,
            I => \N__32463\
        );

    \I__6482\ : Span12Mux_h
    port map (
            O => \N__32463\,
            I => \N__32459\
        );

    \I__6481\ : InMux
    port map (
            O => \N__32462\,
            I => \N__32456\
        );

    \I__6480\ : Odrv12
    port map (
            O => \N__32459\,
            I => pin_oe_4
        );

    \I__6479\ : LocalMux
    port map (
            O => \N__32456\,
            I => pin_oe_4
        );

    \I__6478\ : CascadeMux
    port map (
            O => \N__32451\,
            I => \n11970_cascade_\
        );

    \I__6477\ : IoInMux
    port map (
            O => \N__32448\,
            I => \N__32445\
        );

    \I__6476\ : LocalMux
    port map (
            O => \N__32445\,
            I => \N__32442\
        );

    \I__6475\ : Span12Mux_s4_v
    port map (
            O => \N__32442\,
            I => \N__32439\
        );

    \I__6474\ : Span12Mux_h
    port map (
            O => \N__32439\,
            I => \N__32436\
        );

    \I__6473\ : Span12Mux_v
    port map (
            O => \N__32436\,
            I => \N__32432\
        );

    \I__6472\ : InMux
    port map (
            O => \N__32435\,
            I => \N__32429\
        );

    \I__6471\ : Odrv12
    port map (
            O => \N__32432\,
            I => pin_oe_0
        );

    \I__6470\ : LocalMux
    port map (
            O => \N__32429\,
            I => pin_oe_0
        );

    \I__6469\ : InMux
    port map (
            O => \N__32424\,
            I => \N__32421\
        );

    \I__6468\ : LocalMux
    port map (
            O => \N__32421\,
            I => \N__32418\
        );

    \I__6467\ : Span4Mux_h
    port map (
            O => \N__32418\,
            I => \N__32415\
        );

    \I__6466\ : Odrv4
    port map (
            O => \N__32415\,
            I => n11968
        );

    \I__6465\ : InMux
    port map (
            O => \N__32412\,
            I => \N__32408\
        );

    \I__6464\ : InMux
    port map (
            O => \N__32411\,
            I => \N__32405\
        );

    \I__6463\ : LocalMux
    port map (
            O => \N__32408\,
            I => \N__32400\
        );

    \I__6462\ : LocalMux
    port map (
            O => \N__32405\,
            I => \N__32400\
        );

    \I__6461\ : Span4Mux_h
    port map (
            O => \N__32400\,
            I => \N__32396\
        );

    \I__6460\ : InMux
    port map (
            O => \N__32399\,
            I => \N__32393\
        );

    \I__6459\ : Sp12to4
    port map (
            O => \N__32396\,
            I => \N__32386\
        );

    \I__6458\ : LocalMux
    port map (
            O => \N__32393\,
            I => \N__32386\
        );

    \I__6457\ : InMux
    port map (
            O => \N__32392\,
            I => \N__32383\
        );

    \I__6456\ : InMux
    port map (
            O => \N__32391\,
            I => \N__32380\
        );

    \I__6455\ : Span12Mux_v
    port map (
            O => \N__32386\,
            I => \N__32377\
        );

    \I__6454\ : LocalMux
    port map (
            O => \N__32383\,
            I => \nx.bit_ctr_4\
        );

    \I__6453\ : LocalMux
    port map (
            O => \N__32380\,
            I => \nx.bit_ctr_4\
        );

    \I__6452\ : Odrv12
    port map (
            O => \N__32377\,
            I => \nx.bit_ctr_4\
        );

    \I__6451\ : InMux
    port map (
            O => \N__32370\,
            I => \N__32367\
        );

    \I__6450\ : LocalMux
    port map (
            O => \N__32367\,
            I => \N__32364\
        );

    \I__6449\ : Odrv4
    port map (
            O => \N__32364\,
            I => \nx.n3177\
        );

    \I__6448\ : InMux
    port map (
            O => \N__32361\,
            I => \bfn_13_17_0_\
        );

    \I__6447\ : CascadeMux
    port map (
            O => \N__32358\,
            I => \N__32355\
        );

    \I__6446\ : InMux
    port map (
            O => \N__32355\,
            I => \N__32350\
        );

    \I__6445\ : CascadeMux
    port map (
            O => \N__32354\,
            I => \N__32347\
        );

    \I__6444\ : CascadeMux
    port map (
            O => \N__32353\,
            I => \N__32344\
        );

    \I__6443\ : LocalMux
    port map (
            O => \N__32350\,
            I => \N__32341\
        );

    \I__6442\ : InMux
    port map (
            O => \N__32347\,
            I => \N__32338\
        );

    \I__6441\ : InMux
    port map (
            O => \N__32344\,
            I => \N__32335\
        );

    \I__6440\ : Span4Mux_v
    port map (
            O => \N__32341\,
            I => \N__32332\
        );

    \I__6439\ : LocalMux
    port map (
            O => \N__32338\,
            I => \nx.n3109\
        );

    \I__6438\ : LocalMux
    port map (
            O => \N__32335\,
            I => \nx.n3109\
        );

    \I__6437\ : Odrv4
    port map (
            O => \N__32332\,
            I => \nx.n3109\
        );

    \I__6436\ : InMux
    port map (
            O => \N__32325\,
            I => \N__32322\
        );

    \I__6435\ : LocalMux
    port map (
            O => \N__32322\,
            I => \nx.n3176\
        );

    \I__6434\ : InMux
    port map (
            O => \N__32319\,
            I => \nx.n11079\
        );

    \I__6433\ : CascadeMux
    port map (
            O => \N__32316\,
            I => \nx.n2299_cascade_\
        );

    \I__6432\ : CascadeMux
    port map (
            O => \N__32313\,
            I => \N__32310\
        );

    \I__6431\ : InMux
    port map (
            O => \N__32310\,
            I => \N__32307\
        );

    \I__6430\ : LocalMux
    port map (
            O => \N__32307\,
            I => \nx.n2265\
        );

    \I__6429\ : CascadeMux
    port map (
            O => \N__32304\,
            I => \N__32301\
        );

    \I__6428\ : InMux
    port map (
            O => \N__32301\,
            I => \N__32298\
        );

    \I__6427\ : LocalMux
    port map (
            O => \N__32298\,
            I => \N__32294\
        );

    \I__6426\ : CascadeMux
    port map (
            O => \N__32297\,
            I => \N__32291\
        );

    \I__6425\ : Span4Mux_h
    port map (
            O => \N__32294\,
            I => \N__32287\
        );

    \I__6424\ : InMux
    port map (
            O => \N__32291\,
            I => \N__32284\
        );

    \I__6423\ : InMux
    port map (
            O => \N__32290\,
            I => \N__32281\
        );

    \I__6422\ : Odrv4
    port map (
            O => \N__32287\,
            I => \nx.n2197\
        );

    \I__6421\ : LocalMux
    port map (
            O => \N__32284\,
            I => \nx.n2197\
        );

    \I__6420\ : LocalMux
    port map (
            O => \N__32281\,
            I => \nx.n2197\
        );

    \I__6419\ : CascadeMux
    port map (
            O => \N__32274\,
            I => \N__32271\
        );

    \I__6418\ : InMux
    port map (
            O => \N__32271\,
            I => \N__32267\
        );

    \I__6417\ : InMux
    port map (
            O => \N__32270\,
            I => \N__32264\
        );

    \I__6416\ : LocalMux
    port map (
            O => \N__32267\,
            I => \nx.n2196\
        );

    \I__6415\ : LocalMux
    port map (
            O => \N__32264\,
            I => \nx.n2196\
        );

    \I__6414\ : InMux
    port map (
            O => \N__32259\,
            I => \N__32256\
        );

    \I__6413\ : LocalMux
    port map (
            O => \N__32256\,
            I => \nx.n30_adj_694\
        );

    \I__6412\ : InMux
    port map (
            O => \N__32253\,
            I => \N__32250\
        );

    \I__6411\ : LocalMux
    port map (
            O => \N__32250\,
            I => \N__32247\
        );

    \I__6410\ : Span4Mux_h
    port map (
            O => \N__32247\,
            I => \N__32244\
        );

    \I__6409\ : Odrv4
    port map (
            O => \N__32244\,
            I => \nx.n22_adj_693\
        );

    \I__6408\ : CascadeMux
    port map (
            O => \N__32241\,
            I => \nx.n21_cascade_\
        );

    \I__6407\ : InMux
    port map (
            O => \N__32238\,
            I => \N__32235\
        );

    \I__6406\ : LocalMux
    port map (
            O => \N__32235\,
            I => \nx.n34_adj_695\
        );

    \I__6405\ : InMux
    port map (
            O => \N__32232\,
            I => \N__32229\
        );

    \I__6404\ : LocalMux
    port map (
            O => \N__32229\,
            I => \nx.n2268\
        );

    \I__6403\ : CascadeMux
    port map (
            O => \N__32226\,
            I => \nx.n2225_cascade_\
        );

    \I__6402\ : InMux
    port map (
            O => \N__32223\,
            I => \N__32215\
        );

    \I__6401\ : InMux
    port map (
            O => \N__32222\,
            I => \N__32215\
        );

    \I__6400\ : InMux
    port map (
            O => \N__32221\,
            I => \N__32212\
        );

    \I__6399\ : InMux
    port map (
            O => \N__32220\,
            I => \N__32209\
        );

    \I__6398\ : LocalMux
    port map (
            O => \N__32215\,
            I => \N__32204\
        );

    \I__6397\ : LocalMux
    port map (
            O => \N__32212\,
            I => \N__32204\
        );

    \I__6396\ : LocalMux
    port map (
            O => \N__32209\,
            I => \N__32200\
        );

    \I__6395\ : Sp12to4
    port map (
            O => \N__32204\,
            I => \N__32197\
        );

    \I__6394\ : InMux
    port map (
            O => \N__32203\,
            I => \N__32194\
        );

    \I__6393\ : Span12Mux_s11_h
    port map (
            O => \N__32200\,
            I => \N__32191\
        );

    \I__6392\ : Span12Mux_v
    port map (
            O => \N__32197\,
            I => \N__32188\
        );

    \I__6391\ : LocalMux
    port map (
            O => \N__32194\,
            I => neopxl_color_4
        );

    \I__6390\ : Odrv12
    port map (
            O => \N__32191\,
            I => neopxl_color_4
        );

    \I__6389\ : Odrv12
    port map (
            O => \N__32188\,
            I => neopxl_color_4
        );

    \I__6388\ : SRMux
    port map (
            O => \N__32181\,
            I => \N__32178\
        );

    \I__6387\ : LocalMux
    port map (
            O => \N__32178\,
            I => \N__32175\
        );

    \I__6386\ : Span4Mux_h
    port map (
            O => \N__32175\,
            I => \N__32172\
        );

    \I__6385\ : Span4Mux_v
    port map (
            O => \N__32172\,
            I => \N__32169\
        );

    \I__6384\ : Odrv4
    port map (
            O => \N__32169\,
            I => n22_adj_787
        );

    \I__6383\ : CascadeMux
    port map (
            O => \N__32166\,
            I => \N__32163\
        );

    \I__6382\ : InMux
    port map (
            O => \N__32163\,
            I => \N__32159\
        );

    \I__6381\ : InMux
    port map (
            O => \N__32162\,
            I => \N__32156\
        );

    \I__6380\ : LocalMux
    port map (
            O => \N__32159\,
            I => \N__32153\
        );

    \I__6379\ : LocalMux
    port map (
            O => \N__32156\,
            I => \N__32150\
        );

    \I__6378\ : Span4Mux_h
    port map (
            O => \N__32153\,
            I => \N__32147\
        );

    \I__6377\ : Odrv12
    port map (
            O => \N__32150\,
            I => \nx.n2099\
        );

    \I__6376\ : Odrv4
    port map (
            O => \N__32147\,
            I => \nx.n2099\
        );

    \I__6375\ : InMux
    port map (
            O => \N__32142\,
            I => \N__32139\
        );

    \I__6374\ : LocalMux
    port map (
            O => \N__32139\,
            I => \N__32136\
        );

    \I__6373\ : Odrv4
    port map (
            O => \N__32136\,
            I => \nx.n2166\
        );

    \I__6372\ : InMux
    port map (
            O => \N__32133\,
            I => \N__32129\
        );

    \I__6371\ : InMux
    port map (
            O => \N__32132\,
            I => \N__32125\
        );

    \I__6370\ : LocalMux
    port map (
            O => \N__32129\,
            I => \N__32122\
        );

    \I__6369\ : InMux
    port map (
            O => \N__32128\,
            I => \N__32119\
        );

    \I__6368\ : LocalMux
    port map (
            O => \N__32125\,
            I => \nx.n2198\
        );

    \I__6367\ : Odrv4
    port map (
            O => \N__32122\,
            I => \nx.n2198\
        );

    \I__6366\ : LocalMux
    port map (
            O => \N__32119\,
            I => \nx.n2198\
        );

    \I__6365\ : InMux
    port map (
            O => \N__32112\,
            I => \N__32109\
        );

    \I__6364\ : LocalMux
    port map (
            O => \N__32109\,
            I => \nx.n2274\
        );

    \I__6363\ : CascadeMux
    port map (
            O => \N__32106\,
            I => \N__32102\
        );

    \I__6362\ : InMux
    port map (
            O => \N__32105\,
            I => \N__32099\
        );

    \I__6361\ : InMux
    port map (
            O => \N__32102\,
            I => \N__32096\
        );

    \I__6360\ : LocalMux
    port map (
            O => \N__32099\,
            I => \N__32093\
        );

    \I__6359\ : LocalMux
    port map (
            O => \N__32096\,
            I => \N__32089\
        );

    \I__6358\ : Span4Mux_v
    port map (
            O => \N__32093\,
            I => \N__32086\
        );

    \I__6357\ : InMux
    port map (
            O => \N__32092\,
            I => \N__32083\
        );

    \I__6356\ : Span4Mux_h
    port map (
            O => \N__32089\,
            I => \N__32080\
        );

    \I__6355\ : Odrv4
    port map (
            O => \N__32086\,
            I => \nx.n2207\
        );

    \I__6354\ : LocalMux
    port map (
            O => \N__32083\,
            I => \nx.n2207\
        );

    \I__6353\ : Odrv4
    port map (
            O => \N__32080\,
            I => \nx.n2207\
        );

    \I__6352\ : InMux
    port map (
            O => \N__32073\,
            I => \N__32069\
        );

    \I__6351\ : CascadeMux
    port map (
            O => \N__32072\,
            I => \N__32066\
        );

    \I__6350\ : LocalMux
    port map (
            O => \N__32069\,
            I => \N__32063\
        );

    \I__6349\ : InMux
    port map (
            O => \N__32066\,
            I => \N__32059\
        );

    \I__6348\ : Span4Mux_h
    port map (
            O => \N__32063\,
            I => \N__32056\
        );

    \I__6347\ : InMux
    port map (
            O => \N__32062\,
            I => \N__32053\
        );

    \I__6346\ : LocalMux
    port map (
            O => \N__32059\,
            I => \N__32050\
        );

    \I__6345\ : Odrv4
    port map (
            O => \N__32056\,
            I => \nx.n2208\
        );

    \I__6344\ : LocalMux
    port map (
            O => \N__32053\,
            I => \nx.n2208\
        );

    \I__6343\ : Odrv4
    port map (
            O => \N__32050\,
            I => \nx.n2208\
        );

    \I__6342\ : CascadeMux
    port map (
            O => \N__32043\,
            I => \N__32040\
        );

    \I__6341\ : InMux
    port map (
            O => \N__32040\,
            I => \N__32037\
        );

    \I__6340\ : LocalMux
    port map (
            O => \N__32037\,
            I => \N__32034\
        );

    \I__6339\ : Odrv4
    port map (
            O => \N__32034\,
            I => \nx.n2275\
        );

    \I__6338\ : InMux
    port map (
            O => \N__32031\,
            I => \N__32028\
        );

    \I__6337\ : LocalMux
    port map (
            O => \N__32028\,
            I => \nx.n2272\
        );

    \I__6336\ : CascadeMux
    port map (
            O => \N__32025\,
            I => \N__32021\
        );

    \I__6335\ : InMux
    port map (
            O => \N__32024\,
            I => \N__32018\
        );

    \I__6334\ : InMux
    port map (
            O => \N__32021\,
            I => \N__32015\
        );

    \I__6333\ : LocalMux
    port map (
            O => \N__32018\,
            I => \N__32012\
        );

    \I__6332\ : LocalMux
    port map (
            O => \N__32015\,
            I => \N__32008\
        );

    \I__6331\ : Span4Mux_h
    port map (
            O => \N__32012\,
            I => \N__32005\
        );

    \I__6330\ : InMux
    port map (
            O => \N__32011\,
            I => \N__32002\
        );

    \I__6329\ : Span4Mux_v
    port map (
            O => \N__32008\,
            I => \N__31999\
        );

    \I__6328\ : Odrv4
    port map (
            O => \N__32005\,
            I => \nx.n2205\
        );

    \I__6327\ : LocalMux
    port map (
            O => \N__32002\,
            I => \nx.n2205\
        );

    \I__6326\ : Odrv4
    port map (
            O => \N__31999\,
            I => \nx.n2205\
        );

    \I__6325\ : CascadeMux
    port map (
            O => \N__31992\,
            I => \nx.n2391_cascade_\
        );

    \I__6324\ : CascadeMux
    port map (
            O => \N__31989\,
            I => \nx.n30_adj_696_cascade_\
        );

    \I__6323\ : InMux
    port map (
            O => \N__31986\,
            I => \N__31983\
        );

    \I__6322\ : LocalMux
    port map (
            O => \N__31983\,
            I => \nx.n2266\
        );

    \I__6321\ : CascadeMux
    port map (
            O => \N__31980\,
            I => \N__31976\
        );

    \I__6320\ : InMux
    port map (
            O => \N__31979\,
            I => \N__31973\
        );

    \I__6319\ : InMux
    port map (
            O => \N__31976\,
            I => \N__31970\
        );

    \I__6318\ : LocalMux
    port map (
            O => \N__31973\,
            I => \N__31967\
        );

    \I__6317\ : LocalMux
    port map (
            O => \N__31970\,
            I => \nx.n2199\
        );

    \I__6316\ : Odrv4
    port map (
            O => \N__31967\,
            I => \nx.n2199\
        );

    \I__6315\ : InMux
    port map (
            O => \N__31962\,
            I => \N__31959\
        );

    \I__6314\ : LocalMux
    port map (
            O => \N__31959\,
            I => \nx.n2267\
        );

    \I__6313\ : InMux
    port map (
            O => \N__31956\,
            I => \N__31952\
        );

    \I__6312\ : CascadeMux
    port map (
            O => \N__31955\,
            I => \N__31948\
        );

    \I__6311\ : LocalMux
    port map (
            O => \N__31952\,
            I => \N__31945\
        );

    \I__6310\ : CascadeMux
    port map (
            O => \N__31951\,
            I => \N__31942\
        );

    \I__6309\ : InMux
    port map (
            O => \N__31948\,
            I => \N__31939\
        );

    \I__6308\ : Span4Mux_h
    port map (
            O => \N__31945\,
            I => \N__31936\
        );

    \I__6307\ : InMux
    port map (
            O => \N__31942\,
            I => \N__31933\
        );

    \I__6306\ : LocalMux
    port map (
            O => \N__31939\,
            I => \N__31930\
        );

    \I__6305\ : Odrv4
    port map (
            O => \N__31936\,
            I => \nx.n2204\
        );

    \I__6304\ : LocalMux
    port map (
            O => \N__31933\,
            I => \nx.n2204\
        );

    \I__6303\ : Odrv4
    port map (
            O => \N__31930\,
            I => \nx.n2204\
        );

    \I__6302\ : CascadeMux
    port map (
            O => \N__31923\,
            I => \N__31920\
        );

    \I__6301\ : InMux
    port map (
            O => \N__31920\,
            I => \N__31917\
        );

    \I__6300\ : LocalMux
    port map (
            O => \N__31917\,
            I => \nx.n2271\
        );

    \I__6299\ : CascadeMux
    port map (
            O => \N__31914\,
            I => \nx.n2303_cascade_\
        );

    \I__6298\ : InMux
    port map (
            O => \N__31911\,
            I => \N__31908\
        );

    \I__6297\ : LocalMux
    port map (
            O => \N__31908\,
            I => \nx.n2269\
        );

    \I__6296\ : InMux
    port map (
            O => \N__31905\,
            I => \N__31901\
        );

    \I__6295\ : CascadeMux
    port map (
            O => \N__31904\,
            I => \N__31898\
        );

    \I__6294\ : LocalMux
    port map (
            O => \N__31901\,
            I => \N__31895\
        );

    \I__6293\ : InMux
    port map (
            O => \N__31898\,
            I => \N__31892\
        );

    \I__6292\ : Span4Mux_h
    port map (
            O => \N__31895\,
            I => \N__31887\
        );

    \I__6291\ : LocalMux
    port map (
            O => \N__31892\,
            I => \N__31887\
        );

    \I__6290\ : Odrv4
    port map (
            O => \N__31887\,
            I => \nx.n2202\
        );

    \I__6289\ : InMux
    port map (
            O => \N__31884\,
            I => \N__31880\
        );

    \I__6288\ : CascadeMux
    port map (
            O => \N__31883\,
            I => \N__31877\
        );

    \I__6287\ : LocalMux
    port map (
            O => \N__31880\,
            I => \N__31874\
        );

    \I__6286\ : InMux
    port map (
            O => \N__31877\,
            I => \N__31870\
        );

    \I__6285\ : Span4Mux_v
    port map (
            O => \N__31874\,
            I => \N__31867\
        );

    \I__6284\ : InMux
    port map (
            O => \N__31873\,
            I => \N__31864\
        );

    \I__6283\ : LocalMux
    port map (
            O => \N__31870\,
            I => \N__31861\
        );

    \I__6282\ : Odrv4
    port map (
            O => \N__31867\,
            I => \nx.n2203\
        );

    \I__6281\ : LocalMux
    port map (
            O => \N__31864\,
            I => \nx.n2203\
        );

    \I__6280\ : Odrv12
    port map (
            O => \N__31861\,
            I => \nx.n2203\
        );

    \I__6279\ : CascadeMux
    port map (
            O => \N__31854\,
            I => \N__31851\
        );

    \I__6278\ : InMux
    port map (
            O => \N__31851\,
            I => \N__31848\
        );

    \I__6277\ : LocalMux
    port map (
            O => \N__31848\,
            I => \nx.n2270\
        );

    \I__6276\ : CascadeMux
    port map (
            O => \N__31845\,
            I => \nx.n2302_cascade_\
        );

    \I__6275\ : CascadeMux
    port map (
            O => \N__31842\,
            I => \nx.n2401_cascade_\
        );

    \I__6274\ : InMux
    port map (
            O => \N__31839\,
            I => \N__31836\
        );

    \I__6273\ : LocalMux
    port map (
            O => \N__31836\,
            I => \N__31833\
        );

    \I__6272\ : Odrv4
    port map (
            O => \N__31833\,
            I => \nx.n38\
        );

    \I__6271\ : InMux
    port map (
            O => \N__31830\,
            I => \N__31827\
        );

    \I__6270\ : LocalMux
    port map (
            O => \N__31827\,
            I => \nx.n37\
        );

    \I__6269\ : CascadeMux
    port map (
            O => \N__31824\,
            I => \nx.n39_cascade_\
        );

    \I__6268\ : CascadeMux
    port map (
            O => \N__31821\,
            I => \nx.n2621_cascade_\
        );

    \I__6267\ : CascadeMux
    port map (
            O => \N__31818\,
            I => \N__31815\
        );

    \I__6266\ : InMux
    port map (
            O => \N__31815\,
            I => \N__31810\
        );

    \I__6265\ : InMux
    port map (
            O => \N__31814\,
            I => \N__31807\
        );

    \I__6264\ : InMux
    port map (
            O => \N__31813\,
            I => \N__31804\
        );

    \I__6263\ : LocalMux
    port map (
            O => \N__31810\,
            I => \N__31801\
        );

    \I__6262\ : LocalMux
    port map (
            O => \N__31807\,
            I => \nx.n2707\
        );

    \I__6261\ : LocalMux
    port map (
            O => \N__31804\,
            I => \nx.n2707\
        );

    \I__6260\ : Odrv4
    port map (
            O => \N__31801\,
            I => \nx.n2707\
        );

    \I__6259\ : InMux
    port map (
            O => \N__31794\,
            I => \N__31791\
        );

    \I__6258\ : LocalMux
    port map (
            O => \N__31791\,
            I => \N__31786\
        );

    \I__6257\ : InMux
    port map (
            O => \N__31790\,
            I => \N__31783\
        );

    \I__6256\ : InMux
    port map (
            O => \N__31789\,
            I => \N__31780\
        );

    \I__6255\ : Span4Mux_v
    port map (
            O => \N__31786\,
            I => \N__31775\
        );

    \I__6254\ : LocalMux
    port map (
            O => \N__31783\,
            I => \N__31772\
        );

    \I__6253\ : LocalMux
    port map (
            O => \N__31780\,
            I => \N__31769\
        );

    \I__6252\ : InMux
    port map (
            O => \N__31779\,
            I => \N__31766\
        );

    \I__6251\ : InMux
    port map (
            O => \N__31778\,
            I => \N__31763\
        );

    \I__6250\ : Span4Mux_h
    port map (
            O => \N__31775\,
            I => \N__31760\
        );

    \I__6249\ : Span4Mux_h
    port map (
            O => \N__31772\,
            I => \N__31755\
        );

    \I__6248\ : Span4Mux_v
    port map (
            O => \N__31769\,
            I => \N__31755\
        );

    \I__6247\ : LocalMux
    port map (
            O => \N__31766\,
            I => \nx.bit_ctr_13\
        );

    \I__6246\ : LocalMux
    port map (
            O => \N__31763\,
            I => \nx.bit_ctr_13\
        );

    \I__6245\ : Odrv4
    port map (
            O => \N__31760\,
            I => \nx.bit_ctr_13\
        );

    \I__6244\ : Odrv4
    port map (
            O => \N__31755\,
            I => \nx.bit_ctr_13\
        );

    \I__6243\ : InMux
    port map (
            O => \N__31746\,
            I => \N__31743\
        );

    \I__6242\ : LocalMux
    port map (
            O => \N__31743\,
            I => \nx.n2277\
        );

    \I__6241\ : CascadeMux
    port map (
            O => \N__31740\,
            I => \nx.n2309_cascade_\
        );

    \I__6240\ : CascadeMux
    port map (
            O => \N__31737\,
            I => \nx.n9697_cascade_\
        );

    \I__6239\ : InMux
    port map (
            O => \N__31734\,
            I => \N__31731\
        );

    \I__6238\ : LocalMux
    port map (
            O => \N__31731\,
            I => \nx.n2273\
        );

    \I__6237\ : InMux
    port map (
            O => \N__31728\,
            I => \N__31725\
        );

    \I__6236\ : LocalMux
    port map (
            O => \N__31725\,
            I => \N__31720\
        );

    \I__6235\ : InMux
    port map (
            O => \N__31724\,
            I => \N__31717\
        );

    \I__6234\ : InMux
    port map (
            O => \N__31723\,
            I => \N__31714\
        );

    \I__6233\ : Span4Mux_h
    port map (
            O => \N__31720\,
            I => \N__31709\
        );

    \I__6232\ : LocalMux
    port map (
            O => \N__31717\,
            I => \N__31709\
        );

    \I__6231\ : LocalMux
    port map (
            O => \N__31714\,
            I => \nx.n2206\
        );

    \I__6230\ : Odrv4
    port map (
            O => \N__31709\,
            I => \nx.n2206\
        );

    \I__6229\ : InMux
    port map (
            O => \N__31704\,
            I => \N__31700\
        );

    \I__6228\ : CascadeMux
    port map (
            O => \N__31703\,
            I => \N__31697\
        );

    \I__6227\ : LocalMux
    port map (
            O => \N__31700\,
            I => \N__31693\
        );

    \I__6226\ : InMux
    port map (
            O => \N__31697\,
            I => \N__31690\
        );

    \I__6225\ : InMux
    port map (
            O => \N__31696\,
            I => \N__31687\
        );

    \I__6224\ : Span4Mux_h
    port map (
            O => \N__31693\,
            I => \N__31682\
        );

    \I__6223\ : LocalMux
    port map (
            O => \N__31690\,
            I => \N__31682\
        );

    \I__6222\ : LocalMux
    port map (
            O => \N__31687\,
            I => \nx.n2209\
        );

    \I__6221\ : Odrv4
    port map (
            O => \N__31682\,
            I => \nx.n2209\
        );

    \I__6220\ : CascadeMux
    port map (
            O => \N__31677\,
            I => \N__31674\
        );

    \I__6219\ : InMux
    port map (
            O => \N__31674\,
            I => \N__31671\
        );

    \I__6218\ : LocalMux
    port map (
            O => \N__31671\,
            I => \nx.n2276\
        );

    \I__6217\ : CascadeMux
    port map (
            O => \N__31668\,
            I => \N__31664\
        );

    \I__6216\ : InMux
    port map (
            O => \N__31667\,
            I => \N__31661\
        );

    \I__6215\ : InMux
    port map (
            O => \N__31664\,
            I => \N__31658\
        );

    \I__6214\ : LocalMux
    port map (
            O => \N__31661\,
            I => \N__31654\
        );

    \I__6213\ : LocalMux
    port map (
            O => \N__31658\,
            I => \N__31651\
        );

    \I__6212\ : InMux
    port map (
            O => \N__31657\,
            I => \N__31648\
        );

    \I__6211\ : Odrv4
    port map (
            O => \N__31654\,
            I => \nx.n2695\
        );

    \I__6210\ : Odrv4
    port map (
            O => \N__31651\,
            I => \nx.n2695\
        );

    \I__6209\ : LocalMux
    port map (
            O => \N__31648\,
            I => \nx.n2695\
        );

    \I__6208\ : CascadeMux
    port map (
            O => \N__31641\,
            I => \nx.n2597_cascade_\
        );

    \I__6207\ : CascadeMux
    port map (
            O => \N__31638\,
            I => \N__31634\
        );

    \I__6206\ : InMux
    port map (
            O => \N__31637\,
            I => \N__31631\
        );

    \I__6205\ : InMux
    port map (
            O => \N__31634\,
            I => \N__31628\
        );

    \I__6204\ : LocalMux
    port map (
            O => \N__31631\,
            I => \N__31625\
        );

    \I__6203\ : LocalMux
    port map (
            O => \N__31628\,
            I => \N__31622\
        );

    \I__6202\ : Span4Mux_v
    port map (
            O => \N__31625\,
            I => \N__31619\
        );

    \I__6201\ : Span4Mux_h
    port map (
            O => \N__31622\,
            I => \N__31616\
        );

    \I__6200\ : Odrv4
    port map (
            O => \N__31619\,
            I => \nx.n2691\
        );

    \I__6199\ : Odrv4
    port map (
            O => \N__31616\,
            I => \nx.n2691\
        );

    \I__6198\ : CascadeMux
    port map (
            O => \N__31611\,
            I => \N__31608\
        );

    \I__6197\ : InMux
    port map (
            O => \N__31608\,
            I => \N__31604\
        );

    \I__6196\ : CascadeMux
    port map (
            O => \N__31607\,
            I => \N__31601\
        );

    \I__6195\ : LocalMux
    port map (
            O => \N__31604\,
            I => \N__31598\
        );

    \I__6194\ : InMux
    port map (
            O => \N__31601\,
            I => \N__31595\
        );

    \I__6193\ : Span4Mux_v
    port map (
            O => \N__31598\,
            I => \N__31591\
        );

    \I__6192\ : LocalMux
    port map (
            O => \N__31595\,
            I => \N__31588\
        );

    \I__6191\ : InMux
    port map (
            O => \N__31594\,
            I => \N__31585\
        );

    \I__6190\ : Odrv4
    port map (
            O => \N__31591\,
            I => \nx.n2690\
        );

    \I__6189\ : Odrv4
    port map (
            O => \N__31588\,
            I => \nx.n2690\
        );

    \I__6188\ : LocalMux
    port map (
            O => \N__31585\,
            I => \nx.n2690\
        );

    \I__6187\ : CascadeMux
    port map (
            O => \N__31578\,
            I => \nx.n2691_cascade_\
        );

    \I__6186\ : CascadeMux
    port map (
            O => \N__31575\,
            I => \N__31571\
        );

    \I__6185\ : InMux
    port map (
            O => \N__31574\,
            I => \N__31568\
        );

    \I__6184\ : InMux
    port map (
            O => \N__31571\,
            I => \N__31565\
        );

    \I__6183\ : LocalMux
    port map (
            O => \N__31568\,
            I => \N__31562\
        );

    \I__6182\ : LocalMux
    port map (
            O => \N__31565\,
            I => \N__31559\
        );

    \I__6181\ : Span4Mux_v
    port map (
            O => \N__31562\,
            I => \N__31555\
        );

    \I__6180\ : Span4Mux_v
    port map (
            O => \N__31559\,
            I => \N__31552\
        );

    \I__6179\ : InMux
    port map (
            O => \N__31558\,
            I => \N__31549\
        );

    \I__6178\ : Odrv4
    port map (
            O => \N__31555\,
            I => \nx.n2692\
        );

    \I__6177\ : Odrv4
    port map (
            O => \N__31552\,
            I => \nx.n2692\
        );

    \I__6176\ : LocalMux
    port map (
            O => \N__31549\,
            I => \nx.n2692\
        );

    \I__6175\ : InMux
    port map (
            O => \N__31542\,
            I => \N__31539\
        );

    \I__6174\ : LocalMux
    port map (
            O => \N__31539\,
            I => \nx.n36\
        );

    \I__6173\ : CascadeMux
    port map (
            O => \N__31536\,
            I => \N__31533\
        );

    \I__6172\ : InMux
    port map (
            O => \N__31533\,
            I => \N__31530\
        );

    \I__6171\ : LocalMux
    port map (
            O => \N__31530\,
            I => \N__31525\
        );

    \I__6170\ : InMux
    port map (
            O => \N__31529\,
            I => \N__31522\
        );

    \I__6169\ : InMux
    port map (
            O => \N__31528\,
            I => \N__31519\
        );

    \I__6168\ : Span4Mux_h
    port map (
            O => \N__31525\,
            I => \N__31516\
        );

    \I__6167\ : LocalMux
    port map (
            O => \N__31522\,
            I => \nx.n2700\
        );

    \I__6166\ : LocalMux
    port map (
            O => \N__31519\,
            I => \nx.n2700\
        );

    \I__6165\ : Odrv4
    port map (
            O => \N__31516\,
            I => \nx.n2700\
        );

    \I__6164\ : CascadeMux
    port map (
            O => \N__31509\,
            I => \N__31506\
        );

    \I__6163\ : InMux
    port map (
            O => \N__31506\,
            I => \N__31502\
        );

    \I__6162\ : CascadeMux
    port map (
            O => \N__31505\,
            I => \N__31499\
        );

    \I__6161\ : LocalMux
    port map (
            O => \N__31502\,
            I => \N__31496\
        );

    \I__6160\ : InMux
    port map (
            O => \N__31499\,
            I => \N__31492\
        );

    \I__6159\ : Span4Mux_h
    port map (
            O => \N__31496\,
            I => \N__31489\
        );

    \I__6158\ : InMux
    port map (
            O => \N__31495\,
            I => \N__31486\
        );

    \I__6157\ : LocalMux
    port map (
            O => \N__31492\,
            I => \nx.n2688\
        );

    \I__6156\ : Odrv4
    port map (
            O => \N__31489\,
            I => \nx.n2688\
        );

    \I__6155\ : LocalMux
    port map (
            O => \N__31486\,
            I => \nx.n2688\
        );

    \I__6154\ : CascadeMux
    port map (
            O => \N__31479\,
            I => \N__31475\
        );

    \I__6153\ : CascadeMux
    port map (
            O => \N__31478\,
            I => \N__31472\
        );

    \I__6152\ : InMux
    port map (
            O => \N__31475\,
            I => \N__31469\
        );

    \I__6151\ : InMux
    port map (
            O => \N__31472\,
            I => \N__31466\
        );

    \I__6150\ : LocalMux
    port map (
            O => \N__31469\,
            I => \N__31463\
        );

    \I__6149\ : LocalMux
    port map (
            O => \N__31466\,
            I => \N__31460\
        );

    \I__6148\ : Span4Mux_v
    port map (
            O => \N__31463\,
            I => \N__31456\
        );

    \I__6147\ : Span4Mux_h
    port map (
            O => \N__31460\,
            I => \N__31453\
        );

    \I__6146\ : InMux
    port map (
            O => \N__31459\,
            I => \N__31450\
        );

    \I__6145\ : Odrv4
    port map (
            O => \N__31456\,
            I => \nx.n2689\
        );

    \I__6144\ : Odrv4
    port map (
            O => \N__31453\,
            I => \nx.n2689\
        );

    \I__6143\ : LocalMux
    port map (
            O => \N__31450\,
            I => \nx.n2689\
        );

    \I__6142\ : CascadeMux
    port map (
            O => \N__31443\,
            I => \nx.n34_cascade_\
        );

    \I__6141\ : CascadeMux
    port map (
            O => \N__31440\,
            I => \N__31436\
        );

    \I__6140\ : InMux
    port map (
            O => \N__31439\,
            I => \N__31433\
        );

    \I__6139\ : InMux
    port map (
            O => \N__31436\,
            I => \N__31429\
        );

    \I__6138\ : LocalMux
    port map (
            O => \N__31433\,
            I => \N__31426\
        );

    \I__6137\ : InMux
    port map (
            O => \N__31432\,
            I => \N__31423\
        );

    \I__6136\ : LocalMux
    port map (
            O => \N__31429\,
            I => \N__31420\
        );

    \I__6135\ : Odrv4
    port map (
            O => \N__31426\,
            I => \nx.n2799\
        );

    \I__6134\ : LocalMux
    port map (
            O => \N__31423\,
            I => \nx.n2799\
        );

    \I__6133\ : Odrv4
    port map (
            O => \N__31420\,
            I => \nx.n2799\
        );

    \I__6132\ : InMux
    port map (
            O => \N__31413\,
            I => \N__31410\
        );

    \I__6131\ : LocalMux
    port map (
            O => \N__31410\,
            I => \N__31407\
        );

    \I__6130\ : Span4Mux_v
    port map (
            O => \N__31407\,
            I => \N__31404\
        );

    \I__6129\ : Odrv4
    port map (
            O => \N__31404\,
            I => \nx.n2866\
        );

    \I__6128\ : CascadeMux
    port map (
            O => \N__31401\,
            I => \nx.n2898_cascade_\
        );

    \I__6127\ : InMux
    port map (
            O => \N__31398\,
            I => \N__31394\
        );

    \I__6126\ : InMux
    port map (
            O => \N__31397\,
            I => \N__31391\
        );

    \I__6125\ : LocalMux
    port map (
            O => \N__31394\,
            I => \nx.n2997\
        );

    \I__6124\ : LocalMux
    port map (
            O => \N__31391\,
            I => \nx.n2997\
        );

    \I__6123\ : CascadeMux
    port map (
            O => \N__31386\,
            I => \nx.n2997_cascade_\
        );

    \I__6122\ : InMux
    port map (
            O => \N__31383\,
            I => \N__31380\
        );

    \I__6121\ : LocalMux
    port map (
            O => \N__31380\,
            I => \N__31377\
        );

    \I__6120\ : Span4Mux_h
    port map (
            O => \N__31377\,
            I => \N__31374\
        );

    \I__6119\ : Odrv4
    port map (
            O => \N__31374\,
            I => \nx.n45\
        );

    \I__6118\ : InMux
    port map (
            O => \N__31371\,
            I => \N__31366\
        );

    \I__6117\ : InMux
    port map (
            O => \N__31370\,
            I => \N__31363\
        );

    \I__6116\ : InMux
    port map (
            O => \N__31369\,
            I => \N__31360\
        );

    \I__6115\ : LocalMux
    port map (
            O => \N__31366\,
            I => \nx.n2988\
        );

    \I__6114\ : LocalMux
    port map (
            O => \N__31363\,
            I => \nx.n2988\
        );

    \I__6113\ : LocalMux
    port map (
            O => \N__31360\,
            I => \nx.n2988\
        );

    \I__6112\ : InMux
    port map (
            O => \N__31353\,
            I => \N__31350\
        );

    \I__6111\ : LocalMux
    port map (
            O => \N__31350\,
            I => \N__31347\
        );

    \I__6110\ : Span4Mux_h
    port map (
            O => \N__31347\,
            I => \N__31344\
        );

    \I__6109\ : Odrv4
    port map (
            O => \N__31344\,
            I => \nx.n2855\
        );

    \I__6108\ : CascadeMux
    port map (
            O => \N__31341\,
            I => \N__31338\
        );

    \I__6107\ : InMux
    port map (
            O => \N__31338\,
            I => \N__31335\
        );

    \I__6106\ : LocalMux
    port map (
            O => \N__31335\,
            I => \N__31332\
        );

    \I__6105\ : Span4Mux_h
    port map (
            O => \N__31332\,
            I => \N__31328\
        );

    \I__6104\ : InMux
    port map (
            O => \N__31331\,
            I => \N__31325\
        );

    \I__6103\ : Odrv4
    port map (
            O => \N__31328\,
            I => \nx.n2788\
        );

    \I__6102\ : LocalMux
    port map (
            O => \N__31325\,
            I => \nx.n2788\
        );

    \I__6101\ : InMux
    port map (
            O => \N__31320\,
            I => \N__31317\
        );

    \I__6100\ : LocalMux
    port map (
            O => \N__31317\,
            I => \N__31314\
        );

    \I__6099\ : Span4Mux_v
    port map (
            O => \N__31314\,
            I => \N__31311\
        );

    \I__6098\ : Odrv4
    port map (
            O => \N__31311\,
            I => \nx.n2764\
        );

    \I__6097\ : CascadeMux
    port map (
            O => \N__31308\,
            I => \N__31305\
        );

    \I__6096\ : InMux
    port map (
            O => \N__31305\,
            I => \N__31302\
        );

    \I__6095\ : LocalMux
    port map (
            O => \N__31302\,
            I => \N__31298\
        );

    \I__6094\ : CascadeMux
    port map (
            O => \N__31301\,
            I => \N__31295\
        );

    \I__6093\ : Span4Mux_h
    port map (
            O => \N__31298\,
            I => \N__31291\
        );

    \I__6092\ : InMux
    port map (
            O => \N__31295\,
            I => \N__31288\
        );

    \I__6091\ : InMux
    port map (
            O => \N__31294\,
            I => \N__31285\
        );

    \I__6090\ : Odrv4
    port map (
            O => \N__31291\,
            I => \nx.n2697\
        );

    \I__6089\ : LocalMux
    port map (
            O => \N__31288\,
            I => \nx.n2697\
        );

    \I__6088\ : LocalMux
    port map (
            O => \N__31285\,
            I => \nx.n2697\
        );

    \I__6087\ : CascadeMux
    port map (
            O => \N__31278\,
            I => \N__31271\
        );

    \I__6086\ : CascadeMux
    port map (
            O => \N__31277\,
            I => \N__31265\
        );

    \I__6085\ : CascadeMux
    port map (
            O => \N__31276\,
            I => \N__31262\
        );

    \I__6084\ : CascadeMux
    port map (
            O => \N__31275\,
            I => \N__31256\
        );

    \I__6083\ : InMux
    port map (
            O => \N__31274\,
            I => \N__31249\
        );

    \I__6082\ : InMux
    port map (
            O => \N__31271\,
            I => \N__31244\
        );

    \I__6081\ : InMux
    port map (
            O => \N__31270\,
            I => \N__31244\
        );

    \I__6080\ : InMux
    port map (
            O => \N__31269\,
            I => \N__31231\
        );

    \I__6079\ : InMux
    port map (
            O => \N__31268\,
            I => \N__31231\
        );

    \I__6078\ : InMux
    port map (
            O => \N__31265\,
            I => \N__31231\
        );

    \I__6077\ : InMux
    port map (
            O => \N__31262\,
            I => \N__31231\
        );

    \I__6076\ : InMux
    port map (
            O => \N__31261\,
            I => \N__31231\
        );

    \I__6075\ : InMux
    port map (
            O => \N__31260\,
            I => \N__31231\
        );

    \I__6074\ : CascadeMux
    port map (
            O => \N__31259\,
            I => \N__31227\
        );

    \I__6073\ : InMux
    port map (
            O => \N__31256\,
            I => \N__31223\
        );

    \I__6072\ : CascadeMux
    port map (
            O => \N__31255\,
            I => \N__31217\
        );

    \I__6071\ : CascadeMux
    port map (
            O => \N__31254\,
            I => \N__31213\
        );

    \I__6070\ : CascadeMux
    port map (
            O => \N__31253\,
            I => \N__31209\
        );

    \I__6069\ : CascadeMux
    port map (
            O => \N__31252\,
            I => \N__31206\
        );

    \I__6068\ : LocalMux
    port map (
            O => \N__31249\,
            I => \N__31202\
        );

    \I__6067\ : LocalMux
    port map (
            O => \N__31244\,
            I => \N__31199\
        );

    \I__6066\ : LocalMux
    port map (
            O => \N__31231\,
            I => \N__31196\
        );

    \I__6065\ : InMux
    port map (
            O => \N__31230\,
            I => \N__31189\
        );

    \I__6064\ : InMux
    port map (
            O => \N__31227\,
            I => \N__31189\
        );

    \I__6063\ : InMux
    port map (
            O => \N__31226\,
            I => \N__31189\
        );

    \I__6062\ : LocalMux
    port map (
            O => \N__31223\,
            I => \N__31186\
        );

    \I__6061\ : InMux
    port map (
            O => \N__31222\,
            I => \N__31181\
        );

    \I__6060\ : InMux
    port map (
            O => \N__31221\,
            I => \N__31181\
        );

    \I__6059\ : InMux
    port map (
            O => \N__31220\,
            I => \N__31172\
        );

    \I__6058\ : InMux
    port map (
            O => \N__31217\,
            I => \N__31172\
        );

    \I__6057\ : InMux
    port map (
            O => \N__31216\,
            I => \N__31172\
        );

    \I__6056\ : InMux
    port map (
            O => \N__31213\,
            I => \N__31172\
        );

    \I__6055\ : InMux
    port map (
            O => \N__31212\,
            I => \N__31163\
        );

    \I__6054\ : InMux
    port map (
            O => \N__31209\,
            I => \N__31163\
        );

    \I__6053\ : InMux
    port map (
            O => \N__31206\,
            I => \N__31163\
        );

    \I__6052\ : InMux
    port map (
            O => \N__31205\,
            I => \N__31163\
        );

    \I__6051\ : Span4Mux_v
    port map (
            O => \N__31202\,
            I => \N__31154\
        );

    \I__6050\ : Span4Mux_v
    port map (
            O => \N__31199\,
            I => \N__31154\
        );

    \I__6049\ : Span4Mux_v
    port map (
            O => \N__31196\,
            I => \N__31154\
        );

    \I__6048\ : LocalMux
    port map (
            O => \N__31189\,
            I => \N__31154\
        );

    \I__6047\ : Odrv4
    port map (
            O => \N__31186\,
            I => \nx.n2720\
        );

    \I__6046\ : LocalMux
    port map (
            O => \N__31181\,
            I => \nx.n2720\
        );

    \I__6045\ : LocalMux
    port map (
            O => \N__31172\,
            I => \nx.n2720\
        );

    \I__6044\ : LocalMux
    port map (
            O => \N__31163\,
            I => \nx.n2720\
        );

    \I__6043\ : Odrv4
    port map (
            O => \N__31154\,
            I => \nx.n2720\
        );

    \I__6042\ : CascadeMux
    port map (
            O => \N__31143\,
            I => \N__31140\
        );

    \I__6041\ : InMux
    port map (
            O => \N__31140\,
            I => \N__31135\
        );

    \I__6040\ : CascadeMux
    port map (
            O => \N__31139\,
            I => \N__31132\
        );

    \I__6039\ : InMux
    port map (
            O => \N__31138\,
            I => \N__31129\
        );

    \I__6038\ : LocalMux
    port map (
            O => \N__31135\,
            I => \N__31126\
        );

    \I__6037\ : InMux
    port map (
            O => \N__31132\,
            I => \N__31123\
        );

    \I__6036\ : LocalMux
    port map (
            O => \N__31129\,
            I => \N__31118\
        );

    \I__6035\ : Span4Mux_h
    port map (
            O => \N__31126\,
            I => \N__31118\
        );

    \I__6034\ : LocalMux
    port map (
            O => \N__31123\,
            I => \nx.n2796\
        );

    \I__6033\ : Odrv4
    port map (
            O => \N__31118\,
            I => \nx.n2796\
        );

    \I__6032\ : InMux
    port map (
            O => \N__31113\,
            I => \N__31108\
        );

    \I__6031\ : InMux
    port map (
            O => \N__31112\,
            I => \N__31105\
        );

    \I__6030\ : InMux
    port map (
            O => \N__31111\,
            I => \N__31102\
        );

    \I__6029\ : LocalMux
    port map (
            O => \N__31108\,
            I => \N__31099\
        );

    \I__6028\ : LocalMux
    port map (
            O => \N__31105\,
            I => \nx.n3000\
        );

    \I__6027\ : LocalMux
    port map (
            O => \N__31102\,
            I => \nx.n3000\
        );

    \I__6026\ : Odrv4
    port map (
            O => \N__31099\,
            I => \nx.n3000\
        );

    \I__6025\ : InMux
    port map (
            O => \N__31092\,
            I => \N__31088\
        );

    \I__6024\ : InMux
    port map (
            O => \N__31091\,
            I => \N__31085\
        );

    \I__6023\ : LocalMux
    port map (
            O => \N__31088\,
            I => \nx.n3001\
        );

    \I__6022\ : LocalMux
    port map (
            O => \N__31085\,
            I => \nx.n3001\
        );

    \I__6021\ : CascadeMux
    port map (
            O => \N__31080\,
            I => \nx.n3001_cascade_\
        );

    \I__6020\ : InMux
    port map (
            O => \N__31077\,
            I => \N__31074\
        );

    \I__6019\ : LocalMux
    port map (
            O => \N__31074\,
            I => \N__31071\
        );

    \I__6018\ : Odrv4
    port map (
            O => \N__31071\,
            I => \nx.n44\
        );

    \I__6017\ : InMux
    port map (
            O => \N__31068\,
            I => \N__31063\
        );

    \I__6016\ : InMux
    port map (
            O => \N__31067\,
            I => \N__31060\
        );

    \I__6015\ : InMux
    port map (
            O => \N__31066\,
            I => \N__31057\
        );

    \I__6014\ : LocalMux
    port map (
            O => \N__31063\,
            I => \nx.n3003\
        );

    \I__6013\ : LocalMux
    port map (
            O => \N__31060\,
            I => \nx.n3003\
        );

    \I__6012\ : LocalMux
    port map (
            O => \N__31057\,
            I => \nx.n3003\
        );

    \I__6011\ : InMux
    port map (
            O => \N__31050\,
            I => \N__31045\
        );

    \I__6010\ : InMux
    port map (
            O => \N__31049\,
            I => \N__31042\
        );

    \I__6009\ : InMux
    port map (
            O => \N__31048\,
            I => \N__31039\
        );

    \I__6008\ : LocalMux
    port map (
            O => \N__31045\,
            I => \nx.n3005\
        );

    \I__6007\ : LocalMux
    port map (
            O => \N__31042\,
            I => \nx.n3005\
        );

    \I__6006\ : LocalMux
    port map (
            O => \N__31039\,
            I => \nx.n3005\
        );

    \I__6005\ : CascadeMux
    port map (
            O => \N__31032\,
            I => \N__31029\
        );

    \I__6004\ : InMux
    port map (
            O => \N__31029\,
            I => \N__31026\
        );

    \I__6003\ : LocalMux
    port map (
            O => \N__31026\,
            I => \N__31023\
        );

    \I__6002\ : Span4Mux_v
    port map (
            O => \N__31023\,
            I => \N__31020\
        );

    \I__6001\ : Odrv4
    port map (
            O => \N__31020\,
            I => \nx.n2863\
        );

    \I__6000\ : CascadeMux
    port map (
            O => \N__31017\,
            I => \nx.n2895_cascade_\
        );

    \I__5999\ : CascadeMux
    port map (
            O => \N__31014\,
            I => \N__31009\
        );

    \I__5998\ : InMux
    port map (
            O => \N__31013\,
            I => \N__31006\
        );

    \I__5997\ : InMux
    port map (
            O => \N__31012\,
            I => \N__31003\
        );

    \I__5996\ : InMux
    port map (
            O => \N__31009\,
            I => \N__31000\
        );

    \I__5995\ : LocalMux
    port map (
            O => \N__31006\,
            I => \nx.n2994\
        );

    \I__5994\ : LocalMux
    port map (
            O => \N__31003\,
            I => \nx.n2994\
        );

    \I__5993\ : LocalMux
    port map (
            O => \N__31000\,
            I => \nx.n2994\
        );

    \I__5992\ : CascadeMux
    port map (
            O => \N__30993\,
            I => \nx.n25_adj_748_cascade_\
        );

    \I__5991\ : InMux
    port map (
            O => \N__30990\,
            I => \N__30987\
        );

    \I__5990\ : LocalMux
    port map (
            O => \N__30987\,
            I => \nx.n12785\
        );

    \I__5989\ : InMux
    port map (
            O => \N__30984\,
            I => \N__30981\
        );

    \I__5988\ : LocalMux
    port map (
            O => \N__30981\,
            I => \nx.n19_adj_745\
        );

    \I__5987\ : CascadeMux
    port map (
            O => \N__30978\,
            I => \nx.n12777_cascade_\
        );

    \I__5986\ : InMux
    port map (
            O => \N__30975\,
            I => \N__30972\
        );

    \I__5985\ : LocalMux
    port map (
            O => \N__30972\,
            I => \nx.n12779\
        );

    \I__5984\ : CascadeMux
    port map (
            O => \N__30969\,
            I => \nx.n39_adj_747_cascade_\
        );

    \I__5983\ : InMux
    port map (
            O => \N__30966\,
            I => \N__30963\
        );

    \I__5982\ : LocalMux
    port map (
            O => \N__30963\,
            I => \nx.n12789\
        );

    \I__5981\ : InMux
    port map (
            O => \N__30960\,
            I => \N__30957\
        );

    \I__5980\ : LocalMux
    port map (
            O => \N__30957\,
            I => \N__30954\
        );

    \I__5979\ : Odrv4
    port map (
            O => \N__30954\,
            I => \nx.n12799\
        );

    \I__5978\ : InMux
    port map (
            O => \N__30951\,
            I => \N__30948\
        );

    \I__5977\ : LocalMux
    port map (
            O => \N__30948\,
            I => \nx.n29_adj_746\
        );

    \I__5976\ : InMux
    port map (
            O => \N__30945\,
            I => \N__30942\
        );

    \I__5975\ : LocalMux
    port map (
            O => \N__30942\,
            I => \N__30939\
        );

    \I__5974\ : Span4Mux_h
    port map (
            O => \N__30939\,
            I => \N__30936\
        );

    \I__5973\ : Odrv4
    port map (
            O => \N__30936\,
            I => \nx.n11_adj_751\
        );

    \I__5972\ : InMux
    port map (
            O => \N__30933\,
            I => \N__30930\
        );

    \I__5971\ : LocalMux
    port map (
            O => \N__30930\,
            I => \N__30927\
        );

    \I__5970\ : Odrv4
    port map (
            O => \N__30927\,
            I => \nx.n41_adj_752\
        );

    \I__5969\ : InMux
    port map (
            O => \N__30924\,
            I => \N__30921\
        );

    \I__5968\ : LocalMux
    port map (
            O => \N__30921\,
            I => \N__30916\
        );

    \I__5967\ : InMux
    port map (
            O => \N__30920\,
            I => \N__30913\
        );

    \I__5966\ : InMux
    port map (
            O => \N__30919\,
            I => \N__30910\
        );

    \I__5965\ : Span4Mux_v
    port map (
            O => \N__30916\,
            I => \N__30907\
        );

    \I__5964\ : LocalMux
    port map (
            O => \N__30913\,
            I => \N__30904\
        );

    \I__5963\ : LocalMux
    port map (
            O => \N__30910\,
            I => \N__30901\
        );

    \I__5962\ : Odrv4
    port map (
            O => \N__30907\,
            I => \nx.n2989\
        );

    \I__5961\ : Odrv4
    port map (
            O => \N__30904\,
            I => \nx.n2989\
        );

    \I__5960\ : Odrv4
    port map (
            O => \N__30901\,
            I => \nx.n2989\
        );

    \I__5959\ : CascadeMux
    port map (
            O => \N__30894\,
            I => \N__30891\
        );

    \I__5958\ : InMux
    port map (
            O => \N__30891\,
            I => \N__30888\
        );

    \I__5957\ : LocalMux
    port map (
            O => \N__30888\,
            I => \N__30884\
        );

    \I__5956\ : InMux
    port map (
            O => \N__30887\,
            I => \N__30881\
        );

    \I__5955\ : Span4Mux_v
    port map (
            O => \N__30884\,
            I => \N__30878\
        );

    \I__5954\ : LocalMux
    port map (
            O => \N__30881\,
            I => \nx.n2094\
        );

    \I__5953\ : Odrv4
    port map (
            O => \N__30878\,
            I => \nx.n2094\
        );

    \I__5952\ : InMux
    port map (
            O => \N__30873\,
            I => \N__30870\
        );

    \I__5951\ : LocalMux
    port map (
            O => \N__30870\,
            I => \N__30867\
        );

    \I__5950\ : Odrv4
    port map (
            O => \N__30867\,
            I => \nx.n2161\
        );

    \I__5949\ : InMux
    port map (
            O => \N__30864\,
            I => \bfn_11_31_0_\
        );

    \I__5948\ : InMux
    port map (
            O => \N__30861\,
            I => \N__30858\
        );

    \I__5947\ : LocalMux
    port map (
            O => \N__30858\,
            I => \N__30855\
        );

    \I__5946\ : Span4Mux_v
    port map (
            O => \N__30855\,
            I => \N__30851\
        );

    \I__5945\ : InMux
    port map (
            O => \N__30854\,
            I => \N__30848\
        );

    \I__5944\ : Odrv4
    port map (
            O => \N__30851\,
            I => \nx.n2093\
        );

    \I__5943\ : LocalMux
    port map (
            O => \N__30848\,
            I => \nx.n2093\
        );

    \I__5942\ : InMux
    port map (
            O => \N__30843\,
            I => \nx.n10880\
        );

    \I__5941\ : CascadeMux
    port map (
            O => \N__30840\,
            I => \N__30837\
        );

    \I__5940\ : InMux
    port map (
            O => \N__30837\,
            I => \N__30834\
        );

    \I__5939\ : LocalMux
    port map (
            O => \N__30834\,
            I => \N__30830\
        );

    \I__5938\ : InMux
    port map (
            O => \N__30833\,
            I => \N__30827\
        );

    \I__5937\ : Span4Mux_h
    port map (
            O => \N__30830\,
            I => \N__30822\
        );

    \I__5936\ : LocalMux
    port map (
            O => \N__30827\,
            I => \N__30822\
        );

    \I__5935\ : Odrv4
    port map (
            O => \N__30822\,
            I => \nx.n2192\
        );

    \I__5934\ : CascadeMux
    port map (
            O => \N__30819\,
            I => \nx.n21_adj_750_cascade_\
        );

    \I__5933\ : InMux
    port map (
            O => \N__30816\,
            I => \N__30812\
        );

    \I__5932\ : InMux
    port map (
            O => \N__30815\,
            I => \N__30808\
        );

    \I__5931\ : LocalMux
    port map (
            O => \N__30812\,
            I => \N__30805\
        );

    \I__5930\ : InMux
    port map (
            O => \N__30811\,
            I => \N__30802\
        );

    \I__5929\ : LocalMux
    port map (
            O => \N__30808\,
            I => \N__30799\
        );

    \I__5928\ : Span4Mux_v
    port map (
            O => \N__30805\,
            I => \N__30796\
        );

    \I__5927\ : LocalMux
    port map (
            O => \N__30802\,
            I => \N__30793\
        );

    \I__5926\ : Span4Mux_v
    port map (
            O => \N__30799\,
            I => \N__30788\
        );

    \I__5925\ : Span4Mux_v
    port map (
            O => \N__30796\,
            I => \N__30785\
        );

    \I__5924\ : Span4Mux_v
    port map (
            O => \N__30793\,
            I => \N__30782\
        );

    \I__5923\ : InMux
    port map (
            O => \N__30792\,
            I => \N__30779\
        );

    \I__5922\ : InMux
    port map (
            O => \N__30791\,
            I => \N__30776\
        );

    \I__5921\ : Span4Mux_v
    port map (
            O => \N__30788\,
            I => \N__30771\
        );

    \I__5920\ : Span4Mux_h
    port map (
            O => \N__30785\,
            I => \N__30771\
        );

    \I__5919\ : Odrv4
    port map (
            O => \N__30782\,
            I => \nx.bit_ctr_3\
        );

    \I__5918\ : LocalMux
    port map (
            O => \N__30779\,
            I => \nx.bit_ctr_3\
        );

    \I__5917\ : LocalMux
    port map (
            O => \N__30776\,
            I => \nx.bit_ctr_3\
        );

    \I__5916\ : Odrv4
    port map (
            O => \N__30771\,
            I => \nx.bit_ctr_3\
        );

    \I__5915\ : CascadeMux
    port map (
            O => \N__30762\,
            I => \nx.n12781_cascade_\
        );

    \I__5914\ : InMux
    port map (
            O => \N__30759\,
            I => \N__30756\
        );

    \I__5913\ : LocalMux
    port map (
            O => \N__30756\,
            I => \N__30753\
        );

    \I__5912\ : Odrv4
    port map (
            O => \N__30753\,
            I => \nx.n12801\
        );

    \I__5911\ : CascadeMux
    port map (
            O => \N__30750\,
            I => \nx.n27_adj_744_cascade_\
        );

    \I__5910\ : InMux
    port map (
            O => \N__30747\,
            I => \N__30744\
        );

    \I__5909\ : LocalMux
    port map (
            O => \N__30744\,
            I => \N__30740\
        );

    \I__5908\ : InMux
    port map (
            O => \N__30743\,
            I => \N__30737\
        );

    \I__5907\ : Odrv4
    port map (
            O => \N__30740\,
            I => \nx.n3209\
        );

    \I__5906\ : LocalMux
    port map (
            O => \N__30737\,
            I => \nx.n3209\
        );

    \I__5905\ : InMux
    port map (
            O => \N__30732\,
            I => \bfn_11_30_0_\
        );

    \I__5904\ : InMux
    port map (
            O => \N__30729\,
            I => \nx.n10872\
        );

    \I__5903\ : CascadeMux
    port map (
            O => \N__30726\,
            I => \N__30723\
        );

    \I__5902\ : InMux
    port map (
            O => \N__30723\,
            I => \N__30719\
        );

    \I__5901\ : InMux
    port map (
            O => \N__30722\,
            I => \N__30716\
        );

    \I__5900\ : LocalMux
    port map (
            O => \N__30719\,
            I => \N__30713\
        );

    \I__5899\ : LocalMux
    port map (
            O => \N__30716\,
            I => \N__30709\
        );

    \I__5898\ : Span4Mux_h
    port map (
            O => \N__30713\,
            I => \N__30706\
        );

    \I__5897\ : InMux
    port map (
            O => \N__30712\,
            I => \N__30703\
        );

    \I__5896\ : Odrv4
    port map (
            O => \N__30709\,
            I => \nx.n2100\
        );

    \I__5895\ : Odrv4
    port map (
            O => \N__30706\,
            I => \nx.n2100\
        );

    \I__5894\ : LocalMux
    port map (
            O => \N__30703\,
            I => \nx.n2100\
        );

    \I__5893\ : CascadeMux
    port map (
            O => \N__30696\,
            I => \N__30693\
        );

    \I__5892\ : InMux
    port map (
            O => \N__30693\,
            I => \N__30690\
        );

    \I__5891\ : LocalMux
    port map (
            O => \N__30690\,
            I => \N__30687\
        );

    \I__5890\ : Odrv4
    port map (
            O => \N__30687\,
            I => \nx.n2167\
        );

    \I__5889\ : InMux
    port map (
            O => \N__30684\,
            I => \nx.n10873\
        );

    \I__5888\ : InMux
    port map (
            O => \N__30681\,
            I => \nx.n10874\
        );

    \I__5887\ : CascadeMux
    port map (
            O => \N__30678\,
            I => \N__30675\
        );

    \I__5886\ : InMux
    port map (
            O => \N__30675\,
            I => \N__30672\
        );

    \I__5885\ : LocalMux
    port map (
            O => \N__30672\,
            I => \N__30667\
        );

    \I__5884\ : InMux
    port map (
            O => \N__30671\,
            I => \N__30664\
        );

    \I__5883\ : InMux
    port map (
            O => \N__30670\,
            I => \N__30661\
        );

    \I__5882\ : Span4Mux_s3_v
    port map (
            O => \N__30667\,
            I => \N__30658\
        );

    \I__5881\ : LocalMux
    port map (
            O => \N__30664\,
            I => \N__30655\
        );

    \I__5880\ : LocalMux
    port map (
            O => \N__30661\,
            I => \nx.n2098\
        );

    \I__5879\ : Odrv4
    port map (
            O => \N__30658\,
            I => \nx.n2098\
        );

    \I__5878\ : Odrv4
    port map (
            O => \N__30655\,
            I => \nx.n2098\
        );

    \I__5877\ : InMux
    port map (
            O => \N__30648\,
            I => \N__30645\
        );

    \I__5876\ : LocalMux
    port map (
            O => \N__30645\,
            I => \N__30642\
        );

    \I__5875\ : Odrv4
    port map (
            O => \N__30642\,
            I => \nx.n2165\
        );

    \I__5874\ : InMux
    port map (
            O => \N__30639\,
            I => \nx.n10875\
        );

    \I__5873\ : CascadeMux
    port map (
            O => \N__30636\,
            I => \N__30632\
        );

    \I__5872\ : InMux
    port map (
            O => \N__30635\,
            I => \N__30629\
        );

    \I__5871\ : InMux
    port map (
            O => \N__30632\,
            I => \N__30625\
        );

    \I__5870\ : LocalMux
    port map (
            O => \N__30629\,
            I => \N__30622\
        );

    \I__5869\ : InMux
    port map (
            O => \N__30628\,
            I => \N__30619\
        );

    \I__5868\ : LocalMux
    port map (
            O => \N__30625\,
            I => \nx.n2097\
        );

    \I__5867\ : Odrv4
    port map (
            O => \N__30622\,
            I => \nx.n2097\
        );

    \I__5866\ : LocalMux
    port map (
            O => \N__30619\,
            I => \nx.n2097\
        );

    \I__5865\ : InMux
    port map (
            O => \N__30612\,
            I => \N__30609\
        );

    \I__5864\ : LocalMux
    port map (
            O => \N__30609\,
            I => \N__30606\
        );

    \I__5863\ : Odrv4
    port map (
            O => \N__30606\,
            I => \nx.n2164\
        );

    \I__5862\ : InMux
    port map (
            O => \N__30603\,
            I => \nx.n10876\
        );

    \I__5861\ : CascadeMux
    port map (
            O => \N__30600\,
            I => \N__30597\
        );

    \I__5860\ : InMux
    port map (
            O => \N__30597\,
            I => \N__30593\
        );

    \I__5859\ : InMux
    port map (
            O => \N__30596\,
            I => \N__30590\
        );

    \I__5858\ : LocalMux
    port map (
            O => \N__30593\,
            I => \N__30587\
        );

    \I__5857\ : LocalMux
    port map (
            O => \N__30590\,
            I => \nx.n2096\
        );

    \I__5856\ : Odrv4
    port map (
            O => \N__30587\,
            I => \nx.n2096\
        );

    \I__5855\ : CascadeMux
    port map (
            O => \N__30582\,
            I => \N__30579\
        );

    \I__5854\ : InMux
    port map (
            O => \N__30579\,
            I => \N__30576\
        );

    \I__5853\ : LocalMux
    port map (
            O => \N__30576\,
            I => \nx.n2163\
        );

    \I__5852\ : InMux
    port map (
            O => \N__30573\,
            I => \nx.n10877\
        );

    \I__5851\ : CascadeMux
    port map (
            O => \N__30570\,
            I => \N__30566\
        );

    \I__5850\ : CascadeMux
    port map (
            O => \N__30569\,
            I => \N__30563\
        );

    \I__5849\ : InMux
    port map (
            O => \N__30566\,
            I => \N__30559\
        );

    \I__5848\ : InMux
    port map (
            O => \N__30563\,
            I => \N__30556\
        );

    \I__5847\ : InMux
    port map (
            O => \N__30562\,
            I => \N__30553\
        );

    \I__5846\ : LocalMux
    port map (
            O => \N__30559\,
            I => \nx.n2095\
        );

    \I__5845\ : LocalMux
    port map (
            O => \N__30556\,
            I => \nx.n2095\
        );

    \I__5844\ : LocalMux
    port map (
            O => \N__30553\,
            I => \nx.n2095\
        );

    \I__5843\ : InMux
    port map (
            O => \N__30546\,
            I => \N__30543\
        );

    \I__5842\ : LocalMux
    port map (
            O => \N__30543\,
            I => \N__30540\
        );

    \I__5841\ : Odrv4
    port map (
            O => \N__30540\,
            I => \nx.n2162\
        );

    \I__5840\ : InMux
    port map (
            O => \N__30537\,
            I => \nx.n10878\
        );

    \I__5839\ : CascadeMux
    port map (
            O => \N__30534\,
            I => \N__30529\
        );

    \I__5838\ : InMux
    port map (
            O => \N__30533\,
            I => \N__30525\
        );

    \I__5837\ : InMux
    port map (
            O => \N__30532\,
            I => \N__30522\
        );

    \I__5836\ : InMux
    port map (
            O => \N__30529\,
            I => \N__30519\
        );

    \I__5835\ : InMux
    port map (
            O => \N__30528\,
            I => \N__30516\
        );

    \I__5834\ : LocalMux
    port map (
            O => \N__30525\,
            I => \N__30511\
        );

    \I__5833\ : LocalMux
    port map (
            O => \N__30522\,
            I => \N__30511\
        );

    \I__5832\ : LocalMux
    port map (
            O => \N__30519\,
            I => \N__30507\
        );

    \I__5831\ : LocalMux
    port map (
            O => \N__30516\,
            I => \N__30502\
        );

    \I__5830\ : Span4Mux_v
    port map (
            O => \N__30511\,
            I => \N__30502\
        );

    \I__5829\ : InMux
    port map (
            O => \N__30510\,
            I => \N__30499\
        );

    \I__5828\ : Span4Mux_v
    port map (
            O => \N__30507\,
            I => \N__30496\
        );

    \I__5827\ : Span4Mux_h
    port map (
            O => \N__30502\,
            I => \N__30493\
        );

    \I__5826\ : LocalMux
    port map (
            O => \N__30499\,
            I => \nx.bit_ctr_14\
        );

    \I__5825\ : Odrv4
    port map (
            O => \N__30496\,
            I => \nx.bit_ctr_14\
        );

    \I__5824\ : Odrv4
    port map (
            O => \N__30493\,
            I => \nx.bit_ctr_14\
        );

    \I__5823\ : CascadeMux
    port map (
            O => \N__30486\,
            I => \N__30483\
        );

    \I__5822\ : InMux
    port map (
            O => \N__30483\,
            I => \N__30480\
        );

    \I__5821\ : LocalMux
    port map (
            O => \N__30480\,
            I => \N__30477\
        );

    \I__5820\ : Odrv4
    port map (
            O => \N__30477\,
            I => \nx.n2177\
        );

    \I__5819\ : InMux
    port map (
            O => \N__30474\,
            I => \bfn_11_29_0_\
        );

    \I__5818\ : CascadeMux
    port map (
            O => \N__30471\,
            I => \N__30467\
        );

    \I__5817\ : InMux
    port map (
            O => \N__30470\,
            I => \N__30464\
        );

    \I__5816\ : InMux
    port map (
            O => \N__30467\,
            I => \N__30461\
        );

    \I__5815\ : LocalMux
    port map (
            O => \N__30464\,
            I => \nx.n2109\
        );

    \I__5814\ : LocalMux
    port map (
            O => \N__30461\,
            I => \nx.n2109\
        );

    \I__5813\ : InMux
    port map (
            O => \N__30456\,
            I => \N__30453\
        );

    \I__5812\ : LocalMux
    port map (
            O => \N__30453\,
            I => \nx.n2176\
        );

    \I__5811\ : InMux
    port map (
            O => \N__30450\,
            I => \nx.n10864\
        );

    \I__5810\ : CascadeMux
    port map (
            O => \N__30447\,
            I => \N__30443\
        );

    \I__5809\ : InMux
    port map (
            O => \N__30446\,
            I => \N__30440\
        );

    \I__5808\ : InMux
    port map (
            O => \N__30443\,
            I => \N__30437\
        );

    \I__5807\ : LocalMux
    port map (
            O => \N__30440\,
            I => \nx.n2108\
        );

    \I__5806\ : LocalMux
    port map (
            O => \N__30437\,
            I => \nx.n2108\
        );

    \I__5805\ : InMux
    port map (
            O => \N__30432\,
            I => \N__30429\
        );

    \I__5804\ : LocalMux
    port map (
            O => \N__30429\,
            I => \nx.n2175\
        );

    \I__5803\ : InMux
    port map (
            O => \N__30426\,
            I => \nx.n10865\
        );

    \I__5802\ : CascadeMux
    port map (
            O => \N__30423\,
            I => \N__30419\
        );

    \I__5801\ : InMux
    port map (
            O => \N__30422\,
            I => \N__30416\
        );

    \I__5800\ : InMux
    port map (
            O => \N__30419\,
            I => \N__30413\
        );

    \I__5799\ : LocalMux
    port map (
            O => \N__30416\,
            I => \nx.n2107\
        );

    \I__5798\ : LocalMux
    port map (
            O => \N__30413\,
            I => \nx.n2107\
        );

    \I__5797\ : InMux
    port map (
            O => \N__30408\,
            I => \N__30405\
        );

    \I__5796\ : LocalMux
    port map (
            O => \N__30405\,
            I => \nx.n2174\
        );

    \I__5795\ : InMux
    port map (
            O => \N__30402\,
            I => \nx.n10866\
        );

    \I__5794\ : InMux
    port map (
            O => \N__30399\,
            I => \N__30392\
        );

    \I__5793\ : InMux
    port map (
            O => \N__30398\,
            I => \N__30392\
        );

    \I__5792\ : InMux
    port map (
            O => \N__30397\,
            I => \N__30389\
        );

    \I__5791\ : LocalMux
    port map (
            O => \N__30392\,
            I => \N__30384\
        );

    \I__5790\ : LocalMux
    port map (
            O => \N__30389\,
            I => \N__30384\
        );

    \I__5789\ : Odrv4
    port map (
            O => \N__30384\,
            I => \nx.n2106\
        );

    \I__5788\ : InMux
    port map (
            O => \N__30381\,
            I => \N__30378\
        );

    \I__5787\ : LocalMux
    port map (
            O => \N__30378\,
            I => \nx.n2173\
        );

    \I__5786\ : InMux
    port map (
            O => \N__30375\,
            I => \nx.n10867\
        );

    \I__5785\ : CascadeMux
    port map (
            O => \N__30372\,
            I => \N__30369\
        );

    \I__5784\ : InMux
    port map (
            O => \N__30369\,
            I => \N__30366\
        );

    \I__5783\ : LocalMux
    port map (
            O => \N__30366\,
            I => \N__30362\
        );

    \I__5782\ : InMux
    port map (
            O => \N__30365\,
            I => \N__30359\
        );

    \I__5781\ : Odrv4
    port map (
            O => \N__30362\,
            I => \nx.n2105\
        );

    \I__5780\ : LocalMux
    port map (
            O => \N__30359\,
            I => \nx.n2105\
        );

    \I__5779\ : InMux
    port map (
            O => \N__30354\,
            I => \N__30351\
        );

    \I__5778\ : LocalMux
    port map (
            O => \N__30351\,
            I => \N__30348\
        );

    \I__5777\ : Odrv4
    port map (
            O => \N__30348\,
            I => \nx.n2172\
        );

    \I__5776\ : InMux
    port map (
            O => \N__30345\,
            I => \nx.n10868\
        );

    \I__5775\ : CascadeMux
    port map (
            O => \N__30342\,
            I => \N__30339\
        );

    \I__5774\ : InMux
    port map (
            O => \N__30339\,
            I => \N__30334\
        );

    \I__5773\ : InMux
    port map (
            O => \N__30338\,
            I => \N__30331\
        );

    \I__5772\ : InMux
    port map (
            O => \N__30337\,
            I => \N__30328\
        );

    \I__5771\ : LocalMux
    port map (
            O => \N__30334\,
            I => \N__30325\
        );

    \I__5770\ : LocalMux
    port map (
            O => \N__30331\,
            I => \nx.n2104\
        );

    \I__5769\ : LocalMux
    port map (
            O => \N__30328\,
            I => \nx.n2104\
        );

    \I__5768\ : Odrv4
    port map (
            O => \N__30325\,
            I => \nx.n2104\
        );

    \I__5767\ : InMux
    port map (
            O => \N__30318\,
            I => \N__30315\
        );

    \I__5766\ : LocalMux
    port map (
            O => \N__30315\,
            I => \nx.n2171\
        );

    \I__5765\ : InMux
    port map (
            O => \N__30312\,
            I => \nx.n10869\
        );

    \I__5764\ : CascadeMux
    port map (
            O => \N__30309\,
            I => \N__30306\
        );

    \I__5763\ : InMux
    port map (
            O => \N__30306\,
            I => \N__30302\
        );

    \I__5762\ : InMux
    port map (
            O => \N__30305\,
            I => \N__30299\
        );

    \I__5761\ : LocalMux
    port map (
            O => \N__30302\,
            I => \N__30296\
        );

    \I__5760\ : LocalMux
    port map (
            O => \N__30299\,
            I => \nx.n2103\
        );

    \I__5759\ : Odrv4
    port map (
            O => \N__30296\,
            I => \nx.n2103\
        );

    \I__5758\ : InMux
    port map (
            O => \N__30291\,
            I => \N__30288\
        );

    \I__5757\ : LocalMux
    port map (
            O => \N__30288\,
            I => \nx.n2170\
        );

    \I__5756\ : InMux
    port map (
            O => \N__30285\,
            I => \nx.n10870\
        );

    \I__5755\ : CascadeMux
    port map (
            O => \N__30282\,
            I => \N__30278\
        );

    \I__5754\ : CascadeMux
    port map (
            O => \N__30281\,
            I => \N__30275\
        );

    \I__5753\ : InMux
    port map (
            O => \N__30278\,
            I => \N__30270\
        );

    \I__5752\ : InMux
    port map (
            O => \N__30275\,
            I => \N__30270\
        );

    \I__5751\ : LocalMux
    port map (
            O => \N__30270\,
            I => \N__30267\
        );

    \I__5750\ : Odrv4
    port map (
            O => \N__30267\,
            I => \nx.n2193\
        );

    \I__5749\ : InMux
    port map (
            O => \N__30264\,
            I => \N__30261\
        );

    \I__5748\ : LocalMux
    port map (
            O => \N__30261\,
            I => \nx.n2260\
        );

    \I__5747\ : InMux
    port map (
            O => \N__30258\,
            I => \N__30255\
        );

    \I__5746\ : LocalMux
    port map (
            O => \N__30255\,
            I => \nx.n29\
        );

    \I__5745\ : InMux
    port map (
            O => \N__30252\,
            I => \N__30249\
        );

    \I__5744\ : LocalMux
    port map (
            O => \N__30249\,
            I => \N__30246\
        );

    \I__5743\ : Odrv4
    port map (
            O => \N__30246\,
            I => \nx.n28_adj_686\
        );

    \I__5742\ : CascadeMux
    port map (
            O => \N__30243\,
            I => \N__30240\
        );

    \I__5741\ : InMux
    port map (
            O => \N__30240\,
            I => \N__30237\
        );

    \I__5740\ : LocalMux
    port map (
            O => \N__30237\,
            I => \nx.n27_adj_691\
        );

    \I__5739\ : InMux
    port map (
            O => \N__30234\,
            I => \N__30231\
        );

    \I__5738\ : LocalMux
    port map (
            O => \N__30231\,
            I => \nx.n30_adj_685\
        );

    \I__5737\ : CascadeMux
    port map (
            O => \N__30228\,
            I => \nx.n2126_cascade_\
        );

    \I__5736\ : CascadeMux
    port map (
            O => \N__30225\,
            I => \nx.n2199_cascade_\
        );

    \I__5735\ : CascadeMux
    port map (
            O => \N__30222\,
            I => \nx.n31_cascade_\
        );

    \I__5734\ : InMux
    port map (
            O => \N__30219\,
            I => \N__30216\
        );

    \I__5733\ : LocalMux
    port map (
            O => \N__30216\,
            I => \nx.n28_adj_692\
        );

    \I__5732\ : InMux
    port map (
            O => \N__30213\,
            I => \N__30210\
        );

    \I__5731\ : LocalMux
    port map (
            O => \N__30210\,
            I => \N__30207\
        );

    \I__5730\ : Span4Mux_h
    port map (
            O => \N__30207\,
            I => \N__30204\
        );

    \I__5729\ : Odrv4
    port map (
            O => \N__30204\,
            I => \nx.n2264\
        );

    \I__5728\ : InMux
    port map (
            O => \N__30201\,
            I => \nx.n10893\
        );

    \I__5727\ : InMux
    port map (
            O => \N__30198\,
            I => \nx.n10894\
        );

    \I__5726\ : InMux
    port map (
            O => \N__30195\,
            I => \nx.n10895\
        );

    \I__5725\ : InMux
    port map (
            O => \N__30192\,
            I => \bfn_11_27_0_\
        );

    \I__5724\ : InMux
    port map (
            O => \N__30189\,
            I => \nx.n10897\
        );

    \I__5723\ : InMux
    port map (
            O => \N__30186\,
            I => \nx.n10898\
        );

    \I__5722\ : InMux
    port map (
            O => \N__30183\,
            I => \N__30180\
        );

    \I__5721\ : LocalMux
    port map (
            O => \N__30180\,
            I => \nx.n2263\
        );

    \I__5720\ : CascadeMux
    port map (
            O => \N__30177\,
            I => \nx.n2196_cascade_\
        );

    \I__5719\ : InMux
    port map (
            O => \N__30174\,
            I => \nx.n10884\
        );

    \I__5718\ : InMux
    port map (
            O => \N__30171\,
            I => \nx.n10885\
        );

    \I__5717\ : InMux
    port map (
            O => \N__30168\,
            I => \nx.n10886\
        );

    \I__5716\ : InMux
    port map (
            O => \N__30165\,
            I => \nx.n10887\
        );

    \I__5715\ : InMux
    port map (
            O => \N__30162\,
            I => \bfn_11_26_0_\
        );

    \I__5714\ : InMux
    port map (
            O => \N__30159\,
            I => \nx.n10889\
        );

    \I__5713\ : InMux
    port map (
            O => \N__30156\,
            I => \nx.n10890\
        );

    \I__5712\ : InMux
    port map (
            O => \N__30153\,
            I => \nx.n10891\
        );

    \I__5711\ : InMux
    port map (
            O => \N__30150\,
            I => \nx.n10892\
        );

    \I__5710\ : InMux
    port map (
            O => \N__30147\,
            I => \N__30143\
        );

    \I__5709\ : InMux
    port map (
            O => \N__30146\,
            I => \N__30139\
        );

    \I__5708\ : LocalMux
    port map (
            O => \N__30143\,
            I => \N__30136\
        );

    \I__5707\ : InMux
    port map (
            O => \N__30142\,
            I => \N__30133\
        );

    \I__5706\ : LocalMux
    port map (
            O => \N__30139\,
            I => \N__30129\
        );

    \I__5705\ : Span4Mux_h
    port map (
            O => \N__30136\,
            I => \N__30124\
        );

    \I__5704\ : LocalMux
    port map (
            O => \N__30133\,
            I => \N__30124\
        );

    \I__5703\ : InMux
    port map (
            O => \N__30132\,
            I => \N__30120\
        );

    \I__5702\ : Span4Mux_h
    port map (
            O => \N__30129\,
            I => \N__30115\
        );

    \I__5701\ : Span4Mux_v
    port map (
            O => \N__30124\,
            I => \N__30115\
        );

    \I__5700\ : InMux
    port map (
            O => \N__30123\,
            I => \N__30112\
        );

    \I__5699\ : LocalMux
    port map (
            O => \N__30120\,
            I => \N__30109\
        );

    \I__5698\ : Span4Mux_h
    port map (
            O => \N__30115\,
            I => \N__30106\
        );

    \I__5697\ : LocalMux
    port map (
            O => \N__30112\,
            I => \N__30101\
        );

    \I__5696\ : Span4Mux_h
    port map (
            O => \N__30109\,
            I => \N__30101\
        );

    \I__5695\ : Odrv4
    port map (
            O => \N__30106\,
            I => \nx.bit_ctr_8\
        );

    \I__5694\ : Odrv4
    port map (
            O => \N__30101\,
            I => \nx.bit_ctr_8\
        );

    \I__5693\ : CascadeMux
    port map (
            O => \N__30096\,
            I => \nx.n2698_cascade_\
        );

    \I__5692\ : InMux
    port map (
            O => \N__30093\,
            I => \N__30090\
        );

    \I__5691\ : LocalMux
    port map (
            O => \N__30090\,
            I => \nx.n30\
        );

    \I__5690\ : CascadeMux
    port map (
            O => \N__30087\,
            I => \N__30084\
        );

    \I__5689\ : InMux
    port map (
            O => \N__30084\,
            I => \N__30080\
        );

    \I__5688\ : CascadeMux
    port map (
            O => \N__30083\,
            I => \N__30077\
        );

    \I__5687\ : LocalMux
    port map (
            O => \N__30080\,
            I => \N__30074\
        );

    \I__5686\ : InMux
    port map (
            O => \N__30077\,
            I => \N__30071\
        );

    \I__5685\ : Odrv4
    port map (
            O => \N__30074\,
            I => \nx.n2693\
        );

    \I__5684\ : LocalMux
    port map (
            O => \N__30071\,
            I => \nx.n2693\
        );

    \I__5683\ : CascadeMux
    port map (
            O => \N__30066\,
            I => \N__30063\
        );

    \I__5682\ : InMux
    port map (
            O => \N__30063\,
            I => \N__30059\
        );

    \I__5681\ : CascadeMux
    port map (
            O => \N__30062\,
            I => \N__30056\
        );

    \I__5680\ : LocalMux
    port map (
            O => \N__30059\,
            I => \N__30052\
        );

    \I__5679\ : InMux
    port map (
            O => \N__30056\,
            I => \N__30049\
        );

    \I__5678\ : InMux
    port map (
            O => \N__30055\,
            I => \N__30046\
        );

    \I__5677\ : Odrv4
    port map (
            O => \N__30052\,
            I => \nx.n2694\
        );

    \I__5676\ : LocalMux
    port map (
            O => \N__30049\,
            I => \nx.n2694\
        );

    \I__5675\ : LocalMux
    port map (
            O => \N__30046\,
            I => \nx.n2694\
        );

    \I__5674\ : CascadeMux
    port map (
            O => \N__30039\,
            I => \nx.n2693_cascade_\
        );

    \I__5673\ : CascadeMux
    port map (
            O => \N__30036\,
            I => \N__30032\
        );

    \I__5672\ : InMux
    port map (
            O => \N__30035\,
            I => \N__30028\
        );

    \I__5671\ : InMux
    port map (
            O => \N__30032\,
            I => \N__30025\
        );

    \I__5670\ : InMux
    port map (
            O => \N__30031\,
            I => \N__30022\
        );

    \I__5669\ : LocalMux
    port map (
            O => \N__30028\,
            I => \nx.n2696\
        );

    \I__5668\ : LocalMux
    port map (
            O => \N__30025\,
            I => \nx.n2696\
        );

    \I__5667\ : LocalMux
    port map (
            O => \N__30022\,
            I => \nx.n2696\
        );

    \I__5666\ : InMux
    port map (
            O => \N__30015\,
            I => \N__30012\
        );

    \I__5665\ : LocalMux
    port map (
            O => \N__30012\,
            I => \nx.n37_adj_677\
        );

    \I__5664\ : CascadeMux
    port map (
            O => \N__30009\,
            I => \N__30006\
        );

    \I__5663\ : InMux
    port map (
            O => \N__30006\,
            I => \N__30003\
        );

    \I__5662\ : LocalMux
    port map (
            O => \N__30003\,
            I => \N__30000\
        );

    \I__5661\ : Span4Mux_h
    port map (
            O => \N__30000\,
            I => \N__29996\
        );

    \I__5660\ : CascadeMux
    port map (
            O => \N__29999\,
            I => \N__29992\
        );

    \I__5659\ : Span4Mux_v
    port map (
            O => \N__29996\,
            I => \N__29989\
        );

    \I__5658\ : InMux
    port map (
            O => \N__29995\,
            I => \N__29986\
        );

    \I__5657\ : InMux
    port map (
            O => \N__29992\,
            I => \N__29983\
        );

    \I__5656\ : Odrv4
    port map (
            O => \N__29989\,
            I => \nx.n2709\
        );

    \I__5655\ : LocalMux
    port map (
            O => \N__29986\,
            I => \nx.n2709\
        );

    \I__5654\ : LocalMux
    port map (
            O => \N__29983\,
            I => \nx.n2709\
        );

    \I__5653\ : InMux
    port map (
            O => \N__29976\,
            I => \bfn_11_25_0_\
        );

    \I__5652\ : InMux
    port map (
            O => \N__29973\,
            I => \nx.n10881\
        );

    \I__5651\ : InMux
    port map (
            O => \N__29970\,
            I => \nx.n10882\
        );

    \I__5650\ : InMux
    port map (
            O => \N__29967\,
            I => \nx.n10883\
        );

    \I__5649\ : CascadeMux
    port map (
            O => \N__29964\,
            I => \nx.n2706_cascade_\
        );

    \I__5648\ : InMux
    port map (
            O => \N__29961\,
            I => \N__29958\
        );

    \I__5647\ : LocalMux
    port map (
            O => \N__29958\,
            I => \nx.n40_adj_687\
        );

    \I__5646\ : InMux
    port map (
            O => \N__29955\,
            I => \N__29952\
        );

    \I__5645\ : LocalMux
    port map (
            O => \N__29952\,
            I => \N__29949\
        );

    \I__5644\ : Odrv4
    port map (
            O => \N__29949\,
            I => \nx.n2755\
        );

    \I__5643\ : CascadeMux
    port map (
            O => \N__29946\,
            I => \N__29943\
        );

    \I__5642\ : InMux
    port map (
            O => \N__29943\,
            I => \N__29939\
        );

    \I__5641\ : InMux
    port map (
            O => \N__29942\,
            I => \N__29935\
        );

    \I__5640\ : LocalMux
    port map (
            O => \N__29939\,
            I => \N__29932\
        );

    \I__5639\ : InMux
    port map (
            O => \N__29938\,
            I => \N__29929\
        );

    \I__5638\ : LocalMux
    port map (
            O => \N__29935\,
            I => \nx.n2787\
        );

    \I__5637\ : Odrv4
    port map (
            O => \N__29932\,
            I => \nx.n2787\
        );

    \I__5636\ : LocalMux
    port map (
            O => \N__29929\,
            I => \nx.n2787\
        );

    \I__5635\ : CascadeMux
    port map (
            O => \N__29922\,
            I => \N__29918\
        );

    \I__5634\ : InMux
    port map (
            O => \N__29921\,
            I => \N__29915\
        );

    \I__5633\ : InMux
    port map (
            O => \N__29918\,
            I => \N__29912\
        );

    \I__5632\ : LocalMux
    port map (
            O => \N__29915\,
            I => \nx.n2699\
        );

    \I__5631\ : LocalMux
    port map (
            O => \N__29912\,
            I => \nx.n2699\
        );

    \I__5630\ : InMux
    port map (
            O => \N__29907\,
            I => \N__29904\
        );

    \I__5629\ : LocalMux
    port map (
            O => \N__29904\,
            I => \nx.n2766\
        );

    \I__5628\ : CascadeMux
    port map (
            O => \N__29901\,
            I => \nx.n2699_cascade_\
        );

    \I__5627\ : CascadeMux
    port map (
            O => \N__29898\,
            I => \N__29895\
        );

    \I__5626\ : InMux
    port map (
            O => \N__29895\,
            I => \N__29891\
        );

    \I__5625\ : CascadeMux
    port map (
            O => \N__29894\,
            I => \N__29888\
        );

    \I__5624\ : LocalMux
    port map (
            O => \N__29891\,
            I => \N__29885\
        );

    \I__5623\ : InMux
    port map (
            O => \N__29888\,
            I => \N__29882\
        );

    \I__5622\ : Odrv4
    port map (
            O => \N__29885\,
            I => \nx.n2701\
        );

    \I__5621\ : LocalMux
    port map (
            O => \N__29882\,
            I => \nx.n2701\
        );

    \I__5620\ : CascadeMux
    port map (
            O => \N__29877\,
            I => \nx.n2701_cascade_\
        );

    \I__5619\ : CascadeMux
    port map (
            O => \N__29874\,
            I => \N__29871\
        );

    \I__5618\ : InMux
    port map (
            O => \N__29871\,
            I => \N__29868\
        );

    \I__5617\ : LocalMux
    port map (
            O => \N__29868\,
            I => \N__29865\
        );

    \I__5616\ : Odrv4
    port map (
            O => \N__29865\,
            I => \nx.n42_adj_683\
        );

    \I__5615\ : CascadeMux
    port map (
            O => \N__29862\,
            I => \N__29859\
        );

    \I__5614\ : InMux
    port map (
            O => \N__29859\,
            I => \N__29855\
        );

    \I__5613\ : CascadeMux
    port map (
            O => \N__29858\,
            I => \N__29852\
        );

    \I__5612\ : LocalMux
    port map (
            O => \N__29855\,
            I => \N__29849\
        );

    \I__5611\ : InMux
    port map (
            O => \N__29852\,
            I => \N__29846\
        );

    \I__5610\ : Odrv4
    port map (
            O => \N__29849\,
            I => \nx.n2698\
        );

    \I__5609\ : LocalMux
    port map (
            O => \N__29846\,
            I => \nx.n2698\
        );

    \I__5608\ : InMux
    port map (
            O => \N__29841\,
            I => \N__29838\
        );

    \I__5607\ : LocalMux
    port map (
            O => \N__29838\,
            I => \N__29835\
        );

    \I__5606\ : Odrv4
    port map (
            O => \N__29835\,
            I => \nx.n2765\
        );

    \I__5605\ : InMux
    port map (
            O => \N__29832\,
            I => \N__29829\
        );

    \I__5604\ : LocalMux
    port map (
            O => \N__29829\,
            I => \nx.n41_adj_688\
        );

    \I__5603\ : InMux
    port map (
            O => \N__29826\,
            I => \N__29823\
        );

    \I__5602\ : LocalMux
    port map (
            O => \N__29823\,
            I => \N__29820\
        );

    \I__5601\ : Odrv4
    port map (
            O => \N__29820\,
            I => \nx.n2767\
        );

    \I__5600\ : CascadeMux
    port map (
            O => \N__29817\,
            I => \N__29814\
        );

    \I__5599\ : InMux
    port map (
            O => \N__29814\,
            I => \N__29811\
        );

    \I__5598\ : LocalMux
    port map (
            O => \N__29811\,
            I => \N__29808\
        );

    \I__5597\ : Span4Mux_h
    port map (
            O => \N__29808\,
            I => \N__29805\
        );

    \I__5596\ : Odrv4
    port map (
            O => \N__29805\,
            I => \nx.n2854\
        );

    \I__5595\ : CascadeMux
    port map (
            O => \N__29802\,
            I => \nx.n2886_cascade_\
        );

    \I__5594\ : InMux
    port map (
            O => \N__29799\,
            I => \N__29794\
        );

    \I__5593\ : InMux
    port map (
            O => \N__29798\,
            I => \N__29789\
        );

    \I__5592\ : InMux
    port map (
            O => \N__29797\,
            I => \N__29789\
        );

    \I__5591\ : LocalMux
    port map (
            O => \N__29794\,
            I => \nx.n2985\
        );

    \I__5590\ : LocalMux
    port map (
            O => \N__29789\,
            I => \nx.n2985\
        );

    \I__5589\ : CascadeMux
    port map (
            O => \N__29784\,
            I => \N__29781\
        );

    \I__5588\ : InMux
    port map (
            O => \N__29781\,
            I => \N__29778\
        );

    \I__5587\ : LocalMux
    port map (
            O => \N__29778\,
            I => \nx.n2774\
        );

    \I__5586\ : CascadeMux
    port map (
            O => \N__29775\,
            I => \N__29770\
        );

    \I__5585\ : CascadeMux
    port map (
            O => \N__29774\,
            I => \N__29767\
        );

    \I__5584\ : InMux
    port map (
            O => \N__29773\,
            I => \N__29764\
        );

    \I__5583\ : InMux
    port map (
            O => \N__29770\,
            I => \N__29761\
        );

    \I__5582\ : InMux
    port map (
            O => \N__29767\,
            I => \N__29758\
        );

    \I__5581\ : LocalMux
    port map (
            O => \N__29764\,
            I => \nx.n2800\
        );

    \I__5580\ : LocalMux
    port map (
            O => \N__29761\,
            I => \nx.n2800\
        );

    \I__5579\ : LocalMux
    port map (
            O => \N__29758\,
            I => \nx.n2800\
        );

    \I__5578\ : InMux
    port map (
            O => \N__29751\,
            I => \N__29748\
        );

    \I__5577\ : LocalMux
    port map (
            O => \N__29748\,
            I => \N__29745\
        );

    \I__5576\ : Odrv4
    port map (
            O => \N__29745\,
            I => \nx.n2867\
        );

    \I__5575\ : CascadeMux
    port map (
            O => \N__29742\,
            I => \N__29738\
        );

    \I__5574\ : InMux
    port map (
            O => \N__29741\,
            I => \N__29735\
        );

    \I__5573\ : InMux
    port map (
            O => \N__29738\,
            I => \N__29732\
        );

    \I__5572\ : LocalMux
    port map (
            O => \N__29735\,
            I => \nx.n2706\
        );

    \I__5571\ : LocalMux
    port map (
            O => \N__29732\,
            I => \nx.n2706\
        );

    \I__5570\ : InMux
    port map (
            O => \N__29727\,
            I => \nx.n11074\
        );

    \I__5569\ : InMux
    port map (
            O => \N__29724\,
            I => \N__29720\
        );

    \I__5568\ : InMux
    port map (
            O => \N__29723\,
            I => \N__29717\
        );

    \I__5567\ : LocalMux
    port map (
            O => \N__29720\,
            I => \nx.n2987\
        );

    \I__5566\ : LocalMux
    port map (
            O => \N__29717\,
            I => \nx.n2987\
        );

    \I__5565\ : InMux
    port map (
            O => \N__29712\,
            I => \nx.n11075\
        );

    \I__5564\ : InMux
    port map (
            O => \N__29709\,
            I => \bfn_11_21_0_\
        );

    \I__5563\ : InMux
    port map (
            O => \N__29706\,
            I => \nx.n11077\
        );

    \I__5562\ : CascadeMux
    port map (
            O => \N__29703\,
            I => \N__29698\
        );

    \I__5561\ : CascadeMux
    port map (
            O => \N__29702\,
            I => \N__29695\
        );

    \I__5560\ : CascadeMux
    port map (
            O => \N__29701\,
            I => \N__29692\
        );

    \I__5559\ : InMux
    port map (
            O => \N__29698\,
            I => \N__29666\
        );

    \I__5558\ : InMux
    port map (
            O => \N__29695\,
            I => \N__29661\
        );

    \I__5557\ : InMux
    port map (
            O => \N__29692\,
            I => \N__29661\
        );

    \I__5556\ : CascadeMux
    port map (
            O => \N__29691\,
            I => \N__29658\
        );

    \I__5555\ : CascadeMux
    port map (
            O => \N__29690\,
            I => \N__29655\
        );

    \I__5554\ : CascadeMux
    port map (
            O => \N__29689\,
            I => \N__29652\
        );

    \I__5553\ : CascadeMux
    port map (
            O => \N__29688\,
            I => \N__29649\
        );

    \I__5552\ : CascadeMux
    port map (
            O => \N__29687\,
            I => \N__29646\
        );

    \I__5551\ : CascadeMux
    port map (
            O => \N__29686\,
            I => \N__29643\
        );

    \I__5550\ : CascadeMux
    port map (
            O => \N__29685\,
            I => \N__29640\
        );

    \I__5549\ : CascadeMux
    port map (
            O => \N__29684\,
            I => \N__29637\
        );

    \I__5548\ : CascadeMux
    port map (
            O => \N__29683\,
            I => \N__29634\
        );

    \I__5547\ : CascadeMux
    port map (
            O => \N__29682\,
            I => \N__29631\
        );

    \I__5546\ : CascadeMux
    port map (
            O => \N__29681\,
            I => \N__29628\
        );

    \I__5545\ : CascadeMux
    port map (
            O => \N__29680\,
            I => \N__29625\
        );

    \I__5544\ : CascadeMux
    port map (
            O => \N__29679\,
            I => \N__29622\
        );

    \I__5543\ : CascadeMux
    port map (
            O => \N__29678\,
            I => \N__29619\
        );

    \I__5542\ : CascadeMux
    port map (
            O => \N__29677\,
            I => \N__29616\
        );

    \I__5541\ : CascadeMux
    port map (
            O => \N__29676\,
            I => \N__29613\
        );

    \I__5540\ : CascadeMux
    port map (
            O => \N__29675\,
            I => \N__29610\
        );

    \I__5539\ : CascadeMux
    port map (
            O => \N__29674\,
            I => \N__29607\
        );

    \I__5538\ : CascadeMux
    port map (
            O => \N__29673\,
            I => \N__29604\
        );

    \I__5537\ : CascadeMux
    port map (
            O => \N__29672\,
            I => \N__29601\
        );

    \I__5536\ : CascadeMux
    port map (
            O => \N__29671\,
            I => \N__29598\
        );

    \I__5535\ : CascadeMux
    port map (
            O => \N__29670\,
            I => \N__29595\
        );

    \I__5534\ : InMux
    port map (
            O => \N__29669\,
            I => \N__29592\
        );

    \I__5533\ : LocalMux
    port map (
            O => \N__29666\,
            I => \N__29587\
        );

    \I__5532\ : LocalMux
    port map (
            O => \N__29661\,
            I => \N__29587\
        );

    \I__5531\ : InMux
    port map (
            O => \N__29658\,
            I => \N__29578\
        );

    \I__5530\ : InMux
    port map (
            O => \N__29655\,
            I => \N__29578\
        );

    \I__5529\ : InMux
    port map (
            O => \N__29652\,
            I => \N__29578\
        );

    \I__5528\ : InMux
    port map (
            O => \N__29649\,
            I => \N__29578\
        );

    \I__5527\ : InMux
    port map (
            O => \N__29646\,
            I => \N__29569\
        );

    \I__5526\ : InMux
    port map (
            O => \N__29643\,
            I => \N__29569\
        );

    \I__5525\ : InMux
    port map (
            O => \N__29640\,
            I => \N__29569\
        );

    \I__5524\ : InMux
    port map (
            O => \N__29637\,
            I => \N__29569\
        );

    \I__5523\ : InMux
    port map (
            O => \N__29634\,
            I => \N__29560\
        );

    \I__5522\ : InMux
    port map (
            O => \N__29631\,
            I => \N__29560\
        );

    \I__5521\ : InMux
    port map (
            O => \N__29628\,
            I => \N__29560\
        );

    \I__5520\ : InMux
    port map (
            O => \N__29625\,
            I => \N__29560\
        );

    \I__5519\ : InMux
    port map (
            O => \N__29622\,
            I => \N__29551\
        );

    \I__5518\ : InMux
    port map (
            O => \N__29619\,
            I => \N__29551\
        );

    \I__5517\ : InMux
    port map (
            O => \N__29616\,
            I => \N__29551\
        );

    \I__5516\ : InMux
    port map (
            O => \N__29613\,
            I => \N__29551\
        );

    \I__5515\ : InMux
    port map (
            O => \N__29610\,
            I => \N__29544\
        );

    \I__5514\ : InMux
    port map (
            O => \N__29607\,
            I => \N__29544\
        );

    \I__5513\ : InMux
    port map (
            O => \N__29604\,
            I => \N__29544\
        );

    \I__5512\ : InMux
    port map (
            O => \N__29601\,
            I => \N__29537\
        );

    \I__5511\ : InMux
    port map (
            O => \N__29598\,
            I => \N__29537\
        );

    \I__5510\ : InMux
    port map (
            O => \N__29595\,
            I => \N__29537\
        );

    \I__5509\ : LocalMux
    port map (
            O => \N__29592\,
            I => \N__29534\
        );

    \I__5508\ : Odrv4
    port map (
            O => \N__29587\,
            I => \nx.n3017\
        );

    \I__5507\ : LocalMux
    port map (
            O => \N__29578\,
            I => \nx.n3017\
        );

    \I__5506\ : LocalMux
    port map (
            O => \N__29569\,
            I => \nx.n3017\
        );

    \I__5505\ : LocalMux
    port map (
            O => \N__29560\,
            I => \nx.n3017\
        );

    \I__5504\ : LocalMux
    port map (
            O => \N__29551\,
            I => \nx.n3017\
        );

    \I__5503\ : LocalMux
    port map (
            O => \N__29544\,
            I => \nx.n3017\
        );

    \I__5502\ : LocalMux
    port map (
            O => \N__29537\,
            I => \nx.n3017\
        );

    \I__5501\ : Odrv4
    port map (
            O => \N__29534\,
            I => \nx.n3017\
        );

    \I__5500\ : InMux
    port map (
            O => \N__29517\,
            I => \nx.n11078\
        );

    \I__5499\ : InMux
    port map (
            O => \N__29514\,
            I => \N__29511\
        );

    \I__5498\ : LocalMux
    port map (
            O => \N__29511\,
            I => \N__29508\
        );

    \I__5497\ : Odrv4
    port map (
            O => \N__29508\,
            I => \nx.n40_adj_670\
        );

    \I__5496\ : InMux
    port map (
            O => \N__29505\,
            I => \N__29501\
        );

    \I__5495\ : InMux
    port map (
            O => \N__29504\,
            I => \N__29498\
        );

    \I__5494\ : LocalMux
    port map (
            O => \N__29501\,
            I => \N__29492\
        );

    \I__5493\ : LocalMux
    port map (
            O => \N__29498\,
            I => \N__29492\
        );

    \I__5492\ : InMux
    port map (
            O => \N__29497\,
            I => \N__29489\
        );

    \I__5491\ : Odrv4
    port map (
            O => \N__29492\,
            I => \nx.n2996\
        );

    \I__5490\ : LocalMux
    port map (
            O => \N__29489\,
            I => \nx.n2996\
        );

    \I__5489\ : InMux
    port map (
            O => \N__29484\,
            I => \N__29481\
        );

    \I__5488\ : LocalMux
    port map (
            O => \N__29481\,
            I => \nx.n41_adj_736\
        );

    \I__5487\ : InMux
    port map (
            O => \N__29478\,
            I => \N__29473\
        );

    \I__5486\ : InMux
    port map (
            O => \N__29477\,
            I => \N__29470\
        );

    \I__5485\ : InMux
    port map (
            O => \N__29476\,
            I => \N__29467\
        );

    \I__5484\ : LocalMux
    port map (
            O => \N__29473\,
            I => \N__29462\
        );

    \I__5483\ : LocalMux
    port map (
            O => \N__29470\,
            I => \N__29462\
        );

    \I__5482\ : LocalMux
    port map (
            O => \N__29467\,
            I => \N__29459\
        );

    \I__5481\ : Span4Mux_v
    port map (
            O => \N__29462\,
            I => \N__29454\
        );

    \I__5480\ : Span4Mux_h
    port map (
            O => \N__29459\,
            I => \N__29454\
        );

    \I__5479\ : Odrv4
    port map (
            O => \N__29454\,
            I => \nx.n2998\
        );

    \I__5478\ : InMux
    port map (
            O => \N__29451\,
            I => \nx.n11065\
        );

    \I__5477\ : InMux
    port map (
            O => \N__29448\,
            I => \nx.n11066\
        );

    \I__5476\ : InMux
    port map (
            O => \N__29445\,
            I => \nx.n11067\
        );

    \I__5475\ : InMux
    port map (
            O => \N__29442\,
            I => \bfn_11_20_0_\
        );

    \I__5474\ : InMux
    port map (
            O => \N__29439\,
            I => \nx.n11069\
        );

    \I__5473\ : InMux
    port map (
            O => \N__29436\,
            I => \nx.n11070\
        );

    \I__5472\ : InMux
    port map (
            O => \N__29433\,
            I => \nx.n11071\
        );

    \I__5471\ : InMux
    port map (
            O => \N__29430\,
            I => \nx.n11072\
        );

    \I__5470\ : InMux
    port map (
            O => \N__29427\,
            I => \nx.n11073\
        );

    \I__5469\ : InMux
    port map (
            O => \N__29424\,
            I => \nx.n11056\
        );

    \I__5468\ : InMux
    port map (
            O => \N__29421\,
            I => \nx.n11057\
        );

    \I__5467\ : InMux
    port map (
            O => \N__29418\,
            I => \nx.n11058\
        );

    \I__5466\ : InMux
    port map (
            O => \N__29415\,
            I => \nx.n11059\
        );

    \I__5465\ : InMux
    port map (
            O => \N__29412\,
            I => \bfn_11_19_0_\
        );

    \I__5464\ : InMux
    port map (
            O => \N__29409\,
            I => \nx.n11061\
        );

    \I__5463\ : InMux
    port map (
            O => \N__29406\,
            I => \nx.n11062\
        );

    \I__5462\ : InMux
    port map (
            O => \N__29403\,
            I => \nx.n11063\
        );

    \I__5461\ : InMux
    port map (
            O => \N__29400\,
            I => \nx.n11064\
        );

    \I__5460\ : CascadeMux
    port map (
            O => \N__29397\,
            I => \nx.n42_adj_739_cascade_\
        );

    \I__5459\ : CascadeMux
    port map (
            O => \N__29394\,
            I => \nx.n32_adj_740_cascade_\
        );

    \I__5458\ : InMux
    port map (
            O => \N__29391\,
            I => \N__29388\
        );

    \I__5457\ : LocalMux
    port map (
            O => \N__29388\,
            I => \N__29385\
        );

    \I__5456\ : Span4Mux_h
    port map (
            O => \N__29385\,
            I => \N__29382\
        );

    \I__5455\ : Odrv4
    port map (
            O => \N__29382\,
            I => \nx.n44_adj_741\
        );

    \I__5454\ : InMux
    port map (
            O => \N__29379\,
            I => \N__29376\
        );

    \I__5453\ : LocalMux
    port map (
            O => \N__29376\,
            I => \nx.n50_adj_742\
        );

    \I__5452\ : InMux
    port map (
            O => \N__29373\,
            I => \N__29370\
        );

    \I__5451\ : LocalMux
    port map (
            O => \N__29370\,
            I => \N__29367\
        );

    \I__5450\ : Span4Mux_v
    port map (
            O => \N__29367\,
            I => \N__29364\
        );

    \I__5449\ : Span4Mux_h
    port map (
            O => \N__29364\,
            I => \N__29361\
        );

    \I__5448\ : Odrv4
    port map (
            O => \N__29361\,
            I => \nx.n47\
        );

    \I__5447\ : CascadeMux
    port map (
            O => \N__29358\,
            I => \nx.n49_cascade_\
        );

    \I__5446\ : InMux
    port map (
            O => \N__29355\,
            I => \N__29352\
        );

    \I__5445\ : LocalMux
    port map (
            O => \N__29352\,
            I => \nx.n48\
        );

    \I__5444\ : CascadeMux
    port map (
            O => \N__29349\,
            I => \nx.n3116_cascade_\
        );

    \I__5443\ : InMux
    port map (
            O => \N__29346\,
            I => \N__29342\
        );

    \I__5442\ : InMux
    port map (
            O => \N__29345\,
            I => \N__29339\
        );

    \I__5441\ : LocalMux
    port map (
            O => \N__29342\,
            I => \N__29333\
        );

    \I__5440\ : LocalMux
    port map (
            O => \N__29339\,
            I => \N__29333\
        );

    \I__5439\ : InMux
    port map (
            O => \N__29338\,
            I => \N__29330\
        );

    \I__5438\ : Span4Mux_v
    port map (
            O => \N__29333\,
            I => \N__29325\
        );

    \I__5437\ : LocalMux
    port map (
            O => \N__29330\,
            I => \N__29322\
        );

    \I__5436\ : InMux
    port map (
            O => \N__29329\,
            I => \N__29319\
        );

    \I__5435\ : InMux
    port map (
            O => \N__29328\,
            I => \N__29316\
        );

    \I__5434\ : Span4Mux_h
    port map (
            O => \N__29325\,
            I => \N__29313\
        );

    \I__5433\ : Span4Mux_h
    port map (
            O => \N__29322\,
            I => \N__29310\
        );

    \I__5432\ : LocalMux
    port map (
            O => \N__29319\,
            I => \nx.bit_ctr_5\
        );

    \I__5431\ : LocalMux
    port map (
            O => \N__29316\,
            I => \nx.bit_ctr_5\
        );

    \I__5430\ : Odrv4
    port map (
            O => \N__29313\,
            I => \nx.bit_ctr_5\
        );

    \I__5429\ : Odrv4
    port map (
            O => \N__29310\,
            I => \nx.bit_ctr_5\
        );

    \I__5428\ : InMux
    port map (
            O => \N__29301\,
            I => \bfn_11_18_0_\
        );

    \I__5427\ : InMux
    port map (
            O => \N__29298\,
            I => \N__29294\
        );

    \I__5426\ : InMux
    port map (
            O => \N__29297\,
            I => \N__29291\
        );

    \I__5425\ : LocalMux
    port map (
            O => \N__29294\,
            I => \N__29286\
        );

    \I__5424\ : LocalMux
    port map (
            O => \N__29291\,
            I => \N__29286\
        );

    \I__5423\ : Span4Mux_h
    port map (
            O => \N__29286\,
            I => \N__29283\
        );

    \I__5422\ : Span4Mux_h
    port map (
            O => \N__29283\,
            I => \N__29280\
        );

    \I__5421\ : Odrv4
    port map (
            O => \N__29280\,
            I => \nx.n3009\
        );

    \I__5420\ : CascadeMux
    port map (
            O => \N__29277\,
            I => \N__29273\
        );

    \I__5419\ : CascadeMux
    port map (
            O => \N__29276\,
            I => \N__29270\
        );

    \I__5418\ : InMux
    port map (
            O => \N__29273\,
            I => \N__29267\
        );

    \I__5417\ : InMux
    port map (
            O => \N__29270\,
            I => \N__29264\
        );

    \I__5416\ : LocalMux
    port map (
            O => \N__29267\,
            I => \N__29259\
        );

    \I__5415\ : LocalMux
    port map (
            O => \N__29264\,
            I => \N__29259\
        );

    \I__5414\ : Span4Mux_h
    port map (
            O => \N__29259\,
            I => \N__29256\
        );

    \I__5413\ : Odrv4
    port map (
            O => \N__29256\,
            I => \nx.n13600\
        );

    \I__5412\ : InMux
    port map (
            O => \N__29253\,
            I => \nx.n11053\
        );

    \I__5411\ : InMux
    port map (
            O => \N__29250\,
            I => \N__29245\
        );

    \I__5410\ : InMux
    port map (
            O => \N__29249\,
            I => \N__29242\
        );

    \I__5409\ : InMux
    port map (
            O => \N__29248\,
            I => \N__29239\
        );

    \I__5408\ : LocalMux
    port map (
            O => \N__29245\,
            I => \nx.n3008\
        );

    \I__5407\ : LocalMux
    port map (
            O => \N__29242\,
            I => \nx.n3008\
        );

    \I__5406\ : LocalMux
    port map (
            O => \N__29239\,
            I => \nx.n3008\
        );

    \I__5405\ : InMux
    port map (
            O => \N__29232\,
            I => \nx.n11054\
        );

    \I__5404\ : InMux
    port map (
            O => \N__29229\,
            I => \N__29224\
        );

    \I__5403\ : InMux
    port map (
            O => \N__29228\,
            I => \N__29221\
        );

    \I__5402\ : InMux
    port map (
            O => \N__29227\,
            I => \N__29218\
        );

    \I__5401\ : LocalMux
    port map (
            O => \N__29224\,
            I => \nx.n3007\
        );

    \I__5400\ : LocalMux
    port map (
            O => \N__29221\,
            I => \nx.n3007\
        );

    \I__5399\ : LocalMux
    port map (
            O => \N__29218\,
            I => \nx.n3007\
        );

    \I__5398\ : InMux
    port map (
            O => \N__29211\,
            I => \nx.n11055\
        );

    \I__5397\ : CascadeMux
    port map (
            O => \N__29208\,
            I => \nx.n2193_cascade_\
        );

    \I__5396\ : InMux
    port map (
            O => \N__29205\,
            I => \N__29201\
        );

    \I__5395\ : CascadeMux
    port map (
            O => \N__29204\,
            I => \N__29197\
        );

    \I__5394\ : LocalMux
    port map (
            O => \N__29201\,
            I => \N__29194\
        );

    \I__5393\ : InMux
    port map (
            O => \N__29200\,
            I => \N__29191\
        );

    \I__5392\ : InMux
    port map (
            O => \N__29197\,
            I => \N__29188\
        );

    \I__5391\ : Span4Mux_v
    port map (
            O => \N__29194\,
            I => \N__29181\
        );

    \I__5390\ : LocalMux
    port map (
            O => \N__29191\,
            I => \N__29181\
        );

    \I__5389\ : LocalMux
    port map (
            O => \N__29188\,
            I => \N__29181\
        );

    \I__5388\ : Span4Mux_h
    port map (
            O => \N__29181\,
            I => \N__29178\
        );

    \I__5387\ : Odrv4
    port map (
            O => \N__29178\,
            I => \nx.n2009\
        );

    \I__5386\ : CascadeMux
    port map (
            O => \N__29175\,
            I => \N__29172\
        );

    \I__5385\ : InMux
    port map (
            O => \N__29172\,
            I => \N__29169\
        );

    \I__5384\ : LocalMux
    port map (
            O => \N__29169\,
            I => \N__29166\
        );

    \I__5383\ : Span4Mux_v
    port map (
            O => \N__29166\,
            I => \N__29163\
        );

    \I__5382\ : Odrv4
    port map (
            O => \N__29163\,
            I => \nx.n2076\
        );

    \I__5381\ : CascadeMux
    port map (
            O => \N__29160\,
            I => \nx.n2108_cascade_\
        );

    \I__5380\ : CascadeMux
    port map (
            O => \N__29157\,
            I => \N__29154\
        );

    \I__5379\ : InMux
    port map (
            O => \N__29154\,
            I => \N__29150\
        );

    \I__5378\ : InMux
    port map (
            O => \N__29153\,
            I => \N__29147\
        );

    \I__5377\ : LocalMux
    port map (
            O => \N__29150\,
            I => \N__29144\
        );

    \I__5376\ : LocalMux
    port map (
            O => \N__29147\,
            I => \N__29140\
        );

    \I__5375\ : Span4Mux_h
    port map (
            O => \N__29144\,
            I => \N__29137\
        );

    \I__5374\ : InMux
    port map (
            O => \N__29143\,
            I => \N__29134\
        );

    \I__5373\ : Odrv4
    port map (
            O => \N__29140\,
            I => \nx.n1996\
        );

    \I__5372\ : Odrv4
    port map (
            O => \N__29137\,
            I => \nx.n1996\
        );

    \I__5371\ : LocalMux
    port map (
            O => \N__29134\,
            I => \nx.n1996\
        );

    \I__5370\ : CascadeMux
    port map (
            O => \N__29127\,
            I => \N__29117\
        );

    \I__5369\ : CascadeMux
    port map (
            O => \N__29126\,
            I => \N__29113\
        );

    \I__5368\ : CascadeMux
    port map (
            O => \N__29125\,
            I => \N__29108\
        );

    \I__5367\ : CascadeMux
    port map (
            O => \N__29124\,
            I => \N__29102\
        );

    \I__5366\ : CascadeMux
    port map (
            O => \N__29123\,
            I => \N__29099\
        );

    \I__5365\ : CascadeMux
    port map (
            O => \N__29122\,
            I => \N__29096\
        );

    \I__5364\ : InMux
    port map (
            O => \N__29121\,
            I => \N__29089\
        );

    \I__5363\ : InMux
    port map (
            O => \N__29120\,
            I => \N__29089\
        );

    \I__5362\ : InMux
    port map (
            O => \N__29117\,
            I => \N__29084\
        );

    \I__5361\ : InMux
    port map (
            O => \N__29116\,
            I => \N__29084\
        );

    \I__5360\ : InMux
    port map (
            O => \N__29113\,
            I => \N__29075\
        );

    \I__5359\ : InMux
    port map (
            O => \N__29112\,
            I => \N__29075\
        );

    \I__5358\ : InMux
    port map (
            O => \N__29111\,
            I => \N__29075\
        );

    \I__5357\ : InMux
    port map (
            O => \N__29108\,
            I => \N__29075\
        );

    \I__5356\ : InMux
    port map (
            O => \N__29107\,
            I => \N__29068\
        );

    \I__5355\ : InMux
    port map (
            O => \N__29106\,
            I => \N__29068\
        );

    \I__5354\ : InMux
    port map (
            O => \N__29105\,
            I => \N__29068\
        );

    \I__5353\ : InMux
    port map (
            O => \N__29102\,
            I => \N__29057\
        );

    \I__5352\ : InMux
    port map (
            O => \N__29099\,
            I => \N__29057\
        );

    \I__5351\ : InMux
    port map (
            O => \N__29096\,
            I => \N__29057\
        );

    \I__5350\ : InMux
    port map (
            O => \N__29095\,
            I => \N__29057\
        );

    \I__5349\ : InMux
    port map (
            O => \N__29094\,
            I => \N__29057\
        );

    \I__5348\ : LocalMux
    port map (
            O => \N__29089\,
            I => \N__29048\
        );

    \I__5347\ : LocalMux
    port map (
            O => \N__29084\,
            I => \N__29048\
        );

    \I__5346\ : LocalMux
    port map (
            O => \N__29075\,
            I => \N__29048\
        );

    \I__5345\ : LocalMux
    port map (
            O => \N__29068\,
            I => \N__29048\
        );

    \I__5344\ : LocalMux
    port map (
            O => \N__29057\,
            I => \nx.n2027\
        );

    \I__5343\ : Odrv4
    port map (
            O => \N__29048\,
            I => \nx.n2027\
        );

    \I__5342\ : InMux
    port map (
            O => \N__29043\,
            I => \N__29040\
        );

    \I__5341\ : LocalMux
    port map (
            O => \N__29040\,
            I => \N__29037\
        );

    \I__5340\ : Odrv4
    port map (
            O => \N__29037\,
            I => \nx.n2063\
        );

    \I__5339\ : InMux
    port map (
            O => \N__29034\,
            I => \N__29031\
        );

    \I__5338\ : LocalMux
    port map (
            O => \N__29031\,
            I => \N__29028\
        );

    \I__5337\ : Odrv4
    port map (
            O => \N__29028\,
            I => \nx.n2075\
        );

    \I__5336\ : CascadeMux
    port map (
            O => \N__29025\,
            I => \N__29022\
        );

    \I__5335\ : InMux
    port map (
            O => \N__29022\,
            I => \N__29017\
        );

    \I__5334\ : InMux
    port map (
            O => \N__29021\,
            I => \N__29014\
        );

    \I__5333\ : CascadeMux
    port map (
            O => \N__29020\,
            I => \N__29011\
        );

    \I__5332\ : LocalMux
    port map (
            O => \N__29017\,
            I => \N__29008\
        );

    \I__5331\ : LocalMux
    port map (
            O => \N__29014\,
            I => \N__29005\
        );

    \I__5330\ : InMux
    port map (
            O => \N__29011\,
            I => \N__29002\
        );

    \I__5329\ : Span4Mux_v
    port map (
            O => \N__29008\,
            I => \N__28995\
        );

    \I__5328\ : Span4Mux_h
    port map (
            O => \N__29005\,
            I => \N__28995\
        );

    \I__5327\ : LocalMux
    port map (
            O => \N__29002\,
            I => \N__28995\
        );

    \I__5326\ : Odrv4
    port map (
            O => \N__28995\,
            I => \nx.n2008\
        );

    \I__5325\ : CascadeMux
    port map (
            O => \N__28992\,
            I => \nx.n2107_cascade_\
        );

    \I__5324\ : InMux
    port map (
            O => \N__28989\,
            I => \N__28986\
        );

    \I__5323\ : LocalMux
    port map (
            O => \N__28986\,
            I => \nx.n24_adj_684\
        );

    \I__5322\ : InMux
    port map (
            O => \N__28983\,
            I => \N__28979\
        );

    \I__5321\ : CascadeMux
    port map (
            O => \N__28982\,
            I => \N__28976\
        );

    \I__5320\ : LocalMux
    port map (
            O => \N__28979\,
            I => \N__28973\
        );

    \I__5319\ : InMux
    port map (
            O => \N__28976\,
            I => \N__28970\
        );

    \I__5318\ : Span4Mux_v
    port map (
            O => \N__28973\,
            I => \N__28965\
        );

    \I__5317\ : LocalMux
    port map (
            O => \N__28970\,
            I => \N__28965\
        );

    \I__5316\ : Span4Mux_h
    port map (
            O => \N__28965\,
            I => \N__28961\
        );

    \I__5315\ : InMux
    port map (
            O => \N__28964\,
            I => \N__28958\
        );

    \I__5314\ : Odrv4
    port map (
            O => \N__28961\,
            I => \nx.n1997\
        );

    \I__5313\ : LocalMux
    port map (
            O => \N__28958\,
            I => \nx.n1997\
        );

    \I__5312\ : CascadeMux
    port map (
            O => \N__28953\,
            I => \N__28950\
        );

    \I__5311\ : InMux
    port map (
            O => \N__28950\,
            I => \N__28947\
        );

    \I__5310\ : LocalMux
    port map (
            O => \N__28947\,
            I => \nx.n2064\
        );

    \I__5309\ : CascadeMux
    port map (
            O => \N__28944\,
            I => \nx.n2096_cascade_\
        );

    \I__5308\ : InMux
    port map (
            O => \N__28941\,
            I => \N__28938\
        );

    \I__5307\ : LocalMux
    port map (
            O => \N__28938\,
            I => \N__28933\
        );

    \I__5306\ : InMux
    port map (
            O => \N__28937\,
            I => \N__28930\
        );

    \I__5305\ : InMux
    port map (
            O => \N__28936\,
            I => \N__28926\
        );

    \I__5304\ : Span4Mux_v
    port map (
            O => \N__28933\,
            I => \N__28921\
        );

    \I__5303\ : LocalMux
    port map (
            O => \N__28930\,
            I => \N__28921\
        );

    \I__5302\ : InMux
    port map (
            O => \N__28929\,
            I => \N__28918\
        );

    \I__5301\ : LocalMux
    port map (
            O => \N__28926\,
            I => \N__28914\
        );

    \I__5300\ : Span4Mux_v
    port map (
            O => \N__28921\,
            I => \N__28909\
        );

    \I__5299\ : LocalMux
    port map (
            O => \N__28918\,
            I => \N__28909\
        );

    \I__5298\ : InMux
    port map (
            O => \N__28917\,
            I => \N__28906\
        );

    \I__5297\ : Span4Mux_h
    port map (
            O => \N__28914\,
            I => \N__28903\
        );

    \I__5296\ : Span4Mux_h
    port map (
            O => \N__28909\,
            I => \N__28900\
        );

    \I__5295\ : LocalMux
    port map (
            O => \N__28906\,
            I => \nx.bit_ctr_15\
        );

    \I__5294\ : Odrv4
    port map (
            O => \N__28903\,
            I => \nx.bit_ctr_15\
        );

    \I__5293\ : Odrv4
    port map (
            O => \N__28900\,
            I => \nx.bit_ctr_15\
        );

    \I__5292\ : InMux
    port map (
            O => \N__28893\,
            I => \N__28890\
        );

    \I__5291\ : LocalMux
    port map (
            O => \N__28890\,
            I => \N__28887\
        );

    \I__5290\ : Span4Mux_v
    port map (
            O => \N__28887\,
            I => \N__28884\
        );

    \I__5289\ : Odrv4
    port map (
            O => \N__28884\,
            I => \nx.n2077\
        );

    \I__5288\ : CascadeMux
    port map (
            O => \N__28881\,
            I => \nx.n2109_cascade_\
        );

    \I__5287\ : CascadeMux
    port map (
            O => \N__28878\,
            I => \nx.n2202_cascade_\
        );

    \I__5286\ : InMux
    port map (
            O => \N__28875\,
            I => \N__28872\
        );

    \I__5285\ : LocalMux
    port map (
            O => \N__28872\,
            I => \nx.n18_adj_682\
        );

    \I__5284\ : CascadeMux
    port map (
            O => \N__28869\,
            I => \N__28864\
        );

    \I__5283\ : InMux
    port map (
            O => \N__28868\,
            I => \N__28859\
        );

    \I__5282\ : InMux
    port map (
            O => \N__28867\,
            I => \N__28859\
        );

    \I__5281\ : InMux
    port map (
            O => \N__28864\,
            I => \N__28856\
        );

    \I__5280\ : LocalMux
    port map (
            O => \N__28859\,
            I => \N__28851\
        );

    \I__5279\ : LocalMux
    port map (
            O => \N__28856\,
            I => \N__28851\
        );

    \I__5278\ : Odrv4
    port map (
            O => \N__28851\,
            I => \nx.n2007\
        );

    \I__5277\ : CascadeMux
    port map (
            O => \N__28848\,
            I => \N__28844\
        );

    \I__5276\ : CascadeMux
    port map (
            O => \N__28847\,
            I => \N__28840\
        );

    \I__5275\ : InMux
    port map (
            O => \N__28844\,
            I => \N__28837\
        );

    \I__5274\ : InMux
    port map (
            O => \N__28843\,
            I => \N__28832\
        );

    \I__5273\ : InMux
    port map (
            O => \N__28840\,
            I => \N__28832\
        );

    \I__5272\ : LocalMux
    port map (
            O => \N__28837\,
            I => \N__28827\
        );

    \I__5271\ : LocalMux
    port map (
            O => \N__28832\,
            I => \N__28827\
        );

    \I__5270\ : Span4Mux_h
    port map (
            O => \N__28827\,
            I => \N__28824\
        );

    \I__5269\ : Odrv4
    port map (
            O => \N__28824\,
            I => \nx.n2003\
        );

    \I__5268\ : CascadeMux
    port map (
            O => \N__28821\,
            I => \N__28816\
        );

    \I__5267\ : InMux
    port map (
            O => \N__28820\,
            I => \N__28813\
        );

    \I__5266\ : InMux
    port map (
            O => \N__28819\,
            I => \N__28810\
        );

    \I__5265\ : InMux
    port map (
            O => \N__28816\,
            I => \N__28807\
        );

    \I__5264\ : LocalMux
    port map (
            O => \N__28813\,
            I => \N__28804\
        );

    \I__5263\ : LocalMux
    port map (
            O => \N__28810\,
            I => \nx.n2000\
        );

    \I__5262\ : LocalMux
    port map (
            O => \N__28807\,
            I => \nx.n2000\
        );

    \I__5261\ : Odrv4
    port map (
            O => \N__28804\,
            I => \nx.n2000\
        );

    \I__5260\ : InMux
    port map (
            O => \N__28797\,
            I => \N__28794\
        );

    \I__5259\ : LocalMux
    port map (
            O => \N__28794\,
            I => \nx.n27\
        );

    \I__5258\ : InMux
    port map (
            O => \N__28791\,
            I => \N__28786\
        );

    \I__5257\ : CascadeMux
    port map (
            O => \N__28790\,
            I => \N__28783\
        );

    \I__5256\ : CascadeMux
    port map (
            O => \N__28789\,
            I => \N__28780\
        );

    \I__5255\ : LocalMux
    port map (
            O => \N__28786\,
            I => \N__28777\
        );

    \I__5254\ : InMux
    port map (
            O => \N__28783\,
            I => \N__28774\
        );

    \I__5253\ : InMux
    port map (
            O => \N__28780\,
            I => \N__28771\
        );

    \I__5252\ : Odrv4
    port map (
            O => \N__28777\,
            I => \nx.n2004\
        );

    \I__5251\ : LocalMux
    port map (
            O => \N__28774\,
            I => \nx.n2004\
        );

    \I__5250\ : LocalMux
    port map (
            O => \N__28771\,
            I => \nx.n2004\
        );

    \I__5249\ : InMux
    port map (
            O => \N__28764\,
            I => \N__28761\
        );

    \I__5248\ : LocalMux
    port map (
            O => \N__28761\,
            I => \nx.n2071\
        );

    \I__5247\ : CascadeMux
    port map (
            O => \N__28758\,
            I => \nx.n2103_cascade_\
        );

    \I__5246\ : CascadeMux
    port map (
            O => \N__28755\,
            I => \N__28751\
        );

    \I__5245\ : InMux
    port map (
            O => \N__28754\,
            I => \N__28748\
        );

    \I__5244\ : InMux
    port map (
            O => \N__28751\,
            I => \N__28745\
        );

    \I__5243\ : LocalMux
    port map (
            O => \N__28748\,
            I => \N__28741\
        );

    \I__5242\ : LocalMux
    port map (
            O => \N__28745\,
            I => \N__28738\
        );

    \I__5241\ : InMux
    port map (
            O => \N__28744\,
            I => \N__28735\
        );

    \I__5240\ : Odrv4
    port map (
            O => \N__28741\,
            I => \nx.n1998\
        );

    \I__5239\ : Odrv4
    port map (
            O => \N__28738\,
            I => \nx.n1998\
        );

    \I__5238\ : LocalMux
    port map (
            O => \N__28735\,
            I => \nx.n1998\
        );

    \I__5237\ : InMux
    port map (
            O => \N__28728\,
            I => \N__28725\
        );

    \I__5236\ : LocalMux
    port map (
            O => \N__28725\,
            I => \nx.n2065\
        );

    \I__5235\ : InMux
    port map (
            O => \N__28722\,
            I => \N__28719\
        );

    \I__5234\ : LocalMux
    port map (
            O => \N__28719\,
            I => \nx.n2073\
        );

    \I__5233\ : CascadeMux
    port map (
            O => \N__28716\,
            I => \N__28713\
        );

    \I__5232\ : InMux
    port map (
            O => \N__28713\,
            I => \N__28708\
        );

    \I__5231\ : InMux
    port map (
            O => \N__28712\,
            I => \N__28705\
        );

    \I__5230\ : CascadeMux
    port map (
            O => \N__28711\,
            I => \N__28702\
        );

    \I__5229\ : LocalMux
    port map (
            O => \N__28708\,
            I => \N__28699\
        );

    \I__5228\ : LocalMux
    port map (
            O => \N__28705\,
            I => \N__28696\
        );

    \I__5227\ : InMux
    port map (
            O => \N__28702\,
            I => \N__28693\
        );

    \I__5226\ : Span4Mux_v
    port map (
            O => \N__28699\,
            I => \N__28686\
        );

    \I__5225\ : Span4Mux_h
    port map (
            O => \N__28696\,
            I => \N__28686\
        );

    \I__5224\ : LocalMux
    port map (
            O => \N__28693\,
            I => \N__28686\
        );

    \I__5223\ : Odrv4
    port map (
            O => \N__28686\,
            I => \nx.n2006\
        );

    \I__5222\ : CascadeMux
    port map (
            O => \N__28683\,
            I => \nx.n2105_cascade_\
        );

    \I__5221\ : InMux
    port map (
            O => \N__28680\,
            I => \N__28676\
        );

    \I__5220\ : CascadeMux
    port map (
            O => \N__28679\,
            I => \N__28673\
        );

    \I__5219\ : LocalMux
    port map (
            O => \N__28676\,
            I => \N__28669\
        );

    \I__5218\ : InMux
    port map (
            O => \N__28673\,
            I => \N__28666\
        );

    \I__5217\ : InMux
    port map (
            O => \N__28672\,
            I => \N__28663\
        );

    \I__5216\ : Span4Mux_v
    port map (
            O => \N__28669\,
            I => \N__28656\
        );

    \I__5215\ : LocalMux
    port map (
            O => \N__28666\,
            I => \N__28656\
        );

    \I__5214\ : LocalMux
    port map (
            O => \N__28663\,
            I => \N__28656\
        );

    \I__5213\ : Odrv4
    port map (
            O => \N__28656\,
            I => \nx.n2005\
        );

    \I__5212\ : CascadeMux
    port map (
            O => \N__28653\,
            I => \N__28650\
        );

    \I__5211\ : InMux
    port map (
            O => \N__28650\,
            I => \N__28647\
        );

    \I__5210\ : LocalMux
    port map (
            O => \N__28647\,
            I => \nx.n2072\
        );

    \I__5209\ : CascadeMux
    port map (
            O => \N__28644\,
            I => \N__28640\
        );

    \I__5208\ : InMux
    port map (
            O => \N__28643\,
            I => \N__28637\
        );

    \I__5207\ : InMux
    port map (
            O => \N__28640\,
            I => \N__28633\
        );

    \I__5206\ : LocalMux
    port map (
            O => \N__28637\,
            I => \N__28630\
        );

    \I__5205\ : InMux
    port map (
            O => \N__28636\,
            I => \N__28627\
        );

    \I__5204\ : LocalMux
    port map (
            O => \N__28633\,
            I => \N__28624\
        );

    \I__5203\ : Odrv4
    port map (
            O => \N__28630\,
            I => \nx.n2002\
        );

    \I__5202\ : LocalMux
    port map (
            O => \N__28627\,
            I => \nx.n2002\
        );

    \I__5201\ : Odrv4
    port map (
            O => \N__28624\,
            I => \nx.n2002\
        );

    \I__5200\ : InMux
    port map (
            O => \N__28617\,
            I => \N__28614\
        );

    \I__5199\ : LocalMux
    port map (
            O => \N__28614\,
            I => \nx.n2069\
        );

    \I__5198\ : InMux
    port map (
            O => \N__28611\,
            I => \nx.n11003\
        );

    \I__5197\ : CascadeMux
    port map (
            O => \N__28608\,
            I => \N__28604\
        );

    \I__5196\ : InMux
    port map (
            O => \N__28607\,
            I => \N__28601\
        );

    \I__5195\ : InMux
    port map (
            O => \N__28604\,
            I => \N__28598\
        );

    \I__5194\ : LocalMux
    port map (
            O => \N__28601\,
            I => \N__28595\
        );

    \I__5193\ : LocalMux
    port map (
            O => \N__28598\,
            I => \nx.n2786\
        );

    \I__5192\ : Odrv12
    port map (
            O => \N__28595\,
            I => \nx.n2786\
        );

    \I__5191\ : CascadeMux
    port map (
            O => \N__28590\,
            I => \N__28587\
        );

    \I__5190\ : InMux
    port map (
            O => \N__28587\,
            I => \N__28584\
        );

    \I__5189\ : LocalMux
    port map (
            O => \N__28584\,
            I => \nx.n2070\
        );

    \I__5188\ : CascadeMux
    port map (
            O => \N__28581\,
            I => \nx.n9709_cascade_\
        );

    \I__5187\ : InMux
    port map (
            O => \N__28578\,
            I => \N__28575\
        );

    \I__5186\ : LocalMux
    port map (
            O => \N__28575\,
            I => \N__28572\
        );

    \I__5185\ : Span4Mux_h
    port map (
            O => \N__28572\,
            I => \N__28569\
        );

    \I__5184\ : Odrv4
    port map (
            O => \N__28569\,
            I => \nx.n25\
        );

    \I__5183\ : CascadeMux
    port map (
            O => \N__28566\,
            I => \nx.n26_adj_681_cascade_\
        );

    \I__5182\ : CascadeMux
    port map (
            O => \N__28563\,
            I => \nx.n2027_cascade_\
        );

    \I__5181\ : InMux
    port map (
            O => \N__28560\,
            I => \N__28557\
        );

    \I__5180\ : LocalMux
    port map (
            O => \N__28557\,
            I => \nx.n2074\
        );

    \I__5179\ : CascadeMux
    port map (
            O => \N__28554\,
            I => \N__28550\
        );

    \I__5178\ : InMux
    port map (
            O => \N__28553\,
            I => \N__28547\
        );

    \I__5177\ : InMux
    port map (
            O => \N__28550\,
            I => \N__28544\
        );

    \I__5176\ : LocalMux
    port map (
            O => \N__28547\,
            I => \N__28541\
        );

    \I__5175\ : LocalMux
    port map (
            O => \N__28544\,
            I => \nx.n2001\
        );

    \I__5174\ : Odrv4
    port map (
            O => \N__28541\,
            I => \nx.n2001\
        );

    \I__5173\ : InMux
    port map (
            O => \N__28536\,
            I => \N__28533\
        );

    \I__5172\ : LocalMux
    port map (
            O => \N__28533\,
            I => \nx.n28_adj_680\
        );

    \I__5171\ : CascadeMux
    port map (
            O => \N__28530\,
            I => \N__28527\
        );

    \I__5170\ : InMux
    port map (
            O => \N__28527\,
            I => \N__28524\
        );

    \I__5169\ : LocalMux
    port map (
            O => \N__28524\,
            I => \N__28519\
        );

    \I__5168\ : InMux
    port map (
            O => \N__28523\,
            I => \N__28514\
        );

    \I__5167\ : InMux
    port map (
            O => \N__28522\,
            I => \N__28514\
        );

    \I__5166\ : Odrv4
    port map (
            O => \N__28519\,
            I => \nx.n1999\
        );

    \I__5165\ : LocalMux
    port map (
            O => \N__28514\,
            I => \nx.n1999\
        );

    \I__5164\ : CascadeMux
    port map (
            O => \N__28509\,
            I => \N__28506\
        );

    \I__5163\ : InMux
    port map (
            O => \N__28506\,
            I => \N__28503\
        );

    \I__5162\ : LocalMux
    port map (
            O => \N__28503\,
            I => \nx.n2066\
        );

    \I__5161\ : InMux
    port map (
            O => \N__28500\,
            I => \N__28497\
        );

    \I__5160\ : LocalMux
    port map (
            O => \N__28497\,
            I => \N__28494\
        );

    \I__5159\ : Odrv4
    port map (
            O => \N__28494\,
            I => \nx.n2763\
        );

    \I__5158\ : InMux
    port map (
            O => \N__28491\,
            I => \nx.n10994\
        );

    \I__5157\ : CascadeMux
    port map (
            O => \N__28488\,
            I => \N__28485\
        );

    \I__5156\ : InMux
    port map (
            O => \N__28485\,
            I => \N__28482\
        );

    \I__5155\ : LocalMux
    port map (
            O => \N__28482\,
            I => \nx.n2762\
        );

    \I__5154\ : InMux
    port map (
            O => \N__28479\,
            I => \nx.n10995\
        );

    \I__5153\ : InMux
    port map (
            O => \N__28476\,
            I => \N__28473\
        );

    \I__5152\ : LocalMux
    port map (
            O => \N__28473\,
            I => \nx.n2761\
        );

    \I__5151\ : InMux
    port map (
            O => \N__28470\,
            I => \bfn_10_25_0_\
        );

    \I__5150\ : InMux
    port map (
            O => \N__28467\,
            I => \N__28464\
        );

    \I__5149\ : LocalMux
    port map (
            O => \N__28464\,
            I => \nx.n2760\
        );

    \I__5148\ : InMux
    port map (
            O => \N__28461\,
            I => \nx.n10997\
        );

    \I__5147\ : InMux
    port map (
            O => \N__28458\,
            I => \N__28455\
        );

    \I__5146\ : LocalMux
    port map (
            O => \N__28455\,
            I => \N__28452\
        );

    \I__5145\ : Span4Mux_v
    port map (
            O => \N__28452\,
            I => \N__28449\
        );

    \I__5144\ : Odrv4
    port map (
            O => \N__28449\,
            I => \nx.n2759\
        );

    \I__5143\ : InMux
    port map (
            O => \N__28446\,
            I => \nx.n10998\
        );

    \I__5142\ : InMux
    port map (
            O => \N__28443\,
            I => \N__28440\
        );

    \I__5141\ : LocalMux
    port map (
            O => \N__28440\,
            I => \nx.n2758\
        );

    \I__5140\ : InMux
    port map (
            O => \N__28437\,
            I => \nx.n10999\
        );

    \I__5139\ : InMux
    port map (
            O => \N__28434\,
            I => \N__28431\
        );

    \I__5138\ : LocalMux
    port map (
            O => \N__28431\,
            I => \nx.n2757\
        );

    \I__5137\ : InMux
    port map (
            O => \N__28428\,
            I => \nx.n11000\
        );

    \I__5136\ : InMux
    port map (
            O => \N__28425\,
            I => \N__28422\
        );

    \I__5135\ : LocalMux
    port map (
            O => \N__28422\,
            I => \N__28419\
        );

    \I__5134\ : Odrv4
    port map (
            O => \N__28419\,
            I => \nx.n2756\
        );

    \I__5133\ : InMux
    port map (
            O => \N__28416\,
            I => \nx.n11001\
        );

    \I__5132\ : InMux
    port map (
            O => \N__28413\,
            I => \nx.n11002\
        );

    \I__5131\ : InMux
    port map (
            O => \N__28410\,
            I => \nx.n10985\
        );

    \I__5130\ : InMux
    port map (
            O => \N__28407\,
            I => \N__28404\
        );

    \I__5129\ : LocalMux
    port map (
            O => \N__28404\,
            I => \N__28401\
        );

    \I__5128\ : Odrv12
    port map (
            O => \N__28401\,
            I => \nx.n2771\
        );

    \I__5127\ : InMux
    port map (
            O => \N__28398\,
            I => \nx.n10986\
        );

    \I__5126\ : CascadeMux
    port map (
            O => \N__28395\,
            I => \N__28392\
        );

    \I__5125\ : InMux
    port map (
            O => \N__28392\,
            I => \N__28389\
        );

    \I__5124\ : LocalMux
    port map (
            O => \N__28389\,
            I => \N__28386\
        );

    \I__5123\ : Odrv12
    port map (
            O => \N__28386\,
            I => \nx.n2770\
        );

    \I__5122\ : InMux
    port map (
            O => \N__28383\,
            I => \nx.n10987\
        );

    \I__5121\ : InMux
    port map (
            O => \N__28380\,
            I => \N__28377\
        );

    \I__5120\ : LocalMux
    port map (
            O => \N__28377\,
            I => \nx.n2769\
        );

    \I__5119\ : InMux
    port map (
            O => \N__28374\,
            I => \bfn_10_24_0_\
        );

    \I__5118\ : InMux
    port map (
            O => \N__28371\,
            I => \N__28368\
        );

    \I__5117\ : LocalMux
    port map (
            O => \N__28368\,
            I => \N__28365\
        );

    \I__5116\ : Odrv4
    port map (
            O => \N__28365\,
            I => \nx.n2768\
        );

    \I__5115\ : InMux
    port map (
            O => \N__28362\,
            I => \nx.n10989\
        );

    \I__5114\ : InMux
    port map (
            O => \N__28359\,
            I => \nx.n10990\
        );

    \I__5113\ : InMux
    port map (
            O => \N__28356\,
            I => \nx.n10991\
        );

    \I__5112\ : InMux
    port map (
            O => \N__28353\,
            I => \nx.n10992\
        );

    \I__5111\ : InMux
    port map (
            O => \N__28350\,
            I => \nx.n10993\
        );

    \I__5110\ : CascadeMux
    port map (
            O => \N__28347\,
            I => \nx.n2788_cascade_\
        );

    \I__5109\ : CascadeMux
    port map (
            O => \N__28344\,
            I => \N__28341\
        );

    \I__5108\ : InMux
    port map (
            O => \N__28341\,
            I => \N__28337\
        );

    \I__5107\ : CascadeMux
    port map (
            O => \N__28340\,
            I => \N__28333\
        );

    \I__5106\ : LocalMux
    port map (
            O => \N__28337\,
            I => \N__28330\
        );

    \I__5105\ : InMux
    port map (
            O => \N__28336\,
            I => \N__28327\
        );

    \I__5104\ : InMux
    port map (
            O => \N__28333\,
            I => \N__28324\
        );

    \I__5103\ : Span4Mux_h
    port map (
            O => \N__28330\,
            I => \N__28319\
        );

    \I__5102\ : LocalMux
    port map (
            O => \N__28327\,
            I => \N__28319\
        );

    \I__5101\ : LocalMux
    port map (
            O => \N__28324\,
            I => \nx.n2789\
        );

    \I__5100\ : Odrv4
    port map (
            O => \N__28319\,
            I => \nx.n2789\
        );

    \I__5099\ : CascadeMux
    port map (
            O => \N__28314\,
            I => \nx.n26_adj_706_cascade_\
        );

    \I__5098\ : InMux
    port map (
            O => \N__28311\,
            I => \N__28308\
        );

    \I__5097\ : LocalMux
    port map (
            O => \N__28308\,
            I => \N__28305\
        );

    \I__5096\ : Odrv4
    port map (
            O => \N__28305\,
            I => \nx.n38_adj_713\
        );

    \I__5095\ : InMux
    port map (
            O => \N__28302\,
            I => \N__28299\
        );

    \I__5094\ : LocalMux
    port map (
            O => \N__28299\,
            I => \N__28296\
        );

    \I__5093\ : Odrv4
    port map (
            O => \N__28296\,
            I => \nx.n43_adj_735\
        );

    \I__5092\ : InMux
    port map (
            O => \N__28293\,
            I => \N__28290\
        );

    \I__5091\ : LocalMux
    port map (
            O => \N__28290\,
            I => \N__28287\
        );

    \I__5090\ : Span4Mux_v
    port map (
            O => \N__28287\,
            I => \N__28284\
        );

    \I__5089\ : Odrv4
    port map (
            O => \N__28284\,
            I => \nx.n2777\
        );

    \I__5088\ : InMux
    port map (
            O => \N__28281\,
            I => \bfn_10_23_0_\
        );

    \I__5087\ : InMux
    port map (
            O => \N__28278\,
            I => \N__28275\
        );

    \I__5086\ : LocalMux
    port map (
            O => \N__28275\,
            I => \N__28272\
        );

    \I__5085\ : Span4Mux_v
    port map (
            O => \N__28272\,
            I => \N__28269\
        );

    \I__5084\ : Odrv4
    port map (
            O => \N__28269\,
            I => \nx.n2776\
        );

    \I__5083\ : InMux
    port map (
            O => \N__28266\,
            I => \nx.n10981\
        );

    \I__5082\ : InMux
    port map (
            O => \N__28263\,
            I => \N__28260\
        );

    \I__5081\ : LocalMux
    port map (
            O => \N__28260\,
            I => \N__28257\
        );

    \I__5080\ : Odrv4
    port map (
            O => \N__28257\,
            I => \nx.n2775\
        );

    \I__5079\ : InMux
    port map (
            O => \N__28254\,
            I => \nx.n10982\
        );

    \I__5078\ : InMux
    port map (
            O => \N__28251\,
            I => \nx.n10983\
        );

    \I__5077\ : InMux
    port map (
            O => \N__28248\,
            I => \N__28245\
        );

    \I__5076\ : LocalMux
    port map (
            O => \N__28245\,
            I => \nx.n2773\
        );

    \I__5075\ : InMux
    port map (
            O => \N__28242\,
            I => \nx.n10984\
        );

    \I__5074\ : InMux
    port map (
            O => \N__28239\,
            I => \N__28236\
        );

    \I__5073\ : LocalMux
    port map (
            O => \N__28236\,
            I => \nx.n2772\
        );

    \I__5072\ : InMux
    port map (
            O => \N__28233\,
            I => \N__28230\
        );

    \I__5071\ : LocalMux
    port map (
            O => \N__28230\,
            I => \N__28226\
        );

    \I__5070\ : InMux
    port map (
            O => \N__28229\,
            I => \N__28223\
        );

    \I__5069\ : Odrv4
    port map (
            O => \N__28226\,
            I => \nx.n2809\
        );

    \I__5068\ : LocalMux
    port map (
            O => \N__28223\,
            I => \nx.n2809\
        );

    \I__5067\ : CascadeMux
    port map (
            O => \N__28218\,
            I => \nx.n2809_cascade_\
        );

    \I__5066\ : InMux
    port map (
            O => \N__28215\,
            I => \N__28210\
        );

    \I__5065\ : InMux
    port map (
            O => \N__28214\,
            I => \N__28207\
        );

    \I__5064\ : InMux
    port map (
            O => \N__28213\,
            I => \N__28202\
        );

    \I__5063\ : LocalMux
    port map (
            O => \N__28210\,
            I => \N__28199\
        );

    \I__5062\ : LocalMux
    port map (
            O => \N__28207\,
            I => \N__28196\
        );

    \I__5061\ : InMux
    port map (
            O => \N__28206\,
            I => \N__28193\
        );

    \I__5060\ : InMux
    port map (
            O => \N__28205\,
            I => \N__28190\
        );

    \I__5059\ : LocalMux
    port map (
            O => \N__28202\,
            I => \N__28187\
        );

    \I__5058\ : Span4Mux_v
    port map (
            O => \N__28199\,
            I => \N__28180\
        );

    \I__5057\ : Span4Mux_h
    port map (
            O => \N__28196\,
            I => \N__28180\
        );

    \I__5056\ : LocalMux
    port map (
            O => \N__28193\,
            I => \N__28180\
        );

    \I__5055\ : LocalMux
    port map (
            O => \N__28190\,
            I => \N__28175\
        );

    \I__5054\ : Span4Mux_v
    port map (
            O => \N__28187\,
            I => \N__28175\
        );

    \I__5053\ : Span4Mux_h
    port map (
            O => \N__28180\,
            I => \N__28172\
        );

    \I__5052\ : Odrv4
    port map (
            O => \N__28175\,
            I => \nx.bit_ctr_7\
        );

    \I__5051\ : Odrv4
    port map (
            O => \N__28172\,
            I => \nx.bit_ctr_7\
        );

    \I__5050\ : InMux
    port map (
            O => \N__28167\,
            I => \N__28164\
        );

    \I__5049\ : LocalMux
    port map (
            O => \N__28164\,
            I => \nx.n30_adj_704\
        );

    \I__5048\ : CascadeMux
    port map (
            O => \N__28161\,
            I => \N__28157\
        );

    \I__5047\ : InMux
    port map (
            O => \N__28160\,
            I => \N__28154\
        );

    \I__5046\ : InMux
    port map (
            O => \N__28157\,
            I => \N__28151\
        );

    \I__5045\ : LocalMux
    port map (
            O => \N__28154\,
            I => \nx.n2802\
        );

    \I__5044\ : LocalMux
    port map (
            O => \N__28151\,
            I => \nx.n2802\
        );

    \I__5043\ : InMux
    port map (
            O => \N__28146\,
            I => \N__28143\
        );

    \I__5042\ : LocalMux
    port map (
            O => \N__28143\,
            I => \nx.n2869\
        );

    \I__5041\ : CascadeMux
    port map (
            O => \N__28140\,
            I => \nx.n2802_cascade_\
        );

    \I__5040\ : InMux
    port map (
            O => \N__28137\,
            I => \N__28133\
        );

    \I__5039\ : CascadeMux
    port map (
            O => \N__28136\,
            I => \N__28130\
        );

    \I__5038\ : LocalMux
    port map (
            O => \N__28133\,
            I => \N__28126\
        );

    \I__5037\ : InMux
    port map (
            O => \N__28130\,
            I => \N__28123\
        );

    \I__5036\ : InMux
    port map (
            O => \N__28129\,
            I => \N__28120\
        );

    \I__5035\ : Odrv4
    port map (
            O => \N__28126\,
            I => \nx.n2795\
        );

    \I__5034\ : LocalMux
    port map (
            O => \N__28123\,
            I => \nx.n2795\
        );

    \I__5033\ : LocalMux
    port map (
            O => \N__28120\,
            I => \nx.n2795\
        );

    \I__5032\ : CascadeMux
    port map (
            O => \N__28113\,
            I => \nx.n2720_cascade_\
        );

    \I__5031\ : InMux
    port map (
            O => \N__28110\,
            I => \N__28103\
        );

    \I__5030\ : InMux
    port map (
            O => \N__28109\,
            I => \N__28103\
        );

    \I__5029\ : CascadeMux
    port map (
            O => \N__28108\,
            I => \N__28100\
        );

    \I__5028\ : LocalMux
    port map (
            O => \N__28103\,
            I => \N__28097\
        );

    \I__5027\ : InMux
    port map (
            O => \N__28100\,
            I => \N__28094\
        );

    \I__5026\ : Span4Mux_h
    port map (
            O => \N__28097\,
            I => \N__28091\
        );

    \I__5025\ : LocalMux
    port map (
            O => \N__28094\,
            I => \N__28088\
        );

    \I__5024\ : Odrv4
    port map (
            O => \N__28091\,
            I => \nx.n2801\
        );

    \I__5023\ : Odrv4
    port map (
            O => \N__28088\,
            I => \nx.n2801\
        );

    \I__5022\ : CascadeMux
    port map (
            O => \N__28083\,
            I => \N__28078\
        );

    \I__5021\ : InMux
    port map (
            O => \N__28082\,
            I => \N__28075\
        );

    \I__5020\ : InMux
    port map (
            O => \N__28081\,
            I => \N__28072\
        );

    \I__5019\ : InMux
    port map (
            O => \N__28078\,
            I => \N__28069\
        );

    \I__5018\ : LocalMux
    port map (
            O => \N__28075\,
            I => \nx.n2808\
        );

    \I__5017\ : LocalMux
    port map (
            O => \N__28072\,
            I => \nx.n2808\
        );

    \I__5016\ : LocalMux
    port map (
            O => \N__28069\,
            I => \nx.n2808\
        );

    \I__5015\ : CascadeMux
    port map (
            O => \N__28062\,
            I => \nx.n40_adj_705_cascade_\
        );

    \I__5014\ : CascadeMux
    port map (
            O => \N__28059\,
            I => \nx.n44_adj_721_cascade_\
        );

    \I__5013\ : InMux
    port map (
            O => \N__28056\,
            I => \N__28053\
        );

    \I__5012\ : LocalMux
    port map (
            O => \N__28053\,
            I => \N__28050\
        );

    \I__5011\ : Odrv4
    port map (
            O => \N__28050\,
            I => \nx.n2862\
        );

    \I__5010\ : CascadeMux
    port map (
            O => \N__28047\,
            I => \nx.n2819_cascade_\
        );

    \I__5009\ : InMux
    port map (
            O => \N__28044\,
            I => \N__28041\
        );

    \I__5008\ : LocalMux
    port map (
            O => \N__28041\,
            I => \nx.n2874\
        );

    \I__5007\ : InMux
    port map (
            O => \N__28038\,
            I => \N__28035\
        );

    \I__5006\ : LocalMux
    port map (
            O => \N__28035\,
            I => \nx.n42_adj_730\
        );

    \I__5005\ : CascadeMux
    port map (
            O => \N__28032\,
            I => \N__28028\
        );

    \I__5004\ : CascadeMux
    port map (
            O => \N__28031\,
            I => \N__28024\
        );

    \I__5003\ : InMux
    port map (
            O => \N__28028\,
            I => \N__28019\
        );

    \I__5002\ : InMux
    port map (
            O => \N__28027\,
            I => \N__28019\
        );

    \I__5001\ : InMux
    port map (
            O => \N__28024\,
            I => \N__28016\
        );

    \I__5000\ : LocalMux
    port map (
            O => \N__28019\,
            I => \nx.n2807\
        );

    \I__4999\ : LocalMux
    port map (
            O => \N__28016\,
            I => \nx.n2807\
        );

    \I__4998\ : CascadeMux
    port map (
            O => \N__28011\,
            I => \nx.n2987_cascade_\
        );

    \I__4997\ : CascadeMux
    port map (
            O => \N__28008\,
            I => \nx.n41_cascade_\
        );

    \I__4996\ : InMux
    port map (
            O => \N__28005\,
            I => \N__28002\
        );

    \I__4995\ : LocalMux
    port map (
            O => \N__28002\,
            I => \nx.n39_adj_671\
        );

    \I__4994\ : CascadeMux
    port map (
            O => \N__27999\,
            I => \nx.n50_cascade_\
        );

    \I__4993\ : InMux
    port map (
            O => \N__27996\,
            I => \N__27993\
        );

    \I__4992\ : LocalMux
    port map (
            O => \N__27993\,
            I => \N__27990\
        );

    \I__4991\ : Odrv4
    port map (
            O => \N__27990\,
            I => \nx.n2877\
        );

    \I__4990\ : InMux
    port map (
            O => \N__27987\,
            I => \N__27984\
        );

    \I__4989\ : LocalMux
    port map (
            O => \N__27984\,
            I => \N__27981\
        );

    \I__4988\ : Span4Mux_v
    port map (
            O => \N__27981\,
            I => \N__27978\
        );

    \I__4987\ : Odrv4
    port map (
            O => \N__27978\,
            I => \nx.n2857\
        );

    \I__4986\ : InMux
    port map (
            O => \N__27975\,
            I => \N__27971\
        );

    \I__4985\ : CascadeMux
    port map (
            O => \N__27974\,
            I => \N__27967\
        );

    \I__4984\ : LocalMux
    port map (
            O => \N__27971\,
            I => \N__27964\
        );

    \I__4983\ : CascadeMux
    port map (
            O => \N__27970\,
            I => \N__27961\
        );

    \I__4982\ : InMux
    port map (
            O => \N__27967\,
            I => \N__27958\
        );

    \I__4981\ : Span4Mux_h
    port map (
            O => \N__27964\,
            I => \N__27955\
        );

    \I__4980\ : InMux
    port map (
            O => \N__27961\,
            I => \N__27952\
        );

    \I__4979\ : LocalMux
    port map (
            O => \N__27958\,
            I => \N__27949\
        );

    \I__4978\ : Odrv4
    port map (
            O => \N__27955\,
            I => \nx.n2790\
        );

    \I__4977\ : LocalMux
    port map (
            O => \N__27952\,
            I => \nx.n2790\
        );

    \I__4976\ : Odrv12
    port map (
            O => \N__27949\,
            I => \nx.n2790\
        );

    \I__4975\ : CascadeMux
    port map (
            O => \N__27942\,
            I => \nx.n2889_cascade_\
        );

    \I__4974\ : InMux
    port map (
            O => \N__27939\,
            I => \N__27936\
        );

    \I__4973\ : LocalMux
    port map (
            O => \N__27936\,
            I => \N__27933\
        );

    \I__4972\ : Odrv4
    port map (
            O => \N__27933\,
            I => \nx.n2868\
        );

    \I__4971\ : CascadeMux
    port map (
            O => \N__27930\,
            I => \nx.n12811_cascade_\
        );

    \I__4970\ : CascadeMux
    port map (
            O => \N__27927\,
            I => \nx.n12813_cascade_\
        );

    \I__4969\ : InMux
    port map (
            O => \N__27924\,
            I => \N__27921\
        );

    \I__4968\ : LocalMux
    port map (
            O => \N__27921\,
            I => \nx.n12815\
        );

    \I__4967\ : InMux
    port map (
            O => \N__27918\,
            I => \N__27915\
        );

    \I__4966\ : LocalMux
    port map (
            O => \N__27915\,
            I => \nx.n43_adj_753\
        );

    \I__4965\ : CascadeMux
    port map (
            O => \N__27912\,
            I => \nx.n46_cascade_\
        );

    \I__4964\ : CascadeMux
    port map (
            O => \N__27909\,
            I => \nx.n13_adj_743_cascade_\
        );

    \I__4963\ : InMux
    port map (
            O => \N__27906\,
            I => \N__27903\
        );

    \I__4962\ : LocalMux
    port map (
            O => \N__27903\,
            I => \nx.n12775\
        );

    \I__4961\ : CascadeMux
    port map (
            O => \N__27900\,
            I => \nx.n12787_cascade_\
        );

    \I__4960\ : InMux
    port map (
            O => \N__27897\,
            I => \N__27894\
        );

    \I__4959\ : LocalMux
    port map (
            O => \N__27894\,
            I => \nx.n12803\
        );

    \I__4958\ : InMux
    port map (
            O => \N__27891\,
            I => \N__27888\
        );

    \I__4957\ : LocalMux
    port map (
            O => \N__27888\,
            I => \nx.n35_adj_738\
        );

    \I__4956\ : InMux
    port map (
            O => \N__27885\,
            I => \N__27879\
        );

    \I__4955\ : InMux
    port map (
            O => \N__27884\,
            I => \N__27879\
        );

    \I__4954\ : LocalMux
    port map (
            O => \N__27879\,
            I => \N__27875\
        );

    \I__4953\ : InMux
    port map (
            O => \N__27878\,
            I => \N__27872\
        );

    \I__4952\ : Odrv4
    port map (
            O => \N__27875\,
            I => blink_counter_21
        );

    \I__4951\ : LocalMux
    port map (
            O => \N__27872\,
            I => blink_counter_21
        );

    \I__4950\ : InMux
    port map (
            O => \N__27867\,
            I => n10664
        );

    \I__4949\ : InMux
    port map (
            O => \N__27864\,
            I => \N__27858\
        );

    \I__4948\ : InMux
    port map (
            O => \N__27863\,
            I => \N__27858\
        );

    \I__4947\ : LocalMux
    port map (
            O => \N__27858\,
            I => \N__27854\
        );

    \I__4946\ : InMux
    port map (
            O => \N__27857\,
            I => \N__27851\
        );

    \I__4945\ : Odrv12
    port map (
            O => \N__27854\,
            I => blink_counter_22
        );

    \I__4944\ : LocalMux
    port map (
            O => \N__27851\,
            I => blink_counter_22
        );

    \I__4943\ : InMux
    port map (
            O => \N__27846\,
            I => n10665
        );

    \I__4942\ : CascadeMux
    port map (
            O => \N__27843\,
            I => \N__27839\
        );

    \I__4941\ : InMux
    port map (
            O => \N__27842\,
            I => \N__27834\
        );

    \I__4940\ : InMux
    port map (
            O => \N__27839\,
            I => \N__27834\
        );

    \I__4939\ : LocalMux
    port map (
            O => \N__27834\,
            I => \N__27830\
        );

    \I__4938\ : InMux
    port map (
            O => \N__27833\,
            I => \N__27827\
        );

    \I__4937\ : Odrv4
    port map (
            O => \N__27830\,
            I => blink_counter_23
        );

    \I__4936\ : LocalMux
    port map (
            O => \N__27827\,
            I => blink_counter_23
        );

    \I__4935\ : InMux
    port map (
            O => \N__27822\,
            I => n10666
        );

    \I__4934\ : CascadeMux
    port map (
            O => \N__27819\,
            I => \N__27816\
        );

    \I__4933\ : InMux
    port map (
            O => \N__27816\,
            I => \N__27810\
        );

    \I__4932\ : InMux
    port map (
            O => \N__27815\,
            I => \N__27810\
        );

    \I__4931\ : LocalMux
    port map (
            O => \N__27810\,
            I => \N__27807\
        );

    \I__4930\ : Span4Mux_v
    port map (
            O => \N__27807\,
            I => \N__27803\
        );

    \I__4929\ : InMux
    port map (
            O => \N__27806\,
            I => \N__27800\
        );

    \I__4928\ : Odrv4
    port map (
            O => \N__27803\,
            I => blink_counter_24
        );

    \I__4927\ : LocalMux
    port map (
            O => \N__27800\,
            I => blink_counter_24
        );

    \I__4926\ : InMux
    port map (
            O => \N__27795\,
            I => \bfn_9_32_0_\
        );

    \I__4925\ : InMux
    port map (
            O => \N__27792\,
            I => n10668
        );

    \I__4924\ : InMux
    port map (
            O => \N__27789\,
            I => \N__27786\
        );

    \I__4923\ : LocalMux
    port map (
            O => \N__27786\,
            I => \N__27783\
        );

    \I__4922\ : Span4Mux_v
    port map (
            O => \N__27783\,
            I => \N__27779\
        );

    \I__4921\ : InMux
    port map (
            O => \N__27782\,
            I => \N__27776\
        );

    \I__4920\ : Odrv4
    port map (
            O => \N__27779\,
            I => blink_counter_25
        );

    \I__4919\ : LocalMux
    port map (
            O => \N__27776\,
            I => blink_counter_25
        );

    \I__4918\ : CascadeMux
    port map (
            O => \N__27771\,
            I => \nx.n45_adj_754_cascade_\
        );

    \I__4917\ : CascadeMux
    port map (
            O => \N__27768\,
            I => \nx.n12809_cascade_\
        );

    \I__4916\ : InMux
    port map (
            O => \N__27765\,
            I => \N__27762\
        );

    \I__4915\ : LocalMux
    port map (
            O => \N__27762\,
            I => n13
        );

    \I__4914\ : InMux
    port map (
            O => \N__27759\,
            I => n10656
        );

    \I__4913\ : InMux
    port map (
            O => \N__27756\,
            I => \N__27753\
        );

    \I__4912\ : LocalMux
    port map (
            O => \N__27753\,
            I => n12
        );

    \I__4911\ : InMux
    port map (
            O => \N__27750\,
            I => n10657
        );

    \I__4910\ : InMux
    port map (
            O => \N__27747\,
            I => \N__27744\
        );

    \I__4909\ : LocalMux
    port map (
            O => \N__27744\,
            I => n11
        );

    \I__4908\ : InMux
    port map (
            O => \N__27741\,
            I => n10658
        );

    \I__4907\ : InMux
    port map (
            O => \N__27738\,
            I => \N__27735\
        );

    \I__4906\ : LocalMux
    port map (
            O => \N__27735\,
            I => n10_adj_806
        );

    \I__4905\ : InMux
    port map (
            O => \N__27732\,
            I => \bfn_9_31_0_\
        );

    \I__4904\ : InMux
    port map (
            O => \N__27729\,
            I => \N__27726\
        );

    \I__4903\ : LocalMux
    port map (
            O => \N__27726\,
            I => n9_adj_807
        );

    \I__4902\ : InMux
    port map (
            O => \N__27723\,
            I => n10660
        );

    \I__4901\ : InMux
    port map (
            O => \N__27720\,
            I => \N__27717\
        );

    \I__4900\ : LocalMux
    port map (
            O => \N__27717\,
            I => n8
        );

    \I__4899\ : InMux
    port map (
            O => \N__27714\,
            I => n10661
        );

    \I__4898\ : InMux
    port map (
            O => \N__27711\,
            I => \N__27708\
        );

    \I__4897\ : LocalMux
    port map (
            O => \N__27708\,
            I => n7_adj_808
        );

    \I__4896\ : InMux
    port map (
            O => \N__27705\,
            I => n10662
        );

    \I__4895\ : InMux
    port map (
            O => \N__27702\,
            I => \N__27699\
        );

    \I__4894\ : LocalMux
    port map (
            O => \N__27699\,
            I => n6_adj_809
        );

    \I__4893\ : InMux
    port map (
            O => \N__27696\,
            I => n10663
        );

    \I__4892\ : InMux
    port map (
            O => \N__27693\,
            I => \N__27690\
        );

    \I__4891\ : LocalMux
    port map (
            O => \N__27690\,
            I => n21
        );

    \I__4890\ : InMux
    port map (
            O => \N__27687\,
            I => n10648
        );

    \I__4889\ : InMux
    port map (
            O => \N__27684\,
            I => \N__27681\
        );

    \I__4888\ : LocalMux
    port map (
            O => \N__27681\,
            I => n20
        );

    \I__4887\ : InMux
    port map (
            O => \N__27678\,
            I => n10649
        );

    \I__4886\ : InMux
    port map (
            O => \N__27675\,
            I => \N__27672\
        );

    \I__4885\ : LocalMux
    port map (
            O => \N__27672\,
            I => n19_adj_800
        );

    \I__4884\ : InMux
    port map (
            O => \N__27669\,
            I => n10650
        );

    \I__4883\ : InMux
    port map (
            O => \N__27666\,
            I => \N__27663\
        );

    \I__4882\ : LocalMux
    port map (
            O => \N__27663\,
            I => n18
        );

    \I__4881\ : InMux
    port map (
            O => \N__27660\,
            I => \bfn_9_30_0_\
        );

    \I__4880\ : InMux
    port map (
            O => \N__27657\,
            I => \N__27654\
        );

    \I__4879\ : LocalMux
    port map (
            O => \N__27654\,
            I => n17
        );

    \I__4878\ : InMux
    port map (
            O => \N__27651\,
            I => n10652
        );

    \I__4877\ : InMux
    port map (
            O => \N__27648\,
            I => \N__27645\
        );

    \I__4876\ : LocalMux
    port map (
            O => \N__27645\,
            I => n16
        );

    \I__4875\ : InMux
    port map (
            O => \N__27642\,
            I => n10653
        );

    \I__4874\ : InMux
    port map (
            O => \N__27639\,
            I => \N__27636\
        );

    \I__4873\ : LocalMux
    port map (
            O => \N__27636\,
            I => n15
        );

    \I__4872\ : InMux
    port map (
            O => \N__27633\,
            I => n10654
        );

    \I__4871\ : InMux
    port map (
            O => \N__27630\,
            I => \N__27627\
        );

    \I__4870\ : LocalMux
    port map (
            O => \N__27627\,
            I => n14_adj_802
        );

    \I__4869\ : InMux
    port map (
            O => \N__27624\,
            I => n10655
        );

    \I__4868\ : InMux
    port map (
            O => \N__27621\,
            I => \N__27618\
        );

    \I__4867\ : LocalMux
    port map (
            O => \N__27618\,
            I => \N__27615\
        );

    \I__4866\ : Odrv4
    port map (
            O => \N__27615\,
            I => \nx.n1969\
        );

    \I__4865\ : CascadeMux
    port map (
            O => \N__27612\,
            I => \N__27609\
        );

    \I__4864\ : InMux
    port map (
            O => \N__27609\,
            I => \N__27606\
        );

    \I__4863\ : LocalMux
    port map (
            O => \N__27606\,
            I => \N__27602\
        );

    \I__4862\ : CascadeMux
    port map (
            O => \N__27605\,
            I => \N__27598\
        );

    \I__4861\ : Span4Mux_h
    port map (
            O => \N__27602\,
            I => \N__27595\
        );

    \I__4860\ : InMux
    port map (
            O => \N__27601\,
            I => \N__27592\
        );

    \I__4859\ : InMux
    port map (
            O => \N__27598\,
            I => \N__27589\
        );

    \I__4858\ : Odrv4
    port map (
            O => \N__27595\,
            I => \nx.n1902\
        );

    \I__4857\ : LocalMux
    port map (
            O => \N__27592\,
            I => \nx.n1902\
        );

    \I__4856\ : LocalMux
    port map (
            O => \N__27589\,
            I => \nx.n1902\
        );

    \I__4855\ : CascadeMux
    port map (
            O => \N__27582\,
            I => \N__27577\
        );

    \I__4854\ : CascadeMux
    port map (
            O => \N__27581\,
            I => \N__27573\
        );

    \I__4853\ : CascadeMux
    port map (
            O => \N__27580\,
            I => \N__27569\
        );

    \I__4852\ : InMux
    port map (
            O => \N__27577\,
            I => \N__27558\
        );

    \I__4851\ : InMux
    port map (
            O => \N__27576\,
            I => \N__27558\
        );

    \I__4850\ : InMux
    port map (
            O => \N__27573\,
            I => \N__27558\
        );

    \I__4849\ : InMux
    port map (
            O => \N__27572\,
            I => \N__27558\
        );

    \I__4848\ : InMux
    port map (
            O => \N__27569\,
            I => \N__27553\
        );

    \I__4847\ : InMux
    port map (
            O => \N__27568\,
            I => \N__27553\
        );

    \I__4846\ : CascadeMux
    port map (
            O => \N__27567\,
            I => \N__27547\
        );

    \I__4845\ : LocalMux
    port map (
            O => \N__27558\,
            I => \N__27540\
        );

    \I__4844\ : LocalMux
    port map (
            O => \N__27553\,
            I => \N__27537\
        );

    \I__4843\ : InMux
    port map (
            O => \N__27552\,
            I => \N__27534\
        );

    \I__4842\ : InMux
    port map (
            O => \N__27551\,
            I => \N__27525\
        );

    \I__4841\ : InMux
    port map (
            O => \N__27550\,
            I => \N__27525\
        );

    \I__4840\ : InMux
    port map (
            O => \N__27547\,
            I => \N__27525\
        );

    \I__4839\ : InMux
    port map (
            O => \N__27546\,
            I => \N__27525\
        );

    \I__4838\ : CascadeMux
    port map (
            O => \N__27545\,
            I => \N__27522\
        );

    \I__4837\ : CascadeMux
    port map (
            O => \N__27544\,
            I => \N__27519\
        );

    \I__4836\ : InMux
    port map (
            O => \N__27543\,
            I => \N__27515\
        );

    \I__4835\ : Span4Mux_v
    port map (
            O => \N__27540\,
            I => \N__27510\
        );

    \I__4834\ : Span4Mux_v
    port map (
            O => \N__27537\,
            I => \N__27510\
        );

    \I__4833\ : LocalMux
    port map (
            O => \N__27534\,
            I => \N__27505\
        );

    \I__4832\ : LocalMux
    port map (
            O => \N__27525\,
            I => \N__27505\
        );

    \I__4831\ : InMux
    port map (
            O => \N__27522\,
            I => \N__27498\
        );

    \I__4830\ : InMux
    port map (
            O => \N__27519\,
            I => \N__27498\
        );

    \I__4829\ : InMux
    port map (
            O => \N__27518\,
            I => \N__27498\
        );

    \I__4828\ : LocalMux
    port map (
            O => \N__27515\,
            I => \nx.n1928\
        );

    \I__4827\ : Odrv4
    port map (
            O => \N__27510\,
            I => \nx.n1928\
        );

    \I__4826\ : Odrv4
    port map (
            O => \N__27505\,
            I => \nx.n1928\
        );

    \I__4825\ : LocalMux
    port map (
            O => \N__27498\,
            I => \nx.n1928\
        );

    \I__4824\ : InMux
    port map (
            O => \N__27489\,
            I => \N__27486\
        );

    \I__4823\ : LocalMux
    port map (
            O => \N__27486\,
            I => \nx.n2068\
        );

    \I__4822\ : CascadeMux
    port map (
            O => \N__27483\,
            I => \nx.n2001_cascade_\
        );

    \I__4821\ : InMux
    port map (
            O => \N__27480\,
            I => \N__27477\
        );

    \I__4820\ : LocalMux
    port map (
            O => \N__27477\,
            I => \nx.n2067\
        );

    \I__4819\ : CascadeMux
    port map (
            O => \N__27474\,
            I => \nx.n2099_cascade_\
        );

    \I__4818\ : InMux
    port map (
            O => \N__27471\,
            I => \N__27468\
        );

    \I__4817\ : LocalMux
    port map (
            O => \N__27468\,
            I => n26_adj_798
        );

    \I__4816\ : InMux
    port map (
            O => \N__27465\,
            I => \bfn_9_29_0_\
        );

    \I__4815\ : InMux
    port map (
            O => \N__27462\,
            I => \N__27459\
        );

    \I__4814\ : LocalMux
    port map (
            O => \N__27459\,
            I => n25
        );

    \I__4813\ : InMux
    port map (
            O => \N__27456\,
            I => n10644
        );

    \I__4812\ : InMux
    port map (
            O => \N__27453\,
            I => \N__27450\
        );

    \I__4811\ : LocalMux
    port map (
            O => \N__27450\,
            I => n24
        );

    \I__4810\ : InMux
    port map (
            O => \N__27447\,
            I => n10645
        );

    \I__4809\ : InMux
    port map (
            O => \N__27444\,
            I => \N__27441\
        );

    \I__4808\ : LocalMux
    port map (
            O => \N__27441\,
            I => n23
        );

    \I__4807\ : InMux
    port map (
            O => \N__27438\,
            I => n10646
        );

    \I__4806\ : InMux
    port map (
            O => \N__27435\,
            I => \N__27432\
        );

    \I__4805\ : LocalMux
    port map (
            O => \N__27432\,
            I => n22_adj_799
        );

    \I__4804\ : InMux
    port map (
            O => \N__27429\,
            I => n10647
        );

    \I__4803\ : InMux
    port map (
            O => \N__27426\,
            I => \nx.n10858\
        );

    \I__4802\ : InMux
    port map (
            O => \N__27423\,
            I => \nx.n10859\
        );

    \I__4801\ : InMux
    port map (
            O => \N__27420\,
            I => \nx.n10860\
        );

    \I__4800\ : InMux
    port map (
            O => \N__27417\,
            I => \nx.n10861\
        );

    \I__4799\ : InMux
    port map (
            O => \N__27414\,
            I => \nx.n10862\
        );

    \I__4798\ : InMux
    port map (
            O => \N__27411\,
            I => \N__27408\
        );

    \I__4797\ : LocalMux
    port map (
            O => \N__27408\,
            I => \N__27404\
        );

    \I__4796\ : InMux
    port map (
            O => \N__27407\,
            I => \N__27401\
        );

    \I__4795\ : Odrv4
    port map (
            O => \N__27404\,
            I => \nx.n1994\
        );

    \I__4794\ : LocalMux
    port map (
            O => \N__27401\,
            I => \nx.n1994\
        );

    \I__4793\ : InMux
    port map (
            O => \N__27396\,
            I => \bfn_9_28_0_\
        );

    \I__4792\ : CascadeMux
    port map (
            O => \N__27393\,
            I => \N__27389\
        );

    \I__4791\ : CascadeMux
    port map (
            O => \N__27392\,
            I => \N__27386\
        );

    \I__4790\ : InMux
    port map (
            O => \N__27389\,
            I => \N__27383\
        );

    \I__4789\ : InMux
    port map (
            O => \N__27386\,
            I => \N__27380\
        );

    \I__4788\ : LocalMux
    port map (
            O => \N__27383\,
            I => \N__27375\
        );

    \I__4787\ : LocalMux
    port map (
            O => \N__27380\,
            I => \N__27375\
        );

    \I__4786\ : Span4Mux_v
    port map (
            O => \N__27375\,
            I => \N__27372\
        );

    \I__4785\ : Span4Mux_h
    port map (
            O => \N__27372\,
            I => \N__27369\
        );

    \I__4784\ : Odrv4
    port map (
            O => \N__27369\,
            I => \nx.n1995\
        );

    \I__4783\ : InMux
    port map (
            O => \N__27366\,
            I => \N__27363\
        );

    \I__4782\ : LocalMux
    port map (
            O => \N__27363\,
            I => \nx.n2062\
        );

    \I__4781\ : CascadeMux
    port map (
            O => \N__27360\,
            I => \nx.n2094_cascade_\
        );

    \I__4780\ : InMux
    port map (
            O => \N__27357\,
            I => \N__27352\
        );

    \I__4779\ : CascadeMux
    port map (
            O => \N__27356\,
            I => \N__27349\
        );

    \I__4778\ : InMux
    port map (
            O => \N__27355\,
            I => \N__27346\
        );

    \I__4777\ : LocalMux
    port map (
            O => \N__27352\,
            I => \N__27343\
        );

    \I__4776\ : InMux
    port map (
            O => \N__27349\,
            I => \N__27340\
        );

    \I__4775\ : LocalMux
    port map (
            O => \N__27346\,
            I => \N__27337\
        );

    \I__4774\ : Odrv4
    port map (
            O => \N__27343\,
            I => \nx.n1901\
        );

    \I__4773\ : LocalMux
    port map (
            O => \N__27340\,
            I => \nx.n1901\
        );

    \I__4772\ : Odrv4
    port map (
            O => \N__27337\,
            I => \nx.n1901\
        );

    \I__4771\ : InMux
    port map (
            O => \N__27330\,
            I => \N__27327\
        );

    \I__4770\ : LocalMux
    port map (
            O => \N__27327\,
            I => \N__27324\
        );

    \I__4769\ : Odrv4
    port map (
            O => \N__27324\,
            I => \nx.n1968\
        );

    \I__4768\ : InMux
    port map (
            O => \N__27321\,
            I => \nx.n10849\
        );

    \I__4767\ : InMux
    port map (
            O => \N__27318\,
            I => \nx.n10850\
        );

    \I__4766\ : InMux
    port map (
            O => \N__27315\,
            I => \nx.n10851\
        );

    \I__4765\ : InMux
    port map (
            O => \N__27312\,
            I => \nx.n10852\
        );

    \I__4764\ : InMux
    port map (
            O => \N__27309\,
            I => \nx.n10853\
        );

    \I__4763\ : InMux
    port map (
            O => \N__27306\,
            I => \nx.n10854\
        );

    \I__4762\ : InMux
    port map (
            O => \N__27303\,
            I => \bfn_9_27_0_\
        );

    \I__4761\ : InMux
    port map (
            O => \N__27300\,
            I => \nx.n10856\
        );

    \I__4760\ : InMux
    port map (
            O => \N__27297\,
            I => \nx.n10857\
        );

    \I__4759\ : InMux
    port map (
            O => \N__27294\,
            I => \N__27290\
        );

    \I__4758\ : InMux
    port map (
            O => \N__27293\,
            I => \N__27286\
        );

    \I__4757\ : LocalMux
    port map (
            O => \N__27290\,
            I => \N__27283\
        );

    \I__4756\ : InMux
    port map (
            O => \N__27289\,
            I => \N__27280\
        );

    \I__4755\ : LocalMux
    port map (
            O => \N__27286\,
            I => \N__27275\
        );

    \I__4754\ : Span4Mux_v
    port map (
            O => \N__27283\,
            I => \N__27275\
        );

    \I__4753\ : LocalMux
    port map (
            O => \N__27280\,
            I => \N__27272\
        );

    \I__4752\ : Span4Mux_v
    port map (
            O => \N__27275\,
            I => \N__27267\
        );

    \I__4751\ : Span4Mux_h
    port map (
            O => \N__27272\,
            I => \N__27264\
        );

    \I__4750\ : InMux
    port map (
            O => \N__27271\,
            I => \N__27261\
        );

    \I__4749\ : InMux
    port map (
            O => \N__27270\,
            I => \N__27258\
        );

    \I__4748\ : Span4Mux_h
    port map (
            O => \N__27267\,
            I => \N__27255\
        );

    \I__4747\ : Span4Mux_v
    port map (
            O => \N__27264\,
            I => \N__27252\
        );

    \I__4746\ : LocalMux
    port map (
            O => \N__27261\,
            I => neopxl_color_5
        );

    \I__4745\ : LocalMux
    port map (
            O => \N__27258\,
            I => neopxl_color_5
        );

    \I__4744\ : Odrv4
    port map (
            O => \N__27255\,
            I => neopxl_color_5
        );

    \I__4743\ : Odrv4
    port map (
            O => \N__27252\,
            I => neopxl_color_5
        );

    \I__4742\ : SRMux
    port map (
            O => \N__27243\,
            I => \N__27240\
        );

    \I__4741\ : LocalMux
    port map (
            O => \N__27240\,
            I => \N__27237\
        );

    \I__4740\ : Span4Mux_v
    port map (
            O => \N__27237\,
            I => \N__27234\
        );

    \I__4739\ : Sp12to4
    port map (
            O => \N__27234\,
            I => \N__27231\
        );

    \I__4738\ : Odrv12
    port map (
            O => \N__27231\,
            I => n22
        );

    \I__4737\ : InMux
    port map (
            O => \N__27228\,
            I => \N__27225\
        );

    \I__4736\ : LocalMux
    port map (
            O => \N__27225\,
            I => \N__27222\
        );

    \I__4735\ : Span4Mux_h
    port map (
            O => \N__27222\,
            I => \N__27219\
        );

    \I__4734\ : Odrv4
    port map (
            O => \N__27219\,
            I => \nx.n1966\
        );

    \I__4733\ : InMux
    port map (
            O => \N__27216\,
            I => \N__27213\
        );

    \I__4732\ : LocalMux
    port map (
            O => \N__27213\,
            I => \N__27209\
        );

    \I__4731\ : CascadeMux
    port map (
            O => \N__27212\,
            I => \N__27206\
        );

    \I__4730\ : Span4Mux_h
    port map (
            O => \N__27209\,
            I => \N__27202\
        );

    \I__4729\ : InMux
    port map (
            O => \N__27206\,
            I => \N__27199\
        );

    \I__4728\ : InMux
    port map (
            O => \N__27205\,
            I => \N__27196\
        );

    \I__4727\ : Odrv4
    port map (
            O => \N__27202\,
            I => \nx.n1899\
        );

    \I__4726\ : LocalMux
    port map (
            O => \N__27199\,
            I => \nx.n1899\
        );

    \I__4725\ : LocalMux
    port map (
            O => \N__27196\,
            I => \nx.n1899\
        );

    \I__4724\ : InMux
    port map (
            O => \N__27189\,
            I => \N__27186\
        );

    \I__4723\ : LocalMux
    port map (
            O => \N__27186\,
            I => \N__27183\
        );

    \I__4722\ : Span4Mux_h
    port map (
            O => \N__27183\,
            I => \N__27180\
        );

    \I__4721\ : Odrv4
    port map (
            O => \N__27180\,
            I => \nx.n1967\
        );

    \I__4720\ : CascadeMux
    port map (
            O => \N__27177\,
            I => \N__27174\
        );

    \I__4719\ : InMux
    port map (
            O => \N__27174\,
            I => \N__27171\
        );

    \I__4718\ : LocalMux
    port map (
            O => \N__27171\,
            I => \N__27167\
        );

    \I__4717\ : CascadeMux
    port map (
            O => \N__27170\,
            I => \N__27164\
        );

    \I__4716\ : Span4Mux_h
    port map (
            O => \N__27167\,
            I => \N__27160\
        );

    \I__4715\ : InMux
    port map (
            O => \N__27164\,
            I => \N__27157\
        );

    \I__4714\ : InMux
    port map (
            O => \N__27163\,
            I => \N__27154\
        );

    \I__4713\ : Odrv4
    port map (
            O => \N__27160\,
            I => \nx.n1900\
        );

    \I__4712\ : LocalMux
    port map (
            O => \N__27157\,
            I => \nx.n1900\
        );

    \I__4711\ : LocalMux
    port map (
            O => \N__27154\,
            I => \nx.n1900\
        );

    \I__4710\ : InMux
    port map (
            O => \N__27147\,
            I => \N__27144\
        );

    \I__4709\ : LocalMux
    port map (
            O => \N__27144\,
            I => \N__27141\
        );

    \I__4708\ : Span4Mux_h
    port map (
            O => \N__27141\,
            I => \N__27138\
        );

    \I__4707\ : Odrv4
    port map (
            O => \N__27138\,
            I => \nx.n1970\
        );

    \I__4706\ : InMux
    port map (
            O => \N__27135\,
            I => \N__27132\
        );

    \I__4705\ : LocalMux
    port map (
            O => \N__27132\,
            I => \N__27128\
        );

    \I__4704\ : CascadeMux
    port map (
            O => \N__27131\,
            I => \N__27124\
        );

    \I__4703\ : Span4Mux_h
    port map (
            O => \N__27128\,
            I => \N__27121\
        );

    \I__4702\ : InMux
    port map (
            O => \N__27127\,
            I => \N__27118\
        );

    \I__4701\ : InMux
    port map (
            O => \N__27124\,
            I => \N__27115\
        );

    \I__4700\ : Odrv4
    port map (
            O => \N__27121\,
            I => \nx.n1903\
        );

    \I__4699\ : LocalMux
    port map (
            O => \N__27118\,
            I => \nx.n1903\
        );

    \I__4698\ : LocalMux
    port map (
            O => \N__27115\,
            I => \nx.n1903\
        );

    \I__4697\ : InMux
    port map (
            O => \N__27108\,
            I => \N__27105\
        );

    \I__4696\ : LocalMux
    port map (
            O => \N__27105\,
            I => \N__27102\
        );

    \I__4695\ : Span4Mux_h
    port map (
            O => \N__27102\,
            I => \N__27099\
        );

    \I__4694\ : Odrv4
    port map (
            O => \N__27099\,
            I => \nx.n1972\
        );

    \I__4693\ : CascadeMux
    port map (
            O => \N__27096\,
            I => \N__27093\
        );

    \I__4692\ : InMux
    port map (
            O => \N__27093\,
            I => \N__27090\
        );

    \I__4691\ : LocalMux
    port map (
            O => \N__27090\,
            I => \N__27085\
        );

    \I__4690\ : CascadeMux
    port map (
            O => \N__27089\,
            I => \N__27082\
        );

    \I__4689\ : CascadeMux
    port map (
            O => \N__27088\,
            I => \N__27079\
        );

    \I__4688\ : Span4Mux_h
    port map (
            O => \N__27085\,
            I => \N__27076\
        );

    \I__4687\ : InMux
    port map (
            O => \N__27082\,
            I => \N__27073\
        );

    \I__4686\ : InMux
    port map (
            O => \N__27079\,
            I => \N__27070\
        );

    \I__4685\ : Odrv4
    port map (
            O => \N__27076\,
            I => \nx.n1905\
        );

    \I__4684\ : LocalMux
    port map (
            O => \N__27073\,
            I => \nx.n1905\
        );

    \I__4683\ : LocalMux
    port map (
            O => \N__27070\,
            I => \nx.n1905\
        );

    \I__4682\ : InMux
    port map (
            O => \N__27063\,
            I => \bfn_9_26_0_\
        );

    \I__4681\ : InMux
    port map (
            O => \N__27060\,
            I => \nx.n10848\
        );

    \I__4680\ : InMux
    port map (
            O => \N__27057\,
            I => \nx.n11025\
        );

    \I__4679\ : InMux
    port map (
            O => \N__27054\,
            I => \nx.n11026\
        );

    \I__4678\ : InMux
    port map (
            O => \N__27051\,
            I => \bfn_9_24_0_\
        );

    \I__4677\ : CascadeMux
    port map (
            O => \N__27048\,
            I => \N__27043\
        );

    \I__4676\ : InMux
    port map (
            O => \N__27047\,
            I => \N__27038\
        );

    \I__4675\ : InMux
    port map (
            O => \N__27046\,
            I => \N__27038\
        );

    \I__4674\ : InMux
    port map (
            O => \N__27043\,
            I => \N__27035\
        );

    \I__4673\ : LocalMux
    port map (
            O => \N__27038\,
            I => \N__27032\
        );

    \I__4672\ : LocalMux
    port map (
            O => \N__27035\,
            I => \nx.n2792\
        );

    \I__4671\ : Odrv12
    port map (
            O => \N__27032\,
            I => \nx.n2792\
        );

    \I__4670\ : InMux
    port map (
            O => \N__27027\,
            I => \N__27024\
        );

    \I__4669\ : LocalMux
    port map (
            O => \N__27024\,
            I => \N__27021\
        );

    \I__4668\ : Span12Mux_v
    port map (
            O => \N__27021\,
            I => \N__27018\
        );

    \I__4667\ : Odrv12
    port map (
            O => \N__27018\,
            I => neopxl_color_prev_5
        );

    \I__4666\ : InMux
    port map (
            O => \N__27015\,
            I => \nx.n11016\
        );

    \I__4665\ : InMux
    port map (
            O => \N__27012\,
            I => \nx.n11017\
        );

    \I__4664\ : InMux
    port map (
            O => \N__27009\,
            I => \nx.n11018\
        );

    \I__4663\ : InMux
    port map (
            O => \N__27006\,
            I => \bfn_9_23_0_\
        );

    \I__4662\ : InMux
    port map (
            O => \N__27003\,
            I => \nx.n11020\
        );

    \I__4661\ : InMux
    port map (
            O => \N__27000\,
            I => \N__26997\
        );

    \I__4660\ : LocalMux
    port map (
            O => \N__26997\,
            I => \N__26994\
        );

    \I__4659\ : Odrv4
    port map (
            O => \N__26994\,
            I => \nx.n2859\
        );

    \I__4658\ : InMux
    port map (
            O => \N__26991\,
            I => \nx.n11021\
        );

    \I__4657\ : CascadeMux
    port map (
            O => \N__26988\,
            I => \N__26985\
        );

    \I__4656\ : InMux
    port map (
            O => \N__26985\,
            I => \N__26982\
        );

    \I__4655\ : LocalMux
    port map (
            O => \N__26982\,
            I => \N__26978\
        );

    \I__4654\ : InMux
    port map (
            O => \N__26981\,
            I => \N__26975\
        );

    \I__4653\ : Odrv4
    port map (
            O => \N__26978\,
            I => \nx.n2791\
        );

    \I__4652\ : LocalMux
    port map (
            O => \N__26975\,
            I => \nx.n2791\
        );

    \I__4651\ : InMux
    port map (
            O => \N__26970\,
            I => \N__26967\
        );

    \I__4650\ : LocalMux
    port map (
            O => \N__26967\,
            I => \N__26964\
        );

    \I__4649\ : Odrv4
    port map (
            O => \N__26964\,
            I => \nx.n2858\
        );

    \I__4648\ : InMux
    port map (
            O => \N__26961\,
            I => \nx.n11022\
        );

    \I__4647\ : InMux
    port map (
            O => \N__26958\,
            I => \nx.n11023\
        );

    \I__4646\ : InMux
    port map (
            O => \N__26955\,
            I => \N__26952\
        );

    \I__4645\ : LocalMux
    port map (
            O => \N__26952\,
            I => \N__26949\
        );

    \I__4644\ : Odrv4
    port map (
            O => \N__26949\,
            I => \nx.n2856\
        );

    \I__4643\ : InMux
    port map (
            O => \N__26946\,
            I => \nx.n11024\
        );

    \I__4642\ : InMux
    port map (
            O => \N__26943\,
            I => \nx.n11007\
        );

    \I__4641\ : InMux
    port map (
            O => \N__26940\,
            I => \nx.n11008\
        );

    \I__4640\ : InMux
    port map (
            O => \N__26937\,
            I => \nx.n11009\
        );

    \I__4639\ : InMux
    port map (
            O => \N__26934\,
            I => \nx.n11010\
        );

    \I__4638\ : InMux
    port map (
            O => \N__26931\,
            I => \bfn_9_22_0_\
        );

    \I__4637\ : InMux
    port map (
            O => \N__26928\,
            I => \nx.n11012\
        );

    \I__4636\ : InMux
    port map (
            O => \N__26925\,
            I => \nx.n11013\
        );

    \I__4635\ : InMux
    port map (
            O => \N__26922\,
            I => \nx.n11014\
        );

    \I__4634\ : InMux
    port map (
            O => \N__26919\,
            I => \nx.n11015\
        );

    \I__4633\ : CascadeMux
    port map (
            O => \N__26916\,
            I => \nx.n2791_cascade_\
        );

    \I__4632\ : InMux
    port map (
            O => \N__26913\,
            I => \bfn_9_21_0_\
        );

    \I__4631\ : CascadeMux
    port map (
            O => \N__26910\,
            I => \N__26907\
        );

    \I__4630\ : InMux
    port map (
            O => \N__26907\,
            I => \N__26904\
        );

    \I__4629\ : LocalMux
    port map (
            O => \N__26904\,
            I => \N__26901\
        );

    \I__4628\ : Odrv4
    port map (
            O => \N__26901\,
            I => \nx.n2876\
        );

    \I__4627\ : InMux
    port map (
            O => \N__26898\,
            I => \nx.n11004\
        );

    \I__4626\ : InMux
    port map (
            O => \N__26895\,
            I => \N__26892\
        );

    \I__4625\ : LocalMux
    port map (
            O => \N__26892\,
            I => \N__26889\
        );

    \I__4624\ : Odrv4
    port map (
            O => \N__26889\,
            I => \nx.n2875\
        );

    \I__4623\ : InMux
    port map (
            O => \N__26886\,
            I => \nx.n11005\
        );

    \I__4622\ : InMux
    port map (
            O => \N__26883\,
            I => \nx.n11006\
        );

    \I__4621\ : InMux
    port map (
            O => \N__26880\,
            I => \N__26877\
        );

    \I__4620\ : LocalMux
    port map (
            O => \N__26877\,
            I => \N__26874\
        );

    \I__4619\ : Span4Mux_h
    port map (
            O => \N__26874\,
            I => \N__26871\
        );

    \I__4618\ : Span4Mux_v
    port map (
            O => \N__26871\,
            I => \N__26867\
        );

    \I__4617\ : InMux
    port map (
            O => \N__26870\,
            I => \N__26864\
        );

    \I__4616\ : Odrv4
    port map (
            O => \N__26867\,
            I => \nx.bit_ctr_2\
        );

    \I__4615\ : LocalMux
    port map (
            O => \N__26864\,
            I => \nx.bit_ctr_2\
        );

    \I__4614\ : InMux
    port map (
            O => \N__26859\,
            I => \N__26856\
        );

    \I__4613\ : LocalMux
    port map (
            O => \N__26856\,
            I => \N__26850\
        );

    \I__4612\ : InMux
    port map (
            O => \N__26855\,
            I => \N__26847\
        );

    \I__4611\ : InMux
    port map (
            O => \N__26854\,
            I => \N__26844\
        );

    \I__4610\ : InMux
    port map (
            O => \N__26853\,
            I => \N__26841\
        );

    \I__4609\ : Span4Mux_v
    port map (
            O => \N__26850\,
            I => \N__26838\
        );

    \I__4608\ : LocalMux
    port map (
            O => \N__26847\,
            I => \N__26831\
        );

    \I__4607\ : LocalMux
    port map (
            O => \N__26844\,
            I => \N__26831\
        );

    \I__4606\ : LocalMux
    port map (
            O => \N__26841\,
            I => \N__26831\
        );

    \I__4605\ : Span4Mux_h
    port map (
            O => \N__26838\,
            I => \N__26826\
        );

    \I__4604\ : Span4Mux_v
    port map (
            O => \N__26831\,
            I => \N__26826\
        );

    \I__4603\ : Odrv4
    port map (
            O => \N__26826\,
            I => \state_3_N_448_1\
        );

    \I__4602\ : CascadeMux
    port map (
            O => \N__26823\,
            I => \N__26820\
        );

    \I__4601\ : InMux
    port map (
            O => \N__26820\,
            I => \N__26817\
        );

    \I__4600\ : LocalMux
    port map (
            O => \N__26817\,
            I => \nx.color_bit_N_642_4\
        );

    \I__4599\ : InMux
    port map (
            O => \N__26814\,
            I => \N__26811\
        );

    \I__4598\ : LocalMux
    port map (
            O => \N__26811\,
            I => \N__26808\
        );

    \I__4597\ : Odrv4
    port map (
            O => \N__26808\,
            I => \nx.n13622\
        );

    \I__4596\ : CascadeMux
    port map (
            O => \N__26805\,
            I => \N__26791\
        );

    \I__4595\ : CascadeMux
    port map (
            O => \N__26804\,
            I => \N__26788\
        );

    \I__4594\ : InMux
    port map (
            O => \N__26803\,
            I => \N__26781\
        );

    \I__4593\ : InMux
    port map (
            O => \N__26802\,
            I => \N__26781\
        );

    \I__4592\ : InMux
    port map (
            O => \N__26801\,
            I => \N__26781\
        );

    \I__4591\ : InMux
    port map (
            O => \N__26800\,
            I => \N__26778\
        );

    \I__4590\ : InMux
    port map (
            O => \N__26799\,
            I => \N__26772\
        );

    \I__4589\ : InMux
    port map (
            O => \N__26798\,
            I => \N__26772\
        );

    \I__4588\ : CascadeMux
    port map (
            O => \N__26797\,
            I => \N__26769\
        );

    \I__4587\ : InMux
    port map (
            O => \N__26796\,
            I => \N__26760\
        );

    \I__4586\ : InMux
    port map (
            O => \N__26795\,
            I => \N__26760\
        );

    \I__4585\ : InMux
    port map (
            O => \N__26794\,
            I => \N__26760\
        );

    \I__4584\ : InMux
    port map (
            O => \N__26791\,
            I => \N__26760\
        );

    \I__4583\ : InMux
    port map (
            O => \N__26788\,
            I => \N__26757\
        );

    \I__4582\ : LocalMux
    port map (
            O => \N__26781\,
            I => \N__26754\
        );

    \I__4581\ : LocalMux
    port map (
            O => \N__26778\,
            I => \N__26751\
        );

    \I__4580\ : InMux
    port map (
            O => \N__26777\,
            I => \N__26748\
        );

    \I__4579\ : LocalMux
    port map (
            O => \N__26772\,
            I => \N__26745\
        );

    \I__4578\ : InMux
    port map (
            O => \N__26769\,
            I => \N__26742\
        );

    \I__4577\ : LocalMux
    port map (
            O => \N__26760\,
            I => \N__26737\
        );

    \I__4576\ : LocalMux
    port map (
            O => \N__26757\,
            I => \N__26737\
        );

    \I__4575\ : Span4Mux_v
    port map (
            O => \N__26754\,
            I => \N__26732\
        );

    \I__4574\ : Span4Mux_h
    port map (
            O => \N__26751\,
            I => \N__26732\
        );

    \I__4573\ : LocalMux
    port map (
            O => \N__26748\,
            I => \N__26725\
        );

    \I__4572\ : Span4Mux_v
    port map (
            O => \N__26745\,
            I => \N__26725\
        );

    \I__4571\ : LocalMux
    port map (
            O => \N__26742\,
            I => \N__26725\
        );

    \I__4570\ : Span4Mux_h
    port map (
            O => \N__26737\,
            I => \N__26720\
        );

    \I__4569\ : Span4Mux_h
    port map (
            O => \N__26732\,
            I => \N__26720\
        );

    \I__4568\ : Odrv4
    port map (
            O => \N__26725\,
            I => state_0_adj_792
        );

    \I__4567\ : Odrv4
    port map (
            O => \N__26720\,
            I => state_0_adj_792
        );

    \I__4566\ : CEMux
    port map (
            O => \N__26715\,
            I => \N__26712\
        );

    \I__4565\ : LocalMux
    port map (
            O => \N__26712\,
            I => \N__26709\
        );

    \I__4564\ : Span4Mux_h
    port map (
            O => \N__26709\,
            I => \N__26705\
        );

    \I__4563\ : InMux
    port map (
            O => \N__26708\,
            I => \N__26702\
        );

    \I__4562\ : Odrv4
    port map (
            O => \N__26705\,
            I => n7671
        );

    \I__4561\ : LocalMux
    port map (
            O => \N__26702\,
            I => n7671
        );

    \I__4560\ : SRMux
    port map (
            O => \N__26697\,
            I => \N__26694\
        );

    \I__4559\ : LocalMux
    port map (
            O => \N__26694\,
            I => \N__26691\
        );

    \I__4558\ : Odrv4
    port map (
            O => \N__26691\,
            I => \nx.n7983\
        );

    \I__4557\ : CascadeMux
    port map (
            O => \N__26688\,
            I => \N__26685\
        );

    \I__4556\ : InMux
    port map (
            O => \N__26685\,
            I => \N__26682\
        );

    \I__4555\ : LocalMux
    port map (
            O => \N__26682\,
            I => \nx.n12817\
        );

    \I__4554\ : CascadeMux
    port map (
            O => \N__26679\,
            I => \nx.n12819_cascade_\
        );

    \I__4553\ : InMux
    port map (
            O => \N__26676\,
            I => \N__26673\
        );

    \I__4552\ : LocalMux
    port map (
            O => \N__26673\,
            I => \nx.n12821\
        );

    \I__4551\ : CascadeMux
    port map (
            O => \N__26670\,
            I => \nx.n3009_cascade_\
        );

    \I__4550\ : InMux
    port map (
            O => \N__26667\,
            I => \N__26664\
        );

    \I__4549\ : LocalMux
    port map (
            O => \N__26664\,
            I => \N__26661\
        );

    \I__4548\ : Odrv12
    port map (
            O => \N__26661\,
            I => \nx.n1971\
        );

    \I__4547\ : CascadeMux
    port map (
            O => \N__26658\,
            I => \N__26655\
        );

    \I__4546\ : InMux
    port map (
            O => \N__26655\,
            I => \N__26650\
        );

    \I__4545\ : CascadeMux
    port map (
            O => \N__26654\,
            I => \N__26647\
        );

    \I__4544\ : InMux
    port map (
            O => \N__26653\,
            I => \N__26644\
        );

    \I__4543\ : LocalMux
    port map (
            O => \N__26650\,
            I => \N__26641\
        );

    \I__4542\ : InMux
    port map (
            O => \N__26647\,
            I => \N__26638\
        );

    \I__4541\ : LocalMux
    port map (
            O => \N__26644\,
            I => \N__26635\
        );

    \I__4540\ : Odrv4
    port map (
            O => \N__26641\,
            I => \nx.n1904\
        );

    \I__4539\ : LocalMux
    port map (
            O => \N__26638\,
            I => \nx.n1904\
        );

    \I__4538\ : Odrv4
    port map (
            O => \N__26635\,
            I => \nx.n1904\
        );

    \I__4537\ : InMux
    port map (
            O => \N__26628\,
            I => \N__26625\
        );

    \I__4536\ : LocalMux
    port map (
            O => \N__26625\,
            I => n13360
        );

    \I__4535\ : CascadeMux
    port map (
            O => \N__26622\,
            I => \n13361_cascade_\
        );

    \I__4534\ : IoInMux
    port map (
            O => \N__26619\,
            I => \N__26616\
        );

    \I__4533\ : LocalMux
    port map (
            O => \N__26616\,
            I => \N__26613\
        );

    \I__4532\ : Span12Mux_s1_v
    port map (
            O => \N__26613\,
            I => \N__26610\
        );

    \I__4531\ : Odrv12
    port map (
            O => \N__26610\,
            I => \LED_c\
        );

    \I__4530\ : InMux
    port map (
            O => \N__26607\,
            I => \N__26600\
        );

    \I__4529\ : InMux
    port map (
            O => \N__26606\,
            I => \N__26600\
        );

    \I__4528\ : InMux
    port map (
            O => \N__26605\,
            I => \N__26597\
        );

    \I__4527\ : LocalMux
    port map (
            O => \N__26600\,
            I => \N__26593\
        );

    \I__4526\ : LocalMux
    port map (
            O => \N__26597\,
            I => \N__26590\
        );

    \I__4525\ : InMux
    port map (
            O => \N__26596\,
            I => \N__26587\
        );

    \I__4524\ : Span12Mux_s8_h
    port map (
            O => \N__26593\,
            I => \N__26584\
        );

    \I__4523\ : Span4Mux_h
    port map (
            O => \N__26590\,
            I => \N__26581\
        );

    \I__4522\ : LocalMux
    port map (
            O => \N__26587\,
            I => neopxl_color_12
        );

    \I__4521\ : Odrv12
    port map (
            O => \N__26584\,
            I => neopxl_color_12
        );

    \I__4520\ : Odrv4
    port map (
            O => \N__26581\,
            I => neopxl_color_12
        );

    \I__4519\ : InMux
    port map (
            O => \N__26574\,
            I => \N__26571\
        );

    \I__4518\ : LocalMux
    port map (
            O => \N__26571\,
            I => \nx.n59\
        );

    \I__4517\ : CascadeMux
    port map (
            O => \N__26568\,
            I => \nx.n61_cascade_\
        );

    \I__4516\ : InMux
    port map (
            O => \N__26565\,
            I => \N__26561\
        );

    \I__4515\ : InMux
    port map (
            O => \N__26564\,
            I => \N__26558\
        );

    \I__4514\ : LocalMux
    port map (
            O => \N__26561\,
            I => \N__26555\
        );

    \I__4513\ : LocalMux
    port map (
            O => \N__26558\,
            I => \nx.n11153\
        );

    \I__4512\ : Odrv4
    port map (
            O => \N__26555\,
            I => \nx.n11153\
        );

    \I__4511\ : InMux
    port map (
            O => \N__26550\,
            I => \nx.n10845\
        );

    \I__4510\ : InMux
    port map (
            O => \N__26547\,
            I => \nx.n10846\
        );

    \I__4509\ : CascadeMux
    port map (
            O => \N__26544\,
            I => \N__26540\
        );

    \I__4508\ : InMux
    port map (
            O => \N__26543\,
            I => \N__26537\
        );

    \I__4507\ : InMux
    port map (
            O => \N__26540\,
            I => \N__26534\
        );

    \I__4506\ : LocalMux
    port map (
            O => \N__26537\,
            I => \N__26531\
        );

    \I__4505\ : LocalMux
    port map (
            O => \N__26534\,
            I => \nx.n1895\
        );

    \I__4504\ : Odrv4
    port map (
            O => \N__26531\,
            I => \nx.n1895\
        );

    \I__4503\ : InMux
    port map (
            O => \N__26526\,
            I => \nx.n10847\
        );

    \I__4502\ : InMux
    port map (
            O => \N__26523\,
            I => \N__26520\
        );

    \I__4501\ : LocalMux
    port map (
            O => \N__26520\,
            I => \N__26517\
        );

    \I__4500\ : Odrv4
    port map (
            O => \N__26517\,
            I => \nx.n24\
        );

    \I__4499\ : CascadeMux
    port map (
            O => \N__26514\,
            I => \N__26511\
        );

    \I__4498\ : InMux
    port map (
            O => \N__26511\,
            I => \N__26508\
        );

    \I__4497\ : LocalMux
    port map (
            O => \N__26508\,
            I => \nx.n1963\
        );

    \I__4496\ : CascadeMux
    port map (
            O => \N__26505\,
            I => \N__26501\
        );

    \I__4495\ : CascadeMux
    port map (
            O => \N__26504\,
            I => \N__26497\
        );

    \I__4494\ : InMux
    port map (
            O => \N__26501\,
            I => \N__26494\
        );

    \I__4493\ : InMux
    port map (
            O => \N__26500\,
            I => \N__26491\
        );

    \I__4492\ : InMux
    port map (
            O => \N__26497\,
            I => \N__26488\
        );

    \I__4491\ : LocalMux
    port map (
            O => \N__26494\,
            I => \N__26485\
        );

    \I__4490\ : LocalMux
    port map (
            O => \N__26491\,
            I => \nx.n1896\
        );

    \I__4489\ : LocalMux
    port map (
            O => \N__26488\,
            I => \nx.n1896\
        );

    \I__4488\ : Odrv4
    port map (
            O => \N__26485\,
            I => \nx.n1896\
        );

    \I__4487\ : CascadeMux
    port map (
            O => \N__26478\,
            I => \nx.n1995_cascade_\
        );

    \I__4486\ : InMux
    port map (
            O => \N__26475\,
            I => \N__26472\
        );

    \I__4485\ : LocalMux
    port map (
            O => \N__26472\,
            I => \nx.n1965\
        );

    \I__4484\ : CascadeMux
    port map (
            O => \N__26469\,
            I => \N__26464\
        );

    \I__4483\ : CascadeMux
    port map (
            O => \N__26468\,
            I => \N__26461\
        );

    \I__4482\ : CascadeMux
    port map (
            O => \N__26467\,
            I => \N__26458\
        );

    \I__4481\ : InMux
    port map (
            O => \N__26464\,
            I => \N__26455\
        );

    \I__4480\ : InMux
    port map (
            O => \N__26461\,
            I => \N__26452\
        );

    \I__4479\ : InMux
    port map (
            O => \N__26458\,
            I => \N__26449\
        );

    \I__4478\ : LocalMux
    port map (
            O => \N__26455\,
            I => \nx.n1898\
        );

    \I__4477\ : LocalMux
    port map (
            O => \N__26452\,
            I => \nx.n1898\
        );

    \I__4476\ : LocalMux
    port map (
            O => \N__26449\,
            I => \nx.n1898\
        );

    \I__4475\ : InMux
    port map (
            O => \N__26442\,
            I => \N__26439\
        );

    \I__4474\ : LocalMux
    port map (
            O => \N__26439\,
            I => \nx.n1964\
        );

    \I__4473\ : CascadeMux
    port map (
            O => \N__26436\,
            I => \N__26433\
        );

    \I__4472\ : InMux
    port map (
            O => \N__26433\,
            I => \N__26428\
        );

    \I__4471\ : InMux
    port map (
            O => \N__26432\,
            I => \N__26423\
        );

    \I__4470\ : InMux
    port map (
            O => \N__26431\,
            I => \N__26423\
        );

    \I__4469\ : LocalMux
    port map (
            O => \N__26428\,
            I => \nx.n1897\
        );

    \I__4468\ : LocalMux
    port map (
            O => \N__26423\,
            I => \nx.n1897\
        );

    \I__4467\ : CascadeMux
    port map (
            O => \N__26418\,
            I => \N__26413\
        );

    \I__4466\ : InMux
    port map (
            O => \N__26417\,
            I => \N__26408\
        );

    \I__4465\ : InMux
    port map (
            O => \N__26416\,
            I => \N__26408\
        );

    \I__4464\ : InMux
    port map (
            O => \N__26413\,
            I => \N__26405\
        );

    \I__4463\ : LocalMux
    port map (
            O => \N__26408\,
            I => \nx.n1906\
        );

    \I__4462\ : LocalMux
    port map (
            O => \N__26405\,
            I => \nx.n1906\
        );

    \I__4461\ : InMux
    port map (
            O => \N__26400\,
            I => \N__26397\
        );

    \I__4460\ : LocalMux
    port map (
            O => \N__26397\,
            I => \nx.n1973\
        );

    \I__4459\ : InMux
    port map (
            O => \N__26394\,
            I => \nx.n10836\
        );

    \I__4458\ : InMux
    port map (
            O => \N__26391\,
            I => \nx.n10837\
        );

    \I__4457\ : InMux
    port map (
            O => \N__26388\,
            I => \nx.n10838\
        );

    \I__4456\ : InMux
    port map (
            O => \N__26385\,
            I => \nx.n10839\
        );

    \I__4455\ : InMux
    port map (
            O => \N__26382\,
            I => \bfn_7_28_0_\
        );

    \I__4454\ : InMux
    port map (
            O => \N__26379\,
            I => \nx.n10841\
        );

    \I__4453\ : InMux
    port map (
            O => \N__26376\,
            I => \nx.n10842\
        );

    \I__4452\ : InMux
    port map (
            O => \N__26373\,
            I => \nx.n10843\
        );

    \I__4451\ : InMux
    port map (
            O => \N__26370\,
            I => \nx.n10844\
        );

    \I__4450\ : CascadeMux
    port map (
            O => \N__26367\,
            I => \nx.n28_adj_679_cascade_\
        );

    \I__4449\ : InMux
    port map (
            O => \N__26364\,
            I => \N__26361\
        );

    \I__4448\ : LocalMux
    port map (
            O => \N__26361\,
            I => \nx.n16_adj_678\
        );

    \I__4447\ : CascadeMux
    port map (
            O => \N__26358\,
            I => \nx.n1928_cascade_\
        );

    \I__4446\ : InMux
    port map (
            O => \N__26355\,
            I => \N__26350\
        );

    \I__4445\ : InMux
    port map (
            O => \N__26354\,
            I => \N__26345\
        );

    \I__4444\ : InMux
    port map (
            O => \N__26353\,
            I => \N__26342\
        );

    \I__4443\ : LocalMux
    port map (
            O => \N__26350\,
            I => \N__26339\
        );

    \I__4442\ : InMux
    port map (
            O => \N__26349\,
            I => \N__26334\
        );

    \I__4441\ : InMux
    port map (
            O => \N__26348\,
            I => \N__26334\
        );

    \I__4440\ : LocalMux
    port map (
            O => \N__26345\,
            I => \nx.bit_ctr_16\
        );

    \I__4439\ : LocalMux
    port map (
            O => \N__26342\,
            I => \nx.bit_ctr_16\
        );

    \I__4438\ : Odrv4
    port map (
            O => \N__26339\,
            I => \nx.bit_ctr_16\
        );

    \I__4437\ : LocalMux
    port map (
            O => \N__26334\,
            I => \nx.bit_ctr_16\
        );

    \I__4436\ : InMux
    port map (
            O => \N__26325\,
            I => \N__26322\
        );

    \I__4435\ : LocalMux
    port map (
            O => \N__26322\,
            I => \N__26319\
        );

    \I__4434\ : Odrv4
    port map (
            O => \N__26319\,
            I => \nx.n1977\
        );

    \I__4433\ : InMux
    port map (
            O => \N__26316\,
            I => \bfn_7_27_0_\
        );

    \I__4432\ : CascadeMux
    port map (
            O => \N__26313\,
            I => \N__26310\
        );

    \I__4431\ : InMux
    port map (
            O => \N__26310\,
            I => \N__26305\
        );

    \I__4430\ : CascadeMux
    port map (
            O => \N__26309\,
            I => \N__26302\
        );

    \I__4429\ : InMux
    port map (
            O => \N__26308\,
            I => \N__26299\
        );

    \I__4428\ : LocalMux
    port map (
            O => \N__26305\,
            I => \N__26296\
        );

    \I__4427\ : InMux
    port map (
            O => \N__26302\,
            I => \N__26293\
        );

    \I__4426\ : LocalMux
    port map (
            O => \N__26299\,
            I => \nx.n1909\
        );

    \I__4425\ : Odrv4
    port map (
            O => \N__26296\,
            I => \nx.n1909\
        );

    \I__4424\ : LocalMux
    port map (
            O => \N__26293\,
            I => \nx.n1909\
        );

    \I__4423\ : InMux
    port map (
            O => \N__26286\,
            I => \N__26283\
        );

    \I__4422\ : LocalMux
    port map (
            O => \N__26283\,
            I => \nx.n1976\
        );

    \I__4421\ : InMux
    port map (
            O => \N__26280\,
            I => \nx.n10833\
        );

    \I__4420\ : CascadeMux
    port map (
            O => \N__26277\,
            I => \N__26272\
        );

    \I__4419\ : InMux
    port map (
            O => \N__26276\,
            I => \N__26267\
        );

    \I__4418\ : InMux
    port map (
            O => \N__26275\,
            I => \N__26267\
        );

    \I__4417\ : InMux
    port map (
            O => \N__26272\,
            I => \N__26264\
        );

    \I__4416\ : LocalMux
    port map (
            O => \N__26267\,
            I => \nx.n1908\
        );

    \I__4415\ : LocalMux
    port map (
            O => \N__26264\,
            I => \nx.n1908\
        );

    \I__4414\ : InMux
    port map (
            O => \N__26259\,
            I => \N__26256\
        );

    \I__4413\ : LocalMux
    port map (
            O => \N__26256\,
            I => \nx.n1975\
        );

    \I__4412\ : InMux
    port map (
            O => \N__26253\,
            I => \nx.n10834\
        );

    \I__4411\ : CascadeMux
    port map (
            O => \N__26250\,
            I => \N__26245\
        );

    \I__4410\ : InMux
    port map (
            O => \N__26249\,
            I => \N__26240\
        );

    \I__4409\ : InMux
    port map (
            O => \N__26248\,
            I => \N__26240\
        );

    \I__4408\ : InMux
    port map (
            O => \N__26245\,
            I => \N__26237\
        );

    \I__4407\ : LocalMux
    port map (
            O => \N__26240\,
            I => \nx.n1907\
        );

    \I__4406\ : LocalMux
    port map (
            O => \N__26237\,
            I => \nx.n1907\
        );

    \I__4405\ : CascadeMux
    port map (
            O => \N__26232\,
            I => \N__26229\
        );

    \I__4404\ : InMux
    port map (
            O => \N__26229\,
            I => \N__26226\
        );

    \I__4403\ : LocalMux
    port map (
            O => \N__26226\,
            I => \nx.n1974\
        );

    \I__4402\ : InMux
    port map (
            O => \N__26223\,
            I => \nx.n10835\
        );

    \I__4401\ : CascadeMux
    port map (
            O => \N__26220\,
            I => \N__26216\
        );

    \I__4400\ : InMux
    port map (
            O => \N__26219\,
            I => \N__26213\
        );

    \I__4399\ : InMux
    port map (
            O => \N__26216\,
            I => \N__26210\
        );

    \I__4398\ : LocalMux
    port map (
            O => \N__26213\,
            I => \N__26204\
        );

    \I__4397\ : LocalMux
    port map (
            O => \N__26210\,
            I => \N__26201\
        );

    \I__4396\ : InMux
    port map (
            O => \N__26209\,
            I => \N__26198\
        );

    \I__4395\ : InMux
    port map (
            O => \N__26208\,
            I => \N__26195\
        );

    \I__4394\ : InMux
    port map (
            O => \N__26207\,
            I => \N__26192\
        );

    \I__4393\ : Span4Mux_v
    port map (
            O => \N__26204\,
            I => \N__26187\
        );

    \I__4392\ : Span4Mux_v
    port map (
            O => \N__26201\,
            I => \N__26187\
        );

    \I__4391\ : LocalMux
    port map (
            O => \N__26198\,
            I => \N__26182\
        );

    \I__4390\ : LocalMux
    port map (
            O => \N__26195\,
            I => \N__26182\
        );

    \I__4389\ : LocalMux
    port map (
            O => \N__26192\,
            I => neopxl_color_6
        );

    \I__4388\ : Odrv4
    port map (
            O => \N__26187\,
            I => neopxl_color_6
        );

    \I__4387\ : Odrv12
    port map (
            O => \N__26182\,
            I => neopxl_color_6
        );

    \I__4386\ : CascadeMux
    port map (
            O => \N__26175\,
            I => \N__26171\
        );

    \I__4385\ : InMux
    port map (
            O => \N__26174\,
            I => \N__26167\
        );

    \I__4384\ : InMux
    port map (
            O => \N__26171\,
            I => \N__26162\
        );

    \I__4383\ : InMux
    port map (
            O => \N__26170\,
            I => \N__26162\
        );

    \I__4382\ : LocalMux
    port map (
            O => \N__26167\,
            I => \N__26156\
        );

    \I__4381\ : LocalMux
    port map (
            O => \N__26162\,
            I => \N__26156\
        );

    \I__4380\ : InMux
    port map (
            O => \N__26161\,
            I => \N__26152\
        );

    \I__4379\ : Span4Mux_v
    port map (
            O => \N__26156\,
            I => \N__26149\
        );

    \I__4378\ : InMux
    port map (
            O => \N__26155\,
            I => \N__26146\
        );

    \I__4377\ : LocalMux
    port map (
            O => \N__26152\,
            I => \nx.bit_ctr_0\
        );

    \I__4376\ : Odrv4
    port map (
            O => \N__26149\,
            I => \nx.bit_ctr_0\
        );

    \I__4375\ : LocalMux
    port map (
            O => \N__26146\,
            I => \nx.bit_ctr_0\
        );

    \I__4374\ : InMux
    port map (
            O => \N__26139\,
            I => \N__26136\
        );

    \I__4373\ : LocalMux
    port map (
            O => \N__26136\,
            I => \N__26133\
        );

    \I__4372\ : Odrv12
    port map (
            O => \N__26133\,
            I => \nx.n13373\
        );

    \I__4371\ : InMux
    port map (
            O => \N__26130\,
            I => \N__26123\
        );

    \I__4370\ : InMux
    port map (
            O => \N__26129\,
            I => \N__26114\
        );

    \I__4369\ : InMux
    port map (
            O => \N__26128\,
            I => \N__26114\
        );

    \I__4368\ : InMux
    port map (
            O => \N__26127\,
            I => \N__26114\
        );

    \I__4367\ : InMux
    port map (
            O => \N__26126\,
            I => \N__26114\
        );

    \I__4366\ : LocalMux
    port map (
            O => \N__26123\,
            I => neopxl_color_7
        );

    \I__4365\ : LocalMux
    port map (
            O => \N__26114\,
            I => neopxl_color_7
        );

    \I__4364\ : SRMux
    port map (
            O => \N__26109\,
            I => \N__26106\
        );

    \I__4363\ : LocalMux
    port map (
            O => \N__26106\,
            I => \N__26103\
        );

    \I__4362\ : Odrv12
    port map (
            O => \N__26103\,
            I => n22_adj_793
        );

    \I__4361\ : CascadeMux
    port map (
            O => \N__26100\,
            I => \nx.n26_cascade_\
        );

    \I__4360\ : InMux
    port map (
            O => \N__26097\,
            I => \N__26094\
        );

    \I__4359\ : LocalMux
    port map (
            O => \N__26094\,
            I => \nx.n20\
        );

    \I__4358\ : CascadeMux
    port map (
            O => \N__26091\,
            I => \nx.n11912_cascade_\
        );

    \I__4357\ : InMux
    port map (
            O => \N__26088\,
            I => \N__26085\
        );

    \I__4356\ : LocalMux
    port map (
            O => \N__26085\,
            I => \nx.n58\
        );

    \I__4355\ : CascadeMux
    port map (
            O => \N__26082\,
            I => \N__26078\
        );

    \I__4354\ : InMux
    port map (
            O => \N__26081\,
            I => \N__26075\
        );

    \I__4353\ : InMux
    port map (
            O => \N__26078\,
            I => \N__26070\
        );

    \I__4352\ : LocalMux
    port map (
            O => \N__26075\,
            I => \N__26065\
        );

    \I__4351\ : InMux
    port map (
            O => \N__26074\,
            I => \N__26060\
        );

    \I__4350\ : InMux
    port map (
            O => \N__26073\,
            I => \N__26060\
        );

    \I__4349\ : LocalMux
    port map (
            O => \N__26070\,
            I => \N__26057\
        );

    \I__4348\ : InMux
    port map (
            O => \N__26069\,
            I => \N__26054\
        );

    \I__4347\ : InMux
    port map (
            O => \N__26068\,
            I => \N__26051\
        );

    \I__4346\ : Span4Mux_h
    port map (
            O => \N__26065\,
            I => \N__26046\
        );

    \I__4345\ : LocalMux
    port map (
            O => \N__26060\,
            I => \N__26046\
        );

    \I__4344\ : Sp12to4
    port map (
            O => \N__26057\,
            I => \N__26041\
        );

    \I__4343\ : LocalMux
    port map (
            O => \N__26054\,
            I => \N__26041\
        );

    \I__4342\ : LocalMux
    port map (
            O => \N__26051\,
            I => \nx.bit_ctr_29\
        );

    \I__4341\ : Odrv4
    port map (
            O => \N__26046\,
            I => \nx.bit_ctr_29\
        );

    \I__4340\ : Odrv12
    port map (
            O => \N__26041\,
            I => \nx.bit_ctr_29\
        );

    \I__4339\ : CascadeMux
    port map (
            O => \N__26034\,
            I => \N__26030\
        );

    \I__4338\ : CascadeMux
    port map (
            O => \N__26033\,
            I => \N__26026\
        );

    \I__4337\ : InMux
    port map (
            O => \N__26030\,
            I => \N__26022\
        );

    \I__4336\ : InMux
    port map (
            O => \N__26029\,
            I => \N__26017\
        );

    \I__4335\ : InMux
    port map (
            O => \N__26026\,
            I => \N__26017\
        );

    \I__4334\ : InMux
    port map (
            O => \N__26025\,
            I => \N__26013\
        );

    \I__4333\ : LocalMux
    port map (
            O => \N__26022\,
            I => \N__26010\
        );

    \I__4332\ : LocalMux
    port map (
            O => \N__26017\,
            I => \N__26007\
        );

    \I__4331\ : InMux
    port map (
            O => \N__26016\,
            I => \N__26004\
        );

    \I__4330\ : LocalMux
    port map (
            O => \N__26013\,
            I => \N__26001\
        );

    \I__4329\ : Span4Mux_h
    port map (
            O => \N__26010\,
            I => \N__25996\
        );

    \I__4328\ : Span4Mux_h
    port map (
            O => \N__26007\,
            I => \N__25996\
        );

    \I__4327\ : LocalMux
    port map (
            O => \N__26004\,
            I => \nx.bit_ctr_30\
        );

    \I__4326\ : Odrv12
    port map (
            O => \N__26001\,
            I => \nx.bit_ctr_30\
        );

    \I__4325\ : Odrv4
    port map (
            O => \N__25996\,
            I => \nx.bit_ctr_30\
        );

    \I__4324\ : CascadeMux
    port map (
            O => \N__25989\,
            I => \N__25986\
        );

    \I__4323\ : InMux
    port map (
            O => \N__25986\,
            I => \N__25979\
        );

    \I__4322\ : InMux
    port map (
            O => \N__25985\,
            I => \N__25979\
        );

    \I__4321\ : CascadeMux
    port map (
            O => \N__25984\,
            I => \N__25975\
        );

    \I__4320\ : LocalMux
    port map (
            O => \N__25979\,
            I => \N__25971\
        );

    \I__4319\ : InMux
    port map (
            O => \N__25978\,
            I => \N__25968\
        );

    \I__4318\ : InMux
    port map (
            O => \N__25975\,
            I => \N__25965\
        );

    \I__4317\ : InMux
    port map (
            O => \N__25974\,
            I => \N__25962\
        );

    \I__4316\ : Span4Mux_h
    port map (
            O => \N__25971\,
            I => \N__25959\
        );

    \I__4315\ : LocalMux
    port map (
            O => \N__25968\,
            I => \N__25954\
        );

    \I__4314\ : LocalMux
    port map (
            O => \N__25965\,
            I => \N__25954\
        );

    \I__4313\ : LocalMux
    port map (
            O => \N__25962\,
            I => \nx.bit_ctr_31\
        );

    \I__4312\ : Odrv4
    port map (
            O => \N__25959\,
            I => \nx.bit_ctr_31\
        );

    \I__4311\ : Odrv12
    port map (
            O => \N__25954\,
            I => \nx.bit_ctr_31\
        );

    \I__4310\ : InMux
    port map (
            O => \N__25947\,
            I => \N__25944\
        );

    \I__4309\ : LocalMux
    port map (
            O => \N__25944\,
            I => \nx.n9803\
        );

    \I__4308\ : InMux
    port map (
            O => \N__25941\,
            I => \N__25935\
        );

    \I__4307\ : InMux
    port map (
            O => \N__25940\,
            I => \N__25928\
        );

    \I__4306\ : InMux
    port map (
            O => \N__25939\,
            I => \N__25928\
        );

    \I__4305\ : InMux
    port map (
            O => \N__25938\,
            I => \N__25928\
        );

    \I__4304\ : LocalMux
    port map (
            O => \N__25935\,
            I => \N__25922\
        );

    \I__4303\ : LocalMux
    port map (
            O => \N__25928\,
            I => \N__25919\
        );

    \I__4302\ : InMux
    port map (
            O => \N__25927\,
            I => \N__25914\
        );

    \I__4301\ : InMux
    port map (
            O => \N__25926\,
            I => \N__25914\
        );

    \I__4300\ : InMux
    port map (
            O => \N__25925\,
            I => \N__25911\
        );

    \I__4299\ : Span4Mux_v
    port map (
            O => \N__25922\,
            I => \N__25904\
        );

    \I__4298\ : Span4Mux_v
    port map (
            O => \N__25919\,
            I => \N__25904\
        );

    \I__4297\ : LocalMux
    port map (
            O => \N__25914\,
            I => \N__25904\
        );

    \I__4296\ : LocalMux
    port map (
            O => \N__25911\,
            I => \nx.bit_ctr_27\
        );

    \I__4295\ : Odrv4
    port map (
            O => \N__25904\,
            I => \nx.bit_ctr_27\
        );

    \I__4294\ : InMux
    port map (
            O => \N__25899\,
            I => \N__25890\
        );

    \I__4293\ : InMux
    port map (
            O => \N__25898\,
            I => \N__25885\
        );

    \I__4292\ : InMux
    port map (
            O => \N__25897\,
            I => \N__25885\
        );

    \I__4291\ : InMux
    port map (
            O => \N__25896\,
            I => \N__25878\
        );

    \I__4290\ : InMux
    port map (
            O => \N__25895\,
            I => \N__25878\
        );

    \I__4289\ : InMux
    port map (
            O => \N__25894\,
            I => \N__25878\
        );

    \I__4288\ : InMux
    port map (
            O => \N__25893\,
            I => \N__25875\
        );

    \I__4287\ : LocalMux
    port map (
            O => \N__25890\,
            I => \N__25872\
        );

    \I__4286\ : LocalMux
    port map (
            O => \N__25885\,
            I => \N__25869\
        );

    \I__4285\ : LocalMux
    port map (
            O => \N__25878\,
            I => \N__25866\
        );

    \I__4284\ : LocalMux
    port map (
            O => \N__25875\,
            I => \nx.bit_ctr_28\
        );

    \I__4283\ : Odrv4
    port map (
            O => \N__25872\,
            I => \nx.bit_ctr_28\
        );

    \I__4282\ : Odrv12
    port map (
            O => \N__25869\,
            I => \nx.bit_ctr_28\
        );

    \I__4281\ : Odrv4
    port map (
            O => \N__25866\,
            I => \nx.bit_ctr_28\
        );

    \I__4280\ : CascadeMux
    port map (
            O => \N__25857\,
            I => \N__25852\
        );

    \I__4279\ : CascadeMux
    port map (
            O => \N__25856\,
            I => \N__25849\
        );

    \I__4278\ : CascadeMux
    port map (
            O => \N__25855\,
            I => \N__25846\
        );

    \I__4277\ : InMux
    port map (
            O => \N__25852\,
            I => \N__25843\
        );

    \I__4276\ : InMux
    port map (
            O => \N__25849\,
            I => \N__25840\
        );

    \I__4275\ : InMux
    port map (
            O => \N__25846\,
            I => \N__25837\
        );

    \I__4274\ : LocalMux
    port map (
            O => \N__25843\,
            I => \nx.n11912\
        );

    \I__4273\ : LocalMux
    port map (
            O => \N__25840\,
            I => \nx.n11912\
        );

    \I__4272\ : LocalMux
    port map (
            O => \N__25837\,
            I => \nx.n11912\
        );

    \I__4271\ : InMux
    port map (
            O => \N__25830\,
            I => \N__25824\
        );

    \I__4270\ : InMux
    port map (
            O => \N__25829\,
            I => \N__25819\
        );

    \I__4269\ : InMux
    port map (
            O => \N__25828\,
            I => \N__25819\
        );

    \I__4268\ : InMux
    port map (
            O => \N__25827\,
            I => \N__25816\
        );

    \I__4267\ : LocalMux
    port map (
            O => \N__25824\,
            I => \nx.n708\
        );

    \I__4266\ : LocalMux
    port map (
            O => \N__25819\,
            I => \nx.n708\
        );

    \I__4265\ : LocalMux
    port map (
            O => \N__25816\,
            I => \nx.n708\
        );

    \I__4264\ : CascadeMux
    port map (
            O => \N__25809\,
            I => \N__25804\
        );

    \I__4263\ : InMux
    port map (
            O => \N__25808\,
            I => \N__25801\
        );

    \I__4262\ : InMux
    port map (
            O => \N__25807\,
            I => \N__25796\
        );

    \I__4261\ : InMux
    port map (
            O => \N__25804\,
            I => \N__25796\
        );

    \I__4260\ : LocalMux
    port map (
            O => \N__25801\,
            I => \N__25791\
        );

    \I__4259\ : LocalMux
    port map (
            O => \N__25796\,
            I => \N__25791\
        );

    \I__4258\ : Odrv4
    port map (
            O => \N__25791\,
            I => \nx.n5703\
        );

    \I__4257\ : InMux
    port map (
            O => \N__25788\,
            I => \N__25785\
        );

    \I__4256\ : LocalMux
    port map (
            O => \N__25785\,
            I => \N__25782\
        );

    \I__4255\ : Span4Mux_v
    port map (
            O => \N__25782\,
            I => \N__25779\
        );

    \I__4254\ : Odrv4
    port map (
            O => \N__25779\,
            I => n10_adj_846
        );

    \I__4253\ : InMux
    port map (
            O => \N__25776\,
            I => \N__25773\
        );

    \I__4252\ : LocalMux
    port map (
            O => \N__25773\,
            I => neopxl_color_prev_7
        );

    \I__4251\ : CascadeMux
    port map (
            O => \N__25770\,
            I => \N__25766\
        );

    \I__4250\ : InMux
    port map (
            O => \N__25769\,
            I => \N__25761\
        );

    \I__4249\ : InMux
    port map (
            O => \N__25766\,
            I => \N__25761\
        );

    \I__4248\ : LocalMux
    port map (
            O => \N__25761\,
            I => \N__25758\
        );

    \I__4247\ : Span4Mux_h
    port map (
            O => \N__25758\,
            I => \N__25753\
        );

    \I__4246\ : InMux
    port map (
            O => \N__25757\,
            I => \N__25750\
        );

    \I__4245\ : InMux
    port map (
            O => \N__25756\,
            I => \N__25747\
        );

    \I__4244\ : Span4Mux_v
    port map (
            O => \N__25753\,
            I => \N__25744\
        );

    \I__4243\ : LocalMux
    port map (
            O => \N__25750\,
            I => neopxl_color_15
        );

    \I__4242\ : LocalMux
    port map (
            O => \N__25747\,
            I => neopxl_color_15
        );

    \I__4241\ : Odrv4
    port map (
            O => \N__25744\,
            I => neopxl_color_15
        );

    \I__4240\ : InMux
    port map (
            O => \N__25737\,
            I => \N__25734\
        );

    \I__4239\ : LocalMux
    port map (
            O => \N__25734\,
            I => neopxl_color_prev_15
        );

    \I__4238\ : CascadeMux
    port map (
            O => \N__25731\,
            I => \N__25727\
        );

    \I__4237\ : CascadeMux
    port map (
            O => \N__25730\,
            I => \N__25724\
        );

    \I__4236\ : InMux
    port map (
            O => \N__25727\,
            I => \N__25721\
        );

    \I__4235\ : InMux
    port map (
            O => \N__25724\,
            I => \N__25718\
        );

    \I__4234\ : LocalMux
    port map (
            O => \N__25721\,
            I => \nx.n7497\
        );

    \I__4233\ : LocalMux
    port map (
            O => \N__25718\,
            I => \nx.n7497\
        );

    \I__4232\ : InMux
    port map (
            O => \N__25713\,
            I => \N__25710\
        );

    \I__4231\ : LocalMux
    port map (
            O => \N__25710\,
            I => \nx.n976\
        );

    \I__4230\ : InMux
    port map (
            O => \N__25707\,
            I => \nx.n10738\
        );

    \I__4229\ : CascadeMux
    port map (
            O => \N__25704\,
            I => \N__25701\
        );

    \I__4228\ : InMux
    port map (
            O => \N__25701\,
            I => \N__25698\
        );

    \I__4227\ : LocalMux
    port map (
            O => \N__25698\,
            I => \nx.n7899\
        );

    \I__4226\ : CascadeMux
    port map (
            O => \N__25695\,
            I => \N__25691\
        );

    \I__4225\ : InMux
    port map (
            O => \N__25694\,
            I => \N__25688\
        );

    \I__4224\ : InMux
    port map (
            O => \N__25691\,
            I => \N__25685\
        );

    \I__4223\ : LocalMux
    port map (
            O => \N__25688\,
            I => \nx.n975\
        );

    \I__4222\ : LocalMux
    port map (
            O => \N__25685\,
            I => \nx.n975\
        );

    \I__4221\ : InMux
    port map (
            O => \N__25680\,
            I => \nx.n10739\
        );

    \I__4220\ : InMux
    port map (
            O => \N__25677\,
            I => \N__25671\
        );

    \I__4219\ : InMux
    port map (
            O => \N__25676\,
            I => \N__25671\
        );

    \I__4218\ : LocalMux
    port map (
            O => \N__25671\,
            I => \nx.n974\
        );

    \I__4217\ : InMux
    port map (
            O => \N__25668\,
            I => \nx.n10740\
        );

    \I__4216\ : CascadeMux
    port map (
            O => \N__25665\,
            I => \N__25661\
        );

    \I__4215\ : CascadeMux
    port map (
            O => \N__25664\,
            I => \N__25658\
        );

    \I__4214\ : InMux
    port map (
            O => \N__25661\,
            I => \N__25654\
        );

    \I__4213\ : InMux
    port map (
            O => \N__25658\,
            I => \N__25651\
        );

    \I__4212\ : InMux
    port map (
            O => \N__25657\,
            I => \N__25648\
        );

    \I__4211\ : LocalMux
    port map (
            O => \N__25654\,
            I => \nx.n906\
        );

    \I__4210\ : LocalMux
    port map (
            O => \N__25651\,
            I => \nx.n906\
        );

    \I__4209\ : LocalMux
    port map (
            O => \N__25648\,
            I => \nx.n906\
        );

    \I__4208\ : InMux
    port map (
            O => \N__25641\,
            I => \N__25638\
        );

    \I__4207\ : LocalMux
    port map (
            O => \N__25638\,
            I => \nx.n973\
        );

    \I__4206\ : InMux
    port map (
            O => \N__25635\,
            I => \nx.n10741\
        );

    \I__4205\ : InMux
    port map (
            O => \N__25632\,
            I => \N__25629\
        );

    \I__4204\ : LocalMux
    port map (
            O => \N__25629\,
            I => \nx.n13594\
        );

    \I__4203\ : CascadeMux
    port map (
            O => \N__25626\,
            I => \N__25623\
        );

    \I__4202\ : InMux
    port map (
            O => \N__25623\,
            I => \N__25620\
        );

    \I__4201\ : LocalMux
    port map (
            O => \N__25620\,
            I => \nx.n905\
        );

    \I__4200\ : InMux
    port map (
            O => \N__25617\,
            I => \nx.n10742\
        );

    \I__4199\ : InMux
    port map (
            O => \N__25614\,
            I => \N__25611\
        );

    \I__4198\ : LocalMux
    port map (
            O => \N__25611\,
            I => \N__25607\
        );

    \I__4197\ : InMux
    port map (
            O => \N__25610\,
            I => \N__25604\
        );

    \I__4196\ : Odrv4
    port map (
            O => \N__25607\,
            I => \nx.n4\
        );

    \I__4195\ : LocalMux
    port map (
            O => \N__25604\,
            I => \nx.n4\
        );

    \I__4194\ : CascadeMux
    port map (
            O => \N__25599\,
            I => \N__25596\
        );

    \I__4193\ : InMux
    port map (
            O => \N__25596\,
            I => \N__25589\
        );

    \I__4192\ : InMux
    port map (
            O => \N__25595\,
            I => \N__25589\
        );

    \I__4191\ : InMux
    port map (
            O => \N__25594\,
            I => \N__25586\
        );

    \I__4190\ : LocalMux
    port map (
            O => \N__25589\,
            I => \nx.n807\
        );

    \I__4189\ : LocalMux
    port map (
            O => \N__25586\,
            I => \nx.n807\
        );

    \I__4188\ : CascadeMux
    port map (
            O => \N__25581\,
            I => \N__25576\
        );

    \I__4187\ : InMux
    port map (
            O => \N__25580\,
            I => \N__25571\
        );

    \I__4186\ : InMux
    port map (
            O => \N__25579\,
            I => \N__25571\
        );

    \I__4185\ : InMux
    port map (
            O => \N__25576\,
            I => \N__25568\
        );

    \I__4184\ : LocalMux
    port map (
            O => \N__25571\,
            I => \nx.n11866\
        );

    \I__4183\ : LocalMux
    port map (
            O => \N__25568\,
            I => \nx.n11866\
        );

    \I__4182\ : InMux
    port map (
            O => \N__25563\,
            I => \N__25554\
        );

    \I__4181\ : InMux
    port map (
            O => \N__25562\,
            I => \N__25554\
        );

    \I__4180\ : InMux
    port map (
            O => \N__25561\,
            I => \N__25551\
        );

    \I__4179\ : InMux
    port map (
            O => \N__25560\,
            I => \N__25546\
        );

    \I__4178\ : InMux
    port map (
            O => \N__25559\,
            I => \N__25546\
        );

    \I__4177\ : LocalMux
    port map (
            O => \N__25554\,
            I => \nx.n838\
        );

    \I__4176\ : LocalMux
    port map (
            O => \N__25551\,
            I => \nx.n838\
        );

    \I__4175\ : LocalMux
    port map (
            O => \N__25546\,
            I => \nx.n838\
        );

    \I__4174\ : CascadeMux
    port map (
            O => \N__25539\,
            I => \N__25536\
        );

    \I__4173\ : InMux
    port map (
            O => \N__25536\,
            I => \N__25532\
        );

    \I__4172\ : InMux
    port map (
            O => \N__25535\,
            I => \N__25529\
        );

    \I__4171\ : LocalMux
    port map (
            O => \N__25532\,
            I => \nx.n11868\
        );

    \I__4170\ : LocalMux
    port map (
            O => \N__25529\,
            I => \nx.n11868\
        );

    \I__4169\ : InMux
    port map (
            O => \N__25524\,
            I => \N__25519\
        );

    \I__4168\ : InMux
    port map (
            O => \N__25523\,
            I => \N__25516\
        );

    \I__4167\ : InMux
    port map (
            O => \N__25522\,
            I => \N__25511\
        );

    \I__4166\ : LocalMux
    port map (
            O => \N__25519\,
            I => \N__25506\
        );

    \I__4165\ : LocalMux
    port map (
            O => \N__25516\,
            I => \N__25506\
        );

    \I__4164\ : InMux
    port map (
            O => \N__25515\,
            I => \N__25503\
        );

    \I__4163\ : InMux
    port map (
            O => \N__25514\,
            I => \N__25500\
        );

    \I__4162\ : LocalMux
    port map (
            O => \N__25511\,
            I => \N__25497\
        );

    \I__4161\ : Span4Mux_v
    port map (
            O => \N__25506\,
            I => \N__25494\
        );

    \I__4160\ : LocalMux
    port map (
            O => \N__25503\,
            I => \N__25491\
        );

    \I__4159\ : LocalMux
    port map (
            O => \N__25500\,
            I => \nx.bit_ctr_17\
        );

    \I__4158\ : Odrv4
    port map (
            O => \N__25497\,
            I => \nx.bit_ctr_17\
        );

    \I__4157\ : Odrv4
    port map (
            O => \N__25494\,
            I => \nx.bit_ctr_17\
        );

    \I__4156\ : Odrv12
    port map (
            O => \N__25491\,
            I => \nx.bit_ctr_17\
        );

    \I__4155\ : InMux
    port map (
            O => \N__25482\,
            I => \N__25478\
        );

    \I__4154\ : CascadeMux
    port map (
            O => \N__25481\,
            I => \N__25473\
        );

    \I__4153\ : LocalMux
    port map (
            O => \N__25478\,
            I => \N__25470\
        );

    \I__4152\ : InMux
    port map (
            O => \N__25477\,
            I => \N__25467\
        );

    \I__4151\ : InMux
    port map (
            O => \N__25476\,
            I => \N__25464\
        );

    \I__4150\ : InMux
    port map (
            O => \N__25473\,
            I => \N__25460\
        );

    \I__4149\ : Span4Mux_v
    port map (
            O => \N__25470\,
            I => \N__25455\
        );

    \I__4148\ : LocalMux
    port map (
            O => \N__25467\,
            I => \N__25455\
        );

    \I__4147\ : LocalMux
    port map (
            O => \N__25464\,
            I => \N__25452\
        );

    \I__4146\ : InMux
    port map (
            O => \N__25463\,
            I => \N__25449\
        );

    \I__4145\ : LocalMux
    port map (
            O => \N__25460\,
            I => \N__25446\
        );

    \I__4144\ : Span4Mux_h
    port map (
            O => \N__25455\,
            I => \N__25441\
        );

    \I__4143\ : Span4Mux_h
    port map (
            O => \N__25452\,
            I => \N__25441\
        );

    \I__4142\ : LocalMux
    port map (
            O => \N__25449\,
            I => \nx.bit_ctr_22\
        );

    \I__4141\ : Odrv4
    port map (
            O => \N__25446\,
            I => \nx.bit_ctr_22\
        );

    \I__4140\ : Odrv4
    port map (
            O => \N__25441\,
            I => \nx.bit_ctr_22\
        );

    \I__4139\ : InMux
    port map (
            O => \N__25434\,
            I => \N__25431\
        );

    \I__4138\ : LocalMux
    port map (
            O => \N__25431\,
            I => \N__25428\
        );

    \I__4137\ : Span4Mux_h
    port map (
            O => \N__25428\,
            I => \N__25425\
        );

    \I__4136\ : Odrv4
    port map (
            O => \N__25425\,
            I => \nx.n44_adj_782\
        );

    \I__4135\ : InMux
    port map (
            O => \N__25422\,
            I => \N__25419\
        );

    \I__4134\ : LocalMux
    port map (
            O => \N__25419\,
            I => \nx.n11941\
        );

    \I__4133\ : CascadeMux
    port map (
            O => \N__25416\,
            I => \N__25412\
        );

    \I__4132\ : CascadeMux
    port map (
            O => \N__25415\,
            I => \N__25408\
        );

    \I__4131\ : InMux
    port map (
            O => \N__25412\,
            I => \N__25403\
        );

    \I__4130\ : InMux
    port map (
            O => \N__25411\,
            I => \N__25403\
        );

    \I__4129\ : InMux
    port map (
            O => \N__25408\,
            I => \N__25400\
        );

    \I__4128\ : LocalMux
    port map (
            O => \N__25403\,
            I => \nx.n1008\
        );

    \I__4127\ : LocalMux
    port map (
            O => \N__25400\,
            I => \nx.n1008\
        );

    \I__4126\ : CascadeMux
    port map (
            O => \N__25395\,
            I => \N__25391\
        );

    \I__4125\ : InMux
    port map (
            O => \N__25394\,
            I => \N__25388\
        );

    \I__4124\ : InMux
    port map (
            O => \N__25391\,
            I => \N__25385\
        );

    \I__4123\ : LocalMux
    port map (
            O => \N__25388\,
            I => \nx.n1006\
        );

    \I__4122\ : LocalMux
    port map (
            O => \N__25385\,
            I => \nx.n1006\
        );

    \I__4121\ : CascadeMux
    port map (
            O => \N__25380\,
            I => \nx.n12837_cascade_\
        );

    \I__4120\ : CascadeMux
    port map (
            O => \N__25377\,
            I => \nx.n905_cascade_\
        );

    \I__4119\ : InMux
    port map (
            O => \N__25374\,
            I => \N__25371\
        );

    \I__4118\ : LocalMux
    port map (
            O => \N__25371\,
            I => \nx.n12839\
        );

    \I__4117\ : CascadeMux
    port map (
            O => \N__25368\,
            I => \N__25362\
        );

    \I__4116\ : CascadeMux
    port map (
            O => \N__25367\,
            I => \N__25359\
        );

    \I__4115\ : InMux
    port map (
            O => \N__25366\,
            I => \N__25352\
        );

    \I__4114\ : InMux
    port map (
            O => \N__25365\,
            I => \N__25352\
        );

    \I__4113\ : InMux
    port map (
            O => \N__25362\,
            I => \N__25345\
        );

    \I__4112\ : InMux
    port map (
            O => \N__25359\,
            I => \N__25345\
        );

    \I__4111\ : InMux
    port map (
            O => \N__25358\,
            I => \N__25345\
        );

    \I__4110\ : InMux
    port map (
            O => \N__25357\,
            I => \N__25342\
        );

    \I__4109\ : LocalMux
    port map (
            O => \N__25352\,
            I => \nx.n11174\
        );

    \I__4108\ : LocalMux
    port map (
            O => \N__25345\,
            I => \nx.n11174\
        );

    \I__4107\ : LocalMux
    port map (
            O => \N__25342\,
            I => \nx.n11174\
        );

    \I__4106\ : CascadeMux
    port map (
            O => \N__25335\,
            I => \nx.n11174_cascade_\
        );

    \I__4105\ : CascadeMux
    port map (
            O => \N__25332\,
            I => \N__25329\
        );

    \I__4104\ : InMux
    port map (
            O => \N__25329\,
            I => \N__25323\
        );

    \I__4103\ : InMux
    port map (
            O => \N__25328\,
            I => \N__25320\
        );

    \I__4102\ : InMux
    port map (
            O => \N__25327\,
            I => \N__25317\
        );

    \I__4101\ : InMux
    port map (
            O => \N__25326\,
            I => \N__25314\
        );

    \I__4100\ : LocalMux
    port map (
            O => \N__25323\,
            I => \N__25310\
        );

    \I__4099\ : LocalMux
    port map (
            O => \N__25320\,
            I => \N__25307\
        );

    \I__4098\ : LocalMux
    port map (
            O => \N__25317\,
            I => \N__25302\
        );

    \I__4097\ : LocalMux
    port map (
            O => \N__25314\,
            I => \N__25302\
        );

    \I__4096\ : InMux
    port map (
            O => \N__25313\,
            I => \N__25299\
        );

    \I__4095\ : Span4Mux_h
    port map (
            O => \N__25310\,
            I => \N__25296\
        );

    \I__4094\ : Span4Mux_v
    port map (
            O => \N__25307\,
            I => \N__25291\
        );

    \I__4093\ : Span4Mux_h
    port map (
            O => \N__25302\,
            I => \N__25291\
        );

    \I__4092\ : LocalMux
    port map (
            O => \N__25299\,
            I => \nx.bit_ctr_26\
        );

    \I__4091\ : Odrv4
    port map (
            O => \N__25296\,
            I => \nx.bit_ctr_26\
        );

    \I__4090\ : Odrv4
    port map (
            O => \N__25291\,
            I => \nx.bit_ctr_26\
        );

    \I__4089\ : CascadeMux
    port map (
            O => \N__25284\,
            I => \N__25281\
        );

    \I__4088\ : InMux
    port map (
            O => \N__25281\,
            I => \N__25278\
        );

    \I__4087\ : LocalMux
    port map (
            O => \N__25278\,
            I => \N__25275\
        );

    \I__4086\ : Odrv4
    port map (
            O => \N__25275\,
            I => \nx.n977\
        );

    \I__4085\ : InMux
    port map (
            O => \N__25272\,
            I => \bfn_7_22_0_\
        );

    \I__4084\ : InMux
    port map (
            O => \N__25269\,
            I => \N__25265\
        );

    \I__4083\ : CascadeMux
    port map (
            O => \N__25268\,
            I => \N__25262\
        );

    \I__4082\ : LocalMux
    port map (
            O => \N__25265\,
            I => \N__25259\
        );

    \I__4081\ : InMux
    port map (
            O => \N__25262\,
            I => \N__25255\
        );

    \I__4080\ : Span4Mux_h
    port map (
            O => \N__25259\,
            I => \N__25252\
        );

    \I__4079\ : InMux
    port map (
            O => \N__25258\,
            I => \N__25249\
        );

    \I__4078\ : LocalMux
    port map (
            O => \N__25255\,
            I => \N__25246\
        );

    \I__4077\ : Odrv4
    port map (
            O => \N__25252\,
            I => timer_28
        );

    \I__4076\ : LocalMux
    port map (
            O => \N__25249\,
            I => timer_28
        );

    \I__4075\ : Odrv4
    port map (
            O => \N__25246\,
            I => timer_28
        );

    \I__4074\ : InMux
    port map (
            O => \N__25239\,
            I => \N__25221\
        );

    \I__4073\ : InMux
    port map (
            O => \N__25238\,
            I => \N__25213\
        );

    \I__4072\ : InMux
    port map (
            O => \N__25237\,
            I => \N__25208\
        );

    \I__4071\ : InMux
    port map (
            O => \N__25236\,
            I => \N__25208\
        );

    \I__4070\ : InMux
    port map (
            O => \N__25235\,
            I => \N__25201\
        );

    \I__4069\ : InMux
    port map (
            O => \N__25234\,
            I => \N__25201\
        );

    \I__4068\ : InMux
    port map (
            O => \N__25233\,
            I => \N__25201\
        );

    \I__4067\ : InMux
    port map (
            O => \N__25232\,
            I => \N__25194\
        );

    \I__4066\ : InMux
    port map (
            O => \N__25231\,
            I => \N__25194\
        );

    \I__4065\ : InMux
    port map (
            O => \N__25230\,
            I => \N__25194\
        );

    \I__4064\ : InMux
    port map (
            O => \N__25229\,
            I => \N__25185\
        );

    \I__4063\ : InMux
    port map (
            O => \N__25228\,
            I => \N__25185\
        );

    \I__4062\ : InMux
    port map (
            O => \N__25227\,
            I => \N__25185\
        );

    \I__4061\ : InMux
    port map (
            O => \N__25226\,
            I => \N__25185\
        );

    \I__4060\ : InMux
    port map (
            O => \N__25225\,
            I => \N__25180\
        );

    \I__4059\ : InMux
    port map (
            O => \N__25224\,
            I => \N__25180\
        );

    \I__4058\ : LocalMux
    port map (
            O => \N__25221\,
            I => \N__25173\
        );

    \I__4057\ : InMux
    port map (
            O => \N__25220\,
            I => \N__25170\
        );

    \I__4056\ : InMux
    port map (
            O => \N__25219\,
            I => \N__25167\
        );

    \I__4055\ : InMux
    port map (
            O => \N__25218\,
            I => \N__25158\
        );

    \I__4054\ : InMux
    port map (
            O => \N__25217\,
            I => \N__25158\
        );

    \I__4053\ : InMux
    port map (
            O => \N__25216\,
            I => \N__25158\
        );

    \I__4052\ : LocalMux
    port map (
            O => \N__25213\,
            I => \N__25152\
        );

    \I__4051\ : LocalMux
    port map (
            O => \N__25208\,
            I => \N__25143\
        );

    \I__4050\ : LocalMux
    port map (
            O => \N__25201\,
            I => \N__25143\
        );

    \I__4049\ : LocalMux
    port map (
            O => \N__25194\,
            I => \N__25143\
        );

    \I__4048\ : LocalMux
    port map (
            O => \N__25185\,
            I => \N__25143\
        );

    \I__4047\ : LocalMux
    port map (
            O => \N__25180\,
            I => \N__25140\
        );

    \I__4046\ : InMux
    port map (
            O => \N__25179\,
            I => \N__25131\
        );

    \I__4045\ : InMux
    port map (
            O => \N__25178\,
            I => \N__25131\
        );

    \I__4044\ : InMux
    port map (
            O => \N__25177\,
            I => \N__25131\
        );

    \I__4043\ : InMux
    port map (
            O => \N__25176\,
            I => \N__25131\
        );

    \I__4042\ : Span4Mux_s3_h
    port map (
            O => \N__25173\,
            I => \N__25126\
        );

    \I__4041\ : LocalMux
    port map (
            O => \N__25170\,
            I => \N__25126\
        );

    \I__4040\ : LocalMux
    port map (
            O => \N__25167\,
            I => \N__25123\
        );

    \I__4039\ : InMux
    port map (
            O => \N__25166\,
            I => \N__25118\
        );

    \I__4038\ : InMux
    port map (
            O => \N__25165\,
            I => \N__25118\
        );

    \I__4037\ : LocalMux
    port map (
            O => \N__25158\,
            I => \N__25113\
        );

    \I__4036\ : InMux
    port map (
            O => \N__25157\,
            I => \N__25110\
        );

    \I__4035\ : InMux
    port map (
            O => \N__25156\,
            I => \N__25107\
        );

    \I__4034\ : InMux
    port map (
            O => \N__25155\,
            I => \N__25104\
        );

    \I__4033\ : Span4Mux_v
    port map (
            O => \N__25152\,
            I => \N__25095\
        );

    \I__4032\ : Span4Mux_v
    port map (
            O => \N__25143\,
            I => \N__25095\
        );

    \I__4031\ : Span4Mux_s1_h
    port map (
            O => \N__25140\,
            I => \N__25095\
        );

    \I__4030\ : LocalMux
    port map (
            O => \N__25131\,
            I => \N__25095\
        );

    \I__4029\ : Span4Mux_v
    port map (
            O => \N__25126\,
            I => \N__25088\
        );

    \I__4028\ : Span4Mux_h
    port map (
            O => \N__25123\,
            I => \N__25088\
        );

    \I__4027\ : LocalMux
    port map (
            O => \N__25118\,
            I => \N__25088\
        );

    \I__4026\ : InMux
    port map (
            O => \N__25117\,
            I => \N__25083\
        );

    \I__4025\ : InMux
    port map (
            O => \N__25116\,
            I => \N__25083\
        );

    \I__4024\ : Odrv12
    port map (
            O => \N__25113\,
            I => n11353
        );

    \I__4023\ : LocalMux
    port map (
            O => \N__25110\,
            I => n11353
        );

    \I__4022\ : LocalMux
    port map (
            O => \N__25107\,
            I => n11353
        );

    \I__4021\ : LocalMux
    port map (
            O => \N__25104\,
            I => n11353
        );

    \I__4020\ : Odrv4
    port map (
            O => \N__25095\,
            I => n11353
        );

    \I__4019\ : Odrv4
    port map (
            O => \N__25088\,
            I => n11353
        );

    \I__4018\ : LocalMux
    port map (
            O => \N__25083\,
            I => n11353
        );

    \I__4017\ : InMux
    port map (
            O => \N__25068\,
            I => \N__25064\
        );

    \I__4016\ : InMux
    port map (
            O => \N__25067\,
            I => \N__25061\
        );

    \I__4015\ : LocalMux
    port map (
            O => \N__25064\,
            I => \N__25058\
        );

    \I__4014\ : LocalMux
    port map (
            O => \N__25061\,
            I => neo_pixel_transmitter_t0_28
        );

    \I__4013\ : Odrv4
    port map (
            O => \N__25058\,
            I => neo_pixel_transmitter_t0_28
        );

    \I__4012\ : InMux
    port map (
            O => \N__25053\,
            I => \N__25050\
        );

    \I__4011\ : LocalMux
    port map (
            O => \N__25050\,
            I => n9_adj_847
        );

    \I__4010\ : SRMux
    port map (
            O => \N__25047\,
            I => \N__25044\
        );

    \I__4009\ : LocalMux
    port map (
            O => \N__25044\,
            I => \N__25041\
        );

    \I__4008\ : Span4Mux_v
    port map (
            O => \N__25041\,
            I => \N__25038\
        );

    \I__4007\ : Span4Mux_h
    port map (
            O => \N__25038\,
            I => \N__25035\
        );

    \I__4006\ : Odrv4
    port map (
            O => \N__25035\,
            I => \current_pin_7__N_153\
        );

    \I__4005\ : InMux
    port map (
            O => \N__25032\,
            I => \N__25029\
        );

    \I__4004\ : LocalMux
    port map (
            O => \N__25029\,
            I => neopxl_color_prev_14
        );

    \I__4003\ : CascadeMux
    port map (
            O => \N__25026\,
            I => \N__25020\
        );

    \I__4002\ : InMux
    port map (
            O => \N__25025\,
            I => \N__25017\
        );

    \I__4001\ : InMux
    port map (
            O => \N__25024\,
            I => \N__25010\
        );

    \I__4000\ : InMux
    port map (
            O => \N__25023\,
            I => \N__25010\
        );

    \I__3999\ : InMux
    port map (
            O => \N__25020\,
            I => \N__25010\
        );

    \I__3998\ : LocalMux
    port map (
            O => \N__25017\,
            I => \N__25007\
        );

    \I__3997\ : LocalMux
    port map (
            O => \N__25010\,
            I => neopxl_color_13
        );

    \I__3996\ : Odrv4
    port map (
            O => \N__25007\,
            I => neopxl_color_13
        );

    \I__3995\ : InMux
    port map (
            O => \N__25002\,
            I => \N__24999\
        );

    \I__3994\ : LocalMux
    port map (
            O => \N__24999\,
            I => neopxl_color_prev_13
        );

    \I__3993\ : InMux
    port map (
            O => \N__24996\,
            I => \N__24993\
        );

    \I__3992\ : LocalMux
    port map (
            O => \N__24993\,
            I => n11_adj_845
        );

    \I__3991\ : InMux
    port map (
            O => \N__24990\,
            I => \N__24987\
        );

    \I__3990\ : LocalMux
    port map (
            O => \N__24987\,
            I => neopxl_color_prev_4
        );

    \I__3989\ : InMux
    port map (
            O => \N__24984\,
            I => \N__24980\
        );

    \I__3988\ : CascadeMux
    port map (
            O => \N__24983\,
            I => \N__24975\
        );

    \I__3987\ : LocalMux
    port map (
            O => \N__24980\,
            I => \N__24972\
        );

    \I__3986\ : InMux
    port map (
            O => \N__24979\,
            I => \N__24965\
        );

    \I__3985\ : InMux
    port map (
            O => \N__24978\,
            I => \N__24965\
        );

    \I__3984\ : InMux
    port map (
            O => \N__24975\,
            I => \N__24965\
        );

    \I__3983\ : Span4Mux_h
    port map (
            O => \N__24972\,
            I => \N__24962\
        );

    \I__3982\ : LocalMux
    port map (
            O => \N__24965\,
            I => neopxl_color_14
        );

    \I__3981\ : Odrv4
    port map (
            O => \N__24962\,
            I => neopxl_color_14
        );

    \I__3980\ : CascadeMux
    port map (
            O => \N__24957\,
            I => \N__24952\
        );

    \I__3979\ : CascadeMux
    port map (
            O => \N__24956\,
            I => \N__24949\
        );

    \I__3978\ : InMux
    port map (
            O => \N__24955\,
            I => \N__24946\
        );

    \I__3977\ : InMux
    port map (
            O => \N__24952\,
            I => \N__24937\
        );

    \I__3976\ : InMux
    port map (
            O => \N__24949\,
            I => \N__24934\
        );

    \I__3975\ : LocalMux
    port map (
            O => \N__24946\,
            I => \N__24930\
        );

    \I__3974\ : InMux
    port map (
            O => \N__24945\,
            I => \N__24927\
        );

    \I__3973\ : InMux
    port map (
            O => \N__24944\,
            I => \N__24920\
        );

    \I__3972\ : InMux
    port map (
            O => \N__24943\,
            I => \N__24920\
        );

    \I__3971\ : InMux
    port map (
            O => \N__24942\,
            I => \N__24920\
        );

    \I__3970\ : InMux
    port map (
            O => \N__24941\,
            I => \N__24915\
        );

    \I__3969\ : InMux
    port map (
            O => \N__24940\,
            I => \N__24915\
        );

    \I__3968\ : LocalMux
    port map (
            O => \N__24937\,
            I => \N__24912\
        );

    \I__3967\ : LocalMux
    port map (
            O => \N__24934\,
            I => \N__24909\
        );

    \I__3966\ : InMux
    port map (
            O => \N__24933\,
            I => \N__24904\
        );

    \I__3965\ : Span4Mux_h
    port map (
            O => \N__24930\,
            I => \N__24895\
        );

    \I__3964\ : LocalMux
    port map (
            O => \N__24927\,
            I => \N__24895\
        );

    \I__3963\ : LocalMux
    port map (
            O => \N__24920\,
            I => \N__24895\
        );

    \I__3962\ : LocalMux
    port map (
            O => \N__24915\,
            I => \N__24895\
        );

    \I__3961\ : Span4Mux_h
    port map (
            O => \N__24912\,
            I => \N__24892\
        );

    \I__3960\ : Span4Mux_h
    port map (
            O => \N__24909\,
            I => \N__24889\
        );

    \I__3959\ : InMux
    port map (
            O => \N__24908\,
            I => \N__24884\
        );

    \I__3958\ : InMux
    port map (
            O => \N__24907\,
            I => \N__24884\
        );

    \I__3957\ : LocalMux
    port map (
            O => \N__24904\,
            I => \nx.neo_pixel_transmitter_done\
        );

    \I__3956\ : Odrv4
    port map (
            O => \N__24895\,
            I => \nx.neo_pixel_transmitter_done\
        );

    \I__3955\ : Odrv4
    port map (
            O => \N__24892\,
            I => \nx.neo_pixel_transmitter_done\
        );

    \I__3954\ : Odrv4
    port map (
            O => \N__24889\,
            I => \nx.neo_pixel_transmitter_done\
        );

    \I__3953\ : LocalMux
    port map (
            O => \N__24884\,
            I => \nx.neo_pixel_transmitter_done\
        );

    \I__3952\ : IoInMux
    port map (
            O => \N__24873\,
            I => \N__24870\
        );

    \I__3951\ : LocalMux
    port map (
            O => \N__24870\,
            I => \N__24867\
        );

    \I__3950\ : Odrv12
    port map (
            O => \N__24867\,
            I => \NEOPXL_c\
        );

    \I__3949\ : CEMux
    port map (
            O => \N__24864\,
            I => \N__24861\
        );

    \I__3948\ : LocalMux
    port map (
            O => \N__24861\,
            I => \N__24858\
        );

    \I__3947\ : Odrv12
    port map (
            O => \N__24858\,
            I => \nx.n11988\
        );

    \I__3946\ : SRMux
    port map (
            O => \N__24855\,
            I => \N__24852\
        );

    \I__3945\ : LocalMux
    port map (
            O => \N__24852\,
            I => \N__24849\
        );

    \I__3944\ : Odrv4
    port map (
            O => \N__24849\,
            I => \nx.n12451\
        );

    \I__3943\ : InMux
    port map (
            O => \N__24846\,
            I => \N__24843\
        );

    \I__3942\ : LocalMux
    port map (
            O => \N__24843\,
            I => \N__24839\
        );

    \I__3941\ : InMux
    port map (
            O => \N__24842\,
            I => \N__24836\
        );

    \I__3940\ : Span4Mux_v
    port map (
            O => \N__24839\,
            I => \N__24833\
        );

    \I__3939\ : LocalMux
    port map (
            O => \N__24836\,
            I => \nx.bit_ctr_1\
        );

    \I__3938\ : Odrv4
    port map (
            O => \N__24833\,
            I => \nx.bit_ctr_1\
        );

    \I__3937\ : InMux
    port map (
            O => \N__24828\,
            I => \N__24825\
        );

    \I__3936\ : LocalMux
    port map (
            O => \N__24825\,
            I => \nx.n13364\
        );

    \I__3935\ : CascadeMux
    port map (
            O => \N__24822\,
            I => \nx.n11156_cascade_\
        );

    \I__3934\ : InMux
    port map (
            O => \N__24819\,
            I => \N__24816\
        );

    \I__3933\ : LocalMux
    port map (
            O => \N__24816\,
            I => \nx.n13363\
        );

    \I__3932\ : CascadeMux
    port map (
            O => \N__24813\,
            I => \nx.n13619_cascade_\
        );

    \I__3931\ : InMux
    port map (
            O => \N__24810\,
            I => \N__24807\
        );

    \I__3930\ : LocalMux
    port map (
            O => \N__24807\,
            I => \nx.n11156\
        );

    \I__3929\ : InMux
    port map (
            O => \N__24804\,
            I => \N__24801\
        );

    \I__3928\ : LocalMux
    port map (
            O => \N__24801\,
            I => \N__24798\
        );

    \I__3927\ : Span4Mux_h
    port map (
            O => \N__24798\,
            I => \N__24795\
        );

    \I__3926\ : Odrv4
    port map (
            O => \N__24795\,
            I => n11966
        );

    \I__3925\ : IoInMux
    port map (
            O => \N__24792\,
            I => \N__24789\
        );

    \I__3924\ : LocalMux
    port map (
            O => \N__24789\,
            I => \N__24786\
        );

    \I__3923\ : Span4Mux_s2_h
    port map (
            O => \N__24786\,
            I => \N__24783\
        );

    \I__3922\ : Span4Mux_h
    port map (
            O => \N__24783\,
            I => \N__24779\
        );

    \I__3921\ : InMux
    port map (
            O => \N__24782\,
            I => \N__24776\
        );

    \I__3920\ : Odrv4
    port map (
            O => \N__24779\,
            I => pin_oe_2
        );

    \I__3919\ : LocalMux
    port map (
            O => \N__24776\,
            I => pin_oe_2
        );

    \I__3918\ : InMux
    port map (
            O => \N__24771\,
            I => \N__24768\
        );

    \I__3917\ : LocalMux
    port map (
            O => \N__24768\,
            I => \nx.n13372\
        );

    \I__3916\ : CascadeMux
    port map (
            O => \N__24765\,
            I => \N__24760\
        );

    \I__3915\ : InMux
    port map (
            O => \N__24764\,
            I => \N__24757\
        );

    \I__3914\ : InMux
    port map (
            O => \N__24763\,
            I => \N__24754\
        );

    \I__3913\ : InMux
    port map (
            O => \N__24760\,
            I => \N__24750\
        );

    \I__3912\ : LocalMux
    port map (
            O => \N__24757\,
            I => \N__24747\
        );

    \I__3911\ : LocalMux
    port map (
            O => \N__24754\,
            I => \N__24744\
        );

    \I__3910\ : InMux
    port map (
            O => \N__24753\,
            I => \N__24740\
        );

    \I__3909\ : LocalMux
    port map (
            O => \N__24750\,
            I => \N__24737\
        );

    \I__3908\ : Span12Mux_s5_h
    port map (
            O => \N__24747\,
            I => \N__24734\
        );

    \I__3907\ : Span4Mux_v
    port map (
            O => \N__24744\,
            I => \N__24731\
        );

    \I__3906\ : InMux
    port map (
            O => \N__24743\,
            I => \N__24728\
        );

    \I__3905\ : LocalMux
    port map (
            O => \N__24740\,
            I => \nx.bit_ctr_18\
        );

    \I__3904\ : Odrv12
    port map (
            O => \N__24737\,
            I => \nx.bit_ctr_18\
        );

    \I__3903\ : Odrv12
    port map (
            O => \N__24734\,
            I => \nx.bit_ctr_18\
        );

    \I__3902\ : Odrv4
    port map (
            O => \N__24731\,
            I => \nx.bit_ctr_18\
        );

    \I__3901\ : LocalMux
    port map (
            O => \N__24728\,
            I => \nx.bit_ctr_18\
        );

    \I__3900\ : CascadeMux
    port map (
            O => \N__24717\,
            I => \N__24714\
        );

    \I__3899\ : InMux
    port map (
            O => \N__24714\,
            I => \N__24711\
        );

    \I__3898\ : LocalMux
    port map (
            O => \N__24711\,
            I => \N__24708\
        );

    \I__3897\ : Span4Mux_h
    port map (
            O => \N__24708\,
            I => \N__24705\
        );

    \I__3896\ : Odrv4
    port map (
            O => \N__24705\,
            I => \nx.n48_adj_778\
        );

    \I__3895\ : InMux
    port map (
            O => \N__24702\,
            I => \N__24699\
        );

    \I__3894\ : LocalMux
    port map (
            O => \N__24699\,
            I => \nx.n18_adj_716\
        );

    \I__3893\ : InMux
    port map (
            O => \N__24696\,
            I => \N__24691\
        );

    \I__3892\ : InMux
    port map (
            O => \N__24695\,
            I => \N__24688\
        );

    \I__3891\ : InMux
    port map (
            O => \N__24694\,
            I => \N__24685\
        );

    \I__3890\ : LocalMux
    port map (
            O => \N__24691\,
            I => \nx.n1799\
        );

    \I__3889\ : LocalMux
    port map (
            O => \N__24688\,
            I => \nx.n1799\
        );

    \I__3888\ : LocalMux
    port map (
            O => \N__24685\,
            I => \nx.n1799\
        );

    \I__3887\ : CascadeMux
    port map (
            O => \N__24678\,
            I => \N__24675\
        );

    \I__3886\ : InMux
    port map (
            O => \N__24675\,
            I => \N__24670\
        );

    \I__3885\ : InMux
    port map (
            O => \N__24674\,
            I => \N__24667\
        );

    \I__3884\ : InMux
    port map (
            O => \N__24673\,
            I => \N__24664\
        );

    \I__3883\ : LocalMux
    port map (
            O => \N__24670\,
            I => \N__24661\
        );

    \I__3882\ : LocalMux
    port map (
            O => \N__24667\,
            I => \nx.n1805\
        );

    \I__3881\ : LocalMux
    port map (
            O => \N__24664\,
            I => \nx.n1805\
        );

    \I__3880\ : Odrv4
    port map (
            O => \N__24661\,
            I => \nx.n1805\
        );

    \I__3879\ : InMux
    port map (
            O => \N__24654\,
            I => \N__24651\
        );

    \I__3878\ : LocalMux
    port map (
            O => \N__24651\,
            I => \nx.n24_adj_717\
        );

    \I__3877\ : InMux
    port map (
            O => \N__24648\,
            I => \N__24644\
        );

    \I__3876\ : InMux
    port map (
            O => \N__24647\,
            I => \N__24641\
        );

    \I__3875\ : LocalMux
    port map (
            O => \N__24644\,
            I => \N__24635\
        );

    \I__3874\ : LocalMux
    port map (
            O => \N__24641\,
            I => \N__24635\
        );

    \I__3873\ : InMux
    port map (
            O => \N__24640\,
            I => \N__24632\
        );

    \I__3872\ : Odrv4
    port map (
            O => \N__24635\,
            I => \nx.n1798\
        );

    \I__3871\ : LocalMux
    port map (
            O => \N__24632\,
            I => \nx.n1798\
        );

    \I__3870\ : InMux
    port map (
            O => \N__24627\,
            I => \N__24622\
        );

    \I__3869\ : InMux
    port map (
            O => \N__24626\,
            I => \N__24619\
        );

    \I__3868\ : InMux
    port map (
            O => \N__24625\,
            I => \N__24616\
        );

    \I__3867\ : LocalMux
    port map (
            O => \N__24622\,
            I => \N__24613\
        );

    \I__3866\ : LocalMux
    port map (
            O => \N__24619\,
            I => \nx.n1808\
        );

    \I__3865\ : LocalMux
    port map (
            O => \N__24616\,
            I => \nx.n1808\
        );

    \I__3864\ : Odrv4
    port map (
            O => \N__24613\,
            I => \nx.n1808\
        );

    \I__3863\ : CascadeMux
    port map (
            O => \N__24606\,
            I => \nx.n26_adj_719_cascade_\
        );

    \I__3862\ : InMux
    port map (
            O => \N__24603\,
            I => \N__24598\
        );

    \I__3861\ : InMux
    port map (
            O => \N__24602\,
            I => \N__24595\
        );

    \I__3860\ : InMux
    port map (
            O => \N__24601\,
            I => \N__24592\
        );

    \I__3859\ : LocalMux
    port map (
            O => \N__24598\,
            I => \N__24589\
        );

    \I__3858\ : LocalMux
    port map (
            O => \N__24595\,
            I => \nx.n1809\
        );

    \I__3857\ : LocalMux
    port map (
            O => \N__24592\,
            I => \nx.n1809\
        );

    \I__3856\ : Odrv4
    port map (
            O => \N__24589\,
            I => \nx.n1809\
        );

    \I__3855\ : InMux
    port map (
            O => \N__24582\,
            I => \N__24577\
        );

    \I__3854\ : InMux
    port map (
            O => \N__24581\,
            I => \N__24574\
        );

    \I__3853\ : InMux
    port map (
            O => \N__24580\,
            I => \N__24571\
        );

    \I__3852\ : LocalMux
    port map (
            O => \N__24577\,
            I => \N__24568\
        );

    \I__3851\ : LocalMux
    port map (
            O => \N__24574\,
            I => \nx.n1803\
        );

    \I__3850\ : LocalMux
    port map (
            O => \N__24571\,
            I => \nx.n1803\
        );

    \I__3849\ : Odrv4
    port map (
            O => \N__24568\,
            I => \nx.n1803\
        );

    \I__3848\ : InMux
    port map (
            O => \N__24561\,
            I => \N__24556\
        );

    \I__3847\ : InMux
    port map (
            O => \N__24560\,
            I => \N__24553\
        );

    \I__3846\ : InMux
    port map (
            O => \N__24559\,
            I => \N__24550\
        );

    \I__3845\ : LocalMux
    port map (
            O => \N__24556\,
            I => \nx.n1800\
        );

    \I__3844\ : LocalMux
    port map (
            O => \N__24553\,
            I => \nx.n1800\
        );

    \I__3843\ : LocalMux
    port map (
            O => \N__24550\,
            I => \nx.n1800\
        );

    \I__3842\ : CascadeMux
    port map (
            O => \N__24543\,
            I => \nx.n9717_cascade_\
        );

    \I__3841\ : InMux
    port map (
            O => \N__24540\,
            I => \N__24535\
        );

    \I__3840\ : InMux
    port map (
            O => \N__24539\,
            I => \N__24532\
        );

    \I__3839\ : InMux
    port map (
            O => \N__24538\,
            I => \N__24529\
        );

    \I__3838\ : LocalMux
    port map (
            O => \N__24535\,
            I => \nx.n1796\
        );

    \I__3837\ : LocalMux
    port map (
            O => \N__24532\,
            I => \nx.n1796\
        );

    \I__3836\ : LocalMux
    port map (
            O => \N__24529\,
            I => \nx.n1796\
        );

    \I__3835\ : InMux
    port map (
            O => \N__24522\,
            I => \N__24519\
        );

    \I__3834\ : LocalMux
    port map (
            O => \N__24519\,
            I => \nx.n22_adj_718\
        );

    \I__3833\ : CascadeMux
    port map (
            O => \N__24516\,
            I => \N__24501\
        );

    \I__3832\ : CascadeMux
    port map (
            O => \N__24515\,
            I => \N__24498\
        );

    \I__3831\ : CascadeMux
    port map (
            O => \N__24514\,
            I => \N__24495\
        );

    \I__3830\ : CascadeMux
    port map (
            O => \N__24513\,
            I => \N__24492\
        );

    \I__3829\ : CascadeMux
    port map (
            O => \N__24512\,
            I => \N__24489\
        );

    \I__3828\ : CascadeMux
    port map (
            O => \N__24511\,
            I => \N__24486\
        );

    \I__3827\ : CascadeMux
    port map (
            O => \N__24510\,
            I => \N__24483\
        );

    \I__3826\ : CascadeMux
    port map (
            O => \N__24509\,
            I => \N__24480\
        );

    \I__3825\ : CascadeMux
    port map (
            O => \N__24508\,
            I => \N__24477\
        );

    \I__3824\ : CascadeMux
    port map (
            O => \N__24507\,
            I => \N__24474\
        );

    \I__3823\ : CascadeMux
    port map (
            O => \N__24506\,
            I => \N__24471\
        );

    \I__3822\ : CascadeMux
    port map (
            O => \N__24505\,
            I => \N__24468\
        );

    \I__3821\ : CascadeMux
    port map (
            O => \N__24504\,
            I => \N__24465\
        );

    \I__3820\ : InMux
    port map (
            O => \N__24501\,
            I => \N__24458\
        );

    \I__3819\ : InMux
    port map (
            O => \N__24498\,
            I => \N__24458\
        );

    \I__3818\ : InMux
    port map (
            O => \N__24495\,
            I => \N__24458\
        );

    \I__3817\ : InMux
    port map (
            O => \N__24492\,
            I => \N__24451\
        );

    \I__3816\ : InMux
    port map (
            O => \N__24489\,
            I => \N__24451\
        );

    \I__3815\ : InMux
    port map (
            O => \N__24486\,
            I => \N__24451\
        );

    \I__3814\ : InMux
    port map (
            O => \N__24483\,
            I => \N__24443\
        );

    \I__3813\ : InMux
    port map (
            O => \N__24480\,
            I => \N__24443\
        );

    \I__3812\ : InMux
    port map (
            O => \N__24477\,
            I => \N__24443\
        );

    \I__3811\ : InMux
    port map (
            O => \N__24474\,
            I => \N__24434\
        );

    \I__3810\ : InMux
    port map (
            O => \N__24471\,
            I => \N__24434\
        );

    \I__3809\ : InMux
    port map (
            O => \N__24468\,
            I => \N__24434\
        );

    \I__3808\ : InMux
    port map (
            O => \N__24465\,
            I => \N__24434\
        );

    \I__3807\ : LocalMux
    port map (
            O => \N__24458\,
            I => \N__24429\
        );

    \I__3806\ : LocalMux
    port map (
            O => \N__24451\,
            I => \N__24429\
        );

    \I__3805\ : InMux
    port map (
            O => \N__24450\,
            I => \N__24426\
        );

    \I__3804\ : LocalMux
    port map (
            O => \N__24443\,
            I => \nx.n1829\
        );

    \I__3803\ : LocalMux
    port map (
            O => \N__24434\,
            I => \nx.n1829\
        );

    \I__3802\ : Odrv4
    port map (
            O => \N__24429\,
            I => \nx.n1829\
        );

    \I__3801\ : LocalMux
    port map (
            O => \N__24426\,
            I => \nx.n1829\
        );

    \I__3800\ : CascadeMux
    port map (
            O => \N__24417\,
            I => \N__24413\
        );

    \I__3799\ : CascadeMux
    port map (
            O => \N__24416\,
            I => \N__24410\
        );

    \I__3798\ : InMux
    port map (
            O => \N__24413\,
            I => \N__24407\
        );

    \I__3797\ : InMux
    port map (
            O => \N__24410\,
            I => \N__24404\
        );

    \I__3796\ : LocalMux
    port map (
            O => \N__24407\,
            I => \N__24399\
        );

    \I__3795\ : LocalMux
    port map (
            O => \N__24404\,
            I => \N__24399\
        );

    \I__3794\ : Odrv4
    port map (
            O => \N__24399\,
            I => \nx.n13605\
        );

    \I__3793\ : IoInMux
    port map (
            O => \N__24396\,
            I => \N__24393\
        );

    \I__3792\ : LocalMux
    port map (
            O => \N__24393\,
            I => \N__24390\
        );

    \I__3791\ : Span12Mux_s1_h
    port map (
            O => \N__24390\,
            I => \N__24387\
        );

    \I__3790\ : Span12Mux_h
    port map (
            O => \N__24387\,
            I => \N__24384\
        );

    \I__3789\ : Span12Mux_v
    port map (
            O => \N__24384\,
            I => \N__24380\
        );

    \I__3788\ : InMux
    port map (
            O => \N__24383\,
            I => \N__24377\
        );

    \I__3787\ : Odrv12
    port map (
            O => \N__24380\,
            I => pin_oe_7
        );

    \I__3786\ : LocalMux
    port map (
            O => \N__24377\,
            I => pin_oe_7
        );

    \I__3785\ : InMux
    port map (
            O => \N__24372\,
            I => \N__24367\
        );

    \I__3784\ : InMux
    port map (
            O => \N__24371\,
            I => \N__24364\
        );

    \I__3783\ : InMux
    port map (
            O => \N__24370\,
            I => \N__24361\
        );

    \I__3782\ : LocalMux
    port map (
            O => \N__24367\,
            I => \N__24358\
        );

    \I__3781\ : LocalMux
    port map (
            O => \N__24364\,
            I => \nx.n1804\
        );

    \I__3780\ : LocalMux
    port map (
            O => \N__24361\,
            I => \nx.n1804\
        );

    \I__3779\ : Odrv4
    port map (
            O => \N__24358\,
            I => \nx.n1804\
        );

    \I__3778\ : InMux
    port map (
            O => \N__24351\,
            I => \nx.n10824\
        );

    \I__3777\ : InMux
    port map (
            O => \N__24348\,
            I => \nx.n10825\
        );

    \I__3776\ : InMux
    port map (
            O => \N__24345\,
            I => \N__24340\
        );

    \I__3775\ : InMux
    port map (
            O => \N__24344\,
            I => \N__24337\
        );

    \I__3774\ : InMux
    port map (
            O => \N__24343\,
            I => \N__24334\
        );

    \I__3773\ : LocalMux
    port map (
            O => \N__24340\,
            I => \N__24331\
        );

    \I__3772\ : LocalMux
    port map (
            O => \N__24337\,
            I => \nx.n1802\
        );

    \I__3771\ : LocalMux
    port map (
            O => \N__24334\,
            I => \nx.n1802\
        );

    \I__3770\ : Odrv4
    port map (
            O => \N__24331\,
            I => \nx.n1802\
        );

    \I__3769\ : InMux
    port map (
            O => \N__24324\,
            I => \bfn_6_28_0_\
        );

    \I__3768\ : CascadeMux
    port map (
            O => \N__24321\,
            I => \N__24316\
        );

    \I__3767\ : InMux
    port map (
            O => \N__24320\,
            I => \N__24313\
        );

    \I__3766\ : InMux
    port map (
            O => \N__24319\,
            I => \N__24310\
        );

    \I__3765\ : InMux
    port map (
            O => \N__24316\,
            I => \N__24307\
        );

    \I__3764\ : LocalMux
    port map (
            O => \N__24313\,
            I => \nx.n1801\
        );

    \I__3763\ : LocalMux
    port map (
            O => \N__24310\,
            I => \nx.n1801\
        );

    \I__3762\ : LocalMux
    port map (
            O => \N__24307\,
            I => \nx.n1801\
        );

    \I__3761\ : InMux
    port map (
            O => \N__24300\,
            I => \nx.n10827\
        );

    \I__3760\ : InMux
    port map (
            O => \N__24297\,
            I => \nx.n10828\
        );

    \I__3759\ : InMux
    port map (
            O => \N__24294\,
            I => \nx.n10829\
        );

    \I__3758\ : InMux
    port map (
            O => \N__24291\,
            I => \nx.n10830\
        );

    \I__3757\ : InMux
    port map (
            O => \N__24288\,
            I => \N__24283\
        );

    \I__3756\ : InMux
    port map (
            O => \N__24287\,
            I => \N__24280\
        );

    \I__3755\ : InMux
    port map (
            O => \N__24286\,
            I => \N__24277\
        );

    \I__3754\ : LocalMux
    port map (
            O => \N__24283\,
            I => \nx.n1797\
        );

    \I__3753\ : LocalMux
    port map (
            O => \N__24280\,
            I => \nx.n1797\
        );

    \I__3752\ : LocalMux
    port map (
            O => \N__24277\,
            I => \nx.n1797\
        );

    \I__3751\ : InMux
    port map (
            O => \N__24270\,
            I => \nx.n10831\
        );

    \I__3750\ : InMux
    port map (
            O => \N__24267\,
            I => \nx.n10832\
        );

    \I__3749\ : InMux
    port map (
            O => \N__24264\,
            I => \nx.n10641\
        );

    \I__3748\ : InMux
    port map (
            O => \N__24261\,
            I => \nx.n10642\
        );

    \I__3747\ : InMux
    port map (
            O => \N__24258\,
            I => \nx.n10643\
        );

    \I__3746\ : CEMux
    port map (
            O => \N__24255\,
            I => \N__24251\
        );

    \I__3745\ : CEMux
    port map (
            O => \N__24254\,
            I => \N__24247\
        );

    \I__3744\ : LocalMux
    port map (
            O => \N__24251\,
            I => \N__24244\
        );

    \I__3743\ : CEMux
    port map (
            O => \N__24250\,
            I => \N__24241\
        );

    \I__3742\ : LocalMux
    port map (
            O => \N__24247\,
            I => \N__24237\
        );

    \I__3741\ : Span4Mux_h
    port map (
            O => \N__24244\,
            I => \N__24232\
        );

    \I__3740\ : LocalMux
    port map (
            O => \N__24241\,
            I => \N__24232\
        );

    \I__3739\ : CEMux
    port map (
            O => \N__24240\,
            I => \N__24229\
        );

    \I__3738\ : Span4Mux_v
    port map (
            O => \N__24237\,
            I => \N__24226\
        );

    \I__3737\ : Span4Mux_v
    port map (
            O => \N__24232\,
            I => \N__24223\
        );

    \I__3736\ : LocalMux
    port map (
            O => \N__24229\,
            I => \N__24220\
        );

    \I__3735\ : Odrv4
    port map (
            O => \N__24226\,
            I => \nx.n7657\
        );

    \I__3734\ : Odrv4
    port map (
            O => \N__24223\,
            I => \nx.n7657\
        );

    \I__3733\ : Odrv12
    port map (
            O => \N__24220\,
            I => \nx.n7657\
        );

    \I__3732\ : SRMux
    port map (
            O => \N__24213\,
            I => \N__24209\
        );

    \I__3731\ : SRMux
    port map (
            O => \N__24212\,
            I => \N__24205\
        );

    \I__3730\ : LocalMux
    port map (
            O => \N__24209\,
            I => \N__24201\
        );

    \I__3729\ : SRMux
    port map (
            O => \N__24208\,
            I => \N__24198\
        );

    \I__3728\ : LocalMux
    port map (
            O => \N__24205\,
            I => \N__24195\
        );

    \I__3727\ : SRMux
    port map (
            O => \N__24204\,
            I => \N__24192\
        );

    \I__3726\ : Span4Mux_v
    port map (
            O => \N__24201\,
            I => \N__24189\
        );

    \I__3725\ : LocalMux
    port map (
            O => \N__24198\,
            I => \N__24184\
        );

    \I__3724\ : Span4Mux_v
    port map (
            O => \N__24195\,
            I => \N__24184\
        );

    \I__3723\ : LocalMux
    port map (
            O => \N__24192\,
            I => \N__24181\
        );

    \I__3722\ : Sp12to4
    port map (
            O => \N__24189\,
            I => \N__24178\
        );

    \I__3721\ : Span4Mux_v
    port map (
            O => \N__24184\,
            I => \N__24175\
        );

    \I__3720\ : Odrv12
    port map (
            O => \N__24181\,
            I => \nx.n7994\
        );

    \I__3719\ : Odrv12
    port map (
            O => \N__24178\,
            I => \nx.n7994\
        );

    \I__3718\ : Odrv4
    port map (
            O => \N__24175\,
            I => \nx.n7994\
        );

    \I__3717\ : InMux
    port map (
            O => \N__24168\,
            I => \bfn_6_27_0_\
        );

    \I__3716\ : InMux
    port map (
            O => \N__24165\,
            I => \nx.n10819\
        );

    \I__3715\ : InMux
    port map (
            O => \N__24162\,
            I => \nx.n10820\
        );

    \I__3714\ : InMux
    port map (
            O => \N__24159\,
            I => \N__24154\
        );

    \I__3713\ : InMux
    port map (
            O => \N__24158\,
            I => \N__24151\
        );

    \I__3712\ : InMux
    port map (
            O => \N__24157\,
            I => \N__24148\
        );

    \I__3711\ : LocalMux
    port map (
            O => \N__24154\,
            I => \nx.n1807\
        );

    \I__3710\ : LocalMux
    port map (
            O => \N__24151\,
            I => \nx.n1807\
        );

    \I__3709\ : LocalMux
    port map (
            O => \N__24148\,
            I => \nx.n1807\
        );

    \I__3708\ : InMux
    port map (
            O => \N__24141\,
            I => \nx.n10821\
        );

    \I__3707\ : CascadeMux
    port map (
            O => \N__24138\,
            I => \N__24135\
        );

    \I__3706\ : InMux
    port map (
            O => \N__24135\,
            I => \N__24130\
        );

    \I__3705\ : InMux
    port map (
            O => \N__24134\,
            I => \N__24127\
        );

    \I__3704\ : InMux
    port map (
            O => \N__24133\,
            I => \N__24124\
        );

    \I__3703\ : LocalMux
    port map (
            O => \N__24130\,
            I => \N__24121\
        );

    \I__3702\ : LocalMux
    port map (
            O => \N__24127\,
            I => \nx.n1806\
        );

    \I__3701\ : LocalMux
    port map (
            O => \N__24124\,
            I => \nx.n1806\
        );

    \I__3700\ : Odrv4
    port map (
            O => \N__24121\,
            I => \nx.n1806\
        );

    \I__3699\ : InMux
    port map (
            O => \N__24114\,
            I => \nx.n10822\
        );

    \I__3698\ : InMux
    port map (
            O => \N__24111\,
            I => \nx.n10823\
        );

    \I__3697\ : InMux
    port map (
            O => \N__24108\,
            I => \nx.n10632\
        );

    \I__3696\ : InMux
    port map (
            O => \N__24105\,
            I => \N__24100\
        );

    \I__3695\ : InMux
    port map (
            O => \N__24104\,
            I => \N__24097\
        );

    \I__3694\ : InMux
    port map (
            O => \N__24103\,
            I => \N__24093\
        );

    \I__3693\ : LocalMux
    port map (
            O => \N__24100\,
            I => \N__24087\
        );

    \I__3692\ : LocalMux
    port map (
            O => \N__24097\,
            I => \N__24087\
        );

    \I__3691\ : InMux
    port map (
            O => \N__24096\,
            I => \N__24084\
        );

    \I__3690\ : LocalMux
    port map (
            O => \N__24093\,
            I => \N__24081\
        );

    \I__3689\ : InMux
    port map (
            O => \N__24092\,
            I => \N__24078\
        );

    \I__3688\ : Span4Mux_v
    port map (
            O => \N__24087\,
            I => \N__24075\
        );

    \I__3687\ : LocalMux
    port map (
            O => \N__24084\,
            I => \N__24072\
        );

    \I__3686\ : Span4Mux_h
    port map (
            O => \N__24081\,
            I => \N__24069\
        );

    \I__3685\ : LocalMux
    port map (
            O => \N__24078\,
            I => \nx.bit_ctr_21\
        );

    \I__3684\ : Odrv4
    port map (
            O => \N__24075\,
            I => \nx.bit_ctr_21\
        );

    \I__3683\ : Odrv12
    port map (
            O => \N__24072\,
            I => \nx.bit_ctr_21\
        );

    \I__3682\ : Odrv4
    port map (
            O => \N__24069\,
            I => \nx.bit_ctr_21\
        );

    \I__3681\ : InMux
    port map (
            O => \N__24060\,
            I => \nx.n10633\
        );

    \I__3680\ : InMux
    port map (
            O => \N__24057\,
            I => \nx.n10634\
        );

    \I__3679\ : InMux
    port map (
            O => \N__24054\,
            I => \N__24049\
        );

    \I__3678\ : InMux
    port map (
            O => \N__24053\,
            I => \N__24045\
        );

    \I__3677\ : InMux
    port map (
            O => \N__24052\,
            I => \N__24041\
        );

    \I__3676\ : LocalMux
    port map (
            O => \N__24049\,
            I => \N__24038\
        );

    \I__3675\ : InMux
    port map (
            O => \N__24048\,
            I => \N__24035\
        );

    \I__3674\ : LocalMux
    port map (
            O => \N__24045\,
            I => \N__24032\
        );

    \I__3673\ : InMux
    port map (
            O => \N__24044\,
            I => \N__24029\
        );

    \I__3672\ : LocalMux
    port map (
            O => \N__24041\,
            I => \N__24024\
        );

    \I__3671\ : Span4Mux_h
    port map (
            O => \N__24038\,
            I => \N__24024\
        );

    \I__3670\ : LocalMux
    port map (
            O => \N__24035\,
            I => \N__24021\
        );

    \I__3669\ : Span4Mux_h
    port map (
            O => \N__24032\,
            I => \N__24018\
        );

    \I__3668\ : LocalMux
    port map (
            O => \N__24029\,
            I => \N__24013\
        );

    \I__3667\ : Span4Mux_v
    port map (
            O => \N__24024\,
            I => \N__24013\
        );

    \I__3666\ : Span4Mux_h
    port map (
            O => \N__24021\,
            I => \N__24010\
        );

    \I__3665\ : Odrv4
    port map (
            O => \N__24018\,
            I => \nx.bit_ctr_23\
        );

    \I__3664\ : Odrv4
    port map (
            O => \N__24013\,
            I => \nx.bit_ctr_23\
        );

    \I__3663\ : Odrv4
    port map (
            O => \N__24010\,
            I => \nx.bit_ctr_23\
        );

    \I__3662\ : InMux
    port map (
            O => \N__24003\,
            I => \nx.n10635\
        );

    \I__3661\ : InMux
    port map (
            O => \N__24000\,
            I => \N__23994\
        );

    \I__3660\ : InMux
    port map (
            O => \N__23999\,
            I => \N__23991\
        );

    \I__3659\ : InMux
    port map (
            O => \N__23998\,
            I => \N__23988\
        );

    \I__3658\ : InMux
    port map (
            O => \N__23997\,
            I => \N__23984\
        );

    \I__3657\ : LocalMux
    port map (
            O => \N__23994\,
            I => \N__23981\
        );

    \I__3656\ : LocalMux
    port map (
            O => \N__23991\,
            I => \N__23976\
        );

    \I__3655\ : LocalMux
    port map (
            O => \N__23988\,
            I => \N__23976\
        );

    \I__3654\ : InMux
    port map (
            O => \N__23987\,
            I => \N__23973\
        );

    \I__3653\ : LocalMux
    port map (
            O => \N__23984\,
            I => \N__23970\
        );

    \I__3652\ : Span4Mux_h
    port map (
            O => \N__23981\,
            I => \N__23967\
        );

    \I__3651\ : Span4Mux_v
    port map (
            O => \N__23976\,
            I => \N__23964\
        );

    \I__3650\ : LocalMux
    port map (
            O => \N__23973\,
            I => \nx.bit_ctr_24\
        );

    \I__3649\ : Odrv4
    port map (
            O => \N__23970\,
            I => \nx.bit_ctr_24\
        );

    \I__3648\ : Odrv4
    port map (
            O => \N__23967\,
            I => \nx.bit_ctr_24\
        );

    \I__3647\ : Odrv4
    port map (
            O => \N__23964\,
            I => \nx.bit_ctr_24\
        );

    \I__3646\ : InMux
    port map (
            O => \N__23955\,
            I => \bfn_6_26_0_\
        );

    \I__3645\ : InMux
    port map (
            O => \N__23952\,
            I => \N__23947\
        );

    \I__3644\ : InMux
    port map (
            O => \N__23951\,
            I => \N__23944\
        );

    \I__3643\ : InMux
    port map (
            O => \N__23950\,
            I => \N__23941\
        );

    \I__3642\ : LocalMux
    port map (
            O => \N__23947\,
            I => \N__23936\
        );

    \I__3641\ : LocalMux
    port map (
            O => \N__23944\,
            I => \N__23933\
        );

    \I__3640\ : LocalMux
    port map (
            O => \N__23941\,
            I => \N__23930\
        );

    \I__3639\ : InMux
    port map (
            O => \N__23940\,
            I => \N__23927\
        );

    \I__3638\ : InMux
    port map (
            O => \N__23939\,
            I => \N__23924\
        );

    \I__3637\ : Span4Mux_h
    port map (
            O => \N__23936\,
            I => \N__23921\
        );

    \I__3636\ : Span4Mux_v
    port map (
            O => \N__23933\,
            I => \N__23918\
        );

    \I__3635\ : Span4Mux_v
    port map (
            O => \N__23930\,
            I => \N__23915\
        );

    \I__3634\ : LocalMux
    port map (
            O => \N__23927\,
            I => \N__23912\
        );

    \I__3633\ : LocalMux
    port map (
            O => \N__23924\,
            I => \nx.bit_ctr_25\
        );

    \I__3632\ : Odrv4
    port map (
            O => \N__23921\,
            I => \nx.bit_ctr_25\
        );

    \I__3631\ : Odrv4
    port map (
            O => \N__23918\,
            I => \nx.bit_ctr_25\
        );

    \I__3630\ : Odrv4
    port map (
            O => \N__23915\,
            I => \nx.bit_ctr_25\
        );

    \I__3629\ : Odrv12
    port map (
            O => \N__23912\,
            I => \nx.bit_ctr_25\
        );

    \I__3628\ : InMux
    port map (
            O => \N__23901\,
            I => \nx.n10637\
        );

    \I__3627\ : InMux
    port map (
            O => \N__23898\,
            I => \nx.n10638\
        );

    \I__3626\ : InMux
    port map (
            O => \N__23895\,
            I => \nx.n10639\
        );

    \I__3625\ : InMux
    port map (
            O => \N__23892\,
            I => \nx.n10640\
        );

    \I__3624\ : InMux
    port map (
            O => \N__23889\,
            I => \nx.n10624\
        );

    \I__3623\ : InMux
    port map (
            O => \N__23886\,
            I => \nx.n10625\
        );

    \I__3622\ : InMux
    port map (
            O => \N__23883\,
            I => \nx.n10626\
        );

    \I__3621\ : InMux
    port map (
            O => \N__23880\,
            I => \nx.n10627\
        );

    \I__3620\ : InMux
    port map (
            O => \N__23877\,
            I => \bfn_6_25_0_\
        );

    \I__3619\ : InMux
    port map (
            O => \N__23874\,
            I => \nx.n10629\
        );

    \I__3618\ : InMux
    port map (
            O => \N__23871\,
            I => \nx.n10630\
        );

    \I__3617\ : InMux
    port map (
            O => \N__23868\,
            I => \N__23861\
        );

    \I__3616\ : InMux
    port map (
            O => \N__23867\,
            I => \N__23858\
        );

    \I__3615\ : InMux
    port map (
            O => \N__23866\,
            I => \N__23855\
        );

    \I__3614\ : InMux
    port map (
            O => \N__23865\,
            I => \N__23852\
        );

    \I__3613\ : InMux
    port map (
            O => \N__23864\,
            I => \N__23849\
        );

    \I__3612\ : LocalMux
    port map (
            O => \N__23861\,
            I => \N__23844\
        );

    \I__3611\ : LocalMux
    port map (
            O => \N__23858\,
            I => \N__23844\
        );

    \I__3610\ : LocalMux
    port map (
            O => \N__23855\,
            I => \N__23841\
        );

    \I__3609\ : LocalMux
    port map (
            O => \N__23852\,
            I => \nx.bit_ctr_19\
        );

    \I__3608\ : LocalMux
    port map (
            O => \N__23849\,
            I => \nx.bit_ctr_19\
        );

    \I__3607\ : Odrv4
    port map (
            O => \N__23844\,
            I => \nx.bit_ctr_19\
        );

    \I__3606\ : Odrv4
    port map (
            O => \N__23841\,
            I => \nx.bit_ctr_19\
        );

    \I__3605\ : InMux
    port map (
            O => \N__23832\,
            I => \nx.n10631\
        );

    \I__3604\ : InMux
    port map (
            O => \N__23829\,
            I => \N__23823\
        );

    \I__3603\ : InMux
    port map (
            O => \N__23828\,
            I => \N__23820\
        );

    \I__3602\ : InMux
    port map (
            O => \N__23827\,
            I => \N__23817\
        );

    \I__3601\ : InMux
    port map (
            O => \N__23826\,
            I => \N__23814\
        );

    \I__3600\ : LocalMux
    port map (
            O => \N__23823\,
            I => \N__23810\
        );

    \I__3599\ : LocalMux
    port map (
            O => \N__23820\,
            I => \N__23805\
        );

    \I__3598\ : LocalMux
    port map (
            O => \N__23817\,
            I => \N__23805\
        );

    \I__3597\ : LocalMux
    port map (
            O => \N__23814\,
            I => \N__23802\
        );

    \I__3596\ : InMux
    port map (
            O => \N__23813\,
            I => \N__23799\
        );

    \I__3595\ : Span4Mux_v
    port map (
            O => \N__23810\,
            I => \N__23796\
        );

    \I__3594\ : Span4Mux_v
    port map (
            O => \N__23805\,
            I => \N__23791\
        );

    \I__3593\ : Span4Mux_v
    port map (
            O => \N__23802\,
            I => \N__23791\
        );

    \I__3592\ : LocalMux
    port map (
            O => \N__23799\,
            I => \nx.bit_ctr_20\
        );

    \I__3591\ : Odrv4
    port map (
            O => \N__23796\,
            I => \nx.bit_ctr_20\
        );

    \I__3590\ : Odrv4
    port map (
            O => \N__23791\,
            I => \nx.bit_ctr_20\
        );

    \I__3589\ : InMux
    port map (
            O => \N__23784\,
            I => \nx.n10614\
        );

    \I__3588\ : InMux
    port map (
            O => \N__23781\,
            I => \nx.n10615\
        );

    \I__3587\ : InMux
    port map (
            O => \N__23778\,
            I => \nx.n10616\
        );

    \I__3586\ : InMux
    port map (
            O => \N__23775\,
            I => \nx.n10617\
        );

    \I__3585\ : InMux
    port map (
            O => \N__23772\,
            I => \nx.n10618\
        );

    \I__3584\ : InMux
    port map (
            O => \N__23769\,
            I => \nx.n10619\
        );

    \I__3583\ : InMux
    port map (
            O => \N__23766\,
            I => \bfn_6_24_0_\
        );

    \I__3582\ : InMux
    port map (
            O => \N__23763\,
            I => \nx.n10621\
        );

    \I__3581\ : InMux
    port map (
            O => \N__23760\,
            I => \nx.n10622\
        );

    \I__3580\ : InMux
    port map (
            O => \N__23757\,
            I => \nx.n10623\
        );

    \I__3579\ : CascadeMux
    port map (
            O => \N__23754\,
            I => \nx.n7899_cascade_\
        );

    \I__3578\ : CascadeMux
    port map (
            O => \N__23751\,
            I => \N__23748\
        );

    \I__3577\ : InMux
    port map (
            O => \N__23748\,
            I => \N__23745\
        );

    \I__3576\ : LocalMux
    port map (
            O => \N__23745\,
            I => \nx.n740\
        );

    \I__3575\ : CascadeMux
    port map (
            O => \N__23742\,
            I => \nx.n740_cascade_\
        );

    \I__3574\ : CascadeMux
    port map (
            O => \N__23739\,
            I => \nx.n11866_cascade_\
        );

    \I__3573\ : CascadeMux
    port map (
            O => \N__23736\,
            I => \nx.n838_cascade_\
        );

    \I__3572\ : InMux
    port map (
            O => \N__23733\,
            I => \N__23730\
        );

    \I__3571\ : LocalMux
    port map (
            O => \N__23730\,
            I => \N__23727\
        );

    \I__3570\ : Span4Mux_h
    port map (
            O => \N__23727\,
            I => \N__23724\
        );

    \I__3569\ : Span4Mux_h
    port map (
            O => \N__23724\,
            I => \N__23721\
        );

    \I__3568\ : Odrv4
    port map (
            O => \N__23721\,
            I => n18_adj_815
        );

    \I__3567\ : InMux
    port map (
            O => \N__23718\,
            I => \N__23715\
        );

    \I__3566\ : LocalMux
    port map (
            O => \N__23715\,
            I => \N__23712\
        );

    \I__3565\ : Span4Mux_h
    port map (
            O => \N__23712\,
            I => \N__23708\
        );

    \I__3564\ : InMux
    port map (
            O => \N__23711\,
            I => \N__23705\
        );

    \I__3563\ : Span4Mux_h
    port map (
            O => \N__23708\,
            I => \N__23702\
        );

    \I__3562\ : LocalMux
    port map (
            O => \N__23705\,
            I => delay_counter_31
        );

    \I__3561\ : Odrv4
    port map (
            O => \N__23702\,
            I => delay_counter_31
        );

    \I__3560\ : CascadeMux
    port map (
            O => \N__23697\,
            I => \N__23694\
        );

    \I__3559\ : InMux
    port map (
            O => \N__23694\,
            I => \N__23691\
        );

    \I__3558\ : LocalMux
    port map (
            O => \N__23691\,
            I => \N__23688\
        );

    \I__3557\ : Span4Mux_h
    port map (
            O => \N__23688\,
            I => \N__23685\
        );

    \I__3556\ : Odrv4
    port map (
            O => \N__23685\,
            I => n19_adj_814
        );

    \I__3555\ : InMux
    port map (
            O => \N__23682\,
            I => \N__23679\
        );

    \I__3554\ : LocalMux
    port map (
            O => \N__23679\,
            I => \N__23676\
        );

    \I__3553\ : Span4Mux_h
    port map (
            O => \N__23676\,
            I => \N__23673\
        );

    \I__3552\ : Odrv4
    port map (
            O => \N__23673\,
            I => n17_adj_816
        );

    \I__3551\ : InMux
    port map (
            O => \N__23670\,
            I => \bfn_6_23_0_\
        );

    \I__3550\ : InMux
    port map (
            O => \N__23667\,
            I => \nx.n10613\
        );

    \I__3549\ : InMux
    port map (
            O => \N__23664\,
            I => \N__23661\
        );

    \I__3548\ : LocalMux
    port map (
            O => \N__23661\,
            I => \N__23658\
        );

    \I__3547\ : Span12Mux_s11_v
    port map (
            O => \N__23658\,
            I => \N__23655\
        );

    \I__3546\ : Odrv12
    port map (
            O => \N__23655\,
            I => \nx.n5\
        );

    \I__3545\ : CascadeMux
    port map (
            O => \N__23652\,
            I => \N__23648\
        );

    \I__3544\ : CascadeMux
    port map (
            O => \N__23651\,
            I => \N__23645\
        );

    \I__3543\ : InMux
    port map (
            O => \N__23648\,
            I => \N__23642\
        );

    \I__3542\ : InMux
    port map (
            O => \N__23645\,
            I => \N__23639\
        );

    \I__3541\ : LocalMux
    port map (
            O => \N__23642\,
            I => \nx.n1007\
        );

    \I__3540\ : LocalMux
    port map (
            O => \N__23639\,
            I => \nx.n1007\
        );

    \I__3539\ : InMux
    port map (
            O => \N__23634\,
            I => \N__23631\
        );

    \I__3538\ : LocalMux
    port map (
            O => \N__23631\,
            I => \nx.n1075\
        );

    \I__3537\ : InMux
    port map (
            O => \N__23628\,
            I => \N__23624\
        );

    \I__3536\ : CascadeMux
    port map (
            O => \N__23627\,
            I => \N__23620\
        );

    \I__3535\ : LocalMux
    port map (
            O => \N__23624\,
            I => \N__23617\
        );

    \I__3534\ : InMux
    port map (
            O => \N__23623\,
            I => \N__23614\
        );

    \I__3533\ : InMux
    port map (
            O => \N__23620\,
            I => \N__23611\
        );

    \I__3532\ : Odrv4
    port map (
            O => \N__23617\,
            I => \nx.n1107\
        );

    \I__3531\ : LocalMux
    port map (
            O => \N__23614\,
            I => \nx.n1107\
        );

    \I__3530\ : LocalMux
    port map (
            O => \N__23611\,
            I => \nx.n1107\
        );

    \I__3529\ : CascadeMux
    port map (
            O => \N__23604\,
            I => \N__23600\
        );

    \I__3528\ : CascadeMux
    port map (
            O => \N__23603\,
            I => \N__23597\
        );

    \I__3527\ : InMux
    port map (
            O => \N__23600\,
            I => \N__23594\
        );

    \I__3526\ : InMux
    port map (
            O => \N__23597\,
            I => \N__23591\
        );

    \I__3525\ : LocalMux
    port map (
            O => \N__23594\,
            I => \nx.n1005\
        );

    \I__3524\ : LocalMux
    port map (
            O => \N__23591\,
            I => \nx.n1005\
        );

    \I__3523\ : CascadeMux
    port map (
            O => \N__23586\,
            I => \nx.n1005_cascade_\
        );

    \I__3522\ : CascadeMux
    port map (
            O => \N__23583\,
            I => \N__23578\
        );

    \I__3521\ : InMux
    port map (
            O => \N__23582\,
            I => \N__23575\
        );

    \I__3520\ : InMux
    port map (
            O => \N__23581\,
            I => \N__23572\
        );

    \I__3519\ : InMux
    port map (
            O => \N__23578\,
            I => \N__23569\
        );

    \I__3518\ : LocalMux
    port map (
            O => \N__23575\,
            I => \nx.n1009\
        );

    \I__3517\ : LocalMux
    port map (
            O => \N__23572\,
            I => \nx.n1009\
        );

    \I__3516\ : LocalMux
    port map (
            O => \N__23569\,
            I => \nx.n1009\
        );

    \I__3515\ : CascadeMux
    port map (
            O => \N__23562\,
            I => \nx.n7_adj_690_cascade_\
        );

    \I__3514\ : CascadeMux
    port map (
            O => \N__23559\,
            I => \N__23555\
        );

    \I__3513\ : CascadeMux
    port map (
            O => \N__23558\,
            I => \N__23549\
        );

    \I__3512\ : InMux
    port map (
            O => \N__23555\,
            I => \N__23545\
        );

    \I__3511\ : InMux
    port map (
            O => \N__23554\,
            I => \N__23542\
        );

    \I__3510\ : InMux
    port map (
            O => \N__23553\,
            I => \N__23533\
        );

    \I__3509\ : InMux
    port map (
            O => \N__23552\,
            I => \N__23533\
        );

    \I__3508\ : InMux
    port map (
            O => \N__23549\,
            I => \N__23533\
        );

    \I__3507\ : InMux
    port map (
            O => \N__23548\,
            I => \N__23533\
        );

    \I__3506\ : LocalMux
    port map (
            O => \N__23545\,
            I => \nx.n1037\
        );

    \I__3505\ : LocalMux
    port map (
            O => \N__23542\,
            I => \nx.n1037\
        );

    \I__3504\ : LocalMux
    port map (
            O => \N__23533\,
            I => \nx.n1037\
        );

    \I__3503\ : CascadeMux
    port map (
            O => \N__23526\,
            I => \nx.n1037_cascade_\
        );

    \I__3502\ : InMux
    port map (
            O => \N__23523\,
            I => \N__23520\
        );

    \I__3501\ : LocalMux
    port map (
            O => \N__23520\,
            I => \nx.n1073\
        );

    \I__3500\ : InMux
    port map (
            O => \N__23517\,
            I => \N__23513\
        );

    \I__3499\ : CascadeMux
    port map (
            O => \N__23516\,
            I => \N__23510\
        );

    \I__3498\ : LocalMux
    port map (
            O => \N__23513\,
            I => \N__23506\
        );

    \I__3497\ : InMux
    port map (
            O => \N__23510\,
            I => \N__23503\
        );

    \I__3496\ : InMux
    port map (
            O => \N__23509\,
            I => \N__23500\
        );

    \I__3495\ : Odrv4
    port map (
            O => \N__23506\,
            I => \nx.n1105\
        );

    \I__3494\ : LocalMux
    port map (
            O => \N__23503\,
            I => \nx.n1105\
        );

    \I__3493\ : LocalMux
    port map (
            O => \N__23500\,
            I => \nx.n1105\
        );

    \I__3492\ : InMux
    port map (
            O => \N__23493\,
            I => \N__23489\
        );

    \I__3491\ : InMux
    port map (
            O => \N__23492\,
            I => \N__23486\
        );

    \I__3490\ : LocalMux
    port map (
            O => \N__23489\,
            I => \N__23483\
        );

    \I__3489\ : LocalMux
    port map (
            O => \N__23486\,
            I => \N__23466\
        );

    \I__3488\ : Span4Mux_h
    port map (
            O => \N__23483\,
            I => \N__23463\
        );

    \I__3487\ : InMux
    port map (
            O => \N__23482\,
            I => \N__23458\
        );

    \I__3486\ : InMux
    port map (
            O => \N__23481\,
            I => \N__23458\
        );

    \I__3485\ : InMux
    port map (
            O => \N__23480\,
            I => \N__23453\
        );

    \I__3484\ : InMux
    port map (
            O => \N__23479\,
            I => \N__23453\
        );

    \I__3483\ : InMux
    port map (
            O => \N__23478\,
            I => \N__23450\
        );

    \I__3482\ : InMux
    port map (
            O => \N__23477\,
            I => \N__23445\
        );

    \I__3481\ : InMux
    port map (
            O => \N__23476\,
            I => \N__23445\
        );

    \I__3480\ : InMux
    port map (
            O => \N__23475\,
            I => \N__23440\
        );

    \I__3479\ : InMux
    port map (
            O => \N__23474\,
            I => \N__23440\
        );

    \I__3478\ : InMux
    port map (
            O => \N__23473\,
            I => \N__23433\
        );

    \I__3477\ : InMux
    port map (
            O => \N__23472\,
            I => \N__23433\
        );

    \I__3476\ : InMux
    port map (
            O => \N__23471\,
            I => \N__23433\
        );

    \I__3475\ : InMux
    port map (
            O => \N__23470\,
            I => \N__23428\
        );

    \I__3474\ : InMux
    port map (
            O => \N__23469\,
            I => \N__23428\
        );

    \I__3473\ : Odrv4
    port map (
            O => \N__23466\,
            I => state_1_adj_791
        );

    \I__3472\ : Odrv4
    port map (
            O => \N__23463\,
            I => state_1_adj_791
        );

    \I__3471\ : LocalMux
    port map (
            O => \N__23458\,
            I => state_1_adj_791
        );

    \I__3470\ : LocalMux
    port map (
            O => \N__23453\,
            I => state_1_adj_791
        );

    \I__3469\ : LocalMux
    port map (
            O => \N__23450\,
            I => state_1_adj_791
        );

    \I__3468\ : LocalMux
    port map (
            O => \N__23445\,
            I => state_1_adj_791
        );

    \I__3467\ : LocalMux
    port map (
            O => \N__23440\,
            I => state_1_adj_791
        );

    \I__3466\ : LocalMux
    port map (
            O => \N__23433\,
            I => state_1_adj_791
        );

    \I__3465\ : LocalMux
    port map (
            O => \N__23428\,
            I => state_1_adj_791
        );

    \I__3464\ : CascadeMux
    port map (
            O => \N__23409\,
            I => \nx.n3901_cascade_\
        );

    \I__3463\ : InMux
    port map (
            O => \N__23406\,
            I => \N__23403\
        );

    \I__3462\ : LocalMux
    port map (
            O => \N__23403\,
            I => \N__23400\
        );

    \I__3461\ : Odrv4
    port map (
            O => \N__23400\,
            I => \nx.n13435\
        );

    \I__3460\ : InMux
    port map (
            O => \N__23397\,
            I => \N__23394\
        );

    \I__3459\ : LocalMux
    port map (
            O => \N__23394\,
            I => \nx.n1077\
        );

    \I__3458\ : InMux
    port map (
            O => \N__23391\,
            I => \bfn_6_20_0_\
        );

    \I__3457\ : CascadeMux
    port map (
            O => \N__23388\,
            I => \N__23385\
        );

    \I__3456\ : InMux
    port map (
            O => \N__23385\,
            I => \N__23382\
        );

    \I__3455\ : LocalMux
    port map (
            O => \N__23382\,
            I => \nx.n1076\
        );

    \I__3454\ : InMux
    port map (
            O => \N__23379\,
            I => \nx.n10743\
        );

    \I__3453\ : InMux
    port map (
            O => \N__23376\,
            I => \nx.n10744\
        );

    \I__3452\ : InMux
    port map (
            O => \N__23373\,
            I => \N__23370\
        );

    \I__3451\ : LocalMux
    port map (
            O => \N__23370\,
            I => \nx.n1074\
        );

    \I__3450\ : InMux
    port map (
            O => \N__23367\,
            I => \nx.n10745\
        );

    \I__3449\ : InMux
    port map (
            O => \N__23364\,
            I => \nx.n10746\
        );

    \I__3448\ : InMux
    port map (
            O => \N__23361\,
            I => \N__23358\
        );

    \I__3447\ : LocalMux
    port map (
            O => \N__23358\,
            I => \nx.n1072\
        );

    \I__3446\ : InMux
    port map (
            O => \N__23355\,
            I => \nx.n10747\
        );

    \I__3445\ : InMux
    port map (
            O => \N__23352\,
            I => \nx.n10748\
        );

    \I__3444\ : CascadeMux
    port map (
            O => \N__23349\,
            I => \N__23345\
        );

    \I__3443\ : InMux
    port map (
            O => \N__23348\,
            I => \N__23342\
        );

    \I__3442\ : InMux
    port map (
            O => \N__23345\,
            I => \N__23339\
        );

    \I__3441\ : LocalMux
    port map (
            O => \N__23342\,
            I => \N__23336\
        );

    \I__3440\ : LocalMux
    port map (
            O => \N__23339\,
            I => \nx.n1103\
        );

    \I__3439\ : Odrv4
    port map (
            O => \N__23336\,
            I => \nx.n1103\
        );

    \I__3438\ : InMux
    port map (
            O => \N__23331\,
            I => \N__23328\
        );

    \I__3437\ : LocalMux
    port map (
            O => \N__23328\,
            I => \N__23324\
        );

    \I__3436\ : CascadeMux
    port map (
            O => \N__23327\,
            I => \N__23320\
        );

    \I__3435\ : Span4Mux_h
    port map (
            O => \N__23324\,
            I => \N__23317\
        );

    \I__3434\ : InMux
    port map (
            O => \N__23323\,
            I => \N__23314\
        );

    \I__3433\ : InMux
    port map (
            O => \N__23320\,
            I => \N__23311\
        );

    \I__3432\ : Odrv4
    port map (
            O => \N__23317\,
            I => timer_26
        );

    \I__3431\ : LocalMux
    port map (
            O => \N__23314\,
            I => timer_26
        );

    \I__3430\ : LocalMux
    port map (
            O => \N__23311\,
            I => timer_26
        );

    \I__3429\ : InMux
    port map (
            O => \N__23304\,
            I => \N__23298\
        );

    \I__3428\ : InMux
    port map (
            O => \N__23303\,
            I => \N__23298\
        );

    \I__3427\ : LocalMux
    port map (
            O => \N__23298\,
            I => neo_pixel_transmitter_t0_26
        );

    \I__3426\ : InMux
    port map (
            O => \N__23295\,
            I => \N__23292\
        );

    \I__3425\ : LocalMux
    port map (
            O => \N__23292\,
            I => \N__23289\
        );

    \I__3424\ : Span4Mux_v
    port map (
            O => \N__23289\,
            I => \N__23286\
        );

    \I__3423\ : Odrv4
    port map (
            O => \N__23286\,
            I => \nx.n7\
        );

    \I__3422\ : InMux
    port map (
            O => \N__23283\,
            I => \N__23280\
        );

    \I__3421\ : LocalMux
    port map (
            O => \N__23280\,
            I => \nx.n10_adj_760\
        );

    \I__3420\ : CascadeMux
    port map (
            O => \N__23277\,
            I => \N__23274\
        );

    \I__3419\ : InMux
    port map (
            O => \N__23274\,
            I => \N__23271\
        );

    \I__3418\ : LocalMux
    port map (
            O => \N__23271\,
            I => \N__23268\
        );

    \I__3417\ : Span4Mux_h
    port map (
            O => \N__23268\,
            I => \N__23265\
        );

    \I__3416\ : Odrv4
    port map (
            O => \N__23265\,
            I => n12_adj_844
        );

    \I__3415\ : InMux
    port map (
            O => \N__23262\,
            I => \N__23256\
        );

    \I__3414\ : InMux
    port map (
            O => \N__23261\,
            I => \N__23251\
        );

    \I__3413\ : InMux
    port map (
            O => \N__23260\,
            I => \N__23251\
        );

    \I__3412\ : CascadeMux
    port map (
            O => \N__23259\,
            I => \N__23245\
        );

    \I__3411\ : LocalMux
    port map (
            O => \N__23256\,
            I => \N__23240\
        );

    \I__3410\ : LocalMux
    port map (
            O => \N__23251\,
            I => \N__23237\
        );

    \I__3409\ : InMux
    port map (
            O => \N__23250\,
            I => \N__23234\
        );

    \I__3408\ : InMux
    port map (
            O => \N__23249\,
            I => \N__23231\
        );

    \I__3407\ : InMux
    port map (
            O => \N__23248\,
            I => \N__23222\
        );

    \I__3406\ : InMux
    port map (
            O => \N__23245\,
            I => \N__23222\
        );

    \I__3405\ : InMux
    port map (
            O => \N__23244\,
            I => \N__23222\
        );

    \I__3404\ : InMux
    port map (
            O => \N__23243\,
            I => \N__23222\
        );

    \I__3403\ : Span4Mux_v
    port map (
            O => \N__23240\,
            I => \N__23219\
        );

    \I__3402\ : Span4Mux_h
    port map (
            O => \N__23237\,
            I => \N__23216\
        );

    \I__3401\ : LocalMux
    port map (
            O => \N__23234\,
            I => \nx.start\
        );

    \I__3400\ : LocalMux
    port map (
            O => \N__23231\,
            I => \nx.start\
        );

    \I__3399\ : LocalMux
    port map (
            O => \N__23222\,
            I => \nx.start\
        );

    \I__3398\ : Odrv4
    port map (
            O => \N__23219\,
            I => \nx.start\
        );

    \I__3397\ : Odrv4
    port map (
            O => \N__23216\,
            I => \nx.start\
        );

    \I__3396\ : InMux
    port map (
            O => \N__23205\,
            I => \N__23200\
        );

    \I__3395\ : InMux
    port map (
            O => \N__23204\,
            I => \N__23197\
        );

    \I__3394\ : InMux
    port map (
            O => \N__23203\,
            I => \N__23194\
        );

    \I__3393\ : LocalMux
    port map (
            O => \N__23200\,
            I => \nx.n11908\
        );

    \I__3392\ : LocalMux
    port map (
            O => \N__23197\,
            I => \nx.n11908\
        );

    \I__3391\ : LocalMux
    port map (
            O => \N__23194\,
            I => \nx.n11908\
        );

    \I__3390\ : CascadeMux
    port map (
            O => \N__23187\,
            I => \N__23184\
        );

    \I__3389\ : InMux
    port map (
            O => \N__23184\,
            I => \N__23178\
        );

    \I__3388\ : InMux
    port map (
            O => \N__23183\,
            I => \N__23175\
        );

    \I__3387\ : InMux
    port map (
            O => \N__23182\,
            I => \N__23170\
        );

    \I__3386\ : InMux
    port map (
            O => \N__23181\,
            I => \N__23170\
        );

    \I__3385\ : LocalMux
    port map (
            O => \N__23178\,
            I => \N__23161\
        );

    \I__3384\ : LocalMux
    port map (
            O => \N__23175\,
            I => \N__23161\
        );

    \I__3383\ : LocalMux
    port map (
            O => \N__23170\,
            I => \N__23161\
        );

    \I__3382\ : InMux
    port map (
            O => \N__23169\,
            I => \N__23158\
        );

    \I__3381\ : InMux
    port map (
            O => \N__23168\,
            I => \N__23155\
        );

    \I__3380\ : Span4Mux_h
    port map (
            O => \N__23161\,
            I => \N__23152\
        );

    \I__3379\ : LocalMux
    port map (
            O => \N__23158\,
            I => \N__23149\
        );

    \I__3378\ : LocalMux
    port map (
            O => \N__23155\,
            I => \nx.n7564\
        );

    \I__3377\ : Odrv4
    port map (
            O => \N__23152\,
            I => \nx.n7564\
        );

    \I__3376\ : Odrv12
    port map (
            O => \N__23149\,
            I => \nx.n7564\
        );

    \I__3375\ : InMux
    port map (
            O => \N__23142\,
            I => \N__23138\
        );

    \I__3374\ : InMux
    port map (
            O => \N__23141\,
            I => \N__23135\
        );

    \I__3373\ : LocalMux
    port map (
            O => \N__23138\,
            I => update_color
        );

    \I__3372\ : LocalMux
    port map (
            O => \N__23135\,
            I => update_color
        );

    \I__3371\ : CascadeMux
    port map (
            O => \N__23130\,
            I => \nx.n13436_cascade_\
        );

    \I__3370\ : InMux
    port map (
            O => \N__23127\,
            I => \N__23124\
        );

    \I__3369\ : LocalMux
    port map (
            O => \N__23124\,
            I => \nx.n3901\
        );

    \I__3368\ : InMux
    port map (
            O => \N__23121\,
            I => \N__23118\
        );

    \I__3367\ : LocalMux
    port map (
            O => \N__23118\,
            I => \N__23115\
        );

    \I__3366\ : Odrv4
    port map (
            O => \N__23115\,
            I => \nx.n16_adj_766\
        );

    \I__3365\ : InMux
    port map (
            O => \N__23112\,
            I => \N__23107\
        );

    \I__3364\ : InMux
    port map (
            O => \N__23111\,
            I => \N__23104\
        );

    \I__3363\ : InMux
    port map (
            O => \N__23110\,
            I => \N__23101\
        );

    \I__3362\ : LocalMux
    port map (
            O => \N__23107\,
            I => \N__23094\
        );

    \I__3361\ : LocalMux
    port map (
            O => \N__23104\,
            I => \N__23094\
        );

    \I__3360\ : LocalMux
    port map (
            O => \N__23101\,
            I => \N__23094\
        );

    \I__3359\ : Odrv12
    port map (
            O => \N__23094\,
            I => \nx.n1702\
        );

    \I__3358\ : CascadeMux
    port map (
            O => \N__23091\,
            I => \nx.n22_adj_774_cascade_\
        );

    \I__3357\ : InMux
    port map (
            O => \N__23088\,
            I => \N__23083\
        );

    \I__3356\ : InMux
    port map (
            O => \N__23087\,
            I => \N__23080\
        );

    \I__3355\ : InMux
    port map (
            O => \N__23086\,
            I => \N__23077\
        );

    \I__3354\ : LocalMux
    port map (
            O => \N__23083\,
            I => \N__23074\
        );

    \I__3353\ : LocalMux
    port map (
            O => \N__23080\,
            I => \N__23069\
        );

    \I__3352\ : LocalMux
    port map (
            O => \N__23077\,
            I => \N__23069\
        );

    \I__3351\ : Odrv4
    port map (
            O => \N__23074\,
            I => \nx.n1698\
        );

    \I__3350\ : Odrv4
    port map (
            O => \N__23069\,
            I => \nx.n1698\
        );

    \I__3349\ : InMux
    port map (
            O => \N__23064\,
            I => \N__23059\
        );

    \I__3348\ : InMux
    port map (
            O => \N__23063\,
            I => \N__23056\
        );

    \I__3347\ : InMux
    port map (
            O => \N__23062\,
            I => \N__23053\
        );

    \I__3346\ : LocalMux
    port map (
            O => \N__23059\,
            I => \N__23046\
        );

    \I__3345\ : LocalMux
    port map (
            O => \N__23056\,
            I => \N__23046\
        );

    \I__3344\ : LocalMux
    port map (
            O => \N__23053\,
            I => \N__23046\
        );

    \I__3343\ : Odrv4
    port map (
            O => \N__23046\,
            I => \nx.n1699\
        );

    \I__3342\ : InMux
    port map (
            O => \N__23043\,
            I => \N__23038\
        );

    \I__3341\ : InMux
    port map (
            O => \N__23042\,
            I => \N__23035\
        );

    \I__3340\ : InMux
    port map (
            O => \N__23041\,
            I => \N__23032\
        );

    \I__3339\ : LocalMux
    port map (
            O => \N__23038\,
            I => \N__23029\
        );

    \I__3338\ : LocalMux
    port map (
            O => \N__23035\,
            I => \N__23026\
        );

    \I__3337\ : LocalMux
    port map (
            O => \N__23032\,
            I => \N__23023\
        );

    \I__3336\ : Odrv4
    port map (
            O => \N__23029\,
            I => \nx.n1697\
        );

    \I__3335\ : Odrv12
    port map (
            O => \N__23026\,
            I => \nx.n1697\
        );

    \I__3334\ : Odrv4
    port map (
            O => \N__23023\,
            I => \nx.n1697\
        );

    \I__3333\ : CascadeMux
    port map (
            O => \N__23016\,
            I => \nx.n24_adj_776_cascade_\
        );

    \I__3332\ : InMux
    port map (
            O => \N__23013\,
            I => \N__23010\
        );

    \I__3331\ : LocalMux
    port map (
            O => \N__23010\,
            I => \N__23007\
        );

    \I__3330\ : Odrv4
    port map (
            O => \N__23007\,
            I => \nx.n20_adj_775\
        );

    \I__3329\ : CascadeMux
    port map (
            O => \N__23004\,
            I => \N__22990\
        );

    \I__3328\ : CascadeMux
    port map (
            O => \N__23003\,
            I => \N__22987\
        );

    \I__3327\ : CascadeMux
    port map (
            O => \N__23002\,
            I => \N__22984\
        );

    \I__3326\ : CascadeMux
    port map (
            O => \N__23001\,
            I => \N__22981\
        );

    \I__3325\ : CascadeMux
    port map (
            O => \N__23000\,
            I => \N__22978\
        );

    \I__3324\ : CascadeMux
    port map (
            O => \N__22999\,
            I => \N__22975\
        );

    \I__3323\ : CascadeMux
    port map (
            O => \N__22998\,
            I => \N__22972\
        );

    \I__3322\ : CascadeMux
    port map (
            O => \N__22997\,
            I => \N__22969\
        );

    \I__3321\ : CascadeMux
    port map (
            O => \N__22996\,
            I => \N__22966\
        );

    \I__3320\ : CascadeMux
    port map (
            O => \N__22995\,
            I => \N__22963\
        );

    \I__3319\ : CascadeMux
    port map (
            O => \N__22994\,
            I => \N__22960\
        );

    \I__3318\ : CascadeMux
    port map (
            O => \N__22993\,
            I => \N__22957\
        );

    \I__3317\ : InMux
    port map (
            O => \N__22990\,
            I => \N__22950\
        );

    \I__3316\ : InMux
    port map (
            O => \N__22987\,
            I => \N__22950\
        );

    \I__3315\ : InMux
    port map (
            O => \N__22984\,
            I => \N__22950\
        );

    \I__3314\ : InMux
    port map (
            O => \N__22981\,
            I => \N__22943\
        );

    \I__3313\ : InMux
    port map (
            O => \N__22978\,
            I => \N__22943\
        );

    \I__3312\ : InMux
    port map (
            O => \N__22975\,
            I => \N__22943\
        );

    \I__3311\ : InMux
    port map (
            O => \N__22972\,
            I => \N__22936\
        );

    \I__3310\ : InMux
    port map (
            O => \N__22969\,
            I => \N__22936\
        );

    \I__3309\ : InMux
    port map (
            O => \N__22966\,
            I => \N__22936\
        );

    \I__3308\ : InMux
    port map (
            O => \N__22963\,
            I => \N__22929\
        );

    \I__3307\ : InMux
    port map (
            O => \N__22960\,
            I => \N__22929\
        );

    \I__3306\ : InMux
    port map (
            O => \N__22957\,
            I => \N__22929\
        );

    \I__3305\ : LocalMux
    port map (
            O => \N__22950\,
            I => \N__22924\
        );

    \I__3304\ : LocalMux
    port map (
            O => \N__22943\,
            I => \N__22924\
        );

    \I__3303\ : LocalMux
    port map (
            O => \N__22936\,
            I => \nx.n1730\
        );

    \I__3302\ : LocalMux
    port map (
            O => \N__22929\,
            I => \nx.n1730\
        );

    \I__3301\ : Odrv4
    port map (
            O => \N__22924\,
            I => \nx.n1730\
        );

    \I__3300\ : CascadeMux
    port map (
            O => \N__22917\,
            I => \nx.n1730_cascade_\
        );

    \I__3299\ : CascadeMux
    port map (
            O => \N__22914\,
            I => \N__22910\
        );

    \I__3298\ : CascadeMux
    port map (
            O => \N__22913\,
            I => \N__22907\
        );

    \I__3297\ : InMux
    port map (
            O => \N__22910\,
            I => \N__22904\
        );

    \I__3296\ : InMux
    port map (
            O => \N__22907\,
            I => \N__22901\
        );

    \I__3295\ : LocalMux
    port map (
            O => \N__22904\,
            I => \N__22896\
        );

    \I__3294\ : LocalMux
    port map (
            O => \N__22901\,
            I => \N__22896\
        );

    \I__3293\ : Odrv4
    port map (
            O => \N__22896\,
            I => \nx.n13601\
        );

    \I__3292\ : InMux
    port map (
            O => \N__22893\,
            I => \N__22890\
        );

    \I__3291\ : LocalMux
    port map (
            O => \N__22890\,
            I => n11972
        );

    \I__3290\ : InMux
    port map (
            O => \N__22887\,
            I => \N__22884\
        );

    \I__3289\ : LocalMux
    port map (
            O => \N__22884\,
            I => \nx.n13514\
        );

    \I__3288\ : CascadeMux
    port map (
            O => \N__22881\,
            I => \N__22878\
        );

    \I__3287\ : InMux
    port map (
            O => \N__22878\,
            I => \N__22875\
        );

    \I__3286\ : LocalMux
    port map (
            O => \N__22875\,
            I => \nx.n13513\
        );

    \I__3285\ : InMux
    port map (
            O => \N__22872\,
            I => \N__22869\
        );

    \I__3284\ : LocalMux
    port map (
            O => \N__22869\,
            I => \N__22865\
        );

    \I__3283\ : InMux
    port map (
            O => \N__22868\,
            I => \N__22862\
        );

    \I__3282\ : Odrv4
    port map (
            O => \N__22865\,
            I => \nx.n7598\
        );

    \I__3281\ : LocalMux
    port map (
            O => \N__22862\,
            I => \nx.n7598\
        );

    \I__3280\ : InMux
    port map (
            O => \N__22857\,
            I => \N__22849\
        );

    \I__3279\ : InMux
    port map (
            O => \N__22856\,
            I => \N__22849\
        );

    \I__3278\ : InMux
    port map (
            O => \N__22855\,
            I => \N__22846\
        );

    \I__3277\ : InMux
    port map (
            O => \N__22854\,
            I => \N__22843\
        );

    \I__3276\ : LocalMux
    port map (
            O => \N__22849\,
            I => \nx.n11113\
        );

    \I__3275\ : LocalMux
    port map (
            O => \N__22846\,
            I => \nx.n11113\
        );

    \I__3274\ : LocalMux
    port map (
            O => \N__22843\,
            I => \nx.n11113\
        );

    \I__3273\ : CascadeMux
    port map (
            O => \N__22836\,
            I => \nx.n7598_cascade_\
        );

    \I__3272\ : InMux
    port map (
            O => \N__22833\,
            I => \bfn_5_28_0_\
        );

    \I__3271\ : InMux
    port map (
            O => \N__22830\,
            I => \N__22826\
        );

    \I__3270\ : InMux
    port map (
            O => \N__22829\,
            I => \N__22823\
        );

    \I__3269\ : LocalMux
    port map (
            O => \N__22826\,
            I => \N__22817\
        );

    \I__3268\ : LocalMux
    port map (
            O => \N__22823\,
            I => \N__22817\
        );

    \I__3267\ : InMux
    port map (
            O => \N__22822\,
            I => \N__22814\
        );

    \I__3266\ : Odrv4
    port map (
            O => \N__22817\,
            I => \nx.n1701\
        );

    \I__3265\ : LocalMux
    port map (
            O => \N__22814\,
            I => \nx.n1701\
        );

    \I__3264\ : InMux
    port map (
            O => \N__22809\,
            I => \nx.n10814\
        );

    \I__3263\ : InMux
    port map (
            O => \N__22806\,
            I => \nx.n10815\
        );

    \I__3262\ : InMux
    port map (
            O => \N__22803\,
            I => \nx.n10816\
        );

    \I__3261\ : InMux
    port map (
            O => \N__22800\,
            I => \nx.n10817\
        );

    \I__3260\ : InMux
    port map (
            O => \N__22797\,
            I => \nx.n10818\
        );

    \I__3259\ : InMux
    port map (
            O => \N__22794\,
            I => \N__22791\
        );

    \I__3258\ : LocalMux
    port map (
            O => \N__22791\,
            I => \N__22788\
        );

    \I__3257\ : Span4Mux_v
    port map (
            O => \N__22788\,
            I => \N__22783\
        );

    \I__3256\ : InMux
    port map (
            O => \N__22787\,
            I => \N__22780\
        );

    \I__3255\ : InMux
    port map (
            O => \N__22786\,
            I => \N__22777\
        );

    \I__3254\ : Span4Mux_h
    port map (
            O => \N__22783\,
            I => \N__22772\
        );

    \I__3253\ : LocalMux
    port map (
            O => \N__22780\,
            I => \N__22772\
        );

    \I__3252\ : LocalMux
    port map (
            O => \N__22777\,
            I => \N__22769\
        );

    \I__3251\ : Odrv4
    port map (
            O => \N__22772\,
            I => \nx.n1703\
        );

    \I__3250\ : Odrv12
    port map (
            O => \N__22769\,
            I => \nx.n1703\
        );

    \I__3249\ : InMux
    port map (
            O => \N__22764\,
            I => \N__22759\
        );

    \I__3248\ : InMux
    port map (
            O => \N__22763\,
            I => \N__22756\
        );

    \I__3247\ : InMux
    port map (
            O => \N__22762\,
            I => \N__22753\
        );

    \I__3246\ : LocalMux
    port map (
            O => \N__22759\,
            I => \N__22746\
        );

    \I__3245\ : LocalMux
    port map (
            O => \N__22756\,
            I => \N__22746\
        );

    \I__3244\ : LocalMux
    port map (
            O => \N__22753\,
            I => \N__22746\
        );

    \I__3243\ : Odrv12
    port map (
            O => \N__22746\,
            I => \nx.n1706\
        );

    \I__3242\ : CascadeMux
    port map (
            O => \N__22743\,
            I => \N__22738\
        );

    \I__3241\ : InMux
    port map (
            O => \N__22742\,
            I => \N__22735\
        );

    \I__3240\ : InMux
    port map (
            O => \N__22741\,
            I => \N__22732\
        );

    \I__3239\ : InMux
    port map (
            O => \N__22738\,
            I => \N__22729\
        );

    \I__3238\ : LocalMux
    port map (
            O => \N__22735\,
            I => \N__22724\
        );

    \I__3237\ : LocalMux
    port map (
            O => \N__22732\,
            I => \N__22724\
        );

    \I__3236\ : LocalMux
    port map (
            O => \N__22729\,
            I => \N__22721\
        );

    \I__3235\ : Odrv4
    port map (
            O => \N__22724\,
            I => \nx.n1705\
        );

    \I__3234\ : Odrv12
    port map (
            O => \N__22721\,
            I => \nx.n1705\
        );

    \I__3233\ : InMux
    port map (
            O => \N__22716\,
            I => \N__22711\
        );

    \I__3232\ : InMux
    port map (
            O => \N__22715\,
            I => \N__22708\
        );

    \I__3231\ : InMux
    port map (
            O => \N__22714\,
            I => \N__22705\
        );

    \I__3230\ : LocalMux
    port map (
            O => \N__22711\,
            I => \N__22698\
        );

    \I__3229\ : LocalMux
    port map (
            O => \N__22708\,
            I => \N__22698\
        );

    \I__3228\ : LocalMux
    port map (
            O => \N__22705\,
            I => \N__22698\
        );

    \I__3227\ : Odrv12
    port map (
            O => \N__22698\,
            I => \nx.n1700\
        );

    \I__3226\ : InMux
    port map (
            O => \N__22695\,
            I => \bfn_5_27_0_\
        );

    \I__3225\ : InMux
    port map (
            O => \N__22692\,
            I => \N__22687\
        );

    \I__3224\ : InMux
    port map (
            O => \N__22691\,
            I => \N__22684\
        );

    \I__3223\ : CascadeMux
    port map (
            O => \N__22690\,
            I => \N__22681\
        );

    \I__3222\ : LocalMux
    port map (
            O => \N__22687\,
            I => \N__22676\
        );

    \I__3221\ : LocalMux
    port map (
            O => \N__22684\,
            I => \N__22676\
        );

    \I__3220\ : InMux
    port map (
            O => \N__22681\,
            I => \N__22673\
        );

    \I__3219\ : Odrv12
    port map (
            O => \N__22676\,
            I => \nx.n1709\
        );

    \I__3218\ : LocalMux
    port map (
            O => \N__22673\,
            I => \nx.n1709\
        );

    \I__3217\ : InMux
    port map (
            O => \N__22668\,
            I => \nx.n10806\
        );

    \I__3216\ : InMux
    port map (
            O => \N__22665\,
            I => \N__22662\
        );

    \I__3215\ : LocalMux
    port map (
            O => \N__22662\,
            I => \N__22658\
        );

    \I__3214\ : InMux
    port map (
            O => \N__22661\,
            I => \N__22655\
        );

    \I__3213\ : Span4Mux_h
    port map (
            O => \N__22658\,
            I => \N__22649\
        );

    \I__3212\ : LocalMux
    port map (
            O => \N__22655\,
            I => \N__22649\
        );

    \I__3211\ : InMux
    port map (
            O => \N__22654\,
            I => \N__22646\
        );

    \I__3210\ : Odrv4
    port map (
            O => \N__22649\,
            I => \nx.n1708\
        );

    \I__3209\ : LocalMux
    port map (
            O => \N__22646\,
            I => \nx.n1708\
        );

    \I__3208\ : InMux
    port map (
            O => \N__22641\,
            I => \nx.n10807\
        );

    \I__3207\ : InMux
    port map (
            O => \N__22638\,
            I => \N__22634\
        );

    \I__3206\ : InMux
    port map (
            O => \N__22637\,
            I => \N__22631\
        );

    \I__3205\ : LocalMux
    port map (
            O => \N__22634\,
            I => \N__22625\
        );

    \I__3204\ : LocalMux
    port map (
            O => \N__22631\,
            I => \N__22625\
        );

    \I__3203\ : InMux
    port map (
            O => \N__22630\,
            I => \N__22622\
        );

    \I__3202\ : Odrv4
    port map (
            O => \N__22625\,
            I => \nx.n1707\
        );

    \I__3201\ : LocalMux
    port map (
            O => \N__22622\,
            I => \nx.n1707\
        );

    \I__3200\ : InMux
    port map (
            O => \N__22617\,
            I => \nx.n10808\
        );

    \I__3199\ : InMux
    port map (
            O => \N__22614\,
            I => \nx.n10809\
        );

    \I__3198\ : InMux
    port map (
            O => \N__22611\,
            I => \nx.n10810\
        );

    \I__3197\ : InMux
    port map (
            O => \N__22608\,
            I => \N__22603\
        );

    \I__3196\ : InMux
    port map (
            O => \N__22607\,
            I => \N__22600\
        );

    \I__3195\ : CascadeMux
    port map (
            O => \N__22606\,
            I => \N__22597\
        );

    \I__3194\ : LocalMux
    port map (
            O => \N__22603\,
            I => \N__22592\
        );

    \I__3193\ : LocalMux
    port map (
            O => \N__22600\,
            I => \N__22592\
        );

    \I__3192\ : InMux
    port map (
            O => \N__22597\,
            I => \N__22589\
        );

    \I__3191\ : Odrv4
    port map (
            O => \N__22592\,
            I => \nx.n1704\
        );

    \I__3190\ : LocalMux
    port map (
            O => \N__22589\,
            I => \nx.n1704\
        );

    \I__3189\ : InMux
    port map (
            O => \N__22584\,
            I => \nx.n10811\
        );

    \I__3188\ : InMux
    port map (
            O => \N__22581\,
            I => \nx.n10812\
        );

    \I__3187\ : InMux
    port map (
            O => \N__22578\,
            I => \N__22573\
        );

    \I__3186\ : InMux
    port map (
            O => \N__22577\,
            I => \N__22570\
        );

    \I__3185\ : InMux
    port map (
            O => \N__22576\,
            I => \N__22567\
        );

    \I__3184\ : LocalMux
    port map (
            O => \N__22573\,
            I => \nx.n1605\
        );

    \I__3183\ : LocalMux
    port map (
            O => \N__22570\,
            I => \nx.n1605\
        );

    \I__3182\ : LocalMux
    port map (
            O => \N__22567\,
            I => \nx.n1605\
        );

    \I__3181\ : InMux
    port map (
            O => \N__22560\,
            I => \nx.n10798\
        );

    \I__3180\ : InMux
    port map (
            O => \N__22557\,
            I => \N__22552\
        );

    \I__3179\ : InMux
    port map (
            O => \N__22556\,
            I => \N__22549\
        );

    \I__3178\ : InMux
    port map (
            O => \N__22555\,
            I => \N__22546\
        );

    \I__3177\ : LocalMux
    port map (
            O => \N__22552\,
            I => \nx.n1604\
        );

    \I__3176\ : LocalMux
    port map (
            O => \N__22549\,
            I => \nx.n1604\
        );

    \I__3175\ : LocalMux
    port map (
            O => \N__22546\,
            I => \nx.n1604\
        );

    \I__3174\ : InMux
    port map (
            O => \N__22539\,
            I => \nx.n10799\
        );

    \I__3173\ : CascadeMux
    port map (
            O => \N__22536\,
            I => \N__22531\
        );

    \I__3172\ : InMux
    port map (
            O => \N__22535\,
            I => \N__22528\
        );

    \I__3171\ : InMux
    port map (
            O => \N__22534\,
            I => \N__22525\
        );

    \I__3170\ : InMux
    port map (
            O => \N__22531\,
            I => \N__22522\
        );

    \I__3169\ : LocalMux
    port map (
            O => \N__22528\,
            I => \nx.n1603\
        );

    \I__3168\ : LocalMux
    port map (
            O => \N__22525\,
            I => \nx.n1603\
        );

    \I__3167\ : LocalMux
    port map (
            O => \N__22522\,
            I => \nx.n1603\
        );

    \I__3166\ : InMux
    port map (
            O => \N__22515\,
            I => \nx.n10800\
        );

    \I__3165\ : CascadeMux
    port map (
            O => \N__22512\,
            I => \N__22507\
        );

    \I__3164\ : InMux
    port map (
            O => \N__22511\,
            I => \N__22504\
        );

    \I__3163\ : InMux
    port map (
            O => \N__22510\,
            I => \N__22501\
        );

    \I__3162\ : InMux
    port map (
            O => \N__22507\,
            I => \N__22498\
        );

    \I__3161\ : LocalMux
    port map (
            O => \N__22504\,
            I => \nx.n1602\
        );

    \I__3160\ : LocalMux
    port map (
            O => \N__22501\,
            I => \nx.n1602\
        );

    \I__3159\ : LocalMux
    port map (
            O => \N__22498\,
            I => \nx.n1602\
        );

    \I__3158\ : InMux
    port map (
            O => \N__22491\,
            I => \bfn_5_26_0_\
        );

    \I__3157\ : InMux
    port map (
            O => \N__22488\,
            I => \N__22484\
        );

    \I__3156\ : InMux
    port map (
            O => \N__22487\,
            I => \N__22480\
        );

    \I__3155\ : LocalMux
    port map (
            O => \N__22484\,
            I => \N__22477\
        );

    \I__3154\ : InMux
    port map (
            O => \N__22483\,
            I => \N__22474\
        );

    \I__3153\ : LocalMux
    port map (
            O => \N__22480\,
            I => \nx.n1601\
        );

    \I__3152\ : Odrv4
    port map (
            O => \N__22477\,
            I => \nx.n1601\
        );

    \I__3151\ : LocalMux
    port map (
            O => \N__22474\,
            I => \nx.n1601\
        );

    \I__3150\ : InMux
    port map (
            O => \N__22467\,
            I => \nx.n10802\
        );

    \I__3149\ : InMux
    port map (
            O => \N__22464\,
            I => \N__22459\
        );

    \I__3148\ : InMux
    port map (
            O => \N__22463\,
            I => \N__22456\
        );

    \I__3147\ : CascadeMux
    port map (
            O => \N__22462\,
            I => \N__22453\
        );

    \I__3146\ : LocalMux
    port map (
            O => \N__22459\,
            I => \N__22448\
        );

    \I__3145\ : LocalMux
    port map (
            O => \N__22456\,
            I => \N__22448\
        );

    \I__3144\ : InMux
    port map (
            O => \N__22453\,
            I => \N__22445\
        );

    \I__3143\ : Odrv4
    port map (
            O => \N__22448\,
            I => \nx.n1600\
        );

    \I__3142\ : LocalMux
    port map (
            O => \N__22445\,
            I => \nx.n1600\
        );

    \I__3141\ : InMux
    port map (
            O => \N__22440\,
            I => \nx.n10803\
        );

    \I__3140\ : InMux
    port map (
            O => \N__22437\,
            I => \N__22432\
        );

    \I__3139\ : InMux
    port map (
            O => \N__22436\,
            I => \N__22429\
        );

    \I__3138\ : InMux
    port map (
            O => \N__22435\,
            I => \N__22426\
        );

    \I__3137\ : LocalMux
    port map (
            O => \N__22432\,
            I => \nx.n1599\
        );

    \I__3136\ : LocalMux
    port map (
            O => \N__22429\,
            I => \nx.n1599\
        );

    \I__3135\ : LocalMux
    port map (
            O => \N__22426\,
            I => \nx.n1599\
        );

    \I__3134\ : InMux
    port map (
            O => \N__22419\,
            I => \nx.n10804\
        );

    \I__3133\ : InMux
    port map (
            O => \N__22416\,
            I => \N__22411\
        );

    \I__3132\ : InMux
    port map (
            O => \N__22415\,
            I => \N__22408\
        );

    \I__3131\ : InMux
    port map (
            O => \N__22414\,
            I => \N__22405\
        );

    \I__3130\ : LocalMux
    port map (
            O => \N__22411\,
            I => \N__22402\
        );

    \I__3129\ : LocalMux
    port map (
            O => \N__22408\,
            I => \nx.n1598\
        );

    \I__3128\ : LocalMux
    port map (
            O => \N__22405\,
            I => \nx.n1598\
        );

    \I__3127\ : Odrv4
    port map (
            O => \N__22402\,
            I => \nx.n1598\
        );

    \I__3126\ : CascadeMux
    port map (
            O => \N__22395\,
            I => \N__22382\
        );

    \I__3125\ : CascadeMux
    port map (
            O => \N__22394\,
            I => \N__22379\
        );

    \I__3124\ : CascadeMux
    port map (
            O => \N__22393\,
            I => \N__22376\
        );

    \I__3123\ : CascadeMux
    port map (
            O => \N__22392\,
            I => \N__22373\
        );

    \I__3122\ : CascadeMux
    port map (
            O => \N__22391\,
            I => \N__22370\
        );

    \I__3121\ : CascadeMux
    port map (
            O => \N__22390\,
            I => \N__22367\
        );

    \I__3120\ : CascadeMux
    port map (
            O => \N__22389\,
            I => \N__22364\
        );

    \I__3119\ : CascadeMux
    port map (
            O => \N__22388\,
            I => \N__22361\
        );

    \I__3118\ : CascadeMux
    port map (
            O => \N__22387\,
            I => \N__22358\
        );

    \I__3117\ : CascadeMux
    port map (
            O => \N__22386\,
            I => \N__22355\
        );

    \I__3116\ : CascadeMux
    port map (
            O => \N__22385\,
            I => \N__22352\
        );

    \I__3115\ : InMux
    port map (
            O => \N__22382\,
            I => \N__22347\
        );

    \I__3114\ : InMux
    port map (
            O => \N__22379\,
            I => \N__22347\
        );

    \I__3113\ : InMux
    port map (
            O => \N__22376\,
            I => \N__22340\
        );

    \I__3112\ : InMux
    port map (
            O => \N__22373\,
            I => \N__22340\
        );

    \I__3111\ : InMux
    port map (
            O => \N__22370\,
            I => \N__22340\
        );

    \I__3110\ : InMux
    port map (
            O => \N__22367\,
            I => \N__22333\
        );

    \I__3109\ : InMux
    port map (
            O => \N__22364\,
            I => \N__22333\
        );

    \I__3108\ : InMux
    port map (
            O => \N__22361\,
            I => \N__22333\
        );

    \I__3107\ : InMux
    port map (
            O => \N__22358\,
            I => \N__22326\
        );

    \I__3106\ : InMux
    port map (
            O => \N__22355\,
            I => \N__22326\
        );

    \I__3105\ : InMux
    port map (
            O => \N__22352\,
            I => \N__22326\
        );

    \I__3104\ : LocalMux
    port map (
            O => \N__22347\,
            I => \nx.n1631\
        );

    \I__3103\ : LocalMux
    port map (
            O => \N__22340\,
            I => \nx.n1631\
        );

    \I__3102\ : LocalMux
    port map (
            O => \N__22333\,
            I => \nx.n1631\
        );

    \I__3101\ : LocalMux
    port map (
            O => \N__22326\,
            I => \nx.n1631\
        );

    \I__3100\ : InMux
    port map (
            O => \N__22317\,
            I => \nx.n10805\
        );

    \I__3099\ : CEMux
    port map (
            O => \N__22314\,
            I => \N__22311\
        );

    \I__3098\ : LocalMux
    port map (
            O => \N__22311\,
            I => \N__22307\
        );

    \I__3097\ : CEMux
    port map (
            O => \N__22310\,
            I => \N__22304\
        );

    \I__3096\ : Span4Mux_v
    port map (
            O => \N__22307\,
            I => \N__22297\
        );

    \I__3095\ : LocalMux
    port map (
            O => \N__22304\,
            I => \N__22297\
        );

    \I__3094\ : CEMux
    port map (
            O => \N__22303\,
            I => \N__22294\
        );

    \I__3093\ : CEMux
    port map (
            O => \N__22302\,
            I => \N__22291\
        );

    \I__3092\ : Span4Mux_v
    port map (
            O => \N__22297\,
            I => \N__22286\
        );

    \I__3091\ : LocalMux
    port map (
            O => \N__22294\,
            I => \N__22286\
        );

    \I__3090\ : LocalMux
    port map (
            O => \N__22291\,
            I => \N__22283\
        );

    \I__3089\ : Span4Mux_h
    port map (
            O => \N__22286\,
            I => \N__22280\
        );

    \I__3088\ : Span4Mux_s2_h
    port map (
            O => \N__22283\,
            I => \N__22277\
        );

    \I__3087\ : Odrv4
    port map (
            O => \N__22280\,
            I => n7664
        );

    \I__3086\ : Odrv4
    port map (
            O => \N__22277\,
            I => n7664
        );

    \I__3085\ : CascadeMux
    port map (
            O => \N__22272\,
            I => \nx.n30_adj_777_cascade_\
        );

    \I__3084\ : InMux
    port map (
            O => \N__22269\,
            I => \N__22266\
        );

    \I__3083\ : LocalMux
    port map (
            O => \N__22266\,
            I => \nx.n43_adj_783\
        );

    \I__3082\ : InMux
    port map (
            O => \N__22263\,
            I => \bfn_5_25_0_\
        );

    \I__3081\ : CascadeMux
    port map (
            O => \N__22260\,
            I => \N__22255\
        );

    \I__3080\ : InMux
    port map (
            O => \N__22259\,
            I => \N__22252\
        );

    \I__3079\ : InMux
    port map (
            O => \N__22258\,
            I => \N__22249\
        );

    \I__3078\ : InMux
    port map (
            O => \N__22255\,
            I => \N__22246\
        );

    \I__3077\ : LocalMux
    port map (
            O => \N__22252\,
            I => \nx.n1609\
        );

    \I__3076\ : LocalMux
    port map (
            O => \N__22249\,
            I => \nx.n1609\
        );

    \I__3075\ : LocalMux
    port map (
            O => \N__22246\,
            I => \nx.n1609\
        );

    \I__3074\ : CascadeMux
    port map (
            O => \N__22239\,
            I => \N__22235\
        );

    \I__3073\ : CascadeMux
    port map (
            O => \N__22238\,
            I => \N__22232\
        );

    \I__3072\ : InMux
    port map (
            O => \N__22235\,
            I => \N__22229\
        );

    \I__3071\ : InMux
    port map (
            O => \N__22232\,
            I => \N__22226\
        );

    \I__3070\ : LocalMux
    port map (
            O => \N__22229\,
            I => \nx.n13602\
        );

    \I__3069\ : LocalMux
    port map (
            O => \N__22226\,
            I => \nx.n13602\
        );

    \I__3068\ : InMux
    port map (
            O => \N__22221\,
            I => \nx.n10794\
        );

    \I__3067\ : InMux
    port map (
            O => \N__22218\,
            I => \N__22213\
        );

    \I__3066\ : InMux
    port map (
            O => \N__22217\,
            I => \N__22210\
        );

    \I__3065\ : InMux
    port map (
            O => \N__22216\,
            I => \N__22207\
        );

    \I__3064\ : LocalMux
    port map (
            O => \N__22213\,
            I => \nx.n1608\
        );

    \I__3063\ : LocalMux
    port map (
            O => \N__22210\,
            I => \nx.n1608\
        );

    \I__3062\ : LocalMux
    port map (
            O => \N__22207\,
            I => \nx.n1608\
        );

    \I__3061\ : InMux
    port map (
            O => \N__22200\,
            I => \nx.n10795\
        );

    \I__3060\ : InMux
    port map (
            O => \N__22197\,
            I => \N__22192\
        );

    \I__3059\ : InMux
    port map (
            O => \N__22196\,
            I => \N__22189\
        );

    \I__3058\ : InMux
    port map (
            O => \N__22195\,
            I => \N__22186\
        );

    \I__3057\ : LocalMux
    port map (
            O => \N__22192\,
            I => \nx.n1607\
        );

    \I__3056\ : LocalMux
    port map (
            O => \N__22189\,
            I => \nx.n1607\
        );

    \I__3055\ : LocalMux
    port map (
            O => \N__22186\,
            I => \nx.n1607\
        );

    \I__3054\ : InMux
    port map (
            O => \N__22179\,
            I => \nx.n10796\
        );

    \I__3053\ : InMux
    port map (
            O => \N__22176\,
            I => \N__22171\
        );

    \I__3052\ : InMux
    port map (
            O => \N__22175\,
            I => \N__22168\
        );

    \I__3051\ : InMux
    port map (
            O => \N__22174\,
            I => \N__22165\
        );

    \I__3050\ : LocalMux
    port map (
            O => \N__22171\,
            I => \nx.n1606\
        );

    \I__3049\ : LocalMux
    port map (
            O => \N__22168\,
            I => \nx.n1606\
        );

    \I__3048\ : LocalMux
    port map (
            O => \N__22165\,
            I => \nx.n1606\
        );

    \I__3047\ : InMux
    port map (
            O => \N__22158\,
            I => \nx.n10797\
        );

    \I__3046\ : CascadeMux
    port map (
            O => \N__22155\,
            I => \N__22152\
        );

    \I__3045\ : InMux
    port map (
            O => \N__22152\,
            I => \N__22149\
        );

    \I__3044\ : LocalMux
    port map (
            O => \N__22149\,
            I => \nx.n1273\
        );

    \I__3043\ : InMux
    port map (
            O => \N__22146\,
            I => \nx.n10759\
        );

    \I__3042\ : CascadeMux
    port map (
            O => \N__22143\,
            I => \N__22139\
        );

    \I__3041\ : InMux
    port map (
            O => \N__22142\,
            I => \N__22136\
        );

    \I__3040\ : InMux
    port map (
            O => \N__22139\,
            I => \N__22133\
        );

    \I__3039\ : LocalMux
    port map (
            O => \N__22136\,
            I => \nx.n1205\
        );

    \I__3038\ : LocalMux
    port map (
            O => \N__22133\,
            I => \nx.n1205\
        );

    \I__3037\ : InMux
    port map (
            O => \N__22128\,
            I => \N__22125\
        );

    \I__3036\ : LocalMux
    port map (
            O => \N__22125\,
            I => \nx.n1272\
        );

    \I__3035\ : InMux
    port map (
            O => \N__22122\,
            I => \nx.n10760\
        );

    \I__3034\ : CascadeMux
    port map (
            O => \N__22119\,
            I => \N__22115\
        );

    \I__3033\ : CascadeMux
    port map (
            O => \N__22118\,
            I => \N__22112\
        );

    \I__3032\ : InMux
    port map (
            O => \N__22115\,
            I => \N__22108\
        );

    \I__3031\ : InMux
    port map (
            O => \N__22112\,
            I => \N__22105\
        );

    \I__3030\ : InMux
    port map (
            O => \N__22111\,
            I => \N__22102\
        );

    \I__3029\ : LocalMux
    port map (
            O => \N__22108\,
            I => \nx.n1204\
        );

    \I__3028\ : LocalMux
    port map (
            O => \N__22105\,
            I => \nx.n1204\
        );

    \I__3027\ : LocalMux
    port map (
            O => \N__22102\,
            I => \nx.n1204\
        );

    \I__3026\ : InMux
    port map (
            O => \N__22095\,
            I => \N__22092\
        );

    \I__3025\ : LocalMux
    port map (
            O => \N__22092\,
            I => \N__22089\
        );

    \I__3024\ : Odrv4
    port map (
            O => \N__22089\,
            I => \nx.n1271\
        );

    \I__3023\ : InMux
    port map (
            O => \N__22086\,
            I => \nx.n10761\
        );

    \I__3022\ : InMux
    port map (
            O => \N__22083\,
            I => \nx.n10762\
        );

    \I__3021\ : CascadeMux
    port map (
            O => \N__22080\,
            I => \N__22077\
        );

    \I__3020\ : InMux
    port map (
            O => \N__22077\,
            I => \N__22074\
        );

    \I__3019\ : LocalMux
    port map (
            O => \N__22074\,
            I => \N__22070\
        );

    \I__3018\ : InMux
    port map (
            O => \N__22073\,
            I => \N__22067\
        );

    \I__3017\ : Odrv4
    port map (
            O => \N__22070\,
            I => \nx.n1202\
        );

    \I__3016\ : LocalMux
    port map (
            O => \N__22067\,
            I => \nx.n1202\
        );

    \I__3015\ : InMux
    port map (
            O => \N__22062\,
            I => \bfn_5_23_0_\
        );

    \I__3014\ : CascadeMux
    port map (
            O => \N__22059\,
            I => \N__22055\
        );

    \I__3013\ : CascadeMux
    port map (
            O => \N__22058\,
            I => \N__22052\
        );

    \I__3012\ : InMux
    port map (
            O => \N__22055\,
            I => \N__22047\
        );

    \I__3011\ : InMux
    port map (
            O => \N__22052\,
            I => \N__22047\
        );

    \I__3010\ : LocalMux
    port map (
            O => \N__22047\,
            I => \nx.n1301\
        );

    \I__3009\ : InMux
    port map (
            O => \N__22044\,
            I => \N__22041\
        );

    \I__3008\ : LocalMux
    port map (
            O => \N__22041\,
            I => \N__22037\
        );

    \I__3007\ : InMux
    port map (
            O => \N__22040\,
            I => \N__22034\
        );

    \I__3006\ : Span4Mux_h
    port map (
            O => \N__22037\,
            I => \N__22031\
        );

    \I__3005\ : LocalMux
    port map (
            O => \N__22034\,
            I => delay_counter_19
        );

    \I__3004\ : Odrv4
    port map (
            O => \N__22031\,
            I => delay_counter_19
        );

    \I__3003\ : InMux
    port map (
            O => \N__22026\,
            I => \N__22023\
        );

    \I__3002\ : LocalMux
    port map (
            O => \N__22023\,
            I => \N__22019\
        );

    \I__3001\ : InMux
    port map (
            O => \N__22022\,
            I => \N__22016\
        );

    \I__3000\ : Span4Mux_h
    port map (
            O => \N__22019\,
            I => \N__22013\
        );

    \I__2999\ : LocalMux
    port map (
            O => \N__22016\,
            I => delay_counter_20
        );

    \I__2998\ : Odrv4
    port map (
            O => \N__22013\,
            I => delay_counter_20
        );

    \I__2997\ : InMux
    port map (
            O => \N__22008\,
            I => \N__22005\
        );

    \I__2996\ : LocalMux
    port map (
            O => \N__22005\,
            I => \N__22002\
        );

    \I__2995\ : Odrv12
    port map (
            O => \N__22002\,
            I => n4
        );

    \I__2994\ : CascadeMux
    port map (
            O => \N__21999\,
            I => \N__21995\
        );

    \I__2993\ : InMux
    port map (
            O => \N__21998\,
            I => \N__21992\
        );

    \I__2992\ : InMux
    port map (
            O => \N__21995\,
            I => \N__21989\
        );

    \I__2991\ : LocalMux
    port map (
            O => \N__21992\,
            I => \nx.n1203\
        );

    \I__2990\ : LocalMux
    port map (
            O => \N__21989\,
            I => \nx.n1203\
        );

    \I__2989\ : CascadeMux
    port map (
            O => \N__21984\,
            I => \N__21977\
        );

    \I__2988\ : CascadeMux
    port map (
            O => \N__21983\,
            I => \N__21974\
        );

    \I__2987\ : CascadeMux
    port map (
            O => \N__21982\,
            I => \N__21969\
        );

    \I__2986\ : CascadeMux
    port map (
            O => \N__21981\,
            I => \N__21966\
        );

    \I__2985\ : InMux
    port map (
            O => \N__21980\,
            I => \N__21962\
        );

    \I__2984\ : InMux
    port map (
            O => \N__21977\,
            I => \N__21955\
        );

    \I__2983\ : InMux
    port map (
            O => \N__21974\,
            I => \N__21955\
        );

    \I__2982\ : InMux
    port map (
            O => \N__21973\,
            I => \N__21955\
        );

    \I__2981\ : InMux
    port map (
            O => \N__21972\,
            I => \N__21950\
        );

    \I__2980\ : InMux
    port map (
            O => \N__21969\,
            I => \N__21950\
        );

    \I__2979\ : InMux
    port map (
            O => \N__21966\,
            I => \N__21945\
        );

    \I__2978\ : InMux
    port map (
            O => \N__21965\,
            I => \N__21945\
        );

    \I__2977\ : LocalMux
    port map (
            O => \N__21962\,
            I => \nx.n1235\
        );

    \I__2976\ : LocalMux
    port map (
            O => \N__21955\,
            I => \nx.n1235\
        );

    \I__2975\ : LocalMux
    port map (
            O => \N__21950\,
            I => \nx.n1235\
        );

    \I__2974\ : LocalMux
    port map (
            O => \N__21945\,
            I => \nx.n1235\
        );

    \I__2973\ : InMux
    port map (
            O => \N__21936\,
            I => \N__21933\
        );

    \I__2972\ : LocalMux
    port map (
            O => \N__21933\,
            I => \nx.n1270\
        );

    \I__2971\ : CascadeMux
    port map (
            O => \N__21930\,
            I => \N__21926\
        );

    \I__2970\ : InMux
    port map (
            O => \N__21929\,
            I => \N__21918\
        );

    \I__2969\ : InMux
    port map (
            O => \N__21926\,
            I => \N__21918\
        );

    \I__2968\ : InMux
    port map (
            O => \N__21925\,
            I => \N__21918\
        );

    \I__2967\ : LocalMux
    port map (
            O => \N__21918\,
            I => \nx.n1302\
        );

    \I__2966\ : CascadeMux
    port map (
            O => \N__21915\,
            I => \nx.n49_adj_784_cascade_\
        );

    \I__2965\ : InMux
    port map (
            O => \N__21912\,
            I => \N__21909\
        );

    \I__2964\ : LocalMux
    port map (
            O => \N__21909\,
            I => \N__21906\
        );

    \I__2963\ : Span4Mux_h
    port map (
            O => \N__21906\,
            I => \N__21903\
        );

    \I__2962\ : Odrv4
    port map (
            O => \N__21903\,
            I => \nx.n54\
        );

    \I__2961\ : CascadeMux
    port map (
            O => \N__21900\,
            I => \N__21896\
        );

    \I__2960\ : InMux
    port map (
            O => \N__21899\,
            I => \N__21892\
        );

    \I__2959\ : InMux
    port map (
            O => \N__21896\,
            I => \N__21889\
        );

    \I__2958\ : InMux
    port map (
            O => \N__21895\,
            I => \N__21886\
        );

    \I__2957\ : LocalMux
    port map (
            O => \N__21892\,
            I => \nx.n1106\
        );

    \I__2956\ : LocalMux
    port map (
            O => \N__21889\,
            I => \nx.n1106\
        );

    \I__2955\ : LocalMux
    port map (
            O => \N__21886\,
            I => \nx.n1106\
        );

    \I__2954\ : InMux
    port map (
            O => \N__21879\,
            I => \N__21876\
        );

    \I__2953\ : LocalMux
    port map (
            O => \N__21876\,
            I => \nx.n1173\
        );

    \I__2952\ : InMux
    port map (
            O => \N__21873\,
            I => \nx.n10752\
        );

    \I__2951\ : InMux
    port map (
            O => \N__21870\,
            I => \N__21867\
        );

    \I__2950\ : LocalMux
    port map (
            O => \N__21867\,
            I => \nx.n1172\
        );

    \I__2949\ : InMux
    port map (
            O => \N__21864\,
            I => \nx.n10753\
        );

    \I__2948\ : InMux
    port map (
            O => \N__21861\,
            I => \N__21857\
        );

    \I__2947\ : CascadeMux
    port map (
            O => \N__21860\,
            I => \N__21854\
        );

    \I__2946\ : LocalMux
    port map (
            O => \N__21857\,
            I => \N__21850\
        );

    \I__2945\ : InMux
    port map (
            O => \N__21854\,
            I => \N__21847\
        );

    \I__2944\ : InMux
    port map (
            O => \N__21853\,
            I => \N__21844\
        );

    \I__2943\ : Odrv4
    port map (
            O => \N__21850\,
            I => \nx.n1104\
        );

    \I__2942\ : LocalMux
    port map (
            O => \N__21847\,
            I => \nx.n1104\
        );

    \I__2941\ : LocalMux
    port map (
            O => \N__21844\,
            I => \nx.n1104\
        );

    \I__2940\ : InMux
    port map (
            O => \N__21837\,
            I => \N__21834\
        );

    \I__2939\ : LocalMux
    port map (
            O => \N__21834\,
            I => \nx.n1171\
        );

    \I__2938\ : InMux
    port map (
            O => \N__21831\,
            I => \nx.n10754\
        );

    \I__2937\ : CascadeMux
    port map (
            O => \N__21828\,
            I => \N__21822\
        );

    \I__2936\ : CascadeMux
    port map (
            O => \N__21827\,
            I => \N__21817\
        );

    \I__2935\ : CascadeMux
    port map (
            O => \N__21826\,
            I => \N__21813\
        );

    \I__2934\ : CascadeMux
    port map (
            O => \N__21825\,
            I => \N__21810\
        );

    \I__2933\ : InMux
    port map (
            O => \N__21822\,
            I => \N__21804\
        );

    \I__2932\ : InMux
    port map (
            O => \N__21821\,
            I => \N__21804\
        );

    \I__2931\ : InMux
    port map (
            O => \N__21820\,
            I => \N__21801\
        );

    \I__2930\ : InMux
    port map (
            O => \N__21817\,
            I => \N__21790\
        );

    \I__2929\ : InMux
    port map (
            O => \N__21816\,
            I => \N__21790\
        );

    \I__2928\ : InMux
    port map (
            O => \N__21813\,
            I => \N__21790\
        );

    \I__2927\ : InMux
    port map (
            O => \N__21810\,
            I => \N__21790\
        );

    \I__2926\ : InMux
    port map (
            O => \N__21809\,
            I => \N__21790\
        );

    \I__2925\ : LocalMux
    port map (
            O => \N__21804\,
            I => \N__21787\
        );

    \I__2924\ : LocalMux
    port map (
            O => \N__21801\,
            I => \nx.n1136\
        );

    \I__2923\ : LocalMux
    port map (
            O => \N__21790\,
            I => \nx.n1136\
        );

    \I__2922\ : Odrv4
    port map (
            O => \N__21787\,
            I => \nx.n1136\
        );

    \I__2921\ : InMux
    port map (
            O => \N__21780\,
            I => \nx.n10755\
        );

    \I__2920\ : InMux
    port map (
            O => \N__21777\,
            I => \N__21774\
        );

    \I__2919\ : LocalMux
    port map (
            O => \N__21774\,
            I => \N__21771\
        );

    \I__2918\ : Span4Mux_h
    port map (
            O => \N__21771\,
            I => \N__21768\
        );

    \I__2917\ : Odrv4
    port map (
            O => \N__21768\,
            I => \nx.n1277\
        );

    \I__2916\ : InMux
    port map (
            O => \N__21765\,
            I => \bfn_5_22_0_\
        );

    \I__2915\ : CascadeMux
    port map (
            O => \N__21762\,
            I => \N__21757\
        );

    \I__2914\ : InMux
    port map (
            O => \N__21761\,
            I => \N__21754\
        );

    \I__2913\ : InMux
    port map (
            O => \N__21760\,
            I => \N__21751\
        );

    \I__2912\ : InMux
    port map (
            O => \N__21757\,
            I => \N__21748\
        );

    \I__2911\ : LocalMux
    port map (
            O => \N__21754\,
            I => \nx.n1209\
        );

    \I__2910\ : LocalMux
    port map (
            O => \N__21751\,
            I => \nx.n1209\
        );

    \I__2909\ : LocalMux
    port map (
            O => \N__21748\,
            I => \nx.n1209\
        );

    \I__2908\ : InMux
    port map (
            O => \N__21741\,
            I => \N__21738\
        );

    \I__2907\ : LocalMux
    port map (
            O => \N__21738\,
            I => \N__21735\
        );

    \I__2906\ : Span4Mux_h
    port map (
            O => \N__21735\,
            I => \N__21732\
        );

    \I__2905\ : Odrv4
    port map (
            O => \N__21732\,
            I => \nx.n1276\
        );

    \I__2904\ : InMux
    port map (
            O => \N__21729\,
            I => \nx.n10756\
        );

    \I__2903\ : CascadeMux
    port map (
            O => \N__21726\,
            I => \N__21721\
        );

    \I__2902\ : InMux
    port map (
            O => \N__21725\,
            I => \N__21716\
        );

    \I__2901\ : InMux
    port map (
            O => \N__21724\,
            I => \N__21716\
        );

    \I__2900\ : InMux
    port map (
            O => \N__21721\,
            I => \N__21713\
        );

    \I__2899\ : LocalMux
    port map (
            O => \N__21716\,
            I => \nx.n1208\
        );

    \I__2898\ : LocalMux
    port map (
            O => \N__21713\,
            I => \nx.n1208\
        );

    \I__2897\ : InMux
    port map (
            O => \N__21708\,
            I => \N__21705\
        );

    \I__2896\ : LocalMux
    port map (
            O => \N__21705\,
            I => \nx.n1275\
        );

    \I__2895\ : InMux
    port map (
            O => \N__21702\,
            I => \nx.n10757\
        );

    \I__2894\ : CascadeMux
    port map (
            O => \N__21699\,
            I => \N__21694\
        );

    \I__2893\ : InMux
    port map (
            O => \N__21698\,
            I => \N__21689\
        );

    \I__2892\ : InMux
    port map (
            O => \N__21697\,
            I => \N__21689\
        );

    \I__2891\ : InMux
    port map (
            O => \N__21694\,
            I => \N__21686\
        );

    \I__2890\ : LocalMux
    port map (
            O => \N__21689\,
            I => \nx.n1207\
        );

    \I__2889\ : LocalMux
    port map (
            O => \N__21686\,
            I => \nx.n1207\
        );

    \I__2888\ : InMux
    port map (
            O => \N__21681\,
            I => \N__21678\
        );

    \I__2887\ : LocalMux
    port map (
            O => \N__21678\,
            I => \nx.n1274\
        );

    \I__2886\ : InMux
    port map (
            O => \N__21675\,
            I => \nx.n10758\
        );

    \I__2885\ : CascadeMux
    port map (
            O => \N__21672\,
            I => \N__21667\
        );

    \I__2884\ : InMux
    port map (
            O => \N__21671\,
            I => \N__21662\
        );

    \I__2883\ : InMux
    port map (
            O => \N__21670\,
            I => \N__21662\
        );

    \I__2882\ : InMux
    port map (
            O => \N__21667\,
            I => \N__21659\
        );

    \I__2881\ : LocalMux
    port map (
            O => \N__21662\,
            I => \nx.n1206\
        );

    \I__2880\ : LocalMux
    port map (
            O => \N__21659\,
            I => \nx.n1206\
        );

    \I__2879\ : CascadeMux
    port map (
            O => \N__21654\,
            I => \nx.n1109_cascade_\
        );

    \I__2878\ : CascadeMux
    port map (
            O => \N__21651\,
            I => \nx.n9737_cascade_\
        );

    \I__2877\ : CascadeMux
    port map (
            O => \N__21648\,
            I => \nx.n12_adj_673_cascade_\
        );

    \I__2876\ : InMux
    port map (
            O => \N__21645\,
            I => \N__21642\
        );

    \I__2875\ : LocalMux
    port map (
            O => \N__21642\,
            I => \N__21639\
        );

    \I__2874\ : Odrv4
    port map (
            O => \N__21639\,
            I => \nx.n1177\
        );

    \I__2873\ : InMux
    port map (
            O => \N__21636\,
            I => \bfn_5_21_0_\
        );

    \I__2872\ : CascadeMux
    port map (
            O => \N__21633\,
            I => \N__21629\
        );

    \I__2871\ : InMux
    port map (
            O => \N__21632\,
            I => \N__21626\
        );

    \I__2870\ : InMux
    port map (
            O => \N__21629\,
            I => \N__21623\
        );

    \I__2869\ : LocalMux
    port map (
            O => \N__21626\,
            I => \nx.n1109\
        );

    \I__2868\ : LocalMux
    port map (
            O => \N__21623\,
            I => \nx.n1109\
        );

    \I__2867\ : CascadeMux
    port map (
            O => \N__21618\,
            I => \N__21615\
        );

    \I__2866\ : InMux
    port map (
            O => \N__21615\,
            I => \N__21612\
        );

    \I__2865\ : LocalMux
    port map (
            O => \N__21612\,
            I => \nx.n1176\
        );

    \I__2864\ : InMux
    port map (
            O => \N__21609\,
            I => \nx.n10749\
        );

    \I__2863\ : CascadeMux
    port map (
            O => \N__21606\,
            I => \N__21602\
        );

    \I__2862\ : InMux
    port map (
            O => \N__21605\,
            I => \N__21598\
        );

    \I__2861\ : InMux
    port map (
            O => \N__21602\,
            I => \N__21595\
        );

    \I__2860\ : InMux
    port map (
            O => \N__21601\,
            I => \N__21592\
        );

    \I__2859\ : LocalMux
    port map (
            O => \N__21598\,
            I => \nx.n1108\
        );

    \I__2858\ : LocalMux
    port map (
            O => \N__21595\,
            I => \nx.n1108\
        );

    \I__2857\ : LocalMux
    port map (
            O => \N__21592\,
            I => \nx.n1108\
        );

    \I__2856\ : InMux
    port map (
            O => \N__21585\,
            I => \N__21582\
        );

    \I__2855\ : LocalMux
    port map (
            O => \N__21582\,
            I => \nx.n1175\
        );

    \I__2854\ : InMux
    port map (
            O => \N__21579\,
            I => \nx.n10750\
        );

    \I__2853\ : CascadeMux
    port map (
            O => \N__21576\,
            I => \N__21573\
        );

    \I__2852\ : InMux
    port map (
            O => \N__21573\,
            I => \N__21570\
        );

    \I__2851\ : LocalMux
    port map (
            O => \N__21570\,
            I => \nx.n1174\
        );

    \I__2850\ : InMux
    port map (
            O => \N__21567\,
            I => \nx.n10751\
        );

    \I__2849\ : InMux
    port map (
            O => \N__21564\,
            I => \N__21561\
        );

    \I__2848\ : LocalMux
    port map (
            O => \N__21561\,
            I => \N__21557\
        );

    \I__2847\ : CascadeMux
    port map (
            O => \N__21560\,
            I => \N__21553\
        );

    \I__2846\ : Span4Mux_h
    port map (
            O => \N__21557\,
            I => \N__21550\
        );

    \I__2845\ : InMux
    port map (
            O => \N__21556\,
            I => \N__21547\
        );

    \I__2844\ : InMux
    port map (
            O => \N__21553\,
            I => \N__21544\
        );

    \I__2843\ : Odrv4
    port map (
            O => \N__21550\,
            I => timer_11
        );

    \I__2842\ : LocalMux
    port map (
            O => \N__21547\,
            I => timer_11
        );

    \I__2841\ : LocalMux
    port map (
            O => \N__21544\,
            I => timer_11
        );

    \I__2840\ : InMux
    port map (
            O => \N__21537\,
            I => \N__21534\
        );

    \I__2839\ : LocalMux
    port map (
            O => \N__21534\,
            I => \N__21531\
        );

    \I__2838\ : Sp12to4
    port map (
            O => \N__21531\,
            I => \N__21528\
        );

    \I__2837\ : Span12Mux_v
    port map (
            O => \N__21528\,
            I => \N__21525\
        );

    \I__2836\ : Odrv12
    port map (
            O => \N__21525\,
            I => pin_in_0
        );

    \I__2835\ : InMux
    port map (
            O => \N__21522\,
            I => \N__21519\
        );

    \I__2834\ : LocalMux
    port map (
            O => \N__21519\,
            I => \N__21516\
        );

    \I__2833\ : Span12Mux_h
    port map (
            O => \N__21516\,
            I => \N__21513\
        );

    \I__2832\ : Span12Mux_v
    port map (
            O => \N__21513\,
            I => \N__21510\
        );

    \I__2831\ : Odrv12
    port map (
            O => \N__21510\,
            I => pin_in_1
        );

    \I__2830\ : InMux
    port map (
            O => \N__21507\,
            I => \N__21504\
        );

    \I__2829\ : LocalMux
    port map (
            O => \N__21504\,
            I => \N__21501\
        );

    \I__2828\ : Odrv4
    port map (
            O => \N__21501\,
            I => n13378
        );

    \I__2827\ : InMux
    port map (
            O => \N__21498\,
            I => \N__21495\
        );

    \I__2826\ : LocalMux
    port map (
            O => \N__21495\,
            I => \N__21492\
        );

    \I__2825\ : Span4Mux_h
    port map (
            O => \N__21492\,
            I => \N__21489\
        );

    \I__2824\ : Span4Mux_v
    port map (
            O => \N__21489\,
            I => \N__21486\
        );

    \I__2823\ : Sp12to4
    port map (
            O => \N__21486\,
            I => \N__21483\
        );

    \I__2822\ : Span12Mux_v
    port map (
            O => \N__21483\,
            I => \N__21480\
        );

    \I__2821\ : Odrv12
    port map (
            O => \N__21480\,
            I => pin_in_4
        );

    \I__2820\ : InMux
    port map (
            O => \N__21477\,
            I => \N__21474\
        );

    \I__2819\ : LocalMux
    port map (
            O => \N__21474\,
            I => \N__21471\
        );

    \I__2818\ : Span4Mux_v
    port map (
            O => \N__21471\,
            I => \N__21468\
        );

    \I__2817\ : Span4Mux_v
    port map (
            O => \N__21468\,
            I => \N__21465\
        );

    \I__2816\ : Span4Mux_v
    port map (
            O => \N__21465\,
            I => \N__21462\
        );

    \I__2815\ : Span4Mux_h
    port map (
            O => \N__21462\,
            I => \N__21459\
        );

    \I__2814\ : Odrv4
    port map (
            O => \N__21459\,
            I => pin_in_5
        );

    \I__2813\ : InMux
    port map (
            O => \N__21456\,
            I => \N__21453\
        );

    \I__2812\ : LocalMux
    port map (
            O => \N__21453\,
            I => n13382
        );

    \I__2811\ : CascadeMux
    port map (
            O => \N__21450\,
            I => \n13381_cascade_\
        );

    \I__2810\ : InMux
    port map (
            O => \N__21447\,
            I => \N__21444\
        );

    \I__2809\ : LocalMux
    port map (
            O => \N__21444\,
            I => \N__21441\
        );

    \I__2808\ : Odrv4
    port map (
            O => \N__21441\,
            I => n13613
        );

    \I__2807\ : InMux
    port map (
            O => \N__21438\,
            I => \N__21434\
        );

    \I__2806\ : InMux
    port map (
            O => \N__21437\,
            I => \N__21431\
        );

    \I__2805\ : LocalMux
    port map (
            O => \N__21434\,
            I => neo_pixel_transmitter_t0_11
        );

    \I__2804\ : LocalMux
    port map (
            O => \N__21431\,
            I => neo_pixel_transmitter_t0_11
        );

    \I__2803\ : InMux
    port map (
            O => \N__21426\,
            I => \N__21423\
        );

    \I__2802\ : LocalMux
    port map (
            O => \N__21423\,
            I => \N__21420\
        );

    \I__2801\ : Span4Mux_h
    port map (
            O => \N__21420\,
            I => \N__21417\
        );

    \I__2800\ : Odrv4
    port map (
            O => \N__21417\,
            I => \nx.n22_adj_749\
        );

    \I__2799\ : InMux
    port map (
            O => \N__21414\,
            I => \N__21410\
        );

    \I__2798\ : InMux
    port map (
            O => \N__21413\,
            I => \N__21407\
        );

    \I__2797\ : LocalMux
    port map (
            O => \N__21410\,
            I => neo_pixel_transmitter_t0_19
        );

    \I__2796\ : LocalMux
    port map (
            O => \N__21407\,
            I => neo_pixel_transmitter_t0_19
        );

    \I__2795\ : InMux
    port map (
            O => \N__21402\,
            I => \N__21399\
        );

    \I__2794\ : LocalMux
    port map (
            O => \N__21399\,
            I => \N__21396\
        );

    \I__2793\ : Span4Mux_h
    port map (
            O => \N__21396\,
            I => \N__21393\
        );

    \I__2792\ : Odrv4
    port map (
            O => \N__21393\,
            I => \nx.n14\
        );

    \I__2791\ : InMux
    port map (
            O => \N__21390\,
            I => \N__21387\
        );

    \I__2790\ : LocalMux
    port map (
            O => \N__21387\,
            I => \nx.n13438\
        );

    \I__2789\ : InMux
    port map (
            O => \N__21384\,
            I => \N__21379\
        );

    \I__2788\ : InMux
    port map (
            O => \N__21383\,
            I => \N__21376\
        );

    \I__2787\ : InMux
    port map (
            O => \N__21382\,
            I => \N__21372\
        );

    \I__2786\ : LocalMux
    port map (
            O => \N__21379\,
            I => \N__21367\
        );

    \I__2785\ : LocalMux
    port map (
            O => \N__21376\,
            I => \N__21367\
        );

    \I__2784\ : InMux
    port map (
            O => \N__21375\,
            I => \N__21364\
        );

    \I__2783\ : LocalMux
    port map (
            O => \N__21372\,
            I => \N__21361\
        );

    \I__2782\ : Span4Mux_v
    port map (
            O => \N__21367\,
            I => \N__21356\
        );

    \I__2781\ : LocalMux
    port map (
            O => \N__21364\,
            I => \N__21356\
        );

    \I__2780\ : Odrv4
    port map (
            O => \N__21361\,
            I => \nx.one_wire_N_599_3\
        );

    \I__2779\ : Odrv4
    port map (
            O => \N__21356\,
            I => \nx.one_wire_N_599_3\
        );

    \I__2778\ : CascadeMux
    port map (
            O => \N__21351\,
            I => \nx.n11908_cascade_\
        );

    \I__2777\ : InMux
    port map (
            O => \N__21348\,
            I => \N__21342\
        );

    \I__2776\ : InMux
    port map (
            O => \N__21347\,
            I => \N__21342\
        );

    \I__2775\ : LocalMux
    port map (
            O => \N__21342\,
            I => \nx.n11926\
        );

    \I__2774\ : CascadeMux
    port map (
            O => \N__21339\,
            I => \nx.n11926_cascade_\
        );

    \I__2773\ : CascadeMux
    port map (
            O => \N__21336\,
            I => \n7671_cascade_\
        );

    \I__2772\ : InMux
    port map (
            O => \N__21333\,
            I => \N__21328\
        );

    \I__2771\ : InMux
    port map (
            O => \N__21332\,
            I => \N__21322\
        );

    \I__2770\ : InMux
    port map (
            O => \N__21331\,
            I => \N__21322\
        );

    \I__2769\ : LocalMux
    port map (
            O => \N__21328\,
            I => \N__21319\
        );

    \I__2768\ : InMux
    port map (
            O => \N__21327\,
            I => \N__21316\
        );

    \I__2767\ : LocalMux
    port map (
            O => \N__21322\,
            I => \N__21313\
        );

    \I__2766\ : Span4Mux_v
    port map (
            O => \N__21319\,
            I => \N__21310\
        );

    \I__2765\ : LocalMux
    port map (
            O => \N__21316\,
            I => \N__21307\
        );

    \I__2764\ : Span4Mux_h
    port map (
            O => \N__21313\,
            I => \N__21304\
        );

    \I__2763\ : Odrv4
    port map (
            O => \N__21310\,
            I => \nx.one_wire_N_599_2\
        );

    \I__2762\ : Odrv4
    port map (
            O => \N__21307\,
            I => \nx.one_wire_N_599_2\
        );

    \I__2761\ : Odrv4
    port map (
            O => \N__21304\,
            I => \nx.one_wire_N_599_2\
        );

    \I__2760\ : InMux
    port map (
            O => \N__21297\,
            I => \N__21293\
        );

    \I__2759\ : InMux
    port map (
            O => \N__21296\,
            I => \N__21290\
        );

    \I__2758\ : LocalMux
    port map (
            O => \N__21293\,
            I => \N__21287\
        );

    \I__2757\ : LocalMux
    port map (
            O => \N__21290\,
            I => \N__21284\
        );

    \I__2756\ : Span4Mux_v
    port map (
            O => \N__21287\,
            I => \N__21281\
        );

    \I__2755\ : Odrv4
    port map (
            O => \N__21284\,
            I => \nx.n4_adj_771\
        );

    \I__2754\ : Odrv4
    port map (
            O => \N__21281\,
            I => \nx.n4_adj_771\
        );

    \I__2753\ : CascadeMux
    port map (
            O => \N__21276\,
            I => \N__21273\
        );

    \I__2752\ : InMux
    port map (
            O => \N__21273\,
            I => \N__21270\
        );

    \I__2751\ : LocalMux
    port map (
            O => \N__21270\,
            I => \N__21265\
        );

    \I__2750\ : InMux
    port map (
            O => \N__21269\,
            I => \N__21262\
        );

    \I__2749\ : InMux
    port map (
            O => \N__21268\,
            I => \N__21259\
        );

    \I__2748\ : Span4Mux_v
    port map (
            O => \N__21265\,
            I => \N__21255\
        );

    \I__2747\ : LocalMux
    port map (
            O => \N__21262\,
            I => \N__21250\
        );

    \I__2746\ : LocalMux
    port map (
            O => \N__21259\,
            I => \N__21250\
        );

    \I__2745\ : InMux
    port map (
            O => \N__21258\,
            I => \N__21247\
        );

    \I__2744\ : Odrv4
    port map (
            O => \N__21255\,
            I => \nx.n9747\
        );

    \I__2743\ : Odrv4
    port map (
            O => \N__21250\,
            I => \nx.n9747\
        );

    \I__2742\ : LocalMux
    port map (
            O => \N__21247\,
            I => \nx.n9747\
        );

    \I__2741\ : InMux
    port map (
            O => \N__21240\,
            I => \N__21237\
        );

    \I__2740\ : LocalMux
    port map (
            O => \N__21237\,
            I => \nx.n12381\
        );

    \I__2739\ : InMux
    port map (
            O => \N__21234\,
            I => \N__21231\
        );

    \I__2738\ : LocalMux
    port map (
            O => \N__21231\,
            I => \N__21228\
        );

    \I__2737\ : Span4Mux_v
    port map (
            O => \N__21228\,
            I => \N__21225\
        );

    \I__2736\ : Sp12to4
    port map (
            O => \N__21225\,
            I => \N__21222\
        );

    \I__2735\ : Span12Mux_h
    port map (
            O => \N__21222\,
            I => \N__21219\
        );

    \I__2734\ : Odrv12
    port map (
            O => \N__21219\,
            I => pin_in_10
        );

    \I__2733\ : CascadeMux
    port map (
            O => \N__21216\,
            I => \N__21213\
        );

    \I__2732\ : InMux
    port map (
            O => \N__21213\,
            I => \N__21210\
        );

    \I__2731\ : LocalMux
    port map (
            O => \N__21210\,
            I => \N__21207\
        );

    \I__2730\ : Span4Mux_v
    port map (
            O => \N__21207\,
            I => \N__21204\
        );

    \I__2729\ : Span4Mux_h
    port map (
            O => \N__21204\,
            I => \N__21201\
        );

    \I__2728\ : Span4Mux_v
    port map (
            O => \N__21201\,
            I => \N__21198\
        );

    \I__2727\ : Span4Mux_v
    port map (
            O => \N__21198\,
            I => \N__21195\
        );

    \I__2726\ : Odrv4
    port map (
            O => \N__21195\,
            I => pin_in_11
        );

    \I__2725\ : IoInMux
    port map (
            O => \N__21192\,
            I => \N__21189\
        );

    \I__2724\ : LocalMux
    port map (
            O => \N__21189\,
            I => \N__21186\
        );

    \I__2723\ : IoSpan4Mux
    port map (
            O => \N__21186\,
            I => \N__21183\
        );

    \I__2722\ : Span4Mux_s0_h
    port map (
            O => \N__21183\,
            I => \N__21180\
        );

    \I__2721\ : Sp12to4
    port map (
            O => \N__21180\,
            I => \N__21177\
        );

    \I__2720\ : Span12Mux_v
    port map (
            O => \N__21177\,
            I => \N__21173\
        );

    \I__2719\ : InMux
    port map (
            O => \N__21176\,
            I => \N__21170\
        );

    \I__2718\ : Odrv12
    port map (
            O => \N__21173\,
            I => pin_oe_6
        );

    \I__2717\ : LocalMux
    port map (
            O => \N__21170\,
            I => pin_oe_6
        );

    \I__2716\ : InMux
    port map (
            O => \N__21165\,
            I => \N__21162\
        );

    \I__2715\ : LocalMux
    port map (
            O => \N__21162\,
            I => \N__21159\
        );

    \I__2714\ : Span4Mux_h
    port map (
            O => \N__21159\,
            I => \N__21156\
        );

    \I__2713\ : Sp12to4
    port map (
            O => \N__21156\,
            I => \N__21153\
        );

    \I__2712\ : Span12Mux_v
    port map (
            O => \N__21153\,
            I => \N__21150\
        );

    \I__2711\ : Odrv12
    port map (
            O => \N__21150\,
            I => pin_in_9
        );

    \I__2710\ : CascadeMux
    port map (
            O => \N__21147\,
            I => \N__21144\
        );

    \I__2709\ : InMux
    port map (
            O => \N__21144\,
            I => \N__21141\
        );

    \I__2708\ : LocalMux
    port map (
            O => \N__21141\,
            I => \N__21138\
        );

    \I__2707\ : Span4Mux_h
    port map (
            O => \N__21138\,
            I => \N__21135\
        );

    \I__2706\ : Sp12to4
    port map (
            O => \N__21135\,
            I => \N__21132\
        );

    \I__2705\ : Span12Mux_v
    port map (
            O => \N__21132\,
            I => \N__21129\
        );

    \I__2704\ : Odrv12
    port map (
            O => \N__21129\,
            I => pin_in_8
        );

    \I__2703\ : InMux
    port map (
            O => \N__21126\,
            I => \N__21123\
        );

    \I__2702\ : LocalMux
    port map (
            O => \N__21123\,
            I => n13649
        );

    \I__2701\ : InMux
    port map (
            O => \N__21120\,
            I => \N__21116\
        );

    \I__2700\ : CascadeMux
    port map (
            O => \N__21119\,
            I => \N__21113\
        );

    \I__2699\ : LocalMux
    port map (
            O => \N__21116\,
            I => \N__21110\
        );

    \I__2698\ : InMux
    port map (
            O => \N__21113\,
            I => \N__21106\
        );

    \I__2697\ : Span12Mux_v
    port map (
            O => \N__21110\,
            I => \N__21103\
        );

    \I__2696\ : InMux
    port map (
            O => \N__21109\,
            I => \N__21100\
        );

    \I__2695\ : LocalMux
    port map (
            O => \N__21106\,
            I => \N__21097\
        );

    \I__2694\ : Odrv12
    port map (
            O => \N__21103\,
            I => timer_30
        );

    \I__2693\ : LocalMux
    port map (
            O => \N__21100\,
            I => timer_30
        );

    \I__2692\ : Odrv4
    port map (
            O => \N__21097\,
            I => timer_30
        );

    \I__2691\ : InMux
    port map (
            O => \N__21090\,
            I => \N__21086\
        );

    \I__2690\ : InMux
    port map (
            O => \N__21089\,
            I => \N__21083\
        );

    \I__2689\ : LocalMux
    port map (
            O => \N__21086\,
            I => neo_pixel_transmitter_t0_30
        );

    \I__2688\ : LocalMux
    port map (
            O => \N__21083\,
            I => neo_pixel_transmitter_t0_30
        );

    \I__2687\ : InMux
    port map (
            O => \N__21078\,
            I => \N__21075\
        );

    \I__2686\ : LocalMux
    port map (
            O => \N__21075\,
            I => \nx.n11946\
        );

    \I__2685\ : InMux
    port map (
            O => \N__21072\,
            I => \N__21069\
        );

    \I__2684\ : LocalMux
    port map (
            O => \N__21069\,
            I => \nx.n13445\
        );

    \I__2683\ : CascadeMux
    port map (
            O => \N__21066\,
            I => \nx.n11948_cascade_\
        );

    \I__2682\ : InMux
    port map (
            O => \N__21063\,
            I => \N__21060\
        );

    \I__2681\ : LocalMux
    port map (
            O => \N__21060\,
            I => \N__21057\
        );

    \I__2680\ : Span4Mux_v
    port map (
            O => \N__21057\,
            I => \N__21054\
        );

    \I__2679\ : Span4Mux_h
    port map (
            O => \N__21054\,
            I => \N__21051\
        );

    \I__2678\ : Odrv4
    port map (
            O => \N__21051\,
            I => pin_in_2
        );

    \I__2677\ : InMux
    port map (
            O => \N__21048\,
            I => \N__21045\
        );

    \I__2676\ : LocalMux
    port map (
            O => \N__21045\,
            I => \N__21042\
        );

    \I__2675\ : Span4Mux_v
    port map (
            O => \N__21042\,
            I => \N__21039\
        );

    \I__2674\ : Span4Mux_h
    port map (
            O => \N__21039\,
            I => \N__21036\
        );

    \I__2673\ : Odrv4
    port map (
            O => \N__21036\,
            I => pin_in_3
        );

    \I__2672\ : CascadeMux
    port map (
            O => \N__21033\,
            I => \n13379_cascade_\
        );

    \I__2671\ : InMux
    port map (
            O => \N__21030\,
            I => \N__21025\
        );

    \I__2670\ : InMux
    port map (
            O => \N__21029\,
            I => \N__21022\
        );

    \I__2669\ : InMux
    port map (
            O => \N__21028\,
            I => \N__21019\
        );

    \I__2668\ : LocalMux
    port map (
            O => \N__21025\,
            I => \nx.n1504\
        );

    \I__2667\ : LocalMux
    port map (
            O => \N__21022\,
            I => \nx.n1504\
        );

    \I__2666\ : LocalMux
    port map (
            O => \N__21019\,
            I => \nx.n1504\
        );

    \I__2665\ : InMux
    port map (
            O => \N__21012\,
            I => \nx.n10788\
        );

    \I__2664\ : InMux
    port map (
            O => \N__21009\,
            I => \N__21004\
        );

    \I__2663\ : InMux
    port map (
            O => \N__21008\,
            I => \N__21001\
        );

    \I__2662\ : InMux
    port map (
            O => \N__21007\,
            I => \N__20998\
        );

    \I__2661\ : LocalMux
    port map (
            O => \N__21004\,
            I => \nx.n1503\
        );

    \I__2660\ : LocalMux
    port map (
            O => \N__21001\,
            I => \nx.n1503\
        );

    \I__2659\ : LocalMux
    port map (
            O => \N__20998\,
            I => \nx.n1503\
        );

    \I__2658\ : InMux
    port map (
            O => \N__20991\,
            I => \nx.n10789\
        );

    \I__2657\ : InMux
    port map (
            O => \N__20988\,
            I => \N__20984\
        );

    \I__2656\ : InMux
    port map (
            O => \N__20987\,
            I => \N__20981\
        );

    \I__2655\ : LocalMux
    port map (
            O => \N__20984\,
            I => \N__20976\
        );

    \I__2654\ : LocalMux
    port map (
            O => \N__20981\,
            I => \N__20976\
        );

    \I__2653\ : Odrv4
    port map (
            O => \N__20976\,
            I => \nx.n1502\
        );

    \I__2652\ : InMux
    port map (
            O => \N__20973\,
            I => \bfn_4_27_0_\
        );

    \I__2651\ : InMux
    port map (
            O => \N__20970\,
            I => \N__20966\
        );

    \I__2650\ : InMux
    port map (
            O => \N__20969\,
            I => \N__20963\
        );

    \I__2649\ : LocalMux
    port map (
            O => \N__20966\,
            I => \N__20958\
        );

    \I__2648\ : LocalMux
    port map (
            O => \N__20963\,
            I => \N__20958\
        );

    \I__2647\ : Span4Mux_h
    port map (
            O => \N__20958\,
            I => \N__20954\
        );

    \I__2646\ : InMux
    port map (
            O => \N__20957\,
            I => \N__20951\
        );

    \I__2645\ : Odrv4
    port map (
            O => \N__20954\,
            I => \nx.n1501\
        );

    \I__2644\ : LocalMux
    port map (
            O => \N__20951\,
            I => \nx.n1501\
        );

    \I__2643\ : InMux
    port map (
            O => \N__20946\,
            I => \nx.n10791\
        );

    \I__2642\ : InMux
    port map (
            O => \N__20943\,
            I => \N__20938\
        );

    \I__2641\ : InMux
    port map (
            O => \N__20942\,
            I => \N__20935\
        );

    \I__2640\ : InMux
    port map (
            O => \N__20941\,
            I => \N__20932\
        );

    \I__2639\ : LocalMux
    port map (
            O => \N__20938\,
            I => \nx.n1500\
        );

    \I__2638\ : LocalMux
    port map (
            O => \N__20935\,
            I => \nx.n1500\
        );

    \I__2637\ : LocalMux
    port map (
            O => \N__20932\,
            I => \nx.n1500\
        );

    \I__2636\ : InMux
    port map (
            O => \N__20925\,
            I => \nx.n10792\
        );

    \I__2635\ : InMux
    port map (
            O => \N__20922\,
            I => \N__20918\
        );

    \I__2634\ : InMux
    port map (
            O => \N__20921\,
            I => \N__20915\
        );

    \I__2633\ : LocalMux
    port map (
            O => \N__20918\,
            I => \N__20910\
        );

    \I__2632\ : LocalMux
    port map (
            O => \N__20915\,
            I => \N__20910\
        );

    \I__2631\ : Span4Mux_h
    port map (
            O => \N__20910\,
            I => \N__20906\
        );

    \I__2630\ : InMux
    port map (
            O => \N__20909\,
            I => \N__20903\
        );

    \I__2629\ : Odrv4
    port map (
            O => \N__20906\,
            I => \nx.n1499\
        );

    \I__2628\ : LocalMux
    port map (
            O => \N__20903\,
            I => \nx.n1499\
        );

    \I__2627\ : CascadeMux
    port map (
            O => \N__20898\,
            I => \N__20886\
        );

    \I__2626\ : CascadeMux
    port map (
            O => \N__20897\,
            I => \N__20883\
        );

    \I__2625\ : CascadeMux
    port map (
            O => \N__20896\,
            I => \N__20880\
        );

    \I__2624\ : CascadeMux
    port map (
            O => \N__20895\,
            I => \N__20877\
        );

    \I__2623\ : CascadeMux
    port map (
            O => \N__20894\,
            I => \N__20874\
        );

    \I__2622\ : CascadeMux
    port map (
            O => \N__20893\,
            I => \N__20871\
        );

    \I__2621\ : CascadeMux
    port map (
            O => \N__20892\,
            I => \N__20868\
        );

    \I__2620\ : CascadeMux
    port map (
            O => \N__20891\,
            I => \N__20865\
        );

    \I__2619\ : CascadeMux
    port map (
            O => \N__20890\,
            I => \N__20862\
        );

    \I__2618\ : CascadeMux
    port map (
            O => \N__20889\,
            I => \N__20859\
        );

    \I__2617\ : InMux
    port map (
            O => \N__20886\,
            I => \N__20854\
        );

    \I__2616\ : InMux
    port map (
            O => \N__20883\,
            I => \N__20854\
        );

    \I__2615\ : InMux
    port map (
            O => \N__20880\,
            I => \N__20849\
        );

    \I__2614\ : InMux
    port map (
            O => \N__20877\,
            I => \N__20849\
        );

    \I__2613\ : InMux
    port map (
            O => \N__20874\,
            I => \N__20842\
        );

    \I__2612\ : InMux
    port map (
            O => \N__20871\,
            I => \N__20842\
        );

    \I__2611\ : InMux
    port map (
            O => \N__20868\,
            I => \N__20842\
        );

    \I__2610\ : InMux
    port map (
            O => \N__20865\,
            I => \N__20835\
        );

    \I__2609\ : InMux
    port map (
            O => \N__20862\,
            I => \N__20835\
        );

    \I__2608\ : InMux
    port map (
            O => \N__20859\,
            I => \N__20835\
        );

    \I__2607\ : LocalMux
    port map (
            O => \N__20854\,
            I => \nx.n1532\
        );

    \I__2606\ : LocalMux
    port map (
            O => \N__20849\,
            I => \nx.n1532\
        );

    \I__2605\ : LocalMux
    port map (
            O => \N__20842\,
            I => \nx.n1532\
        );

    \I__2604\ : LocalMux
    port map (
            O => \N__20835\,
            I => \nx.n1532\
        );

    \I__2603\ : InMux
    port map (
            O => \N__20826\,
            I => \nx.n10793\
        );

    \I__2602\ : InMux
    port map (
            O => \N__20823\,
            I => \N__20820\
        );

    \I__2601\ : LocalMux
    port map (
            O => \N__20820\,
            I => \nx.n45_adj_781\
        );

    \I__2600\ : InMux
    port map (
            O => \N__20817\,
            I => \N__20814\
        );

    \I__2599\ : LocalMux
    port map (
            O => \N__20814\,
            I => \N__20811\
        );

    \I__2598\ : Odrv4
    port map (
            O => \N__20811\,
            I => \nx.n19\
        );

    \I__2597\ : InMux
    port map (
            O => \N__20808\,
            I => \N__20805\
        );

    \I__2596\ : LocalMux
    port map (
            O => \N__20805\,
            I => \N__20802\
        );

    \I__2595\ : Odrv4
    port map (
            O => \N__20802\,
            I => \nx.n47_adj_780\
        );

    \I__2594\ : InMux
    port map (
            O => \N__20799\,
            I => \N__20796\
        );

    \I__2593\ : LocalMux
    port map (
            O => \N__20796\,
            I => \nx.n18\
        );

    \I__2592\ : InMux
    port map (
            O => \N__20793\,
            I => \N__20789\
        );

    \I__2591\ : InMux
    port map (
            O => \N__20792\,
            I => \N__20786\
        );

    \I__2590\ : LocalMux
    port map (
            O => \N__20789\,
            I => \N__20783\
        );

    \I__2589\ : LocalMux
    port map (
            O => \N__20786\,
            I => delay_counter_28
        );

    \I__2588\ : Odrv4
    port map (
            O => \N__20783\,
            I => delay_counter_28
        );

    \I__2587\ : InMux
    port map (
            O => \N__20778\,
            I => \N__20774\
        );

    \I__2586\ : InMux
    port map (
            O => \N__20777\,
            I => \N__20771\
        );

    \I__2585\ : LocalMux
    port map (
            O => \N__20774\,
            I => \N__20768\
        );

    \I__2584\ : LocalMux
    port map (
            O => \N__20771\,
            I => delay_counter_24
        );

    \I__2583\ : Odrv4
    port map (
            O => \N__20768\,
            I => delay_counter_24
        );

    \I__2582\ : CascadeMux
    port map (
            O => \N__20763\,
            I => \N__20760\
        );

    \I__2581\ : InMux
    port map (
            O => \N__20760\,
            I => \N__20757\
        );

    \I__2580\ : LocalMux
    port map (
            O => \N__20757\,
            I => \N__20753\
        );

    \I__2579\ : InMux
    port map (
            O => \N__20756\,
            I => \N__20750\
        );

    \I__2578\ : Span4Mux_h
    port map (
            O => \N__20753\,
            I => \N__20747\
        );

    \I__2577\ : LocalMux
    port map (
            O => \N__20750\,
            I => delay_counter_22
        );

    \I__2576\ : Odrv4
    port map (
            O => \N__20747\,
            I => delay_counter_22
        );

    \I__2575\ : InMux
    port map (
            O => \N__20742\,
            I => \N__20738\
        );

    \I__2574\ : InMux
    port map (
            O => \N__20741\,
            I => \N__20735\
        );

    \I__2573\ : LocalMux
    port map (
            O => \N__20738\,
            I => \N__20732\
        );

    \I__2572\ : LocalMux
    port map (
            O => \N__20735\,
            I => delay_counter_26
        );

    \I__2571\ : Odrv4
    port map (
            O => \N__20732\,
            I => delay_counter_26
        );

    \I__2570\ : InMux
    port map (
            O => \N__20727\,
            I => \bfn_4_26_0_\
        );

    \I__2569\ : InMux
    port map (
            O => \N__20724\,
            I => \N__20720\
        );

    \I__2568\ : InMux
    port map (
            O => \N__20723\,
            I => \N__20717\
        );

    \I__2567\ : LocalMux
    port map (
            O => \N__20720\,
            I => \nx.n1509\
        );

    \I__2566\ : LocalMux
    port map (
            O => \N__20717\,
            I => \nx.n1509\
        );

    \I__2565\ : CascadeMux
    port map (
            O => \N__20712\,
            I => \N__20708\
        );

    \I__2564\ : CascadeMux
    port map (
            O => \N__20711\,
            I => \N__20705\
        );

    \I__2563\ : InMux
    port map (
            O => \N__20708\,
            I => \N__20702\
        );

    \I__2562\ : InMux
    port map (
            O => \N__20705\,
            I => \N__20699\
        );

    \I__2561\ : LocalMux
    port map (
            O => \N__20702\,
            I => \nx.n13604\
        );

    \I__2560\ : LocalMux
    port map (
            O => \N__20699\,
            I => \nx.n13604\
        );

    \I__2559\ : InMux
    port map (
            O => \N__20694\,
            I => \nx.n10783\
        );

    \I__2558\ : InMux
    port map (
            O => \N__20691\,
            I => \N__20686\
        );

    \I__2557\ : InMux
    port map (
            O => \N__20690\,
            I => \N__20683\
        );

    \I__2556\ : InMux
    port map (
            O => \N__20689\,
            I => \N__20680\
        );

    \I__2555\ : LocalMux
    port map (
            O => \N__20686\,
            I => \nx.n1508\
        );

    \I__2554\ : LocalMux
    port map (
            O => \N__20683\,
            I => \nx.n1508\
        );

    \I__2553\ : LocalMux
    port map (
            O => \N__20680\,
            I => \nx.n1508\
        );

    \I__2552\ : InMux
    port map (
            O => \N__20673\,
            I => \nx.n10784\
        );

    \I__2551\ : InMux
    port map (
            O => \N__20670\,
            I => \N__20666\
        );

    \I__2550\ : InMux
    port map (
            O => \N__20669\,
            I => \N__20663\
        );

    \I__2549\ : LocalMux
    port map (
            O => \N__20666\,
            I => \nx.n1507\
        );

    \I__2548\ : LocalMux
    port map (
            O => \N__20663\,
            I => \nx.n1507\
        );

    \I__2547\ : InMux
    port map (
            O => \N__20658\,
            I => \nx.n10785\
        );

    \I__2546\ : InMux
    port map (
            O => \N__20655\,
            I => \N__20650\
        );

    \I__2545\ : InMux
    port map (
            O => \N__20654\,
            I => \N__20647\
        );

    \I__2544\ : InMux
    port map (
            O => \N__20653\,
            I => \N__20644\
        );

    \I__2543\ : LocalMux
    port map (
            O => \N__20650\,
            I => \nx.n1506\
        );

    \I__2542\ : LocalMux
    port map (
            O => \N__20647\,
            I => \nx.n1506\
        );

    \I__2541\ : LocalMux
    port map (
            O => \N__20644\,
            I => \nx.n1506\
        );

    \I__2540\ : InMux
    port map (
            O => \N__20637\,
            I => \nx.n10786\
        );

    \I__2539\ : InMux
    port map (
            O => \N__20634\,
            I => \N__20629\
        );

    \I__2538\ : InMux
    port map (
            O => \N__20633\,
            I => \N__20626\
        );

    \I__2537\ : InMux
    port map (
            O => \N__20632\,
            I => \N__20623\
        );

    \I__2536\ : LocalMux
    port map (
            O => \N__20629\,
            I => \nx.n1505\
        );

    \I__2535\ : LocalMux
    port map (
            O => \N__20626\,
            I => \nx.n1505\
        );

    \I__2534\ : LocalMux
    port map (
            O => \N__20623\,
            I => \nx.n1505\
        );

    \I__2533\ : InMux
    port map (
            O => \N__20616\,
            I => \nx.n10787\
        );

    \I__2532\ : InMux
    port map (
            O => \N__20613\,
            I => \N__20609\
        );

    \I__2531\ : InMux
    port map (
            O => \N__20612\,
            I => \N__20606\
        );

    \I__2530\ : LocalMux
    port map (
            O => \N__20609\,
            I => \N__20603\
        );

    \I__2529\ : LocalMux
    port map (
            O => \N__20606\,
            I => delay_counter_18
        );

    \I__2528\ : Odrv4
    port map (
            O => \N__20603\,
            I => delay_counter_18
        );

    \I__2527\ : InMux
    port map (
            O => \N__20598\,
            I => \N__20594\
        );

    \I__2526\ : InMux
    port map (
            O => \N__20597\,
            I => \N__20591\
        );

    \I__2525\ : LocalMux
    port map (
            O => \N__20594\,
            I => \N__20588\
        );

    \I__2524\ : LocalMux
    port map (
            O => \N__20591\,
            I => delay_counter_16
        );

    \I__2523\ : Odrv4
    port map (
            O => \N__20588\,
            I => delay_counter_16
        );

    \I__2522\ : InMux
    port map (
            O => \N__20583\,
            I => \N__20580\
        );

    \I__2521\ : LocalMux
    port map (
            O => \N__20580\,
            I => \N__20577\
        );

    \I__2520\ : Odrv4
    port map (
            O => \N__20577\,
            I => n6_adj_843
        );

    \I__2519\ : CascadeMux
    port map (
            O => \N__20574\,
            I => \N__20569\
        );

    \I__2518\ : InMux
    port map (
            O => \N__20573\,
            I => \N__20566\
        );

    \I__2517\ : InMux
    port map (
            O => \N__20572\,
            I => \N__20563\
        );

    \I__2516\ : InMux
    port map (
            O => \N__20569\,
            I => \N__20560\
        );

    \I__2515\ : LocalMux
    port map (
            O => \N__20566\,
            I => \N__20555\
        );

    \I__2514\ : LocalMux
    port map (
            O => \N__20563\,
            I => \N__20555\
        );

    \I__2513\ : LocalMux
    port map (
            O => \N__20560\,
            I => \nx.n1304\
        );

    \I__2512\ : Odrv4
    port map (
            O => \N__20555\,
            I => \nx.n1304\
        );

    \I__2511\ : CascadeMux
    port map (
            O => \N__20550\,
            I => \N__20546\
        );

    \I__2510\ : CascadeMux
    port map (
            O => \N__20549\,
            I => \N__20542\
        );

    \I__2509\ : InMux
    port map (
            O => \N__20546\,
            I => \N__20539\
        );

    \I__2508\ : InMux
    port map (
            O => \N__20545\,
            I => \N__20536\
        );

    \I__2507\ : InMux
    port map (
            O => \N__20542\,
            I => \N__20533\
        );

    \I__2506\ : LocalMux
    port map (
            O => \N__20539\,
            I => \N__20528\
        );

    \I__2505\ : LocalMux
    port map (
            O => \N__20536\,
            I => \N__20528\
        );

    \I__2504\ : LocalMux
    port map (
            O => \N__20533\,
            I => \nx.n1305\
        );

    \I__2503\ : Odrv4
    port map (
            O => \N__20528\,
            I => \nx.n1305\
        );

    \I__2502\ : CascadeMux
    port map (
            O => \N__20523\,
            I => \nx.n10_adj_668_cascade_\
        );

    \I__2501\ : CascadeMux
    port map (
            O => \N__20520\,
            I => \N__20515\
        );

    \I__2500\ : InMux
    port map (
            O => \N__20519\,
            I => \N__20512\
        );

    \I__2499\ : InMux
    port map (
            O => \N__20518\,
            I => \N__20509\
        );

    \I__2498\ : InMux
    port map (
            O => \N__20515\,
            I => \N__20506\
        );

    \I__2497\ : LocalMux
    port map (
            O => \N__20512\,
            I => \N__20501\
        );

    \I__2496\ : LocalMux
    port map (
            O => \N__20509\,
            I => \N__20501\
        );

    \I__2495\ : LocalMux
    port map (
            O => \N__20506\,
            I => \nx.n1307\
        );

    \I__2494\ : Odrv4
    port map (
            O => \N__20501\,
            I => \nx.n1307\
        );

    \I__2493\ : InMux
    port map (
            O => \N__20496\,
            I => \N__20493\
        );

    \I__2492\ : LocalMux
    port map (
            O => \N__20493\,
            I => \nx.n16\
        );

    \I__2491\ : CascadeMux
    port map (
            O => \N__20490\,
            I => \N__20487\
        );

    \I__2490\ : InMux
    port map (
            O => \N__20487\,
            I => \N__20484\
        );

    \I__2489\ : LocalMux
    port map (
            O => \N__20484\,
            I => \nx.n1369\
        );

    \I__2488\ : CascadeMux
    port map (
            O => \N__20481\,
            I => \N__20477\
        );

    \I__2487\ : CascadeMux
    port map (
            O => \N__20480\,
            I => \N__20471\
        );

    \I__2486\ : InMux
    port map (
            O => \N__20477\,
            I => \N__20462\
        );

    \I__2485\ : InMux
    port map (
            O => \N__20476\,
            I => \N__20462\
        );

    \I__2484\ : InMux
    port map (
            O => \N__20475\,
            I => \N__20453\
        );

    \I__2483\ : InMux
    port map (
            O => \N__20474\,
            I => \N__20453\
        );

    \I__2482\ : InMux
    port map (
            O => \N__20471\,
            I => \N__20453\
        );

    \I__2481\ : InMux
    port map (
            O => \N__20470\,
            I => \N__20453\
        );

    \I__2480\ : InMux
    port map (
            O => \N__20469\,
            I => \N__20448\
        );

    \I__2479\ : InMux
    port map (
            O => \N__20468\,
            I => \N__20448\
        );

    \I__2478\ : InMux
    port map (
            O => \N__20467\,
            I => \N__20445\
        );

    \I__2477\ : LocalMux
    port map (
            O => \N__20462\,
            I => \nx.n1334\
        );

    \I__2476\ : LocalMux
    port map (
            O => \N__20453\,
            I => \nx.n1334\
        );

    \I__2475\ : LocalMux
    port map (
            O => \N__20448\,
            I => \nx.n1334\
        );

    \I__2474\ : LocalMux
    port map (
            O => \N__20445\,
            I => \nx.n1334\
        );

    \I__2473\ : CascadeMux
    port map (
            O => \N__20436\,
            I => \N__20433\
        );

    \I__2472\ : InMux
    port map (
            O => \N__20433\,
            I => \N__20429\
        );

    \I__2471\ : InMux
    port map (
            O => \N__20432\,
            I => \N__20426\
        );

    \I__2470\ : LocalMux
    port map (
            O => \N__20429\,
            I => \N__20423\
        );

    \I__2469\ : LocalMux
    port map (
            O => \N__20426\,
            I => \N__20419\
        );

    \I__2468\ : Span4Mux_s3_h
    port map (
            O => \N__20423\,
            I => \N__20416\
        );

    \I__2467\ : InMux
    port map (
            O => \N__20422\,
            I => \N__20413\
        );

    \I__2466\ : Odrv4
    port map (
            O => \N__20419\,
            I => \nx.n1401\
        );

    \I__2465\ : Odrv4
    port map (
            O => \N__20416\,
            I => \nx.n1401\
        );

    \I__2464\ : LocalMux
    port map (
            O => \N__20413\,
            I => \nx.n1401\
        );

    \I__2463\ : SRMux
    port map (
            O => \N__20406\,
            I => \N__20403\
        );

    \I__2462\ : LocalMux
    port map (
            O => \N__20403\,
            I => \N__20400\
        );

    \I__2461\ : Sp12to4
    port map (
            O => \N__20400\,
            I => \N__20397\
        );

    \I__2460\ : Odrv12
    port map (
            O => \N__20397\,
            I => n22_adj_795
        );

    \I__2459\ : CascadeMux
    port map (
            O => \N__20394\,
            I => \nx.n1631_cascade_\
        );

    \I__2458\ : CascadeMux
    port map (
            O => \N__20391\,
            I => \nx.n15_adj_676_cascade_\
        );

    \I__2457\ : InMux
    port map (
            O => \N__20388\,
            I => \N__20385\
        );

    \I__2456\ : LocalMux
    port map (
            O => \N__20385\,
            I => \nx.n22\
        );

    \I__2455\ : CascadeMux
    port map (
            O => \N__20382\,
            I => \N__20378\
        );

    \I__2454\ : InMux
    port map (
            O => \N__20381\,
            I => \N__20375\
        );

    \I__2453\ : InMux
    port map (
            O => \N__20378\,
            I => \N__20372\
        );

    \I__2452\ : LocalMux
    port map (
            O => \N__20375\,
            I => \nx.n1308\
        );

    \I__2451\ : LocalMux
    port map (
            O => \N__20372\,
            I => \nx.n1308\
        );

    \I__2450\ : InMux
    port map (
            O => \N__20367\,
            I => \N__20364\
        );

    \I__2449\ : LocalMux
    port map (
            O => \N__20364\,
            I => \N__20361\
        );

    \I__2448\ : Span4Mux_s3_h
    port map (
            O => \N__20361\,
            I => \N__20358\
        );

    \I__2447\ : Odrv4
    port map (
            O => \N__20358\,
            I => \nx.n1375\
        );

    \I__2446\ : InMux
    port map (
            O => \N__20355\,
            I => \nx.n10765\
        );

    \I__2445\ : InMux
    port map (
            O => \N__20352\,
            I => \N__20349\
        );

    \I__2444\ : LocalMux
    port map (
            O => \N__20349\,
            I => \nx.n1374\
        );

    \I__2443\ : InMux
    port map (
            O => \N__20346\,
            I => \nx.n10766\
        );

    \I__2442\ : CascadeMux
    port map (
            O => \N__20343\,
            I => \N__20338\
        );

    \I__2441\ : InMux
    port map (
            O => \N__20342\,
            I => \N__20333\
        );

    \I__2440\ : InMux
    port map (
            O => \N__20341\,
            I => \N__20333\
        );

    \I__2439\ : InMux
    port map (
            O => \N__20338\,
            I => \N__20330\
        );

    \I__2438\ : LocalMux
    port map (
            O => \N__20333\,
            I => \nx.n1306\
        );

    \I__2437\ : LocalMux
    port map (
            O => \N__20330\,
            I => \nx.n1306\
        );

    \I__2436\ : CascadeMux
    port map (
            O => \N__20325\,
            I => \N__20322\
        );

    \I__2435\ : InMux
    port map (
            O => \N__20322\,
            I => \N__20319\
        );

    \I__2434\ : LocalMux
    port map (
            O => \N__20319\,
            I => \nx.n1373\
        );

    \I__2433\ : InMux
    port map (
            O => \N__20316\,
            I => \nx.n10767\
        );

    \I__2432\ : InMux
    port map (
            O => \N__20313\,
            I => \N__20310\
        );

    \I__2431\ : LocalMux
    port map (
            O => \N__20310\,
            I => \nx.n1372\
        );

    \I__2430\ : InMux
    port map (
            O => \N__20307\,
            I => \nx.n10768\
        );

    \I__2429\ : CascadeMux
    port map (
            O => \N__20304\,
            I => \N__20301\
        );

    \I__2428\ : InMux
    port map (
            O => \N__20301\,
            I => \N__20298\
        );

    \I__2427\ : LocalMux
    port map (
            O => \N__20298\,
            I => \nx.n1371\
        );

    \I__2426\ : InMux
    port map (
            O => \N__20295\,
            I => \nx.n10769\
        );

    \I__2425\ : CascadeMux
    port map (
            O => \N__20292\,
            I => \N__20287\
        );

    \I__2424\ : InMux
    port map (
            O => \N__20291\,
            I => \N__20282\
        );

    \I__2423\ : InMux
    port map (
            O => \N__20290\,
            I => \N__20282\
        );

    \I__2422\ : InMux
    port map (
            O => \N__20287\,
            I => \N__20279\
        );

    \I__2421\ : LocalMux
    port map (
            O => \N__20282\,
            I => \nx.n1303\
        );

    \I__2420\ : LocalMux
    port map (
            O => \N__20279\,
            I => \nx.n1303\
        );

    \I__2419\ : InMux
    port map (
            O => \N__20274\,
            I => \N__20271\
        );

    \I__2418\ : LocalMux
    port map (
            O => \N__20271\,
            I => \nx.n1370\
        );

    \I__2417\ : InMux
    port map (
            O => \N__20268\,
            I => \nx.n10770\
        );

    \I__2416\ : InMux
    port map (
            O => \N__20265\,
            I => \bfn_4_24_0_\
        );

    \I__2415\ : InMux
    port map (
            O => \N__20262\,
            I => \nx.n10772\
        );

    \I__2414\ : InMux
    port map (
            O => \N__20259\,
            I => \N__20256\
        );

    \I__2413\ : LocalMux
    port map (
            O => \N__20256\,
            I => \N__20253\
        );

    \I__2412\ : Span4Mux_s3_h
    port map (
            O => \N__20253\,
            I => \N__20249\
        );

    \I__2411\ : InMux
    port map (
            O => \N__20252\,
            I => \N__20246\
        );

    \I__2410\ : Odrv4
    port map (
            O => \N__20249\,
            I => \nx.n1400\
        );

    \I__2409\ : LocalMux
    port map (
            O => \N__20246\,
            I => \nx.n1400\
        );

    \I__2408\ : CascadeMux
    port map (
            O => \N__20241\,
            I => \nx.n1235_cascade_\
        );

    \I__2407\ : CascadeMux
    port map (
            O => \N__20238\,
            I => \nx.n1203_cascade_\
        );

    \I__2406\ : CascadeMux
    port map (
            O => \N__20235\,
            I => \N__20232\
        );

    \I__2405\ : InMux
    port map (
            O => \N__20232\,
            I => \N__20229\
        );

    \I__2404\ : LocalMux
    port map (
            O => \N__20229\,
            I => \nx.n13_adj_675\
        );

    \I__2403\ : InMux
    port map (
            O => \N__20226\,
            I => \N__20223\
        );

    \I__2402\ : LocalMux
    port map (
            O => \N__20223\,
            I => \N__20220\
        );

    \I__2401\ : Span4Mux_s3_h
    port map (
            O => \N__20220\,
            I => \N__20217\
        );

    \I__2400\ : Odrv4
    port map (
            O => \N__20217\,
            I => \nx.n1377\
        );

    \I__2399\ : InMux
    port map (
            O => \N__20214\,
            I => \bfn_4_23_0_\
        );

    \I__2398\ : CascadeMux
    port map (
            O => \N__20211\,
            I => \N__20207\
        );

    \I__2397\ : InMux
    port map (
            O => \N__20210\,
            I => \N__20204\
        );

    \I__2396\ : InMux
    port map (
            O => \N__20207\,
            I => \N__20201\
        );

    \I__2395\ : LocalMux
    port map (
            O => \N__20204\,
            I => \nx.n1309\
        );

    \I__2394\ : LocalMux
    port map (
            O => \N__20201\,
            I => \nx.n1309\
        );

    \I__2393\ : CascadeMux
    port map (
            O => \N__20196\,
            I => \N__20193\
        );

    \I__2392\ : InMux
    port map (
            O => \N__20193\,
            I => \N__20190\
        );

    \I__2391\ : LocalMux
    port map (
            O => \N__20190\,
            I => \nx.n1376\
        );

    \I__2390\ : InMux
    port map (
            O => \N__20187\,
            I => \nx.n10764\
        );

    \I__2389\ : CascadeMux
    port map (
            O => \N__20184\,
            I => \N__20181\
        );

    \I__2388\ : InMux
    port map (
            O => \N__20181\,
            I => \N__20178\
        );

    \I__2387\ : LocalMux
    port map (
            O => \N__20178\,
            I => \N__20173\
        );

    \I__2386\ : InMux
    port map (
            O => \N__20177\,
            I => \N__20170\
        );

    \I__2385\ : InMux
    port map (
            O => \N__20176\,
            I => \N__20167\
        );

    \I__2384\ : Span4Mux_v
    port map (
            O => \N__20173\,
            I => \N__20164\
        );

    \I__2383\ : LocalMux
    port map (
            O => \N__20170\,
            I => timer_29
        );

    \I__2382\ : LocalMux
    port map (
            O => \N__20167\,
            I => timer_29
        );

    \I__2381\ : Odrv4
    port map (
            O => \N__20164\,
            I => timer_29
        );

    \I__2380\ : InMux
    port map (
            O => \N__20157\,
            I => \N__20154\
        );

    \I__2379\ : LocalMux
    port map (
            O => \N__20154\,
            I => \N__20150\
        );

    \I__2378\ : InMux
    port map (
            O => \N__20153\,
            I => \N__20147\
        );

    \I__2377\ : Span4Mux_h
    port map (
            O => \N__20150\,
            I => \N__20144\
        );

    \I__2376\ : LocalMux
    port map (
            O => \N__20147\,
            I => neo_pixel_transmitter_t0_29
        );

    \I__2375\ : Odrv4
    port map (
            O => \N__20144\,
            I => neo_pixel_transmitter_t0_29
        );

    \I__2374\ : InMux
    port map (
            O => \N__20139\,
            I => \N__20135\
        );

    \I__2373\ : InMux
    port map (
            O => \N__20138\,
            I => \N__20132\
        );

    \I__2372\ : LocalMux
    port map (
            O => \N__20135\,
            I => neo_pixel_transmitter_t0_25
        );

    \I__2371\ : LocalMux
    port map (
            O => \N__20132\,
            I => neo_pixel_transmitter_t0_25
        );

    \I__2370\ : CascadeMux
    port map (
            O => \N__20127\,
            I => \N__20124\
        );

    \I__2369\ : InMux
    port map (
            O => \N__20124\,
            I => \N__20121\
        );

    \I__2368\ : LocalMux
    port map (
            O => \N__20121\,
            I => \N__20118\
        );

    \I__2367\ : Span4Mux_s3_h
    port map (
            O => \N__20118\,
            I => \N__20115\
        );

    \I__2366\ : Odrv4
    port map (
            O => \N__20115\,
            I => \nx.n8\
        );

    \I__2365\ : CascadeMux
    port map (
            O => \N__20112\,
            I => \nx.n1205_cascade_\
        );

    \I__2364\ : InMux
    port map (
            O => \N__20109\,
            I => \N__20106\
        );

    \I__2363\ : LocalMux
    port map (
            O => \N__20106\,
            I => \nx.n11_adj_674\
        );

    \I__2362\ : CascadeMux
    port map (
            O => \N__20103\,
            I => \nx.n6_adj_786_cascade_\
        );

    \I__2361\ : InMux
    port map (
            O => \N__20100\,
            I => \N__20096\
        );

    \I__2360\ : InMux
    port map (
            O => \N__20099\,
            I => \N__20093\
        );

    \I__2359\ : LocalMux
    port map (
            O => \N__20096\,
            I => \N__20090\
        );

    \I__2358\ : LocalMux
    port map (
            O => \N__20093\,
            I => \N__20087\
        );

    \I__2357\ : Span4Mux_h
    port map (
            O => \N__20090\,
            I => \N__20084\
        );

    \I__2356\ : Odrv4
    port map (
            O => \N__20087\,
            I => \nx.one_wire_N_599_5\
        );

    \I__2355\ : Odrv4
    port map (
            O => \N__20084\,
            I => \nx.one_wire_N_599_5\
        );

    \I__2354\ : CEMux
    port map (
            O => \N__20079\,
            I => \N__20076\
        );

    \I__2353\ : LocalMux
    port map (
            O => \N__20076\,
            I => \N__20073\
        );

    \I__2352\ : Span4Mux_v
    port map (
            O => \N__20073\,
            I => \N__20070\
        );

    \I__2351\ : Odrv4
    port map (
            O => \N__20070\,
            I => \nx.n13659\
        );

    \I__2350\ : InMux
    port map (
            O => \N__20067\,
            I => \N__20064\
        );

    \I__2349\ : LocalMux
    port map (
            O => \N__20064\,
            I => \N__20060\
        );

    \I__2348\ : InMux
    port map (
            O => \N__20063\,
            I => \N__20057\
        );

    \I__2347\ : Span4Mux_v
    port map (
            O => \N__20060\,
            I => \N__20052\
        );

    \I__2346\ : LocalMux
    port map (
            O => \N__20057\,
            I => \N__20052\
        );

    \I__2345\ : Odrv4
    port map (
            O => \N__20052\,
            I => \nx.one_wire_N_599_7\
        );

    \I__2344\ : InMux
    port map (
            O => \N__20049\,
            I => \N__20040\
        );

    \I__2343\ : InMux
    port map (
            O => \N__20048\,
            I => \N__20040\
        );

    \I__2342\ : InMux
    port map (
            O => \N__20047\,
            I => \N__20040\
        );

    \I__2341\ : LocalMux
    port map (
            O => \N__20040\,
            I => \N__20037\
        );

    \I__2340\ : Span4Mux_v
    port map (
            O => \N__20037\,
            I => \N__20034\
        );

    \I__2339\ : Odrv4
    port map (
            O => \N__20034\,
            I => \nx.one_wire_N_599_8\
        );

    \I__2338\ : CascadeMux
    port map (
            O => \N__20031\,
            I => \N__20027\
        );

    \I__2337\ : InMux
    port map (
            O => \N__20030\,
            I => \N__20022\
        );

    \I__2336\ : InMux
    port map (
            O => \N__20027\,
            I => \N__20022\
        );

    \I__2335\ : LocalMux
    port map (
            O => \N__20022\,
            I => \N__20019\
        );

    \I__2334\ : Odrv4
    port map (
            O => \N__20019\,
            I => \nx.one_wire_N_599_6\
        );

    \I__2333\ : InMux
    port map (
            O => \N__20016\,
            I => \N__20013\
        );

    \I__2332\ : LocalMux
    port map (
            O => \N__20013\,
            I => \nx.n13211\
        );

    \I__2331\ : CascadeMux
    port map (
            O => \N__20010\,
            I => \N__20006\
        );

    \I__2330\ : InMux
    port map (
            O => \N__20009\,
            I => \N__19998\
        );

    \I__2329\ : InMux
    port map (
            O => \N__20006\,
            I => \N__19998\
        );

    \I__2328\ : InMux
    port map (
            O => \N__20005\,
            I => \N__19998\
        );

    \I__2327\ : LocalMux
    port map (
            O => \N__19998\,
            I => \N__19995\
        );

    \I__2326\ : Span4Mux_h
    port map (
            O => \N__19995\,
            I => \N__19992\
        );

    \I__2325\ : Odrv4
    port map (
            O => \N__19992\,
            I => \nx.one_wire_N_599_10\
        );

    \I__2324\ : InMux
    port map (
            O => \N__19989\,
            I => \N__19984\
        );

    \I__2323\ : InMux
    port map (
            O => \N__19988\,
            I => \N__19979\
        );

    \I__2322\ : InMux
    port map (
            O => \N__19987\,
            I => \N__19979\
        );

    \I__2321\ : LocalMux
    port map (
            O => \N__19984\,
            I => \N__19976\
        );

    \I__2320\ : LocalMux
    port map (
            O => \N__19979\,
            I => \N__19973\
        );

    \I__2319\ : Span4Mux_v
    port map (
            O => \N__19976\,
            I => \N__19968\
        );

    \I__2318\ : Span4Mux_v
    port map (
            O => \N__19973\,
            I => \N__19968\
        );

    \I__2317\ : Odrv4
    port map (
            O => \N__19968\,
            I => \nx.one_wire_N_599_9\
        );

    \I__2316\ : CascadeMux
    port map (
            O => \N__19965\,
            I => \nx.n13217_cascade_\
        );

    \I__2315\ : InMux
    port map (
            O => \N__19962\,
            I => \N__19953\
        );

    \I__2314\ : InMux
    port map (
            O => \N__19961\,
            I => \N__19953\
        );

    \I__2313\ : InMux
    port map (
            O => \N__19960\,
            I => \N__19953\
        );

    \I__2312\ : LocalMux
    port map (
            O => \N__19953\,
            I => \N__19950\
        );

    \I__2311\ : Span4Mux_h
    port map (
            O => \N__19950\,
            I => \N__19947\
        );

    \I__2310\ : Odrv4
    port map (
            O => \N__19947\,
            I => \nx.n7608\
        );

    \I__2309\ : InMux
    port map (
            O => \N__19944\,
            I => \N__19941\
        );

    \I__2308\ : LocalMux
    port map (
            O => \N__19941\,
            I => \N__19938\
        );

    \I__2307\ : Span4Mux_s3_h
    port map (
            O => \N__19938\,
            I => \N__19935\
        );

    \I__2306\ : Odrv4
    port map (
            O => \N__19935\,
            I => \nx.n20_adj_726\
        );

    \I__2305\ : CascadeMux
    port map (
            O => \N__19932\,
            I => \N__19929\
        );

    \I__2304\ : InMux
    port map (
            O => \N__19929\,
            I => \N__19924\
        );

    \I__2303\ : InMux
    port map (
            O => \N__19928\,
            I => \N__19921\
        );

    \I__2302\ : InMux
    port map (
            O => \N__19927\,
            I => \N__19918\
        );

    \I__2301\ : LocalMux
    port map (
            O => \N__19924\,
            I => \N__19915\
        );

    \I__2300\ : LocalMux
    port map (
            O => \N__19921\,
            I => timer_13
        );

    \I__2299\ : LocalMux
    port map (
            O => \N__19918\,
            I => timer_13
        );

    \I__2298\ : Odrv4
    port map (
            O => \N__19915\,
            I => timer_13
        );

    \I__2297\ : InMux
    port map (
            O => \N__19908\,
            I => \N__19902\
        );

    \I__2296\ : InMux
    port map (
            O => \N__19907\,
            I => \N__19902\
        );

    \I__2295\ : LocalMux
    port map (
            O => \N__19902\,
            I => neo_pixel_transmitter_t0_13
        );

    \I__2294\ : InMux
    port map (
            O => \N__19899\,
            I => \N__19894\
        );

    \I__2293\ : InMux
    port map (
            O => \N__19898\,
            I => \N__19891\
        );

    \I__2292\ : InMux
    port map (
            O => \N__19897\,
            I => \N__19888\
        );

    \I__2291\ : LocalMux
    port map (
            O => \N__19894\,
            I => timer_25
        );

    \I__2290\ : LocalMux
    port map (
            O => \N__19891\,
            I => timer_25
        );

    \I__2289\ : LocalMux
    port map (
            O => \N__19888\,
            I => timer_25
        );

    \I__2288\ : CascadeMux
    port map (
            O => \N__19881\,
            I => \N__19876\
        );

    \I__2287\ : InMux
    port map (
            O => \N__19880\,
            I => \N__19873\
        );

    \I__2286\ : InMux
    port map (
            O => \N__19879\,
            I => \N__19870\
        );

    \I__2285\ : InMux
    port map (
            O => \N__19876\,
            I => \N__19867\
        );

    \I__2284\ : LocalMux
    port map (
            O => \N__19873\,
            I => timer_19
        );

    \I__2283\ : LocalMux
    port map (
            O => \N__19870\,
            I => timer_19
        );

    \I__2282\ : LocalMux
    port map (
            O => \N__19867\,
            I => timer_19
        );

    \I__2281\ : InMux
    port map (
            O => \N__19860\,
            I => \N__19857\
        );

    \I__2280\ : LocalMux
    port map (
            O => \N__19857\,
            I => \N__19854\
        );

    \I__2279\ : Span4Mux_h
    port map (
            O => \N__19854\,
            I => \N__19851\
        );

    \I__2278\ : Span4Mux_v
    port map (
            O => \N__19851\,
            I => \N__19848\
        );

    \I__2277\ : Span4Mux_v
    port map (
            O => \N__19848\,
            I => \N__19845\
        );

    \I__2276\ : Odrv4
    port map (
            O => \N__19845\,
            I => pin_in_7
        );

    \I__2275\ : InMux
    port map (
            O => \N__19842\,
            I => \N__19839\
        );

    \I__2274\ : LocalMux
    port map (
            O => \N__19839\,
            I => \N__19836\
        );

    \I__2273\ : Span12Mux_v
    port map (
            O => \N__19836\,
            I => \N__19833\
        );

    \I__2272\ : Odrv12
    port map (
            O => \N__19833\,
            I => pin_in_6
        );

    \I__2271\ : InMux
    port map (
            O => \N__19830\,
            I => \N__19827\
        );

    \I__2270\ : LocalMux
    port map (
            O => \N__19827\,
            I => \nx.n103\
        );

    \I__2269\ : CascadeMux
    port map (
            O => \N__19824\,
            I => \N__19821\
        );

    \I__2268\ : InMux
    port map (
            O => \N__19821\,
            I => \N__19818\
        );

    \I__2267\ : LocalMux
    port map (
            O => \N__19818\,
            I => \nx.n11892\
        );

    \I__2266\ : InMux
    port map (
            O => \N__19815\,
            I => \N__19812\
        );

    \I__2265\ : LocalMux
    port map (
            O => \N__19812\,
            I => \N__19809\
        );

    \I__2264\ : Span4Mux_s3_h
    port map (
            O => \N__19809\,
            I => \N__19806\
        );

    \I__2263\ : Odrv4
    port map (
            O => \N__19806\,
            I => \nx.n30_adj_712\
        );

    \I__2262\ : InMux
    port map (
            O => \N__19803\,
            I => \N__19800\
        );

    \I__2261\ : LocalMux
    port map (
            O => \N__19800\,
            I => \N__19797\
        );

    \I__2260\ : Span4Mux_s3_h
    port map (
            O => \N__19797\,
            I => \N__19794\
        );

    \I__2259\ : Odrv4
    port map (
            O => \N__19794\,
            I => \nx.n32\
        );

    \I__2258\ : CascadeMux
    port map (
            O => \N__19791\,
            I => \N__19788\
        );

    \I__2257\ : InMux
    port map (
            O => \N__19788\,
            I => \N__19785\
        );

    \I__2256\ : LocalMux
    port map (
            O => \N__19785\,
            I => \N__19782\
        );

    \I__2255\ : Span4Mux_v
    port map (
            O => \N__19782\,
            I => \N__19779\
        );

    \I__2254\ : Sp12to4
    port map (
            O => \N__19779\,
            I => \N__19776\
        );

    \I__2253\ : Odrv12
    port map (
            O => \N__19776\,
            I => \nx.n28_adj_715\
        );

    \I__2252\ : InMux
    port map (
            O => \N__19773\,
            I => \N__19768\
        );

    \I__2251\ : InMux
    port map (
            O => \N__19772\,
            I => \N__19765\
        );

    \I__2250\ : InMux
    port map (
            O => \N__19771\,
            I => \N__19762\
        );

    \I__2249\ : LocalMux
    port map (
            O => \N__19768\,
            I => timer_5
        );

    \I__2248\ : LocalMux
    port map (
            O => \N__19765\,
            I => timer_5
        );

    \I__2247\ : LocalMux
    port map (
            O => \N__19762\,
            I => timer_5
        );

    \I__2246\ : CascadeMux
    port map (
            O => \N__19755\,
            I => \N__19752\
        );

    \I__2245\ : InMux
    port map (
            O => \N__19752\,
            I => \N__19746\
        );

    \I__2244\ : InMux
    port map (
            O => \N__19751\,
            I => \N__19746\
        );

    \I__2243\ : LocalMux
    port map (
            O => \N__19746\,
            I => neo_pixel_transmitter_t0_5
        );

    \I__2242\ : CascadeMux
    port map (
            O => \N__19743\,
            I => \N__19738\
        );

    \I__2241\ : InMux
    port map (
            O => \N__19742\,
            I => \N__19735\
        );

    \I__2240\ : InMux
    port map (
            O => \N__19741\,
            I => \N__19732\
        );

    \I__2239\ : InMux
    port map (
            O => \N__19738\,
            I => \N__19729\
        );

    \I__2238\ : LocalMux
    port map (
            O => \N__19735\,
            I => timer_1
        );

    \I__2237\ : LocalMux
    port map (
            O => \N__19732\,
            I => timer_1
        );

    \I__2236\ : LocalMux
    port map (
            O => \N__19729\,
            I => timer_1
        );

    \I__2235\ : CascadeMux
    port map (
            O => \N__19722\,
            I => \N__19719\
        );

    \I__2234\ : InMux
    port map (
            O => \N__19719\,
            I => \N__19713\
        );

    \I__2233\ : InMux
    port map (
            O => \N__19718\,
            I => \N__19713\
        );

    \I__2232\ : LocalMux
    port map (
            O => \N__19713\,
            I => neo_pixel_transmitter_t0_1
        );

    \I__2231\ : CascadeMux
    port map (
            O => \N__19710\,
            I => \N__19705\
        );

    \I__2230\ : InMux
    port map (
            O => \N__19709\,
            I => \N__19702\
        );

    \I__2229\ : InMux
    port map (
            O => \N__19708\,
            I => \N__19699\
        );

    \I__2228\ : InMux
    port map (
            O => \N__19705\,
            I => \N__19696\
        );

    \I__2227\ : LocalMux
    port map (
            O => \N__19702\,
            I => timer_3
        );

    \I__2226\ : LocalMux
    port map (
            O => \N__19699\,
            I => timer_3
        );

    \I__2225\ : LocalMux
    port map (
            O => \N__19696\,
            I => timer_3
        );

    \I__2224\ : InMux
    port map (
            O => \N__19689\,
            I => \N__19685\
        );

    \I__2223\ : InMux
    port map (
            O => \N__19688\,
            I => \N__19682\
        );

    \I__2222\ : LocalMux
    port map (
            O => \N__19685\,
            I => neo_pixel_transmitter_t0_3
        );

    \I__2221\ : LocalMux
    port map (
            O => \N__19682\,
            I => neo_pixel_transmitter_t0_3
        );

    \I__2220\ : InMux
    port map (
            O => \N__19677\,
            I => \N__19674\
        );

    \I__2219\ : LocalMux
    port map (
            O => \N__19674\,
            I => \nx.n16_adj_785\
        );

    \I__2218\ : CascadeMux
    port map (
            O => \N__19671\,
            I => \N__19667\
        );

    \I__2217\ : InMux
    port map (
            O => \N__19670\,
            I => \N__19664\
        );

    \I__2216\ : InMux
    port map (
            O => \N__19667\,
            I => \N__19661\
        );

    \I__2215\ : LocalMux
    port map (
            O => \N__19664\,
            I => \N__19658\
        );

    \I__2214\ : LocalMux
    port map (
            O => \N__19661\,
            I => \N__19655\
        );

    \I__2213\ : Span4Mux_h
    port map (
            O => \N__19658\,
            I => \N__19652\
        );

    \I__2212\ : Odrv4
    port map (
            O => \N__19655\,
            I => \nx.one_wire_N_599_4\
        );

    \I__2211\ : Odrv4
    port map (
            O => \N__19652\,
            I => \nx.one_wire_N_599_4\
        );

    \I__2210\ : InMux
    port map (
            O => \N__19647\,
            I => \N__19644\
        );

    \I__2209\ : LocalMux
    port map (
            O => \N__19644\,
            I => \nx.n46_adj_779\
        );

    \I__2208\ : InMux
    port map (
            O => \N__19641\,
            I => \N__19638\
        );

    \I__2207\ : LocalMux
    port map (
            O => \N__19638\,
            I => \N__19635\
        );

    \I__2206\ : Span4Mux_v
    port map (
            O => \N__19635\,
            I => \N__19632\
        );

    \I__2205\ : Span4Mux_v
    port map (
            O => \N__19632\,
            I => \N__19629\
        );

    \I__2204\ : Odrv4
    port map (
            O => \N__19629\,
            I => \nx.n3\
        );

    \I__2203\ : CascadeMux
    port map (
            O => \N__19626\,
            I => \nx.n7_adj_764_cascade_\
        );

    \I__2202\ : CascadeMux
    port map (
            O => \N__19623\,
            I => \nx.n11864_cascade_\
        );

    \I__2201\ : CEMux
    port map (
            O => \N__19620\,
            I => \N__19617\
        );

    \I__2200\ : LocalMux
    port map (
            O => \N__19617\,
            I => \nx.n7_adj_667\
        );

    \I__2199\ : InMux
    port map (
            O => \N__19614\,
            I => \N__19611\
        );

    \I__2198\ : LocalMux
    port map (
            O => \N__19611\,
            I => \nx.n1476\
        );

    \I__2197\ : CascadeMux
    port map (
            O => \N__19608\,
            I => \N__19604\
        );

    \I__2196\ : InMux
    port map (
            O => \N__19607\,
            I => \N__19600\
        );

    \I__2195\ : InMux
    port map (
            O => \N__19604\,
            I => \N__19597\
        );

    \I__2194\ : InMux
    port map (
            O => \N__19603\,
            I => \N__19594\
        );

    \I__2193\ : LocalMux
    port map (
            O => \N__19600\,
            I => \nx.n1409\
        );

    \I__2192\ : LocalMux
    port map (
            O => \N__19597\,
            I => \nx.n1409\
        );

    \I__2191\ : LocalMux
    port map (
            O => \N__19594\,
            I => \nx.n1409\
        );

    \I__2190\ : CascadeMux
    port map (
            O => \N__19587\,
            I => \N__19584\
        );

    \I__2189\ : InMux
    port map (
            O => \N__19584\,
            I => \N__19581\
        );

    \I__2188\ : LocalMux
    port map (
            O => \N__19581\,
            I => \nx.n1468\
        );

    \I__2187\ : InMux
    port map (
            O => \N__19578\,
            I => \N__19575\
        );

    \I__2186\ : LocalMux
    port map (
            O => \N__19575\,
            I => \nx.n1475\
        );

    \I__2185\ : InMux
    port map (
            O => \N__19572\,
            I => \N__19568\
        );

    \I__2184\ : CascadeMux
    port map (
            O => \N__19571\,
            I => \N__19565\
        );

    \I__2183\ : LocalMux
    port map (
            O => \N__19568\,
            I => \N__19561\
        );

    \I__2182\ : InMux
    port map (
            O => \N__19565\,
            I => \N__19558\
        );

    \I__2181\ : InMux
    port map (
            O => \N__19564\,
            I => \N__19555\
        );

    \I__2180\ : Odrv4
    port map (
            O => \N__19561\,
            I => \nx.n1408\
        );

    \I__2179\ : LocalMux
    port map (
            O => \N__19558\,
            I => \nx.n1408\
        );

    \I__2178\ : LocalMux
    port map (
            O => \N__19555\,
            I => \nx.n1408\
        );

    \I__2177\ : CascadeMux
    port map (
            O => \N__19548\,
            I => \nx.n1507_cascade_\
        );

    \I__2176\ : CascadeMux
    port map (
            O => \N__19545\,
            I => \nx.n18_adj_731_cascade_\
        );

    \I__2175\ : CascadeMux
    port map (
            O => \N__19542\,
            I => \nx.n20_adj_733_cascade_\
        );

    \I__2174\ : InMux
    port map (
            O => \N__19539\,
            I => \N__19536\
        );

    \I__2173\ : LocalMux
    port map (
            O => \N__19536\,
            I => \nx.n16_adj_732\
        );

    \I__2172\ : CascadeMux
    port map (
            O => \N__19533\,
            I => \nx.n1532_cascade_\
        );

    \I__2171\ : InMux
    port map (
            O => \N__19530\,
            I => \N__19527\
        );

    \I__2170\ : LocalMux
    port map (
            O => \N__19527\,
            I => \N__19524\
        );

    \I__2169\ : Odrv4
    port map (
            O => \N__19524\,
            I => \nx.n1477\
        );

    \I__2168\ : CascadeMux
    port map (
            O => \N__19521\,
            I => \N__19515\
        );

    \I__2167\ : CascadeMux
    port map (
            O => \N__19520\,
            I => \N__19510\
        );

    \I__2166\ : CascadeMux
    port map (
            O => \N__19519\,
            I => \N__19506\
        );

    \I__2165\ : CascadeMux
    port map (
            O => \N__19518\,
            I => \N__19502\
        );

    \I__2164\ : InMux
    port map (
            O => \N__19515\,
            I => \N__19495\
        );

    \I__2163\ : InMux
    port map (
            O => \N__19514\,
            I => \N__19495\
        );

    \I__2162\ : InMux
    port map (
            O => \N__19513\,
            I => \N__19484\
        );

    \I__2161\ : InMux
    port map (
            O => \N__19510\,
            I => \N__19484\
        );

    \I__2160\ : InMux
    port map (
            O => \N__19509\,
            I => \N__19484\
        );

    \I__2159\ : InMux
    port map (
            O => \N__19506\,
            I => \N__19484\
        );

    \I__2158\ : InMux
    port map (
            O => \N__19505\,
            I => \N__19484\
        );

    \I__2157\ : InMux
    port map (
            O => \N__19502\,
            I => \N__19477\
        );

    \I__2156\ : InMux
    port map (
            O => \N__19501\,
            I => \N__19477\
        );

    \I__2155\ : InMux
    port map (
            O => \N__19500\,
            I => \N__19477\
        );

    \I__2154\ : LocalMux
    port map (
            O => \N__19495\,
            I => \nx.n1433\
        );

    \I__2153\ : LocalMux
    port map (
            O => \N__19484\,
            I => \nx.n1433\
        );

    \I__2152\ : LocalMux
    port map (
            O => \N__19477\,
            I => \nx.n1433\
        );

    \I__2151\ : CascadeMux
    port map (
            O => \N__19470\,
            I => \nx.n1509_cascade_\
        );

    \I__2150\ : InMux
    port map (
            O => \N__19467\,
            I => \N__19464\
        );

    \I__2149\ : LocalMux
    port map (
            O => \N__19464\,
            I => \nx.n9729\
        );

    \I__2148\ : CascadeMux
    port map (
            O => \N__19461\,
            I => \nx.n16_adj_727_cascade_\
        );

    \I__2147\ : CascadeMux
    port map (
            O => \N__19458\,
            I => \N__19455\
        );

    \I__2146\ : InMux
    port map (
            O => \N__19455\,
            I => \N__19452\
        );

    \I__2145\ : LocalMux
    port map (
            O => \N__19452\,
            I => \nx.n1471\
        );

    \I__2144\ : InMux
    port map (
            O => \N__19449\,
            I => \N__19446\
        );

    \I__2143\ : LocalMux
    port map (
            O => \N__19446\,
            I => \nx.n1473\
        );

    \I__2142\ : CascadeMux
    port map (
            O => \N__19443\,
            I => \N__19439\
        );

    \I__2141\ : InMux
    port map (
            O => \N__19442\,
            I => \N__19435\
        );

    \I__2140\ : InMux
    port map (
            O => \N__19439\,
            I => \N__19432\
        );

    \I__2139\ : InMux
    port map (
            O => \N__19438\,
            I => \N__19429\
        );

    \I__2138\ : LocalMux
    port map (
            O => \N__19435\,
            I => \nx.n1406\
        );

    \I__2137\ : LocalMux
    port map (
            O => \N__19432\,
            I => \nx.n1406\
        );

    \I__2136\ : LocalMux
    port map (
            O => \N__19429\,
            I => \nx.n1406\
        );

    \I__2135\ : CascadeMux
    port map (
            O => \N__19422\,
            I => \N__19419\
        );

    \I__2134\ : InMux
    port map (
            O => \N__19419\,
            I => \N__19414\
        );

    \I__2133\ : InMux
    port map (
            O => \N__19418\,
            I => \N__19409\
        );

    \I__2132\ : InMux
    port map (
            O => \N__19417\,
            I => \N__19409\
        );

    \I__2131\ : LocalMux
    port map (
            O => \N__19414\,
            I => \nx.n1404\
        );

    \I__2130\ : LocalMux
    port map (
            O => \N__19409\,
            I => \nx.n1404\
        );

    \I__2129\ : CascadeMux
    port map (
            O => \N__19404\,
            I => \N__19401\
        );

    \I__2128\ : InMux
    port map (
            O => \N__19401\,
            I => \N__19398\
        );

    \I__2127\ : LocalMux
    port map (
            O => \N__19398\,
            I => \nx.n13_adj_729\
        );

    \I__2126\ : InMux
    port map (
            O => \N__19395\,
            I => \N__19392\
        );

    \I__2125\ : LocalMux
    port map (
            O => \N__19392\,
            I => \nx.n18_adj_728\
        );

    \I__2124\ : InMux
    port map (
            O => \N__19389\,
            I => \N__19384\
        );

    \I__2123\ : InMux
    port map (
            O => \N__19388\,
            I => \N__19381\
        );

    \I__2122\ : CascadeMux
    port map (
            O => \N__19387\,
            I => \N__19378\
        );

    \I__2121\ : LocalMux
    port map (
            O => \N__19384\,
            I => \N__19373\
        );

    \I__2120\ : LocalMux
    port map (
            O => \N__19381\,
            I => \N__19373\
        );

    \I__2119\ : InMux
    port map (
            O => \N__19378\,
            I => \N__19370\
        );

    \I__2118\ : Odrv4
    port map (
            O => \N__19373\,
            I => \nx.n1405\
        );

    \I__2117\ : LocalMux
    port map (
            O => \N__19370\,
            I => \nx.n1405\
        );

    \I__2116\ : CascadeMux
    port map (
            O => \N__19365\,
            I => \nx.n1433_cascade_\
        );

    \I__2115\ : InMux
    port map (
            O => \N__19362\,
            I => \N__19359\
        );

    \I__2114\ : LocalMux
    port map (
            O => \N__19359\,
            I => \nx.n1472\
        );

    \I__2113\ : InMux
    port map (
            O => \N__19356\,
            I => \N__19353\
        );

    \I__2112\ : LocalMux
    port map (
            O => \N__19353\,
            I => \nx.n1470\
        );

    \I__2111\ : CascadeMux
    port map (
            O => \N__19350\,
            I => \N__19346\
        );

    \I__2110\ : CascadeMux
    port map (
            O => \N__19349\,
            I => \N__19343\
        );

    \I__2109\ : InMux
    port map (
            O => \N__19346\,
            I => \N__19340\
        );

    \I__2108\ : InMux
    port map (
            O => \N__19343\,
            I => \N__19337\
        );

    \I__2107\ : LocalMux
    port map (
            O => \N__19340\,
            I => \nx.n1403\
        );

    \I__2106\ : LocalMux
    port map (
            O => \N__19337\,
            I => \nx.n1403\
        );

    \I__2105\ : CascadeMux
    port map (
            O => \N__19332\,
            I => \nx.n1502_cascade_\
        );

    \I__2104\ : InMux
    port map (
            O => \N__19329\,
            I => \N__19326\
        );

    \I__2103\ : LocalMux
    port map (
            O => \N__19326\,
            I => \nx.n1474\
        );

    \I__2102\ : CascadeMux
    port map (
            O => \N__19323\,
            I => \N__19319\
        );

    \I__2101\ : CascadeMux
    port map (
            O => \N__19322\,
            I => \N__19315\
        );

    \I__2100\ : InMux
    port map (
            O => \N__19319\,
            I => \N__19310\
        );

    \I__2099\ : InMux
    port map (
            O => \N__19318\,
            I => \N__19310\
        );

    \I__2098\ : InMux
    port map (
            O => \N__19315\,
            I => \N__19307\
        );

    \I__2097\ : LocalMux
    port map (
            O => \N__19310\,
            I => \nx.n1407\
        );

    \I__2096\ : LocalMux
    port map (
            O => \N__19307\,
            I => \nx.n1407\
        );

    \I__2095\ : InMux
    port map (
            O => \N__19302\,
            I => \N__19299\
        );

    \I__2094\ : LocalMux
    port map (
            O => \N__19299\,
            I => \N__19295\
        );

    \I__2093\ : InMux
    port map (
            O => \N__19298\,
            I => \N__19292\
        );

    \I__2092\ : Span4Mux_h
    port map (
            O => \N__19295\,
            I => \N__19289\
        );

    \I__2091\ : LocalMux
    port map (
            O => \N__19292\,
            I => delay_counter_21
        );

    \I__2090\ : Odrv4
    port map (
            O => \N__19289\,
            I => delay_counter_21
        );

    \I__2089\ : CascadeMux
    port map (
            O => \N__19284\,
            I => \N__19281\
        );

    \I__2088\ : InMux
    port map (
            O => \N__19281\,
            I => \N__19278\
        );

    \I__2087\ : LocalMux
    port map (
            O => \N__19278\,
            I => \N__19274\
        );

    \I__2086\ : InMux
    port map (
            O => \N__19277\,
            I => \N__19271\
        );

    \I__2085\ : Span4Mux_h
    port map (
            O => \N__19274\,
            I => \N__19268\
        );

    \I__2084\ : LocalMux
    port map (
            O => \N__19271\,
            I => delay_counter_29
        );

    \I__2083\ : Odrv4
    port map (
            O => \N__19268\,
            I => delay_counter_29
        );

    \I__2082\ : InMux
    port map (
            O => \N__19263\,
            I => \N__19260\
        );

    \I__2081\ : LocalMux
    port map (
            O => \N__19260\,
            I => n12379
        );

    \I__2080\ : InMux
    port map (
            O => \N__19257\,
            I => \N__19254\
        );

    \I__2079\ : LocalMux
    port map (
            O => \N__19254\,
            I => \nx.n12_adj_669\
        );

    \I__2078\ : CascadeMux
    port map (
            O => \N__19251\,
            I => \nx.n1308_cascade_\
        );

    \I__2077\ : CascadeMux
    port map (
            O => \N__19248\,
            I => \nx.n1334_cascade_\
        );

    \I__2076\ : CascadeMux
    port map (
            O => \N__19245\,
            I => \nx.n1403_cascade_\
        );

    \I__2075\ : CascadeMux
    port map (
            O => \N__19242\,
            I => \N__19239\
        );

    \I__2074\ : InMux
    port map (
            O => \N__19239\,
            I => \N__19233\
        );

    \I__2073\ : InMux
    port map (
            O => \N__19238\,
            I => \N__19233\
        );

    \I__2072\ : LocalMux
    port map (
            O => \N__19233\,
            I => \N__19229\
        );

    \I__2071\ : InMux
    port map (
            O => \N__19232\,
            I => \N__19226\
        );

    \I__2070\ : Odrv4
    port map (
            O => \N__19229\,
            I => \nx.n1402\
        );

    \I__2069\ : LocalMux
    port map (
            O => \N__19226\,
            I => \nx.n1402\
        );

    \I__2068\ : InMux
    port map (
            O => \N__19221\,
            I => \N__19218\
        );

    \I__2067\ : LocalMux
    port map (
            O => \N__19218\,
            I => \N__19214\
        );

    \I__2066\ : InMux
    port map (
            O => \N__19217\,
            I => \N__19211\
        );

    \I__2065\ : Span4Mux_h
    port map (
            O => \N__19214\,
            I => \N__19208\
        );

    \I__2064\ : LocalMux
    port map (
            O => \N__19211\,
            I => delay_counter_17
        );

    \I__2063\ : Odrv4
    port map (
            O => \N__19208\,
            I => delay_counter_17
        );

    \I__2062\ : CascadeMux
    port map (
            O => \N__19203\,
            I => \N__19200\
        );

    \I__2061\ : InMux
    port map (
            O => \N__19200\,
            I => \N__19197\
        );

    \I__2060\ : LocalMux
    port map (
            O => \N__19197\,
            I => \N__19193\
        );

    \I__2059\ : InMux
    port map (
            O => \N__19196\,
            I => \N__19190\
        );

    \I__2058\ : Span4Mux_h
    port map (
            O => \N__19193\,
            I => \N__19187\
        );

    \I__2057\ : LocalMux
    port map (
            O => \N__19190\,
            I => delay_counter_15
        );

    \I__2056\ : Odrv4
    port map (
            O => \N__19187\,
            I => delay_counter_15
        );

    \I__2055\ : InMux
    port map (
            O => \N__19182\,
            I => \N__19179\
        );

    \I__2054\ : LocalMux
    port map (
            O => \N__19179\,
            I => \N__19176\
        );

    \I__2053\ : Span4Mux_h
    port map (
            O => \N__19176\,
            I => \N__19173\
        );

    \I__2052\ : Odrv4
    port map (
            O => \N__19173\,
            I => n12382
        );

    \I__2051\ : CascadeMux
    port map (
            O => \N__19170\,
            I => \n11828_cascade_\
        );

    \I__2050\ : IoInMux
    port map (
            O => \N__19167\,
            I => \N__19164\
        );

    \I__2049\ : LocalMux
    port map (
            O => \N__19164\,
            I => \N__19161\
        );

    \I__2048\ : Span4Mux_s0_h
    port map (
            O => \N__19161\,
            I => \N__19158\
        );

    \I__2047\ : Span4Mux_v
    port map (
            O => \N__19158\,
            I => \N__19155\
        );

    \I__2046\ : Span4Mux_v
    port map (
            O => \N__19155\,
            I => \N__19151\
        );

    \I__2045\ : InMux
    port map (
            O => \N__19154\,
            I => \N__19148\
        );

    \I__2044\ : Odrv4
    port map (
            O => \N__19151\,
            I => pin_oe_5
        );

    \I__2043\ : LocalMux
    port map (
            O => \N__19148\,
            I => pin_oe_5
        );

    \I__2042\ : InMux
    port map (
            O => \N__19143\,
            I => \N__19140\
        );

    \I__2041\ : LocalMux
    port map (
            O => \N__19140\,
            I => \N__19135\
        );

    \I__2040\ : InMux
    port map (
            O => \N__19139\,
            I => \N__19132\
        );

    \I__2039\ : InMux
    port map (
            O => \N__19138\,
            I => \N__19129\
        );

    \I__2038\ : Odrv4
    port map (
            O => \N__19135\,
            I => timer_16
        );

    \I__2037\ : LocalMux
    port map (
            O => \N__19132\,
            I => timer_16
        );

    \I__2036\ : LocalMux
    port map (
            O => \N__19129\,
            I => timer_16
        );

    \I__2035\ : InMux
    port map (
            O => \N__19122\,
            I => \N__19118\
        );

    \I__2034\ : InMux
    port map (
            O => \N__19121\,
            I => \N__19115\
        );

    \I__2033\ : LocalMux
    port map (
            O => \N__19118\,
            I => neo_pixel_transmitter_t0_16
        );

    \I__2032\ : LocalMux
    port map (
            O => \N__19115\,
            I => neo_pixel_transmitter_t0_16
        );

    \I__2031\ : CascadeMux
    port map (
            O => \N__19110\,
            I => \N__19107\
        );

    \I__2030\ : InMux
    port map (
            O => \N__19107\,
            I => \N__19104\
        );

    \I__2029\ : LocalMux
    port map (
            O => \N__19104\,
            I => \N__19101\
        );

    \I__2028\ : Odrv4
    port map (
            O => \N__19101\,
            I => \nx.n17\
        );

    \I__2027\ : CascadeMux
    port map (
            O => \N__19098\,
            I => \nx.n1309_cascade_\
        );

    \I__2026\ : InMux
    port map (
            O => \N__19095\,
            I => \nx.n10731\
        );

    \I__2025\ : InMux
    port map (
            O => \N__19092\,
            I => \nx.n10732\
        );

    \I__2024\ : CascadeMux
    port map (
            O => \N__19089\,
            I => \N__19085\
        );

    \I__2023\ : InMux
    port map (
            O => \N__19088\,
            I => \N__19081\
        );

    \I__2022\ : InMux
    port map (
            O => \N__19085\,
            I => \N__19078\
        );

    \I__2021\ : InMux
    port map (
            O => \N__19084\,
            I => \N__19075\
        );

    \I__2020\ : LocalMux
    port map (
            O => \N__19081\,
            I => \N__19070\
        );

    \I__2019\ : LocalMux
    port map (
            O => \N__19078\,
            I => \N__19070\
        );

    \I__2018\ : LocalMux
    port map (
            O => \N__19075\,
            I => \N__19065\
        );

    \I__2017\ : Span4Mux_v
    port map (
            O => \N__19070\,
            I => \N__19065\
        );

    \I__2016\ : Odrv4
    port map (
            O => \N__19065\,
            I => timer_27
        );

    \I__2015\ : InMux
    port map (
            O => \N__19062\,
            I => \nx.n10733\
        );

    \I__2014\ : InMux
    port map (
            O => \N__19059\,
            I => \nx.n10734\
        );

    \I__2013\ : InMux
    port map (
            O => \N__19056\,
            I => \nx.n10735\
        );

    \I__2012\ : InMux
    port map (
            O => \N__19053\,
            I => \nx.n10736\
        );

    \I__2011\ : InMux
    port map (
            O => \N__19050\,
            I => \nx.n10737\
        );

    \I__2010\ : InMux
    port map (
            O => \N__19047\,
            I => \N__19042\
        );

    \I__2009\ : InMux
    port map (
            O => \N__19046\,
            I => \N__19039\
        );

    \I__2008\ : InMux
    port map (
            O => \N__19045\,
            I => \N__19036\
        );

    \I__2007\ : LocalMux
    port map (
            O => \N__19042\,
            I => \N__19033\
        );

    \I__2006\ : LocalMux
    port map (
            O => \N__19039\,
            I => \N__19030\
        );

    \I__2005\ : LocalMux
    port map (
            O => \N__19036\,
            I => timer_31
        );

    \I__2004\ : Odrv12
    port map (
            O => \N__19033\,
            I => timer_31
        );

    \I__2003\ : Odrv4
    port map (
            O => \N__19030\,
            I => timer_31
        );

    \I__2002\ : CascadeMux
    port map (
            O => \N__19023\,
            I => \n11826_cascade_\
        );

    \I__2001\ : IoInMux
    port map (
            O => \N__19020\,
            I => \N__19017\
        );

    \I__2000\ : LocalMux
    port map (
            O => \N__19017\,
            I => \N__19014\
        );

    \I__1999\ : Span4Mux_s2_v
    port map (
            O => \N__19014\,
            I => \N__19011\
        );

    \I__1998\ : Span4Mux_v
    port map (
            O => \N__19011\,
            I => \N__19008\
        );

    \I__1997\ : Span4Mux_v
    port map (
            O => \N__19008\,
            I => \N__19004\
        );

    \I__1996\ : InMux
    port map (
            O => \N__19007\,
            I => \N__19001\
        );

    \I__1995\ : Odrv4
    port map (
            O => \N__19004\,
            I => pin_oe_1
        );

    \I__1994\ : LocalMux
    port map (
            O => \N__19001\,
            I => pin_oe_1
        );

    \I__1993\ : InMux
    port map (
            O => \N__18996\,
            I => \bfn_3_20_0_\
        );

    \I__1992\ : InMux
    port map (
            O => \N__18993\,
            I => \N__18989\
        );

    \I__1991\ : CascadeMux
    port map (
            O => \N__18992\,
            I => \N__18985\
        );

    \I__1990\ : LocalMux
    port map (
            O => \N__18989\,
            I => \N__18982\
        );

    \I__1989\ : InMux
    port map (
            O => \N__18988\,
            I => \N__18979\
        );

    \I__1988\ : InMux
    port map (
            O => \N__18985\,
            I => \N__18976\
        );

    \I__1987\ : Odrv4
    port map (
            O => \N__18982\,
            I => timer_17
        );

    \I__1986\ : LocalMux
    port map (
            O => \N__18979\,
            I => timer_17
        );

    \I__1985\ : LocalMux
    port map (
            O => \N__18976\,
            I => timer_17
        );

    \I__1984\ : InMux
    port map (
            O => \N__18969\,
            I => \nx.n10723\
        );

    \I__1983\ : InMux
    port map (
            O => \N__18966\,
            I => \N__18962\
        );

    \I__1982\ : CascadeMux
    port map (
            O => \N__18965\,
            I => \N__18959\
        );

    \I__1981\ : LocalMux
    port map (
            O => \N__18962\,
            I => \N__18955\
        );

    \I__1980\ : InMux
    port map (
            O => \N__18959\,
            I => \N__18952\
        );

    \I__1979\ : InMux
    port map (
            O => \N__18958\,
            I => \N__18949\
        );

    \I__1978\ : Span4Mux_s2_h
    port map (
            O => \N__18955\,
            I => \N__18944\
        );

    \I__1977\ : LocalMux
    port map (
            O => \N__18952\,
            I => \N__18944\
        );

    \I__1976\ : LocalMux
    port map (
            O => \N__18949\,
            I => timer_18
        );

    \I__1975\ : Odrv4
    port map (
            O => \N__18944\,
            I => timer_18
        );

    \I__1974\ : InMux
    port map (
            O => \N__18939\,
            I => \nx.n10724\
        );

    \I__1973\ : InMux
    port map (
            O => \N__18936\,
            I => \nx.n10725\
        );

    \I__1972\ : InMux
    port map (
            O => \N__18933\,
            I => \N__18930\
        );

    \I__1971\ : LocalMux
    port map (
            O => \N__18930\,
            I => \N__18927\
        );

    \I__1970\ : Span4Mux_s2_h
    port map (
            O => \N__18927\,
            I => \N__18922\
        );

    \I__1969\ : InMux
    port map (
            O => \N__18926\,
            I => \N__18919\
        );

    \I__1968\ : InMux
    port map (
            O => \N__18925\,
            I => \N__18916\
        );

    \I__1967\ : Odrv4
    port map (
            O => \N__18922\,
            I => timer_20
        );

    \I__1966\ : LocalMux
    port map (
            O => \N__18919\,
            I => timer_20
        );

    \I__1965\ : LocalMux
    port map (
            O => \N__18916\,
            I => timer_20
        );

    \I__1964\ : InMux
    port map (
            O => \N__18909\,
            I => \nx.n10726\
        );

    \I__1963\ : InMux
    port map (
            O => \N__18906\,
            I => \N__18903\
        );

    \I__1962\ : LocalMux
    port map (
            O => \N__18903\,
            I => \N__18899\
        );

    \I__1961\ : InMux
    port map (
            O => \N__18902\,
            I => \N__18895\
        );

    \I__1960\ : Span4Mux_v
    port map (
            O => \N__18899\,
            I => \N__18892\
        );

    \I__1959\ : InMux
    port map (
            O => \N__18898\,
            I => \N__18889\
        );

    \I__1958\ : LocalMux
    port map (
            O => \N__18895\,
            I => \N__18886\
        );

    \I__1957\ : Odrv4
    port map (
            O => \N__18892\,
            I => timer_21
        );

    \I__1956\ : LocalMux
    port map (
            O => \N__18889\,
            I => timer_21
        );

    \I__1955\ : Odrv4
    port map (
            O => \N__18886\,
            I => timer_21
        );

    \I__1954\ : InMux
    port map (
            O => \N__18879\,
            I => \nx.n10727\
        );

    \I__1953\ : InMux
    port map (
            O => \N__18876\,
            I => \N__18872\
        );

    \I__1952\ : CascadeMux
    port map (
            O => \N__18875\,
            I => \N__18869\
        );

    \I__1951\ : LocalMux
    port map (
            O => \N__18872\,
            I => \N__18865\
        );

    \I__1950\ : InMux
    port map (
            O => \N__18869\,
            I => \N__18862\
        );

    \I__1949\ : InMux
    port map (
            O => \N__18868\,
            I => \N__18859\
        );

    \I__1948\ : Span4Mux_v
    port map (
            O => \N__18865\,
            I => \N__18854\
        );

    \I__1947\ : LocalMux
    port map (
            O => \N__18862\,
            I => \N__18854\
        );

    \I__1946\ : LocalMux
    port map (
            O => \N__18859\,
            I => timer_22
        );

    \I__1945\ : Odrv4
    port map (
            O => \N__18854\,
            I => timer_22
        );

    \I__1944\ : InMux
    port map (
            O => \N__18849\,
            I => \nx.n10728\
        );

    \I__1943\ : InMux
    port map (
            O => \N__18846\,
            I => \N__18843\
        );

    \I__1942\ : LocalMux
    port map (
            O => \N__18843\,
            I => \N__18838\
        );

    \I__1941\ : InMux
    port map (
            O => \N__18842\,
            I => \N__18835\
        );

    \I__1940\ : InMux
    port map (
            O => \N__18841\,
            I => \N__18832\
        );

    \I__1939\ : Span4Mux_v
    port map (
            O => \N__18838\,
            I => \N__18827\
        );

    \I__1938\ : LocalMux
    port map (
            O => \N__18835\,
            I => \N__18827\
        );

    \I__1937\ : LocalMux
    port map (
            O => \N__18832\,
            I => timer_23
        );

    \I__1936\ : Odrv4
    port map (
            O => \N__18827\,
            I => timer_23
        );

    \I__1935\ : InMux
    port map (
            O => \N__18822\,
            I => \nx.n10729\
        );

    \I__1934\ : InMux
    port map (
            O => \N__18819\,
            I => \N__18815\
        );

    \I__1933\ : CascadeMux
    port map (
            O => \N__18818\,
            I => \N__18811\
        );

    \I__1932\ : LocalMux
    port map (
            O => \N__18815\,
            I => \N__18808\
        );

    \I__1931\ : InMux
    port map (
            O => \N__18814\,
            I => \N__18805\
        );

    \I__1930\ : InMux
    port map (
            O => \N__18811\,
            I => \N__18802\
        );

    \I__1929\ : Odrv4
    port map (
            O => \N__18808\,
            I => timer_24
        );

    \I__1928\ : LocalMux
    port map (
            O => \N__18805\,
            I => timer_24
        );

    \I__1927\ : LocalMux
    port map (
            O => \N__18802\,
            I => timer_24
        );

    \I__1926\ : InMux
    port map (
            O => \N__18795\,
            I => \bfn_3_21_0_\
        );

    \I__1925\ : InMux
    port map (
            O => \N__18792\,
            I => \N__18789\
        );

    \I__1924\ : LocalMux
    port map (
            O => \N__18789\,
            I => \N__18784\
        );

    \I__1923\ : InMux
    port map (
            O => \N__18788\,
            I => \N__18781\
        );

    \I__1922\ : InMux
    port map (
            O => \N__18787\,
            I => \N__18778\
        );

    \I__1921\ : Odrv4
    port map (
            O => \N__18784\,
            I => timer_8
        );

    \I__1920\ : LocalMux
    port map (
            O => \N__18781\,
            I => timer_8
        );

    \I__1919\ : LocalMux
    port map (
            O => \N__18778\,
            I => timer_8
        );

    \I__1918\ : InMux
    port map (
            O => \N__18771\,
            I => \bfn_3_19_0_\
        );

    \I__1917\ : InMux
    port map (
            O => \N__18768\,
            I => \N__18765\
        );

    \I__1916\ : LocalMux
    port map (
            O => \N__18765\,
            I => \N__18760\
        );

    \I__1915\ : InMux
    port map (
            O => \N__18764\,
            I => \N__18757\
        );

    \I__1914\ : InMux
    port map (
            O => \N__18763\,
            I => \N__18754\
        );

    \I__1913\ : Odrv4
    port map (
            O => \N__18760\,
            I => timer_9
        );

    \I__1912\ : LocalMux
    port map (
            O => \N__18757\,
            I => timer_9
        );

    \I__1911\ : LocalMux
    port map (
            O => \N__18754\,
            I => timer_9
        );

    \I__1910\ : InMux
    port map (
            O => \N__18747\,
            I => \nx.n10715\
        );

    \I__1909\ : InMux
    port map (
            O => \N__18744\,
            I => \N__18740\
        );

    \I__1908\ : CascadeMux
    port map (
            O => \N__18743\,
            I => \N__18736\
        );

    \I__1907\ : LocalMux
    port map (
            O => \N__18740\,
            I => \N__18733\
        );

    \I__1906\ : InMux
    port map (
            O => \N__18739\,
            I => \N__18730\
        );

    \I__1905\ : InMux
    port map (
            O => \N__18736\,
            I => \N__18727\
        );

    \I__1904\ : Odrv4
    port map (
            O => \N__18733\,
            I => timer_10
        );

    \I__1903\ : LocalMux
    port map (
            O => \N__18730\,
            I => timer_10
        );

    \I__1902\ : LocalMux
    port map (
            O => \N__18727\,
            I => timer_10
        );

    \I__1901\ : InMux
    port map (
            O => \N__18720\,
            I => \nx.n10716\
        );

    \I__1900\ : InMux
    port map (
            O => \N__18717\,
            I => \nx.n10717\
        );

    \I__1899\ : InMux
    port map (
            O => \N__18714\,
            I => \N__18711\
        );

    \I__1898\ : LocalMux
    port map (
            O => \N__18711\,
            I => \N__18707\
        );

    \I__1897\ : CascadeMux
    port map (
            O => \N__18710\,
            I => \N__18703\
        );

    \I__1896\ : Span4Mux_s2_h
    port map (
            O => \N__18707\,
            I => \N__18700\
        );

    \I__1895\ : InMux
    port map (
            O => \N__18706\,
            I => \N__18697\
        );

    \I__1894\ : InMux
    port map (
            O => \N__18703\,
            I => \N__18694\
        );

    \I__1893\ : Odrv4
    port map (
            O => \N__18700\,
            I => timer_12
        );

    \I__1892\ : LocalMux
    port map (
            O => \N__18697\,
            I => timer_12
        );

    \I__1891\ : LocalMux
    port map (
            O => \N__18694\,
            I => timer_12
        );

    \I__1890\ : InMux
    port map (
            O => \N__18687\,
            I => \nx.n10718\
        );

    \I__1889\ : InMux
    port map (
            O => \N__18684\,
            I => \nx.n10719\
        );

    \I__1888\ : InMux
    port map (
            O => \N__18681\,
            I => \N__18677\
        );

    \I__1887\ : CascadeMux
    port map (
            O => \N__18680\,
            I => \N__18673\
        );

    \I__1886\ : LocalMux
    port map (
            O => \N__18677\,
            I => \N__18670\
        );

    \I__1885\ : InMux
    port map (
            O => \N__18676\,
            I => \N__18667\
        );

    \I__1884\ : InMux
    port map (
            O => \N__18673\,
            I => \N__18664\
        );

    \I__1883\ : Odrv12
    port map (
            O => \N__18670\,
            I => timer_14
        );

    \I__1882\ : LocalMux
    port map (
            O => \N__18667\,
            I => timer_14
        );

    \I__1881\ : LocalMux
    port map (
            O => \N__18664\,
            I => timer_14
        );

    \I__1880\ : InMux
    port map (
            O => \N__18657\,
            I => \nx.n10720\
        );

    \I__1879\ : InMux
    port map (
            O => \N__18654\,
            I => \N__18651\
        );

    \I__1878\ : LocalMux
    port map (
            O => \N__18651\,
            I => \N__18646\
        );

    \I__1877\ : InMux
    port map (
            O => \N__18650\,
            I => \N__18643\
        );

    \I__1876\ : InMux
    port map (
            O => \N__18649\,
            I => \N__18640\
        );

    \I__1875\ : Span4Mux_v
    port map (
            O => \N__18646\,
            I => \N__18635\
        );

    \I__1874\ : LocalMux
    port map (
            O => \N__18643\,
            I => \N__18635\
        );

    \I__1873\ : LocalMux
    port map (
            O => \N__18640\,
            I => timer_15
        );

    \I__1872\ : Odrv4
    port map (
            O => \N__18635\,
            I => timer_15
        );

    \I__1871\ : InMux
    port map (
            O => \N__18630\,
            I => \nx.n10721\
        );

    \I__1870\ : CascadeMux
    port map (
            O => \N__18627\,
            I => \nx.n11834_cascade_\
        );

    \I__1869\ : InMux
    port map (
            O => \N__18624\,
            I => \N__18621\
        );

    \I__1868\ : LocalMux
    port map (
            O => \N__18621\,
            I => \N__18617\
        );

    \I__1867\ : CascadeMux
    port map (
            O => \N__18620\,
            I => \N__18613\
        );

    \I__1866\ : Span4Mux_v
    port map (
            O => \N__18617\,
            I => \N__18610\
        );

    \I__1865\ : InMux
    port map (
            O => \N__18616\,
            I => \N__18607\
        );

    \I__1864\ : InMux
    port map (
            O => \N__18613\,
            I => \N__18604\
        );

    \I__1863\ : Odrv4
    port map (
            O => \N__18610\,
            I => timer_0
        );

    \I__1862\ : LocalMux
    port map (
            O => \N__18607\,
            I => timer_0
        );

    \I__1861\ : LocalMux
    port map (
            O => \N__18604\,
            I => timer_0
        );

    \I__1860\ : InMux
    port map (
            O => \N__18597\,
            I => \bfn_3_18_0_\
        );

    \I__1859\ : InMux
    port map (
            O => \N__18594\,
            I => \nx.n10707\
        );

    \I__1858\ : CascadeMux
    port map (
            O => \N__18591\,
            I => \N__18586\
        );

    \I__1857\ : InMux
    port map (
            O => \N__18590\,
            I => \N__18583\
        );

    \I__1856\ : InMux
    port map (
            O => \N__18589\,
            I => \N__18580\
        );

    \I__1855\ : InMux
    port map (
            O => \N__18586\,
            I => \N__18577\
        );

    \I__1854\ : LocalMux
    port map (
            O => \N__18583\,
            I => timer_2
        );

    \I__1853\ : LocalMux
    port map (
            O => \N__18580\,
            I => timer_2
        );

    \I__1852\ : LocalMux
    port map (
            O => \N__18577\,
            I => timer_2
        );

    \I__1851\ : InMux
    port map (
            O => \N__18570\,
            I => \nx.n10708\
        );

    \I__1850\ : InMux
    port map (
            O => \N__18567\,
            I => \nx.n10709\
        );

    \I__1849\ : InMux
    port map (
            O => \N__18564\,
            I => \N__18560\
        );

    \I__1848\ : CascadeMux
    port map (
            O => \N__18563\,
            I => \N__18556\
        );

    \I__1847\ : LocalMux
    port map (
            O => \N__18560\,
            I => \N__18553\
        );

    \I__1846\ : InMux
    port map (
            O => \N__18559\,
            I => \N__18550\
        );

    \I__1845\ : InMux
    port map (
            O => \N__18556\,
            I => \N__18547\
        );

    \I__1844\ : Odrv4
    port map (
            O => \N__18553\,
            I => timer_4
        );

    \I__1843\ : LocalMux
    port map (
            O => \N__18550\,
            I => timer_4
        );

    \I__1842\ : LocalMux
    port map (
            O => \N__18547\,
            I => timer_4
        );

    \I__1841\ : InMux
    port map (
            O => \N__18540\,
            I => \nx.n10710\
        );

    \I__1840\ : InMux
    port map (
            O => \N__18537\,
            I => \nx.n10711\
        );

    \I__1839\ : CascadeMux
    port map (
            O => \N__18534\,
            I => \N__18529\
        );

    \I__1838\ : InMux
    port map (
            O => \N__18533\,
            I => \N__18526\
        );

    \I__1837\ : InMux
    port map (
            O => \N__18532\,
            I => \N__18523\
        );

    \I__1836\ : InMux
    port map (
            O => \N__18529\,
            I => \N__18520\
        );

    \I__1835\ : LocalMux
    port map (
            O => \N__18526\,
            I => timer_6
        );

    \I__1834\ : LocalMux
    port map (
            O => \N__18523\,
            I => timer_6
        );

    \I__1833\ : LocalMux
    port map (
            O => \N__18520\,
            I => timer_6
        );

    \I__1832\ : InMux
    port map (
            O => \N__18513\,
            I => \nx.n10712\
        );

    \I__1831\ : InMux
    port map (
            O => \N__18510\,
            I => \N__18506\
        );

    \I__1830\ : CascadeMux
    port map (
            O => \N__18509\,
            I => \N__18502\
        );

    \I__1829\ : LocalMux
    port map (
            O => \N__18506\,
            I => \N__18499\
        );

    \I__1828\ : InMux
    port map (
            O => \N__18505\,
            I => \N__18496\
        );

    \I__1827\ : InMux
    port map (
            O => \N__18502\,
            I => \N__18493\
        );

    \I__1826\ : Odrv4
    port map (
            O => \N__18499\,
            I => timer_7
        );

    \I__1825\ : LocalMux
    port map (
            O => \N__18496\,
            I => timer_7
        );

    \I__1824\ : LocalMux
    port map (
            O => \N__18493\,
            I => timer_7
        );

    \I__1823\ : InMux
    port map (
            O => \N__18486\,
            I => \nx.n10713\
        );

    \I__1822\ : InMux
    port map (
            O => \N__18483\,
            I => \bfn_2_26_0_\
        );

    \I__1821\ : InMux
    port map (
            O => \N__18480\,
            I => \nx.n10781\
        );

    \I__1820\ : InMux
    port map (
            O => \N__18477\,
            I => \nx.n10782\
        );

    \I__1819\ : InMux
    port map (
            O => \N__18474\,
            I => \N__18471\
        );

    \I__1818\ : LocalMux
    port map (
            O => \N__18471\,
            I => \nx.n1469\
        );

    \I__1817\ : InMux
    port map (
            O => \N__18468\,
            I => \N__18462\
        );

    \I__1816\ : InMux
    port map (
            O => \N__18467\,
            I => \N__18462\
        );

    \I__1815\ : LocalMux
    port map (
            O => \N__18462\,
            I => neo_pixel_transmitter_t0_14
        );

    \I__1814\ : InMux
    port map (
            O => \N__18459\,
            I => \N__18456\
        );

    \I__1813\ : LocalMux
    port map (
            O => \N__18456\,
            I => \N__18453\
        );

    \I__1812\ : Span4Mux_v
    port map (
            O => \N__18453\,
            I => \N__18450\
        );

    \I__1811\ : Odrv4
    port map (
            O => \N__18450\,
            I => \nx.n19_adj_725\
        );

    \I__1810\ : InMux
    port map (
            O => \N__18447\,
            I => \bfn_2_25_0_\
        );

    \I__1809\ : InMux
    port map (
            O => \N__18444\,
            I => \nx.n10773\
        );

    \I__1808\ : InMux
    port map (
            O => \N__18441\,
            I => \nx.n10774\
        );

    \I__1807\ : InMux
    port map (
            O => \N__18438\,
            I => \nx.n10775\
        );

    \I__1806\ : InMux
    port map (
            O => \N__18435\,
            I => \nx.n10776\
        );

    \I__1805\ : InMux
    port map (
            O => \N__18432\,
            I => \nx.n10777\
        );

    \I__1804\ : InMux
    port map (
            O => \N__18429\,
            I => \nx.n10778\
        );

    \I__1803\ : InMux
    port map (
            O => \N__18426\,
            I => \nx.n10779\
        );

    \I__1802\ : InMux
    port map (
            O => \N__18423\,
            I => \N__18420\
        );

    \I__1801\ : LocalMux
    port map (
            O => \N__18420\,
            I => \nx.n13201\
        );

    \I__1800\ : InMux
    port map (
            O => \N__18417\,
            I => \bfn_2_23_0_\
        );

    \I__1799\ : InMux
    port map (
            O => \N__18414\,
            I => \N__18411\
        );

    \I__1798\ : LocalMux
    port map (
            O => \N__18411\,
            I => \nx.n13203\
        );

    \I__1797\ : InMux
    port map (
            O => \N__18408\,
            I => \nx.n10696\
        );

    \I__1796\ : InMux
    port map (
            O => \N__18405\,
            I => \N__18402\
        );

    \I__1795\ : LocalMux
    port map (
            O => \N__18402\,
            I => \nx.n13205\
        );

    \I__1794\ : InMux
    port map (
            O => \N__18399\,
            I => \N__18396\
        );

    \I__1793\ : LocalMux
    port map (
            O => \N__18396\,
            I => \N__18393\
        );

    \I__1792\ : Span4Mux_v
    port map (
            O => \N__18393\,
            I => \N__18390\
        );

    \I__1791\ : Odrv4
    port map (
            O => \N__18390\,
            I => \nx.n4_adj_710\
        );

    \I__1790\ : InMux
    port map (
            O => \N__18387\,
            I => \nx.n10697\
        );

    \I__1789\ : InMux
    port map (
            O => \N__18384\,
            I => \N__18381\
        );

    \I__1788\ : LocalMux
    port map (
            O => \N__18381\,
            I => \nx.n13207\
        );

    \I__1787\ : InMux
    port map (
            O => \N__18378\,
            I => \nx.n10698\
        );

    \I__1786\ : InMux
    port map (
            O => \N__18375\,
            I => \N__18372\
        );

    \I__1785\ : LocalMux
    port map (
            O => \N__18372\,
            I => \N__18369\
        );

    \I__1784\ : Odrv4
    port map (
            O => \N__18369\,
            I => \nx.n2\
        );

    \I__1783\ : CascadeMux
    port map (
            O => \N__18366\,
            I => \N__18363\
        );

    \I__1782\ : InMux
    port map (
            O => \N__18363\,
            I => \N__18360\
        );

    \I__1781\ : LocalMux
    port map (
            O => \N__18360\,
            I => \nx.n13209\
        );

    \I__1780\ : InMux
    port map (
            O => \N__18357\,
            I => \nx.n10699\
        );

    \I__1779\ : InMux
    port map (
            O => \N__18354\,
            I => \N__18351\
        );

    \I__1778\ : LocalMux
    port map (
            O => \N__18351\,
            I => \nx.n6\
        );

    \I__1777\ : InMux
    port map (
            O => \N__18348\,
            I => \N__18342\
        );

    \I__1776\ : InMux
    port map (
            O => \N__18347\,
            I => \N__18342\
        );

    \I__1775\ : LocalMux
    port map (
            O => \N__18342\,
            I => neo_pixel_transmitter_t0_27
        );

    \I__1774\ : InMux
    port map (
            O => \N__18339\,
            I => \N__18336\
        );

    \I__1773\ : LocalMux
    port map (
            O => \N__18336\,
            I => \nx.n13189\
        );

    \I__1772\ : CascadeMux
    port map (
            O => \N__18333\,
            I => \N__18330\
        );

    \I__1771\ : InMux
    port map (
            O => \N__18330\,
            I => \N__18327\
        );

    \I__1770\ : LocalMux
    port map (
            O => \N__18327\,
            I => \N__18324\
        );

    \I__1769\ : Span4Mux_v
    port map (
            O => \N__18324\,
            I => \N__18321\
        );

    \I__1768\ : Odrv4
    port map (
            O => \N__18321\,
            I => \nx.n12\
        );

    \I__1767\ : InMux
    port map (
            O => \N__18318\,
            I => \bfn_2_22_0_\
        );

    \I__1766\ : InMux
    port map (
            O => \N__18315\,
            I => \N__18312\
        );

    \I__1765\ : LocalMux
    port map (
            O => \N__18312\,
            I => \nx.n13191\
        );

    \I__1764\ : InMux
    port map (
            O => \N__18309\,
            I => \N__18306\
        );

    \I__1763\ : LocalMux
    port map (
            O => \N__18306\,
            I => \N__18303\
        );

    \I__1762\ : Odrv12
    port map (
            O => \N__18303\,
            I => \nx.n11\
        );

    \I__1761\ : InMux
    port map (
            O => \N__18300\,
            I => \nx.n10690\
        );

    \I__1760\ : InMux
    port map (
            O => \N__18297\,
            I => \N__18294\
        );

    \I__1759\ : LocalMux
    port map (
            O => \N__18294\,
            I => \nx.n13193\
        );

    \I__1758\ : CascadeMux
    port map (
            O => \N__18291\,
            I => \N__18288\
        );

    \I__1757\ : InMux
    port map (
            O => \N__18288\,
            I => \N__18285\
        );

    \I__1756\ : LocalMux
    port map (
            O => \N__18285\,
            I => \N__18282\
        );

    \I__1755\ : Odrv12
    port map (
            O => \N__18282\,
            I => \nx.n10\
        );

    \I__1754\ : InMux
    port map (
            O => \N__18279\,
            I => \nx.n10691\
        );

    \I__1753\ : InMux
    port map (
            O => \N__18276\,
            I => \N__18273\
        );

    \I__1752\ : LocalMux
    port map (
            O => \N__18273\,
            I => \N__18270\
        );

    \I__1751\ : Odrv4
    port map (
            O => \N__18270\,
            I => \nx.n13195\
        );

    \I__1750\ : InMux
    port map (
            O => \N__18267\,
            I => \N__18264\
        );

    \I__1749\ : LocalMux
    port map (
            O => \N__18264\,
            I => \nx.n9\
        );

    \I__1748\ : InMux
    port map (
            O => \N__18261\,
            I => \nx.n10692\
        );

    \I__1747\ : InMux
    port map (
            O => \N__18258\,
            I => \N__18255\
        );

    \I__1746\ : LocalMux
    port map (
            O => \N__18255\,
            I => \N__18252\
        );

    \I__1745\ : Odrv4
    port map (
            O => \N__18252\,
            I => \nx.n13197\
        );

    \I__1744\ : InMux
    port map (
            O => \N__18249\,
            I => \nx.n10693\
        );

    \I__1743\ : InMux
    port map (
            O => \N__18246\,
            I => \N__18243\
        );

    \I__1742\ : LocalMux
    port map (
            O => \N__18243\,
            I => \N__18240\
        );

    \I__1741\ : Odrv4
    port map (
            O => \N__18240\,
            I => \nx.n13199\
        );

    \I__1740\ : InMux
    port map (
            O => \N__18237\,
            I => \nx.n10694\
        );

    \I__1739\ : InMux
    port map (
            O => \N__18234\,
            I => \N__18231\
        );

    \I__1738\ : LocalMux
    port map (
            O => \N__18231\,
            I => \nx.n13177\
        );

    \I__1737\ : CascadeMux
    port map (
            O => \N__18228\,
            I => \N__18225\
        );

    \I__1736\ : InMux
    port map (
            O => \N__18225\,
            I => \N__18222\
        );

    \I__1735\ : LocalMux
    port map (
            O => \N__18222\,
            I => \N__18219\
        );

    \I__1734\ : Odrv12
    port map (
            O => \N__18219\,
            I => \nx.n18_adj_723\
        );

    \I__1733\ : InMux
    port map (
            O => \N__18216\,
            I => \bfn_2_21_0_\
        );

    \I__1732\ : InMux
    port map (
            O => \N__18213\,
            I => \N__18210\
        );

    \I__1731\ : LocalMux
    port map (
            O => \N__18210\,
            I => \nx.n13179\
        );

    \I__1730\ : InMux
    port map (
            O => \N__18207\,
            I => \nx.n10684\
        );

    \I__1729\ : InMux
    port map (
            O => \N__18204\,
            I => \N__18201\
        );

    \I__1728\ : LocalMux
    port map (
            O => \N__18201\,
            I => \nx.n13181\
        );

    \I__1727\ : InMux
    port map (
            O => \N__18198\,
            I => \N__18195\
        );

    \I__1726\ : LocalMux
    port map (
            O => \N__18195\,
            I => \N__18192\
        );

    \I__1725\ : Odrv4
    port map (
            O => \N__18192\,
            I => \nx.n16_adj_672\
        );

    \I__1724\ : InMux
    port map (
            O => \N__18189\,
            I => \nx.n10685\
        );

    \I__1723\ : InMux
    port map (
            O => \N__18186\,
            I => \N__18183\
        );

    \I__1722\ : LocalMux
    port map (
            O => \N__18183\,
            I => \N__18180\
        );

    \I__1721\ : Odrv4
    port map (
            O => \N__18180\,
            I => \nx.n13183\
        );

    \I__1720\ : InMux
    port map (
            O => \N__18177\,
            I => \N__18174\
        );

    \I__1719\ : LocalMux
    port map (
            O => \N__18174\,
            I => \nx.n15\
        );

    \I__1718\ : InMux
    port map (
            O => \N__18171\,
            I => \nx.n10686\
        );

    \I__1717\ : InMux
    port map (
            O => \N__18168\,
            I => \N__18165\
        );

    \I__1716\ : LocalMux
    port map (
            O => \N__18165\,
            I => \nx.n13185\
        );

    \I__1715\ : InMux
    port map (
            O => \N__18162\,
            I => \nx.n10687\
        );

    \I__1714\ : InMux
    port map (
            O => \N__18159\,
            I => \N__18156\
        );

    \I__1713\ : LocalMux
    port map (
            O => \N__18156\,
            I => \N__18153\
        );

    \I__1712\ : Odrv4
    port map (
            O => \N__18153\,
            I => \nx.n13187\
        );

    \I__1711\ : CascadeMux
    port map (
            O => \N__18150\,
            I => \N__18147\
        );

    \I__1710\ : InMux
    port map (
            O => \N__18147\,
            I => \N__18144\
        );

    \I__1709\ : LocalMux
    port map (
            O => \N__18144\,
            I => \nx.n13\
        );

    \I__1708\ : InMux
    port map (
            O => \N__18141\,
            I => \nx.n10688\
        );

    \I__1707\ : InMux
    port map (
            O => \N__18138\,
            I => \N__18135\
        );

    \I__1706\ : LocalMux
    port map (
            O => \N__18135\,
            I => \nx.n26_adj_722\
        );

    \I__1705\ : InMux
    port map (
            O => \N__18132\,
            I => \nx.n10675\
        );

    \I__1704\ : CascadeMux
    port map (
            O => \N__18129\,
            I => \N__18126\
        );

    \I__1703\ : InMux
    port map (
            O => \N__18126\,
            I => \N__18123\
        );

    \I__1702\ : LocalMux
    port map (
            O => \N__18123\,
            I => \N__18120\
        );

    \I__1701\ : Odrv12
    port map (
            O => \N__18120\,
            I => \nx.n25_adj_724\
        );

    \I__1700\ : InMux
    port map (
            O => \N__18117\,
            I => \bfn_2_20_0_\
        );

    \I__1699\ : CascadeMux
    port map (
            O => \N__18114\,
            I => \N__18111\
        );

    \I__1698\ : InMux
    port map (
            O => \N__18111\,
            I => \N__18108\
        );

    \I__1697\ : LocalMux
    port map (
            O => \N__18108\,
            I => \nx.n24_adj_734\
        );

    \I__1696\ : InMux
    port map (
            O => \N__18105\,
            I => \nx.n10677\
        );

    \I__1695\ : InMux
    port map (
            O => \N__18102\,
            I => \N__18099\
        );

    \I__1694\ : LocalMux
    port map (
            O => \N__18099\,
            I => \N__18096\
        );

    \I__1693\ : Odrv4
    port map (
            O => \N__18096\,
            I => \nx.n23\
        );

    \I__1692\ : InMux
    port map (
            O => \N__18093\,
            I => \nx.n10678\
        );

    \I__1691\ : InMux
    port map (
            O => \N__18090\,
            I => \nx.n10679\
        );

    \I__1690\ : InMux
    port map (
            O => \N__18087\,
            I => \N__18084\
        );

    \I__1689\ : LocalMux
    port map (
            O => \N__18084\,
            I => \nx.one_wire_N_599_11\
        );

    \I__1688\ : InMux
    port map (
            O => \N__18081\,
            I => \N__18078\
        );

    \I__1687\ : LocalMux
    port map (
            O => \N__18078\,
            I => \N__18075\
        );

    \I__1686\ : Span4Mux_h
    port map (
            O => \N__18075\,
            I => \N__18072\
        );

    \I__1685\ : Odrv4
    port map (
            O => \N__18072\,
            I => \nx.n21_adj_737\
        );

    \I__1684\ : InMux
    port map (
            O => \N__18069\,
            I => \nx.n10680\
        );

    \I__1683\ : InMux
    port map (
            O => \N__18066\,
            I => \N__18063\
        );

    \I__1682\ : LocalMux
    port map (
            O => \N__18063\,
            I => \nx.n13173\
        );

    \I__1681\ : InMux
    port map (
            O => \N__18060\,
            I => \nx.n10681\
        );

    \I__1680\ : InMux
    port map (
            O => \N__18057\,
            I => \N__18054\
        );

    \I__1679\ : LocalMux
    port map (
            O => \N__18054\,
            I => \nx.n13175\
        );

    \I__1678\ : InMux
    port map (
            O => \N__18051\,
            I => \nx.n10682\
        );

    \I__1677\ : InMux
    port map (
            O => \N__18048\,
            I => \N__18042\
        );

    \I__1676\ : InMux
    port map (
            O => \N__18047\,
            I => \N__18042\
        );

    \I__1675\ : LocalMux
    port map (
            O => \N__18042\,
            I => neo_pixel_transmitter_t0_22
        );

    \I__1674\ : InMux
    port map (
            O => \N__18039\,
            I => \N__18033\
        );

    \I__1673\ : InMux
    port map (
            O => \N__18038\,
            I => \N__18033\
        );

    \I__1672\ : LocalMux
    port map (
            O => \N__18033\,
            I => neo_pixel_transmitter_t0_10
        );

    \I__1671\ : InMux
    port map (
            O => \N__18030\,
            I => \N__18027\
        );

    \I__1670\ : LocalMux
    port map (
            O => \N__18027\,
            I => \N__18024\
        );

    \I__1669\ : Odrv4
    port map (
            O => \N__18024\,
            I => \nx.n33\
        );

    \I__1668\ : InMux
    port map (
            O => \N__18021\,
            I => \nx.n10669\
        );

    \I__1667\ : InMux
    port map (
            O => \N__18018\,
            I => \N__18015\
        );

    \I__1666\ : LocalMux
    port map (
            O => \N__18015\,
            I => \N__18012\
        );

    \I__1665\ : Odrv4
    port map (
            O => \N__18012\,
            I => \nx.n31_adj_711\
        );

    \I__1664\ : InMux
    port map (
            O => \N__18009\,
            I => \nx.n10670\
        );

    \I__1663\ : InMux
    port map (
            O => \N__18006\,
            I => \nx.n10671\
        );

    \I__1662\ : InMux
    port map (
            O => \N__18003\,
            I => \N__18000\
        );

    \I__1661\ : LocalMux
    port map (
            O => \N__18000\,
            I => \nx.n29_adj_714\
        );

    \I__1660\ : InMux
    port map (
            O => \N__17997\,
            I => \nx.n10672\
        );

    \I__1659\ : InMux
    port map (
            O => \N__17994\,
            I => \nx.n10673\
        );

    \I__1658\ : InMux
    port map (
            O => \N__17991\,
            I => \N__17988\
        );

    \I__1657\ : LocalMux
    port map (
            O => \N__17988\,
            I => \nx.n27_adj_720\
        );

    \I__1656\ : InMux
    port map (
            O => \N__17985\,
            I => \nx.n10674\
        );

    \I__1655\ : InMux
    port map (
            O => \N__17982\,
            I => \N__17976\
        );

    \I__1654\ : InMux
    port map (
            O => \N__17981\,
            I => \N__17976\
        );

    \I__1653\ : LocalMux
    port map (
            O => \N__17976\,
            I => neo_pixel_transmitter_t0_23
        );

    \I__1652\ : InMux
    port map (
            O => \N__17973\,
            I => \N__17967\
        );

    \I__1651\ : InMux
    port map (
            O => \N__17972\,
            I => \N__17967\
        );

    \I__1650\ : LocalMux
    port map (
            O => \N__17967\,
            I => neo_pixel_transmitter_t0_15
        );

    \I__1649\ : InMux
    port map (
            O => \N__17964\,
            I => \N__17958\
        );

    \I__1648\ : InMux
    port map (
            O => \N__17963\,
            I => \N__17958\
        );

    \I__1647\ : LocalMux
    port map (
            O => \N__17958\,
            I => neo_pixel_transmitter_t0_8
        );

    \I__1646\ : InMux
    port map (
            O => \N__17955\,
            I => \N__17949\
        );

    \I__1645\ : InMux
    port map (
            O => \N__17954\,
            I => \N__17949\
        );

    \I__1644\ : LocalMux
    port map (
            O => \N__17949\,
            I => neo_pixel_transmitter_t0_2
        );

    \I__1643\ : InMux
    port map (
            O => \N__17946\,
            I => \N__17942\
        );

    \I__1642\ : InMux
    port map (
            O => \N__17945\,
            I => \N__17939\
        );

    \I__1641\ : LocalMux
    port map (
            O => \N__17942\,
            I => neo_pixel_transmitter_t0_6
        );

    \I__1640\ : LocalMux
    port map (
            O => \N__17939\,
            I => neo_pixel_transmitter_t0_6
        );

    \I__1639\ : InMux
    port map (
            O => \N__17934\,
            I => \N__17928\
        );

    \I__1638\ : InMux
    port map (
            O => \N__17933\,
            I => \N__17928\
        );

    \I__1637\ : LocalMux
    port map (
            O => \N__17928\,
            I => neo_pixel_transmitter_t0_17
        );

    \I__1636\ : InMux
    port map (
            O => \N__17925\,
            I => \N__17921\
        );

    \I__1635\ : InMux
    port map (
            O => \N__17924\,
            I => \N__17918\
        );

    \I__1634\ : LocalMux
    port map (
            O => \N__17921\,
            I => \N__17915\
        );

    \I__1633\ : LocalMux
    port map (
            O => \N__17918\,
            I => delay_counter_27
        );

    \I__1632\ : Odrv12
    port map (
            O => \N__17915\,
            I => delay_counter_27
        );

    \I__1631\ : InMux
    port map (
            O => \N__17910\,
            I => n10608
        );

    \I__1630\ : InMux
    port map (
            O => \N__17907\,
            I => n10609
        );

    \I__1629\ : InMux
    port map (
            O => \N__17904\,
            I => n10610
        );

    \I__1628\ : InMux
    port map (
            O => \N__17901\,
            I => \N__17897\
        );

    \I__1627\ : InMux
    port map (
            O => \N__17900\,
            I => \N__17894\
        );

    \I__1626\ : LocalMux
    port map (
            O => \N__17897\,
            I => \N__17891\
        );

    \I__1625\ : LocalMux
    port map (
            O => \N__17894\,
            I => delay_counter_30
        );

    \I__1624\ : Odrv12
    port map (
            O => \N__17891\,
            I => delay_counter_30
        );

    \I__1623\ : InMux
    port map (
            O => \N__17886\,
            I => n10611
        );

    \I__1622\ : InMux
    port map (
            O => \N__17883\,
            I => n10612
        );

    \I__1621\ : InMux
    port map (
            O => \N__17880\,
            I => n10599
        );

    \I__1620\ : InMux
    port map (
            O => \N__17877\,
            I => n10600
        );

    \I__1619\ : InMux
    port map (
            O => \N__17874\,
            I => n10601
        );

    \I__1618\ : InMux
    port map (
            O => \N__17871\,
            I => n10602
        );

    \I__1617\ : InMux
    port map (
            O => \N__17868\,
            I => n10603
        );

    \I__1616\ : CascadeMux
    port map (
            O => \N__17865\,
            I => \N__17862\
        );

    \I__1615\ : InMux
    port map (
            O => \N__17862\,
            I => \N__17858\
        );

    \I__1614\ : InMux
    port map (
            O => \N__17861\,
            I => \N__17855\
        );

    \I__1613\ : LocalMux
    port map (
            O => \N__17858\,
            I => \N__17852\
        );

    \I__1612\ : LocalMux
    port map (
            O => \N__17855\,
            I => delay_counter_23
        );

    \I__1611\ : Odrv12
    port map (
            O => \N__17852\,
            I => delay_counter_23
        );

    \I__1610\ : InMux
    port map (
            O => \N__17847\,
            I => n10604
        );

    \I__1609\ : InMux
    port map (
            O => \N__17844\,
            I => \bfn_1_25_0_\
        );

    \I__1608\ : InMux
    port map (
            O => \N__17841\,
            I => \N__17837\
        );

    \I__1607\ : InMux
    port map (
            O => \N__17840\,
            I => \N__17834\
        );

    \I__1606\ : LocalMux
    port map (
            O => \N__17837\,
            I => \N__17831\
        );

    \I__1605\ : LocalMux
    port map (
            O => \N__17834\,
            I => delay_counter_25
        );

    \I__1604\ : Odrv12
    port map (
            O => \N__17831\,
            I => delay_counter_25
        );

    \I__1603\ : InMux
    port map (
            O => \N__17826\,
            I => n10606
        );

    \I__1602\ : InMux
    port map (
            O => \N__17823\,
            I => n10607
        );

    \I__1601\ : CascadeMux
    port map (
            O => \N__17820\,
            I => \N__17817\
        );

    \I__1600\ : InMux
    port map (
            O => \N__17817\,
            I => \N__17813\
        );

    \I__1599\ : InMux
    port map (
            O => \N__17816\,
            I => \N__17810\
        );

    \I__1598\ : LocalMux
    port map (
            O => \N__17813\,
            I => \N__17807\
        );

    \I__1597\ : LocalMux
    port map (
            O => \N__17810\,
            I => delay_counter_9
        );

    \I__1596\ : Odrv4
    port map (
            O => \N__17807\,
            I => delay_counter_9
        );

    \I__1595\ : InMux
    port map (
            O => \N__17802\,
            I => n10590
        );

    \I__1594\ : InMux
    port map (
            O => \N__17799\,
            I => \N__17795\
        );

    \I__1593\ : InMux
    port map (
            O => \N__17798\,
            I => \N__17792\
        );

    \I__1592\ : LocalMux
    port map (
            O => \N__17795\,
            I => \N__17789\
        );

    \I__1591\ : LocalMux
    port map (
            O => \N__17792\,
            I => delay_counter_10
        );

    \I__1590\ : Odrv4
    port map (
            O => \N__17789\,
            I => delay_counter_10
        );

    \I__1589\ : InMux
    port map (
            O => \N__17784\,
            I => n10591
        );

    \I__1588\ : InMux
    port map (
            O => \N__17781\,
            I => \N__17777\
        );

    \I__1587\ : InMux
    port map (
            O => \N__17780\,
            I => \N__17774\
        );

    \I__1586\ : LocalMux
    port map (
            O => \N__17777\,
            I => \N__17771\
        );

    \I__1585\ : LocalMux
    port map (
            O => \N__17774\,
            I => delay_counter_11
        );

    \I__1584\ : Odrv4
    port map (
            O => \N__17771\,
            I => delay_counter_11
        );

    \I__1583\ : InMux
    port map (
            O => \N__17766\,
            I => n10592
        );

    \I__1582\ : InMux
    port map (
            O => \N__17763\,
            I => \N__17759\
        );

    \I__1581\ : InMux
    port map (
            O => \N__17762\,
            I => \N__17756\
        );

    \I__1580\ : LocalMux
    port map (
            O => \N__17759\,
            I => \N__17753\
        );

    \I__1579\ : LocalMux
    port map (
            O => \N__17756\,
            I => delay_counter_12
        );

    \I__1578\ : Odrv4
    port map (
            O => \N__17753\,
            I => delay_counter_12
        );

    \I__1577\ : InMux
    port map (
            O => \N__17748\,
            I => n10593
        );

    \I__1576\ : InMux
    port map (
            O => \N__17745\,
            I => \N__17741\
        );

    \I__1575\ : InMux
    port map (
            O => \N__17744\,
            I => \N__17738\
        );

    \I__1574\ : LocalMux
    port map (
            O => \N__17741\,
            I => \N__17735\
        );

    \I__1573\ : LocalMux
    port map (
            O => \N__17738\,
            I => delay_counter_13
        );

    \I__1572\ : Odrv4
    port map (
            O => \N__17735\,
            I => delay_counter_13
        );

    \I__1571\ : InMux
    port map (
            O => \N__17730\,
            I => n10594
        );

    \I__1570\ : InMux
    port map (
            O => \N__17727\,
            I => \N__17723\
        );

    \I__1569\ : InMux
    port map (
            O => \N__17726\,
            I => \N__17720\
        );

    \I__1568\ : LocalMux
    port map (
            O => \N__17723\,
            I => \N__17717\
        );

    \I__1567\ : LocalMux
    port map (
            O => \N__17720\,
            I => delay_counter_14
        );

    \I__1566\ : Odrv12
    port map (
            O => \N__17717\,
            I => delay_counter_14
        );

    \I__1565\ : InMux
    port map (
            O => \N__17712\,
            I => n10595
        );

    \I__1564\ : InMux
    port map (
            O => \N__17709\,
            I => n10596
        );

    \I__1563\ : InMux
    port map (
            O => \N__17706\,
            I => \bfn_1_24_0_\
        );

    \I__1562\ : InMux
    port map (
            O => \N__17703\,
            I => n10598
        );

    \I__1561\ : InMux
    port map (
            O => \N__17700\,
            I => \N__17696\
        );

    \I__1560\ : InMux
    port map (
            O => \N__17699\,
            I => \N__17693\
        );

    \I__1559\ : LocalMux
    port map (
            O => \N__17696\,
            I => delay_counter_1
        );

    \I__1558\ : LocalMux
    port map (
            O => \N__17693\,
            I => delay_counter_1
        );

    \I__1557\ : InMux
    port map (
            O => \N__17688\,
            I => n10582
        );

    \I__1556\ : CascadeMux
    port map (
            O => \N__17685\,
            I => \N__17681\
        );

    \I__1555\ : InMux
    port map (
            O => \N__17684\,
            I => \N__17678\
        );

    \I__1554\ : InMux
    port map (
            O => \N__17681\,
            I => \N__17675\
        );

    \I__1553\ : LocalMux
    port map (
            O => \N__17678\,
            I => delay_counter_2
        );

    \I__1552\ : LocalMux
    port map (
            O => \N__17675\,
            I => delay_counter_2
        );

    \I__1551\ : InMux
    port map (
            O => \N__17670\,
            I => n10583
        );

    \I__1550\ : InMux
    port map (
            O => \N__17667\,
            I => \N__17663\
        );

    \I__1549\ : InMux
    port map (
            O => \N__17666\,
            I => \N__17660\
        );

    \I__1548\ : LocalMux
    port map (
            O => \N__17663\,
            I => delay_counter_3
        );

    \I__1547\ : LocalMux
    port map (
            O => \N__17660\,
            I => delay_counter_3
        );

    \I__1546\ : InMux
    port map (
            O => \N__17655\,
            I => n10584
        );

    \I__1545\ : InMux
    port map (
            O => \N__17652\,
            I => \N__17648\
        );

    \I__1544\ : InMux
    port map (
            O => \N__17651\,
            I => \N__17645\
        );

    \I__1543\ : LocalMux
    port map (
            O => \N__17648\,
            I => delay_counter_4
        );

    \I__1542\ : LocalMux
    port map (
            O => \N__17645\,
            I => delay_counter_4
        );

    \I__1541\ : InMux
    port map (
            O => \N__17640\,
            I => n10585
        );

    \I__1540\ : InMux
    port map (
            O => \N__17637\,
            I => \N__17633\
        );

    \I__1539\ : InMux
    port map (
            O => \N__17636\,
            I => \N__17630\
        );

    \I__1538\ : LocalMux
    port map (
            O => \N__17633\,
            I => delay_counter_5
        );

    \I__1537\ : LocalMux
    port map (
            O => \N__17630\,
            I => delay_counter_5
        );

    \I__1536\ : InMux
    port map (
            O => \N__17625\,
            I => n10586
        );

    \I__1535\ : InMux
    port map (
            O => \N__17622\,
            I => \N__17618\
        );

    \I__1534\ : InMux
    port map (
            O => \N__17621\,
            I => \N__17615\
        );

    \I__1533\ : LocalMux
    port map (
            O => \N__17618\,
            I => delay_counter_6
        );

    \I__1532\ : LocalMux
    port map (
            O => \N__17615\,
            I => delay_counter_6
        );

    \I__1531\ : InMux
    port map (
            O => \N__17610\,
            I => n10587
        );

    \I__1530\ : CascadeMux
    port map (
            O => \N__17607\,
            I => \N__17604\
        );

    \I__1529\ : InMux
    port map (
            O => \N__17604\,
            I => \N__17600\
        );

    \I__1528\ : InMux
    port map (
            O => \N__17603\,
            I => \N__17597\
        );

    \I__1527\ : LocalMux
    port map (
            O => \N__17600\,
            I => \N__17594\
        );

    \I__1526\ : LocalMux
    port map (
            O => \N__17597\,
            I => delay_counter_7
        );

    \I__1525\ : Odrv4
    port map (
            O => \N__17594\,
            I => delay_counter_7
        );

    \I__1524\ : InMux
    port map (
            O => \N__17589\,
            I => n10588
        );

    \I__1523\ : InMux
    port map (
            O => \N__17586\,
            I => \N__17582\
        );

    \I__1522\ : InMux
    port map (
            O => \N__17585\,
            I => \N__17579\
        );

    \I__1521\ : LocalMux
    port map (
            O => \N__17582\,
            I => \N__17576\
        );

    \I__1520\ : LocalMux
    port map (
            O => \N__17579\,
            I => delay_counter_8
        );

    \I__1519\ : Odrv4
    port map (
            O => \N__17576\,
            I => delay_counter_8
        );

    \I__1518\ : InMux
    port map (
            O => \N__17571\,
            I => \bfn_1_23_0_\
        );

    \I__1517\ : InMux
    port map (
            O => \N__17568\,
            I => \N__17564\
        );

    \I__1516\ : InMux
    port map (
            O => \N__17567\,
            I => \N__17561\
        );

    \I__1515\ : LocalMux
    port map (
            O => \N__17564\,
            I => neo_pixel_transmitter_t0_18
        );

    \I__1514\ : LocalMux
    port map (
            O => \N__17561\,
            I => neo_pixel_transmitter_t0_18
        );

    \I__1513\ : InMux
    port map (
            O => \N__17556\,
            I => \N__17552\
        );

    \I__1512\ : InMux
    port map (
            O => \N__17555\,
            I => \N__17549\
        );

    \I__1511\ : LocalMux
    port map (
            O => \N__17552\,
            I => neo_pixel_transmitter_t0_20
        );

    \I__1510\ : LocalMux
    port map (
            O => \N__17549\,
            I => neo_pixel_transmitter_t0_20
        );

    \I__1509\ : InMux
    port map (
            O => \N__17544\,
            I => \N__17538\
        );

    \I__1508\ : InMux
    port map (
            O => \N__17543\,
            I => \N__17538\
        );

    \I__1507\ : LocalMux
    port map (
            O => \N__17538\,
            I => neo_pixel_transmitter_t0_24
        );

    \I__1506\ : InMux
    port map (
            O => \N__17535\,
            I => \N__17529\
        );

    \I__1505\ : InMux
    port map (
            O => \N__17534\,
            I => \N__17529\
        );

    \I__1504\ : LocalMux
    port map (
            O => \N__17529\,
            I => neo_pixel_transmitter_t0_31
        );

    \I__1503\ : InMux
    port map (
            O => \N__17526\,
            I => \N__17523\
        );

    \I__1502\ : LocalMux
    port map (
            O => \N__17523\,
            I => n15_adj_841
        );

    \I__1501\ : InMux
    port map (
            O => \N__17520\,
            I => \N__17517\
        );

    \I__1500\ : LocalMux
    port map (
            O => \N__17517\,
            I => n14_adj_842
        );

    \I__1499\ : InMux
    port map (
            O => \N__17514\,
            I => \N__17510\
        );

    \I__1498\ : InMux
    port map (
            O => \N__17513\,
            I => \N__17507\
        );

    \I__1497\ : LocalMux
    port map (
            O => \N__17510\,
            I => \N__17504\
        );

    \I__1496\ : LocalMux
    port map (
            O => \N__17507\,
            I => delay_counter_0
        );

    \I__1495\ : Odrv4
    port map (
            O => \N__17504\,
            I => delay_counter_0
        );

    \I__1494\ : InMux
    port map (
            O => \N__17499\,
            I => \bfn_1_22_0_\
        );

    \I__1493\ : InMux
    port map (
            O => \N__17496\,
            I => \N__17490\
        );

    \I__1492\ : InMux
    port map (
            O => \N__17495\,
            I => \N__17490\
        );

    \I__1491\ : LocalMux
    port map (
            O => \N__17490\,
            I => neo_pixel_transmitter_t0_9
        );

    \I__1490\ : InMux
    port map (
            O => \N__17487\,
            I => \N__17484\
        );

    \I__1489\ : LocalMux
    port map (
            O => \N__17484\,
            I => neopxl_color_prev_12
        );

    \I__1488\ : CascadeMux
    port map (
            O => \N__17481\,
            I => \n24_adj_801_cascade_\
        );

    \I__1487\ : InMux
    port map (
            O => \N__17478\,
            I => \N__17475\
        );

    \I__1486\ : LocalMux
    port map (
            O => \N__17475\,
            I => n12414
        );

    \I__1485\ : InMux
    port map (
            O => \N__17472\,
            I => \N__17469\
        );

    \I__1484\ : LocalMux
    port map (
            O => \N__17469\,
            I => \N__17466\
        );

    \I__1483\ : Odrv4
    port map (
            O => \N__17466\,
            I => neopxl_color_prev_6
        );

    \I__1482\ : InMux
    port map (
            O => \N__17463\,
            I => \N__17457\
        );

    \I__1481\ : InMux
    port map (
            O => \N__17462\,
            I => \N__17457\
        );

    \I__1480\ : LocalMux
    port map (
            O => \N__17457\,
            I => neo_pixel_transmitter_t0_21
        );

    \I__1479\ : InMux
    port map (
            O => \N__17454\,
            I => \N__17448\
        );

    \I__1478\ : InMux
    port map (
            O => \N__17453\,
            I => \N__17448\
        );

    \I__1477\ : LocalMux
    port map (
            O => \N__17448\,
            I => neo_pixel_transmitter_t0_7
        );

    \I__1476\ : InMux
    port map (
            O => \N__17445\,
            I => \N__17439\
        );

    \I__1475\ : InMux
    port map (
            O => \N__17444\,
            I => \N__17439\
        );

    \I__1474\ : LocalMux
    port map (
            O => \N__17439\,
            I => neo_pixel_transmitter_t0_12
        );

    \I__1473\ : InMux
    port map (
            O => \N__17436\,
            I => \N__17430\
        );

    \I__1472\ : InMux
    port map (
            O => \N__17435\,
            I => \N__17430\
        );

    \I__1471\ : LocalMux
    port map (
            O => \N__17430\,
            I => neo_pixel_transmitter_t0_4
        );

    \I__1470\ : InMux
    port map (
            O => \N__17427\,
            I => \N__17421\
        );

    \I__1469\ : InMux
    port map (
            O => \N__17426\,
            I => \N__17421\
        );

    \I__1468\ : LocalMux
    port map (
            O => \N__17421\,
            I => neo_pixel_transmitter_t0_0
        );

    \I__1467\ : IoInMux
    port map (
            O => \N__17418\,
            I => \N__17415\
        );

    \I__1466\ : LocalMux
    port map (
            O => \N__17415\,
            I => \N__17412\
        );

    \I__1465\ : IoSpan4Mux
    port map (
            O => \N__17412\,
            I => \N__17409\
        );

    \I__1464\ : IoSpan4Mux
    port map (
            O => \N__17409\,
            I => \N__17406\
        );

    \I__1463\ : IoSpan4Mux
    port map (
            O => \N__17406\,
            I => \N__17403\
        );

    \I__1462\ : Odrv4
    port map (
            O => \N__17403\,
            I => \CLK_pad_gb_input\
        );

    \IN_MUX_bfv_2_19_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_2_19_0_\
        );

    \IN_MUX_bfv_2_20_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \nx.n10676\,
            carryinitout => \bfn_2_20_0_\
        );

    \IN_MUX_bfv_2_21_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \nx.n10683_THRU_CRY_0_THRU_CO\,
            carryinitout => \bfn_2_21_0_\
        );

    \IN_MUX_bfv_2_22_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \nx.n10689_THRU_CRY_1_THRU_CO\,
            carryinitout => \bfn_2_22_0_\
        );

    \IN_MUX_bfv_2_23_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \nx.n10695_THRU_CRY_1_THRU_CO\,
            carryinitout => \bfn_2_23_0_\
        );

    \IN_MUX_bfv_3_18_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_3_18_0_\
        );

    \IN_MUX_bfv_3_19_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \nx.n10714\,
            carryinitout => \bfn_3_19_0_\
        );

    \IN_MUX_bfv_3_20_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \nx.n10722\,
            carryinitout => \bfn_3_20_0_\
        );

    \IN_MUX_bfv_3_21_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \nx.n10730\,
            carryinitout => \bfn_3_21_0_\
        );

    \IN_MUX_bfv_4_23_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_4_23_0_\
        );

    \IN_MUX_bfv_4_24_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \nx.n10771\,
            carryinitout => \bfn_4_24_0_\
        );

    \IN_MUX_bfv_5_22_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_5_22_0_\
        );

    \IN_MUX_bfv_5_23_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \nx.n10763\,
            carryinitout => \bfn_5_23_0_\
        );

    \IN_MUX_bfv_5_21_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_5_21_0_\
        );

    \IN_MUX_bfv_6_20_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_6_20_0_\
        );

    \IN_MUX_bfv_7_22_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_7_22_0_\
        );

    \IN_MUX_bfv_13_17_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_13_17_0_\
        );

    \IN_MUX_bfv_13_18_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \nx.n11086\,
            carryinitout => \bfn_13_18_0_\
        );

    \IN_MUX_bfv_13_19_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \nx.n11094\,
            carryinitout => \bfn_13_19_0_\
        );

    \IN_MUX_bfv_13_20_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \nx.n11102\,
            carryinitout => \bfn_13_20_0_\
        );

    \IN_MUX_bfv_11_18_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_11_18_0_\
        );

    \IN_MUX_bfv_11_19_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \nx.n11060\,
            carryinitout => \bfn_11_19_0_\
        );

    \IN_MUX_bfv_11_20_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \nx.n11068\,
            carryinitout => \bfn_11_20_0_\
        );

    \IN_MUX_bfv_11_21_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \nx.n11076\,
            carryinitout => \bfn_11_21_0_\
        );

    \IN_MUX_bfv_14_19_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_14_19_0_\
        );

    \IN_MUX_bfv_14_20_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \nx.n11035\,
            carryinitout => \bfn_14_20_0_\
        );

    \IN_MUX_bfv_14_21_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \nx.n11043\,
            carryinitout => \bfn_14_21_0_\
        );

    \IN_MUX_bfv_14_22_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \nx.n11051\,
            carryinitout => \bfn_14_22_0_\
        );

    \IN_MUX_bfv_9_21_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_9_21_0_\
        );

    \IN_MUX_bfv_9_22_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \nx.n11011\,
            carryinitout => \bfn_9_22_0_\
        );

    \IN_MUX_bfv_9_23_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \nx.n11019\,
            carryinitout => \bfn_9_23_0_\
        );

    \IN_MUX_bfv_9_24_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \nx.n11027\,
            carryinitout => \bfn_9_24_0_\
        );

    \IN_MUX_bfv_10_23_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_10_23_0_\
        );

    \IN_MUX_bfv_10_24_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \nx.n10988\,
            carryinitout => \bfn_10_24_0_\
        );

    \IN_MUX_bfv_10_25_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \nx.n10996\,
            carryinitout => \bfn_10_25_0_\
        );

    \IN_MUX_bfv_16_21_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_16_21_0_\
        );

    \IN_MUX_bfv_16_22_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \nx.n10966\,
            carryinitout => \bfn_16_22_0_\
        );

    \IN_MUX_bfv_16_23_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \nx.n10974\,
            carryinitout => \bfn_16_23_0_\
        );

    \IN_MUX_bfv_16_24_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_16_24_0_\
        );

    \IN_MUX_bfv_16_25_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \nx.n10945\,
            carryinitout => \bfn_16_25_0_\
        );

    \IN_MUX_bfv_16_26_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \nx.n10953\,
            carryinitout => \bfn_16_26_0_\
        );

    \IN_MUX_bfv_14_24_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_14_24_0_\
        );

    \IN_MUX_bfv_14_25_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \nx.n10925\,
            carryinitout => \bfn_14_25_0_\
        );

    \IN_MUX_bfv_14_26_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \nx.n10933\,
            carryinitout => \bfn_14_26_0_\
        );

    \IN_MUX_bfv_13_26_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_13_26_0_\
        );

    \IN_MUX_bfv_13_27_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \nx.n10906\,
            carryinitout => \bfn_13_27_0_\
        );

    \IN_MUX_bfv_13_28_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \nx.n10914\,
            carryinitout => \bfn_13_28_0_\
        );

    \IN_MUX_bfv_11_25_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_11_25_0_\
        );

    \IN_MUX_bfv_11_26_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \nx.n10888\,
            carryinitout => \bfn_11_26_0_\
        );

    \IN_MUX_bfv_11_27_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \nx.n10896\,
            carryinitout => \bfn_11_27_0_\
        );

    \IN_MUX_bfv_11_29_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_11_29_0_\
        );

    \IN_MUX_bfv_11_30_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \nx.n10871\,
            carryinitout => \bfn_11_30_0_\
        );

    \IN_MUX_bfv_11_31_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \nx.n10879\,
            carryinitout => \bfn_11_31_0_\
        );

    \IN_MUX_bfv_9_26_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_9_26_0_\
        );

    \IN_MUX_bfv_9_27_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \nx.n10855\,
            carryinitout => \bfn_9_27_0_\
        );

    \IN_MUX_bfv_9_28_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \nx.n10863\,
            carryinitout => \bfn_9_28_0_\
        );

    \IN_MUX_bfv_7_27_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_7_27_0_\
        );

    \IN_MUX_bfv_7_28_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \nx.n10840\,
            carryinitout => \bfn_7_28_0_\
        );

    \IN_MUX_bfv_6_27_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_6_27_0_\
        );

    \IN_MUX_bfv_6_28_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \nx.n10826\,
            carryinitout => \bfn_6_28_0_\
        );

    \IN_MUX_bfv_5_27_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_5_27_0_\
        );

    \IN_MUX_bfv_5_28_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \nx.n10813\,
            carryinitout => \bfn_5_28_0_\
        );

    \IN_MUX_bfv_5_25_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_5_25_0_\
        );

    \IN_MUX_bfv_5_26_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \nx.n10801\,
            carryinitout => \bfn_5_26_0_\
        );

    \IN_MUX_bfv_4_26_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_4_26_0_\
        );

    \IN_MUX_bfv_4_27_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \nx.n10790\,
            carryinitout => \bfn_4_27_0_\
        );

    \IN_MUX_bfv_2_25_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_2_25_0_\
        );

    \IN_MUX_bfv_2_26_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \nx.n10780\,
            carryinitout => \bfn_2_26_0_\
        );

    \IN_MUX_bfv_6_23_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_6_23_0_\
        );

    \IN_MUX_bfv_6_24_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \nx.n10620\,
            carryinitout => \bfn_6_24_0_\
        );

    \IN_MUX_bfv_6_25_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \nx.n10628\,
            carryinitout => \bfn_6_25_0_\
        );

    \IN_MUX_bfv_6_26_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \nx.n10636\,
            carryinitout => \bfn_6_26_0_\
        );

    \IN_MUX_bfv_1_22_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_1_22_0_\
        );

    \IN_MUX_bfv_1_23_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n10589,
            carryinitout => \bfn_1_23_0_\
        );

    \IN_MUX_bfv_1_24_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n10597,
            carryinitout => \bfn_1_24_0_\
        );

    \IN_MUX_bfv_1_25_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n10605,
            carryinitout => \bfn_1_25_0_\
        );

    \IN_MUX_bfv_17_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_17_15_0_\
        );

    \IN_MUX_bfv_9_29_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_9_29_0_\
        );

    \IN_MUX_bfv_9_30_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n10651,
            carryinitout => \bfn_9_30_0_\
        );

    \IN_MUX_bfv_9_31_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n10659,
            carryinitout => \bfn_9_31_0_\
        );

    \IN_MUX_bfv_9_32_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n10667,
            carryinitout => \bfn_9_32_0_\
        );

    \IN_MUX_bfv_17_17_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_17_17_0_\
        );

    \CLK_pad_gb\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__17418\,
            GLOBALBUFFEROUTPUT => \CLK_c\
        );

    \VCC\ : VCC
    port map (
            Y => \VCCG0\
        );

    \GND\ : GND
    port map (
            Y => \GNDG0\
        );

    \GND_Inst\ : GND
    port map (
            Y => \_gnd_net_\
        );

    \nx.neo_pixel_transmitter_t0_i0_i0_LC_1_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__18624\,
            in1 => \N__17427\,
            in2 => \_gnd_net_\,
            in3 => \N__25224\,
            lcout => neo_pixel_transmitter_t0_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46839\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.sub_14_inv_0_i22_1_lut_LC_1_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__17462\,
            lcout => \nx.n12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.sub_14_inv_0_i1_1_lut_LC_1_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__17426\,
            lcout => \nx.n33\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.neo_pixel_transmitter_t0_i0_i21_LC_1_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__25225\,
            in1 => \N__18906\,
            in2 => \_gnd_net_\,
            in3 => \N__17463\,
            lcout => neo_pixel_transmitter_t0_21,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46839\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.neo_pixel_transmitter_t0_i0_i12_LC_1_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__25230\,
            in1 => \N__18714\,
            in2 => \_gnd_net_\,
            in3 => \N__17445\,
            lcout => neo_pixel_transmitter_t0_12,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46841\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.sub_14_inv_0_i8_1_lut_LC_1_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__17453\,
            lcout => \nx.n26_adj_722\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.sub_14_inv_0_i5_1_lut_LC_1_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__17435\,
            lcout => \nx.n29_adj_714\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.neo_pixel_transmitter_t0_i0_i7_LC_1_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__25232\,
            in1 => \N__18510\,
            in2 => \_gnd_net_\,
            in3 => \N__17454\,
            lcout => neo_pixel_transmitter_t0_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46841\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.sub_14_inv_0_i7_1_lut_LC_1_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__17945\,
            lcout => \nx.n27_adj_720\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.sub_14_inv_0_i13_1_lut_LC_1_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__17444\,
            lcout => \nx.n21_adj_737\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.neo_pixel_transmitter_t0_i0_i4_LC_1_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__18564\,
            in1 => \N__17436\,
            in2 => \_gnd_net_\,
            in3 => \N__25231\,
            lcout => neo_pixel_transmitter_t0_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46841\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.neo_pixel_transmitter_t0_i0_i20_LC_1_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__25234\,
            in1 => \N__18933\,
            in2 => \_gnd_net_\,
            in3 => \N__17556\,
            lcout => neo_pixel_transmitter_t0_20,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46843\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.neo_pixel_transmitter_t0_i0_i9_LC_1_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__17496\,
            in1 => \N__18768\,
            in2 => \_gnd_net_\,
            in3 => \N__25235\,
            lcout => neo_pixel_transmitter_t0_9,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46843\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i4_4_lut_adj_169_LC_1_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111101111011110"
        )
    port map (
            in0 => \N__17472\,
            in1 => \N__26606\,
            in2 => \N__26220\,
            in3 => \N__17487\,
            lcout => n12_adj_844,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.sub_14_inv_0_i10_1_lut_LC_1_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__17495\,
            lcout => \nx.n24_adj_734\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \neopxl_color_prev_i12_LC_1_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26607\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => neopxl_color_prev_12,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46843\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.sub_14_inv_0_i30_1_lut_LC_1_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20157\,
            lcout => \nx.n4_adj_710\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.neo_pixel_transmitter_t0_i0_i18_LC_1_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__18966\,
            in1 => \N__17568\,
            in2 => \_gnd_net_\,
            in3 => \N__25233\,
            lcout => neo_pixel_transmitter_t0_18,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46843\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i820_4_lut_LC_1_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100100010001000"
        )
    port map (
            in0 => \N__17799\,
            in1 => \N__17781\,
            in2 => \N__17820\,
            in3 => \N__17478\,
            lcout => OPEN,
            ltout => \n24_adj_801_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i2_4_lut_LC_1_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010100000000000"
        )
    port map (
            in0 => \N__17745\,
            in1 => \N__17763\,
            in2 => \N__17481\,
            in3 => \N__17727\,
            lcout => n12382,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i8_4_lut_LC_1_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__17514\,
            in1 => \N__17520\,
            in2 => \N__17607\,
            in3 => \N__17526\,
            lcout => n12414,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \neopxl_color_prev_i6_LC_1_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26219\,
            lcout => neopxl_color_prev_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46845\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.sub_14_inv_0_i19_1_lut_LC_1_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__17567\,
            lcout => \nx.n15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.sub_14_inv_0_i21_1_lut_LC_1_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17555\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \nx.n13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.neo_pixel_transmitter_t0_i0_i31_LC_1_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__19047\,
            in1 => \N__17535\,
            in2 => \_gnd_net_\,
            in3 => \N__25237\,
            lcout => neo_pixel_transmitter_t0_31,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46848\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.neo_pixel_transmitter_t0_i0_i24_LC_1_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__25236\,
            in1 => \N__18819\,
            in2 => \_gnd_net_\,
            in3 => \N__17544\,
            lcout => neo_pixel_transmitter_t0_24,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46848\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i7_4_lut_LC_1_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__17841\,
            in1 => \N__17925\,
            in2 => \N__17865\,
            in3 => \N__17901\,
            lcout => n18_adj_815,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.sub_14_inv_0_i25_1_lut_LC_1_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__17543\,
            lcout => \nx.n9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.sub_14_inv_0_i32_1_lut_LC_1_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__17534\,
            lcout => \nx.n2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i6_4_lut_LC_1_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__17699\,
            in1 => \N__17621\,
            in2 => \N__17685\,
            in3 => \N__17586\,
            lcout => n15_adj_841,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i5_3_lut_LC_1_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101110"
        )
    port map (
            in0 => \N__17651\,
            in1 => \N__17636\,
            in2 => \_gnd_net_\,
            in3 => \N__17666\,
            lcout => n14_adj_842,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_counter_634__i0_LC_1_22_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17513\,
            in2 => \_gnd_net_\,
            in3 => \N__17499\,
            lcout => delay_counter_0,
            ltout => OPEN,
            carryin => \bfn_1_22_0_\,
            carryout => n10582,
            clk => \N__46852\,
            ce => \N__22314\,
            sr => \N__43506\
        );

    \delay_counter_634__i1_LC_1_22_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17700\,
            in2 => \_gnd_net_\,
            in3 => \N__17688\,
            lcout => delay_counter_1,
            ltout => OPEN,
            carryin => n10582,
            carryout => n10583,
            clk => \N__46852\,
            ce => \N__22314\,
            sr => \N__43506\
        );

    \delay_counter_634__i2_LC_1_22_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17684\,
            in2 => \_gnd_net_\,
            in3 => \N__17670\,
            lcout => delay_counter_2,
            ltout => OPEN,
            carryin => n10583,
            carryout => n10584,
            clk => \N__46852\,
            ce => \N__22314\,
            sr => \N__43506\
        );

    \delay_counter_634__i3_LC_1_22_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17667\,
            in2 => \_gnd_net_\,
            in3 => \N__17655\,
            lcout => delay_counter_3,
            ltout => OPEN,
            carryin => n10584,
            carryout => n10585,
            clk => \N__46852\,
            ce => \N__22314\,
            sr => \N__43506\
        );

    \delay_counter_634__i4_LC_1_22_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17652\,
            in2 => \_gnd_net_\,
            in3 => \N__17640\,
            lcout => delay_counter_4,
            ltout => OPEN,
            carryin => n10585,
            carryout => n10586,
            clk => \N__46852\,
            ce => \N__22314\,
            sr => \N__43506\
        );

    \delay_counter_634__i5_LC_1_22_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17637\,
            in2 => \_gnd_net_\,
            in3 => \N__17625\,
            lcout => delay_counter_5,
            ltout => OPEN,
            carryin => n10586,
            carryout => n10587,
            clk => \N__46852\,
            ce => \N__22314\,
            sr => \N__43506\
        );

    \delay_counter_634__i6_LC_1_22_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17622\,
            in2 => \_gnd_net_\,
            in3 => \N__17610\,
            lcout => delay_counter_6,
            ltout => OPEN,
            carryin => n10587,
            carryout => n10588,
            clk => \N__46852\,
            ce => \N__22314\,
            sr => \N__43506\
        );

    \delay_counter_634__i7_LC_1_22_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17603\,
            in2 => \_gnd_net_\,
            in3 => \N__17589\,
            lcout => delay_counter_7,
            ltout => OPEN,
            carryin => n10588,
            carryout => n10589,
            clk => \N__46852\,
            ce => \N__22314\,
            sr => \N__43506\
        );

    \delay_counter_634__i8_LC_1_23_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17585\,
            in2 => \_gnd_net_\,
            in3 => \N__17571\,
            lcout => delay_counter_8,
            ltout => OPEN,
            carryin => \bfn_1_23_0_\,
            carryout => n10590,
            clk => \N__46858\,
            ce => \N__22303\,
            sr => \N__43491\
        );

    \delay_counter_634__i9_LC_1_23_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17816\,
            in2 => \_gnd_net_\,
            in3 => \N__17802\,
            lcout => delay_counter_9,
            ltout => OPEN,
            carryin => n10590,
            carryout => n10591,
            clk => \N__46858\,
            ce => \N__22303\,
            sr => \N__43491\
        );

    \delay_counter_634__i10_LC_1_23_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17798\,
            in2 => \_gnd_net_\,
            in3 => \N__17784\,
            lcout => delay_counter_10,
            ltout => OPEN,
            carryin => n10591,
            carryout => n10592,
            clk => \N__46858\,
            ce => \N__22303\,
            sr => \N__43491\
        );

    \delay_counter_634__i11_LC_1_23_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17780\,
            in2 => \_gnd_net_\,
            in3 => \N__17766\,
            lcout => delay_counter_11,
            ltout => OPEN,
            carryin => n10592,
            carryout => n10593,
            clk => \N__46858\,
            ce => \N__22303\,
            sr => \N__43491\
        );

    \delay_counter_634__i12_LC_1_23_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17762\,
            in2 => \_gnd_net_\,
            in3 => \N__17748\,
            lcout => delay_counter_12,
            ltout => OPEN,
            carryin => n10593,
            carryout => n10594,
            clk => \N__46858\,
            ce => \N__22303\,
            sr => \N__43491\
        );

    \delay_counter_634__i13_LC_1_23_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17744\,
            in2 => \_gnd_net_\,
            in3 => \N__17730\,
            lcout => delay_counter_13,
            ltout => OPEN,
            carryin => n10594,
            carryout => n10595,
            clk => \N__46858\,
            ce => \N__22303\,
            sr => \N__43491\
        );

    \delay_counter_634__i14_LC_1_23_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17726\,
            in2 => \_gnd_net_\,
            in3 => \N__17712\,
            lcout => delay_counter_14,
            ltout => OPEN,
            carryin => n10595,
            carryout => n10596,
            clk => \N__46858\,
            ce => \N__22303\,
            sr => \N__43491\
        );

    \delay_counter_634__i15_LC_1_23_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19196\,
            in2 => \_gnd_net_\,
            in3 => \N__17709\,
            lcout => delay_counter_15,
            ltout => OPEN,
            carryin => n10596,
            carryout => n10597,
            clk => \N__46858\,
            ce => \N__22303\,
            sr => \N__43491\
        );

    \delay_counter_634__i16_LC_1_24_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20597\,
            in2 => \_gnd_net_\,
            in3 => \N__17706\,
            lcout => delay_counter_16,
            ltout => OPEN,
            carryin => \bfn_1_24_0_\,
            carryout => n10598,
            clk => \N__46863\,
            ce => \N__22302\,
            sr => \N__43505\
        );

    \delay_counter_634__i17_LC_1_24_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19217\,
            in2 => \_gnd_net_\,
            in3 => \N__17703\,
            lcout => delay_counter_17,
            ltout => OPEN,
            carryin => n10598,
            carryout => n10599,
            clk => \N__46863\,
            ce => \N__22302\,
            sr => \N__43505\
        );

    \delay_counter_634__i18_LC_1_24_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20612\,
            in2 => \_gnd_net_\,
            in3 => \N__17880\,
            lcout => delay_counter_18,
            ltout => OPEN,
            carryin => n10599,
            carryout => n10600,
            clk => \N__46863\,
            ce => \N__22302\,
            sr => \N__43505\
        );

    \delay_counter_634__i19_LC_1_24_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22040\,
            in2 => \_gnd_net_\,
            in3 => \N__17877\,
            lcout => delay_counter_19,
            ltout => OPEN,
            carryin => n10600,
            carryout => n10601,
            clk => \N__46863\,
            ce => \N__22302\,
            sr => \N__43505\
        );

    \delay_counter_634__i20_LC_1_24_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22022\,
            in2 => \_gnd_net_\,
            in3 => \N__17874\,
            lcout => delay_counter_20,
            ltout => OPEN,
            carryin => n10601,
            carryout => n10602,
            clk => \N__46863\,
            ce => \N__22302\,
            sr => \N__43505\
        );

    \delay_counter_634__i21_LC_1_24_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19298\,
            in2 => \_gnd_net_\,
            in3 => \N__17871\,
            lcout => delay_counter_21,
            ltout => OPEN,
            carryin => n10602,
            carryout => n10603,
            clk => \N__46863\,
            ce => \N__22302\,
            sr => \N__43505\
        );

    \delay_counter_634__i22_LC_1_24_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20756\,
            in2 => \_gnd_net_\,
            in3 => \N__17868\,
            lcout => delay_counter_22,
            ltout => OPEN,
            carryin => n10603,
            carryout => n10604,
            clk => \N__46863\,
            ce => \N__22302\,
            sr => \N__43505\
        );

    \delay_counter_634__i23_LC_1_24_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17861\,
            in2 => \_gnd_net_\,
            in3 => \N__17847\,
            lcout => delay_counter_23,
            ltout => OPEN,
            carryin => n10604,
            carryout => n10605,
            clk => \N__46863\,
            ce => \N__22302\,
            sr => \N__43505\
        );

    \delay_counter_634__i24_LC_1_25_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20777\,
            in2 => \_gnd_net_\,
            in3 => \N__17844\,
            lcout => delay_counter_24,
            ltout => OPEN,
            carryin => \bfn_1_25_0_\,
            carryout => n10606,
            clk => \N__46870\,
            ce => \N__22310\,
            sr => \N__43492\
        );

    \delay_counter_634__i25_LC_1_25_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17840\,
            in2 => \_gnd_net_\,
            in3 => \N__17826\,
            lcout => delay_counter_25,
            ltout => OPEN,
            carryin => n10606,
            carryout => n10607,
            clk => \N__46870\,
            ce => \N__22310\,
            sr => \N__43492\
        );

    \delay_counter_634__i26_LC_1_25_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20741\,
            in2 => \_gnd_net_\,
            in3 => \N__17823\,
            lcout => delay_counter_26,
            ltout => OPEN,
            carryin => n10607,
            carryout => n10608,
            clk => \N__46870\,
            ce => \N__22310\,
            sr => \N__43492\
        );

    \delay_counter_634__i27_LC_1_25_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17924\,
            in2 => \_gnd_net_\,
            in3 => \N__17910\,
            lcout => delay_counter_27,
            ltout => OPEN,
            carryin => n10608,
            carryout => n10609,
            clk => \N__46870\,
            ce => \N__22310\,
            sr => \N__43492\
        );

    \delay_counter_634__i28_LC_1_25_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20792\,
            in2 => \_gnd_net_\,
            in3 => \N__17907\,
            lcout => delay_counter_28,
            ltout => OPEN,
            carryin => n10609,
            carryout => n10610,
            clk => \N__46870\,
            ce => \N__22310\,
            sr => \N__43492\
        );

    \delay_counter_634__i29_LC_1_25_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19277\,
            in2 => \_gnd_net_\,
            in3 => \N__17904\,
            lcout => delay_counter_29,
            ltout => OPEN,
            carryin => n10610,
            carryout => n10611,
            clk => \N__46870\,
            ce => \N__22310\,
            sr => \N__43492\
        );

    \delay_counter_634__i30_LC_1_25_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17900\,
            in2 => \_gnd_net_\,
            in3 => \N__17886\,
            lcout => delay_counter_30,
            ltout => OPEN,
            carryin => n10611,
            carryout => n10612,
            clk => \N__46870\,
            ce => \N__22310\,
            sr => \N__43492\
        );

    \delay_counter_634__i31_LC_1_25_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23711\,
            in2 => \_gnd_net_\,
            in3 => \N__17883\,
            lcout => delay_counter_31,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46870\,
            ce => \N__22310\,
            sr => \N__43492\
        );

    \nx.sub_14_inv_0_i9_1_lut_LC_2_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__17963\,
            lcout => \nx.n25_adj_724\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.sub_14_inv_0_i3_1_lut_LC_2_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__17954\,
            lcout => \nx.n31_adj_711\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.neo_pixel_transmitter_t0_i0_i15_LC_2_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__17973\,
            in1 => \N__18654\,
            in2 => \_gnd_net_\,
            in3 => \N__25176\,
            lcout => neo_pixel_transmitter_t0_15,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46840\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.sub_14_inv_0_i24_1_lut_LC_2_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__17981\,
            lcout => \nx.n10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.neo_pixel_transmitter_t0_i0_i23_LC_2_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__17982\,
            in1 => \N__18846\,
            in2 => \_gnd_net_\,
            in3 => \N__25177\,
            lcout => neo_pixel_transmitter_t0_23,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46840\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.sub_14_inv_0_i16_1_lut_LC_2_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__17972\,
            lcout => \nx.n18_adj_723\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.neo_pixel_transmitter_t0_i0_i8_LC_2_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__18792\,
            in1 => \N__17964\,
            in2 => \_gnd_net_\,
            in3 => \N__25179\,
            lcout => neo_pixel_transmitter_t0_8,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46840\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.neo_pixel_transmitter_t0_i0_i2_LC_2_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__25178\,
            in1 => \N__18590\,
            in2 => \_gnd_net_\,
            in3 => \N__17955\,
            lcout => neo_pixel_transmitter_t0_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46840\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.neo_pixel_transmitter_t0_i0_i6_LC_2_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__25229\,
            in1 => \N__18533\,
            in2 => \_gnd_net_\,
            in3 => \N__17946\,
            lcout => neo_pixel_transmitter_t0_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46844\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.sub_14_inv_0_i23_1_lut_LC_2_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18047\,
            lcout => \nx.n11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.neo_pixel_transmitter_t0_i0_i17_LC_2_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__25227\,
            in1 => \N__18993\,
            in2 => \_gnd_net_\,
            in3 => \N__17934\,
            lcout => neo_pixel_transmitter_t0_17,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46844\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.neo_pixel_transmitter_t0_i0_i10_LC_2_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__18744\,
            in1 => \N__18039\,
            in2 => \_gnd_net_\,
            in3 => \N__25226\,
            lcout => neo_pixel_transmitter_t0_10,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46844\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.sub_14_inv_0_i18_1_lut_LC_2_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__17933\,
            lcout => \nx.n16_adj_672\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.neo_pixel_transmitter_t0_i0_i22_LC_2_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__18876\,
            in1 => \N__18048\,
            in2 => \_gnd_net_\,
            in3 => \N__25228\,
            lcout => neo_pixel_transmitter_t0_22,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46844\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.sub_14_inv_0_i11_1_lut_LC_2_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18038\,
            lcout => \nx.n23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.sub_14_add_2_2_LC_2_19_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18030\,
            in2 => \N__18620\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_2_19_0_\,
            carryout => \nx.n10669\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.sub_14_add_2_3_lut_LC_2_19_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__21375\,
            in1 => \N__19803\,
            in2 => \N__19743\,
            in3 => \N__18021\,
            lcout => \nx.n4_adj_771\,
            ltout => OPEN,
            carryin => \nx.n10669\,
            carryout => \nx.n10670\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.sub_14_add_2_4_lut_LC_2_19_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18018\,
            in2 => \N__18591\,
            in3 => \N__18009\,
            lcout => \nx.one_wire_N_599_2\,
            ltout => OPEN,
            carryin => \nx.n10670\,
            carryout => \nx.n10671\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.sub_14_add_2_5_lut_LC_2_19_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19815\,
            in2 => \N__19710\,
            in3 => \N__18006\,
            lcout => \nx.one_wire_N_599_3\,
            ltout => OPEN,
            carryin => \nx.n10671\,
            carryout => \nx.n10672\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.sub_14_add_2_6_lut_LC_2_19_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18003\,
            in2 => \N__18563\,
            in3 => \N__17997\,
            lcout => \nx.one_wire_N_599_4\,
            ltout => OPEN,
            carryin => \nx.n10672\,
            carryout => \nx.n10673\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.sub_14_add_2_7_lut_LC_2_19_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19771\,
            in2 => \N__19791\,
            in3 => \N__17994\,
            lcout => \nx.one_wire_N_599_5\,
            ltout => OPEN,
            carryin => \nx.n10673\,
            carryout => \nx.n10674\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.sub_14_add_2_8_lut_LC_2_19_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17991\,
            in2 => \N__18534\,
            in3 => \N__17985\,
            lcout => \nx.one_wire_N_599_6\,
            ltout => OPEN,
            carryin => \nx.n10674\,
            carryout => \nx.n10675\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.sub_14_add_2_9_lut_LC_2_19_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18138\,
            in2 => \N__18509\,
            in3 => \N__18132\,
            lcout => \nx.one_wire_N_599_7\,
            ltout => OPEN,
            carryin => \nx.n10675\,
            carryout => \nx.n10676\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.sub_14_add_2_10_lut_LC_2_20_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18787\,
            in2 => \N__18129\,
            in3 => \N__18117\,
            lcout => \nx.one_wire_N_599_8\,
            ltout => OPEN,
            carryin => \bfn_2_20_0_\,
            carryout => \nx.n10677\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.sub_14_add_2_11_lut_LC_2_20_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18763\,
            in2 => \N__18114\,
            in3 => \N__18105\,
            lcout => \nx.one_wire_N_599_9\,
            ltout => OPEN,
            carryin => \nx.n10677\,
            carryout => \nx.n10678\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.sub_14_add_2_12_lut_LC_2_20_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18102\,
            in2 => \N__18743\,
            in3 => \N__18093\,
            lcout => \nx.one_wire_N_599_10\,
            ltout => OPEN,
            carryin => \nx.n10678\,
            carryout => \nx.n10679\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.sub_14_add_2_13_lut_LC_2_20_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21426\,
            in2 => \N__21560\,
            in3 => \N__18090\,
            lcout => \nx.one_wire_N_599_11\,
            ltout => OPEN,
            carryin => \nx.n10679\,
            carryout => \nx.n10680\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.sub_14_add_2_14_lut_LC_2_20_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101110111110"
        )
    port map (
            in0 => \N__18087\,
            in1 => \N__18081\,
            in2 => \N__18710\,
            in3 => \N__18069\,
            lcout => \nx.n13173\,
            ltout => OPEN,
            carryin => \nx.n10680\,
            carryout => \nx.n10681\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.sub_14_add_2_15_lut_LC_2_20_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101110111110"
        )
    port map (
            in0 => \N__18066\,
            in1 => \N__19944\,
            in2 => \N__19932\,
            in3 => \N__18060\,
            lcout => \nx.n13175\,
            ltout => OPEN,
            carryin => \nx.n10681\,
            carryout => \nx.n10682\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.sub_14_add_2_16_lut_LC_2_20_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101110111110"
        )
    port map (
            in0 => \N__18057\,
            in1 => \N__18459\,
            in2 => \N__18680\,
            in3 => \N__18051\,
            lcout => \nx.n13177\,
            ltout => OPEN,
            carryin => \nx.n10682\,
            carryout => \nx.n10683\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.sub_14_add_2_16_THRU_CRY_0_LC_2_20_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42223\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \nx.n10683\,
            carryout => \nx.n10683_THRU_CRY_0_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.sub_14_add_2_17_lut_LC_2_21_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101110111110"
        )
    port map (
            in0 => \N__18234\,
            in1 => \N__18650\,
            in2 => \N__18228\,
            in3 => \N__18216\,
            lcout => \nx.n13179\,
            ltout => OPEN,
            carryin => \bfn_2_21_0_\,
            carryout => \nx.n10684\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.sub_14_add_2_18_lut_LC_2_21_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101110111110"
        )
    port map (
            in0 => \N__18213\,
            in1 => \N__19138\,
            in2 => \N__19110\,
            in3 => \N__18207\,
            lcout => \nx.n13181\,
            ltout => OPEN,
            carryin => \nx.n10684\,
            carryout => \nx.n10685\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.sub_14_add_2_19_lut_LC_2_21_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101110111110"
        )
    port map (
            in0 => \N__18204\,
            in1 => \N__18198\,
            in2 => \N__18992\,
            in3 => \N__18189\,
            lcout => \nx.n13183\,
            ltout => OPEN,
            carryin => \nx.n10685\,
            carryout => \nx.n10686\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.sub_14_add_2_20_lut_LC_2_21_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101110111110"
        )
    port map (
            in0 => \N__18186\,
            in1 => \N__18177\,
            in2 => \N__18965\,
            in3 => \N__18171\,
            lcout => \nx.n13185\,
            ltout => OPEN,
            carryin => \nx.n10686\,
            carryout => \nx.n10687\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.sub_14_add_2_21_lut_LC_2_21_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101110111110"
        )
    port map (
            in0 => \N__18168\,
            in1 => \N__21402\,
            in2 => \N__19881\,
            in3 => \N__18162\,
            lcout => \nx.n13187\,
            ltout => OPEN,
            carryin => \nx.n10687\,
            carryout => \nx.n10688\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.sub_14_add_2_22_lut_LC_2_21_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101110111110"
        )
    port map (
            in0 => \N__18159\,
            in1 => \N__18925\,
            in2 => \N__18150\,
            in3 => \N__18141\,
            lcout => \nx.n13189\,
            ltout => OPEN,
            carryin => \nx.n10688\,
            carryout => \nx.n10689\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.sub_14_add_2_22_THRU_CRY_0_LC_2_21_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42225\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \nx.n10689\,
            carryout => \nx.n10689_THRU_CRY_0_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.sub_14_add_2_22_THRU_CRY_1_LC_2_21_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \GNDG0\,
            in2 => \N__42281\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \nx.n10689_THRU_CRY_0_THRU_CO\,
            carryout => \nx.n10689_THRU_CRY_1_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.sub_14_add_2_23_lut_LC_2_22_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101110111110"
        )
    port map (
            in0 => \N__18339\,
            in1 => \N__18902\,
            in2 => \N__18333\,
            in3 => \N__18318\,
            lcout => \nx.n13191\,
            ltout => OPEN,
            carryin => \bfn_2_22_0_\,
            carryout => \nx.n10690\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.sub_14_add_2_24_lut_LC_2_22_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101110111110"
        )
    port map (
            in0 => \N__18315\,
            in1 => \N__18309\,
            in2 => \N__18875\,
            in3 => \N__18300\,
            lcout => \nx.n13193\,
            ltout => OPEN,
            carryin => \nx.n10690\,
            carryout => \nx.n10691\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.sub_14_add_2_25_lut_LC_2_22_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101110111110"
        )
    port map (
            in0 => \N__18297\,
            in1 => \N__18842\,
            in2 => \N__18291\,
            in3 => \N__18279\,
            lcout => \nx.n13195\,
            ltout => OPEN,
            carryin => \nx.n10691\,
            carryout => \nx.n10692\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.sub_14_add_2_26_lut_LC_2_22_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101110111110"
        )
    port map (
            in0 => \N__18276\,
            in1 => \N__18267\,
            in2 => \N__18818\,
            in3 => \N__18261\,
            lcout => \nx.n13197\,
            ltout => OPEN,
            carryin => \nx.n10692\,
            carryout => \nx.n10693\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.sub_14_add_2_27_lut_LC_2_22_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101110111110"
        )
    port map (
            in0 => \N__18258\,
            in1 => \N__19897\,
            in2 => \N__20127\,
            in3 => \N__18249\,
            lcout => \nx.n13199\,
            ltout => OPEN,
            carryin => \nx.n10693\,
            carryout => \nx.n10694\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.sub_14_add_2_28_lut_LC_2_22_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101110111110"
        )
    port map (
            in0 => \N__18246\,
            in1 => \N__23295\,
            in2 => \N__23327\,
            in3 => \N__18237\,
            lcout => \nx.n13201\,
            ltout => OPEN,
            carryin => \nx.n10694\,
            carryout => \nx.n10695\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.sub_14_add_2_28_THRU_CRY_0_LC_2_22_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42229\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \nx.n10695\,
            carryout => \nx.n10695_THRU_CRY_0_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.sub_14_add_2_28_THRU_CRY_1_LC_2_22_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42224\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \nx.n10695_THRU_CRY_0_THRU_CO\,
            carryout => \nx.n10695_THRU_CRY_1_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.sub_14_add_2_29_lut_LC_2_23_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101110111110"
        )
    port map (
            in0 => \N__18423\,
            in1 => \N__18354\,
            in2 => \N__19089\,
            in3 => \N__18417\,
            lcout => \nx.n13203\,
            ltout => OPEN,
            carryin => \bfn_2_23_0_\,
            carryout => \nx.n10696\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.sub_14_add_2_30_lut_LC_2_23_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101110111110"
        )
    port map (
            in0 => \N__18414\,
            in1 => \N__23664\,
            in2 => \N__25268\,
            in3 => \N__18408\,
            lcout => \nx.n13205\,
            ltout => OPEN,
            carryin => \nx.n10696\,
            carryout => \nx.n10697\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.sub_14_add_2_31_lut_LC_2_23_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101110111110"
        )
    port map (
            in0 => \N__18405\,
            in1 => \N__18399\,
            in2 => \N__20184\,
            in3 => \N__18387\,
            lcout => \nx.n13207\,
            ltout => OPEN,
            carryin => \nx.n10697\,
            carryout => \nx.n10698\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.sub_14_add_2_32_lut_LC_2_23_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101110111110"
        )
    port map (
            in0 => \N__18384\,
            in1 => \N__19641\,
            in2 => \N__21119\,
            in3 => \N__18378\,
            lcout => \nx.n13209\,
            ltout => OPEN,
            carryin => \nx.n10698\,
            carryout => \nx.n10699\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.sub_14_add_2_33_lut_LC_2_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100111110110"
        )
    port map (
            in0 => \N__18375\,
            in1 => \N__19046\,
            in2 => \N__18366\,
            in3 => \N__18357\,
            lcout => \nx.n7608\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.sub_14_inv_0_i28_1_lut_LC_2_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18347\,
            lcout => \nx.n6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.neo_pixel_transmitter_t0_i0_i27_LC_2_23_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__18348\,
            in1 => \N__19088\,
            in2 => \_gnd_net_\,
            in3 => \N__25239\,
            lcout => neo_pixel_transmitter_t0_27,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46864\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \neopxl_color_i6_LC_2_24_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0101010101000000"
        )
    port map (
            in0 => \N__43675\,
            in1 => \N__43955\,
            in2 => \N__47697\,
            in3 => \N__26207\,
            lcout => neopxl_color_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46871\,
            ce => 'H',
            sr => \N__20406\
        );

    \nx.mod_5_i946_3_lut_LC_2_24_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20367\,
            in2 => \N__20481\,
            in3 => \N__20381\,
            lcout => \nx.n1407\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i948_3_lut_LC_2_24_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__20226\,
            in1 => \N__25482\,
            in2 => \_gnd_net_\,
            in3 => \N__20476\,
            lcout => \nx.n1409\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1004_2_lut_LC_2_25_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24096\,
            in2 => \_gnd_net_\,
            in3 => \N__18447\,
            lcout => \nx.n1477\,
            ltout => OPEN,
            carryin => \bfn_2_25_0_\,
            carryout => \nx.n10773\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1004_3_lut_LC_2_25_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__19608\,
            in3 => \N__18444\,
            lcout => \nx.n1476\,
            ltout => OPEN,
            carryin => \nx.n10773\,
            carryout => \nx.n10774\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1004_4_lut_LC_2_25_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42282\,
            in2 => \N__19571\,
            in3 => \N__18441\,
            lcout => \nx.n1475\,
            ltout => OPEN,
            carryin => \nx.n10774\,
            carryout => \nx.n10775\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1004_5_lut_LC_2_25_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42288\,
            in2 => \N__19322\,
            in3 => \N__18438\,
            lcout => \nx.n1474\,
            ltout => OPEN,
            carryin => \nx.n10775\,
            carryout => \nx.n10776\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1004_6_lut_LC_2_25_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42283\,
            in2 => \N__19443\,
            in3 => \N__18435\,
            lcout => \nx.n1473\,
            ltout => OPEN,
            carryin => \nx.n10776\,
            carryout => \nx.n10777\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1004_7_lut_LC_2_25_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19388\,
            in2 => \N__42299\,
            in3 => \N__18432\,
            lcout => \nx.n1472\,
            ltout => OPEN,
            carryin => \nx.n10777\,
            carryout => \nx.n10778\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1004_8_lut_LC_2_25_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42287\,
            in2 => \N__19422\,
            in3 => \N__18429\,
            lcout => \nx.n1471\,
            ltout => OPEN,
            carryin => \nx.n10778\,
            carryout => \nx.n10779\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1004_9_lut_LC_2_25_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42289\,
            in2 => \N__19349\,
            in3 => \N__18426\,
            lcout => \nx.n1470\,
            ltout => OPEN,
            carryin => \nx.n10779\,
            carryout => \nx.n10780\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1004_10_lut_LC_2_26_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19238\,
            in2 => \N__42300\,
            in3 => \N__18483\,
            lcout => \nx.n1469\,
            ltout => OPEN,
            carryin => \bfn_2_26_0_\,
            carryout => \nx.n10781\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1004_11_lut_LC_2_26_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42293\,
            in2 => \N__20436\,
            in3 => \N__18480\,
            lcout => \nx.n1468\,
            ltout => OPEN,
            carryin => \nx.n10781\,
            carryout => \nx.n10782\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1004_12_lut_LC_2_26_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001000001100000"
        )
    port map (
            in0 => \N__42294\,
            in1 => \N__20259\,
            in2 => \N__19521\,
            in3 => \N__18477\,
            lcout => \nx.n1499\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i18_4_lut_adj_134_LC_2_26_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__24105\,
            in1 => \N__23829\,
            in2 => \N__30534\,
            in3 => \N__36060\,
            lcout => \nx.n46_adj_779\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1008_3_lut_LC_2_26_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18474\,
            in2 => \N__19242\,
            in3 => \N__19514\,
            lcout => \nx.n1501\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.neo_pixel_transmitter_t0_i0_i14_LC_3_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__18681\,
            in1 => \N__18468\,
            in2 => \_gnd_net_\,
            in3 => \N__25156\,
            lcout => neo_pixel_transmitter_t0_14,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46846\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.sub_14_inv_0_i15_1_lut_LC_3_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18467\,
            lcout => \nx.n19_adj_725\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.neo_pixel_transmitter_done_104_LC_3_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101000010001"
        )
    port map (
            in0 => \N__24908\,
            in1 => \N__23250\,
            in2 => \_gnd_net_\,
            in3 => \N__23493\,
            lcout => \nx.neo_pixel_transmitter_done\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46842\,
            ce => \N__20079\,
            sr => \_gnd_net_\
        );

    \nx.i9152_2_lut_LC_3_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26800\,
            in2 => \_gnd_net_\,
            in3 => \N__24907\,
            lcout => OPEN,
            ltout => \nx.n11834_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i1_4_lut_adj_151_LC_3_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000111110001"
        )
    port map (
            in0 => \N__21327\,
            in1 => \N__21382\,
            in2 => \N__18627\,
            in3 => \N__21296\,
            lcout => \nx.n103\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.timer_632__i0_LC_3_18_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18616\,
            in2 => \_gnd_net_\,
            in3 => \N__18597\,
            lcout => timer_0,
            ltout => OPEN,
            carryin => \bfn_3_18_0_\,
            carryout => \nx.n10707\,
            clk => \N__46847\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.timer_632__i1_LC_3_18_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19741\,
            in2 => \_gnd_net_\,
            in3 => \N__18594\,
            lcout => timer_1,
            ltout => OPEN,
            carryin => \nx.n10707\,
            carryout => \nx.n10708\,
            clk => \N__46847\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.timer_632__i2_LC_3_18_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18589\,
            in2 => \_gnd_net_\,
            in3 => \N__18570\,
            lcout => timer_2,
            ltout => OPEN,
            carryin => \nx.n10708\,
            carryout => \nx.n10709\,
            clk => \N__46847\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.timer_632__i3_LC_3_18_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19708\,
            in2 => \_gnd_net_\,
            in3 => \N__18567\,
            lcout => timer_3,
            ltout => OPEN,
            carryin => \nx.n10709\,
            carryout => \nx.n10710\,
            clk => \N__46847\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.timer_632__i4_LC_3_18_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18559\,
            in2 => \_gnd_net_\,
            in3 => \N__18540\,
            lcout => timer_4,
            ltout => OPEN,
            carryin => \nx.n10710\,
            carryout => \nx.n10711\,
            clk => \N__46847\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.timer_632__i5_LC_3_18_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19772\,
            in2 => \_gnd_net_\,
            in3 => \N__18537\,
            lcout => timer_5,
            ltout => OPEN,
            carryin => \nx.n10711\,
            carryout => \nx.n10712\,
            clk => \N__46847\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.timer_632__i6_LC_3_18_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18532\,
            in2 => \_gnd_net_\,
            in3 => \N__18513\,
            lcout => timer_6,
            ltout => OPEN,
            carryin => \nx.n10712\,
            carryout => \nx.n10713\,
            clk => \N__46847\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.timer_632__i7_LC_3_18_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18505\,
            in2 => \_gnd_net_\,
            in3 => \N__18486\,
            lcout => timer_7,
            ltout => OPEN,
            carryin => \nx.n10713\,
            carryout => \nx.n10714\,
            clk => \N__46847\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.timer_632__i8_LC_3_19_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18788\,
            in2 => \_gnd_net_\,
            in3 => \N__18771\,
            lcout => timer_8,
            ltout => OPEN,
            carryin => \bfn_3_19_0_\,
            carryout => \nx.n10715\,
            clk => \N__46849\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.timer_632__i9_LC_3_19_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18764\,
            in2 => \_gnd_net_\,
            in3 => \N__18747\,
            lcout => timer_9,
            ltout => OPEN,
            carryin => \nx.n10715\,
            carryout => \nx.n10716\,
            clk => \N__46849\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.timer_632__i10_LC_3_19_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18739\,
            in2 => \_gnd_net_\,
            in3 => \N__18720\,
            lcout => timer_10,
            ltout => OPEN,
            carryin => \nx.n10716\,
            carryout => \nx.n10717\,
            clk => \N__46849\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.timer_632__i11_LC_3_19_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21556\,
            in2 => \_gnd_net_\,
            in3 => \N__18717\,
            lcout => timer_11,
            ltout => OPEN,
            carryin => \nx.n10717\,
            carryout => \nx.n10718\,
            clk => \N__46849\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.timer_632__i12_LC_3_19_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18706\,
            in2 => \_gnd_net_\,
            in3 => \N__18687\,
            lcout => timer_12,
            ltout => OPEN,
            carryin => \nx.n10718\,
            carryout => \nx.n10719\,
            clk => \N__46849\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.timer_632__i13_LC_3_19_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19927\,
            in2 => \_gnd_net_\,
            in3 => \N__18684\,
            lcout => timer_13,
            ltout => OPEN,
            carryin => \nx.n10719\,
            carryout => \nx.n10720\,
            clk => \N__46849\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.timer_632__i14_LC_3_19_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18676\,
            in2 => \_gnd_net_\,
            in3 => \N__18657\,
            lcout => timer_14,
            ltout => OPEN,
            carryin => \nx.n10720\,
            carryout => \nx.n10721\,
            clk => \N__46849\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.timer_632__i15_LC_3_19_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18649\,
            in2 => \_gnd_net_\,
            in3 => \N__18630\,
            lcout => timer_15,
            ltout => OPEN,
            carryin => \nx.n10721\,
            carryout => \nx.n10722\,
            clk => \N__46849\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.timer_632__i16_LC_3_20_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19139\,
            in2 => \_gnd_net_\,
            in3 => \N__18996\,
            lcout => timer_16,
            ltout => OPEN,
            carryin => \bfn_3_20_0_\,
            carryout => \nx.n10723\,
            clk => \N__46853\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.timer_632__i17_LC_3_20_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18988\,
            in2 => \_gnd_net_\,
            in3 => \N__18969\,
            lcout => timer_17,
            ltout => OPEN,
            carryin => \nx.n10723\,
            carryout => \nx.n10724\,
            clk => \N__46853\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.timer_632__i18_LC_3_20_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18958\,
            in2 => \_gnd_net_\,
            in3 => \N__18939\,
            lcout => timer_18,
            ltout => OPEN,
            carryin => \nx.n10724\,
            carryout => \nx.n10725\,
            clk => \N__46853\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.timer_632__i19_LC_3_20_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19879\,
            in2 => \_gnd_net_\,
            in3 => \N__18936\,
            lcout => timer_19,
            ltout => OPEN,
            carryin => \nx.n10725\,
            carryout => \nx.n10726\,
            clk => \N__46853\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.timer_632__i20_LC_3_20_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18926\,
            in2 => \_gnd_net_\,
            in3 => \N__18909\,
            lcout => timer_20,
            ltout => OPEN,
            carryin => \nx.n10726\,
            carryout => \nx.n10727\,
            clk => \N__46853\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.timer_632__i21_LC_3_20_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18898\,
            in2 => \_gnd_net_\,
            in3 => \N__18879\,
            lcout => timer_21,
            ltout => OPEN,
            carryin => \nx.n10727\,
            carryout => \nx.n10728\,
            clk => \N__46853\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.timer_632__i22_LC_3_20_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18868\,
            in2 => \_gnd_net_\,
            in3 => \N__18849\,
            lcout => timer_22,
            ltout => OPEN,
            carryin => \nx.n10728\,
            carryout => \nx.n10729\,
            clk => \N__46853\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.timer_632__i23_LC_3_20_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18841\,
            in2 => \_gnd_net_\,
            in3 => \N__18822\,
            lcout => timer_23,
            ltout => OPEN,
            carryin => \nx.n10729\,
            carryout => \nx.n10730\,
            clk => \N__46853\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.timer_632__i24_LC_3_21_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18814\,
            in2 => \_gnd_net_\,
            in3 => \N__18795\,
            lcout => timer_24,
            ltout => OPEN,
            carryin => \bfn_3_21_0_\,
            carryout => \nx.n10731\,
            clk => \N__46859\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.timer_632__i25_LC_3_21_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19898\,
            in2 => \_gnd_net_\,
            in3 => \N__19095\,
            lcout => timer_25,
            ltout => OPEN,
            carryin => \nx.n10731\,
            carryout => \nx.n10732\,
            clk => \N__46859\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.timer_632__i26_LC_3_21_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23323\,
            in2 => \_gnd_net_\,
            in3 => \N__19092\,
            lcout => timer_26,
            ltout => OPEN,
            carryin => \nx.n10732\,
            carryout => \nx.n10733\,
            clk => \N__46859\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.timer_632__i27_LC_3_21_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19084\,
            in2 => \_gnd_net_\,
            in3 => \N__19062\,
            lcout => timer_27,
            ltout => OPEN,
            carryin => \nx.n10733\,
            carryout => \nx.n10734\,
            clk => \N__46859\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.timer_632__i28_LC_3_21_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25258\,
            in2 => \_gnd_net_\,
            in3 => \N__19059\,
            lcout => timer_28,
            ltout => OPEN,
            carryin => \nx.n10734\,
            carryout => \nx.n10735\,
            clk => \N__46859\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.timer_632__i29_LC_3_21_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20176\,
            in2 => \_gnd_net_\,
            in3 => \N__19056\,
            lcout => timer_29,
            ltout => OPEN,
            carryin => \nx.n10735\,
            carryout => \nx.n10736\,
            clk => \N__46859\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.timer_632__i30_LC_3_21_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21109\,
            in2 => \_gnd_net_\,
            in3 => \N__19053\,
            lcout => timer_30,
            ltout => OPEN,
            carryin => \nx.n10736\,
            carryout => \nx.n10737\,
            clk => \N__46859\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.timer_632__i31_LC_3_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19045\,
            in2 => \_gnd_net_\,
            in3 => \N__19050\,
            lcout => timer_31,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46859\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_2_lut_3_lut_4_lut_4_lut_adj_184_LC_3_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011001000"
        )
    port map (
            in0 => \N__45020\,
            in1 => \N__47667\,
            in2 => \N__45695\,
            in3 => \N__42639\,
            lcout => OPEN,
            ltout => \n11826_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pin_output_enable__i1_LC_3_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100111011000100"
        )
    port map (
            in0 => \N__47125\,
            in1 => \N__19007\,
            in2 => \N__19023\,
            in3 => \N__47672\,
            lcout => pin_oe_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46865\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i4_4_lut_LC_3_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__19221\,
            in1 => \N__20583\,
            in2 => \N__19203\,
            in3 => \N__19182\,
            lcout => n12379,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_2_lut_3_lut_4_lut_4_lut_adj_187_LC_3_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010001010"
        )
    port map (
            in0 => \N__47666\,
            in1 => \N__42635\,
            in2 => \N__45696\,
            in3 => \N__45021\,
            lcout => OPEN,
            ltout => \n11828_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pin_output_enable__i5_LC_3_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010110010101010"
        )
    port map (
            in0 => \N__19154\,
            in1 => \N__47668\,
            in2 => \N__19170\,
            in3 => \N__47126\,
            lcout => pin_oe_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46865\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.neo_pixel_transmitter_t0_i0_i16_LC_3_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__19143\,
            in1 => \N__19122\,
            in2 => \_gnd_net_\,
            in3 => \N__25220\,
            lcout => neo_pixel_transmitter_t0_16,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46865\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i874_3_lut_LC_3_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22095\,
            in2 => \N__22119\,
            in3 => \N__21980\,
            lcout => \nx.n1303\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i944_3_lut_LC_3_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010101010"
        )
    port map (
            in0 => \N__20342\,
            in1 => \_gnd_net_\,
            in2 => \N__20325\,
            in3 => \N__20467\,
            lcout => \nx.n1405\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.sub_14_inv_0_i17_1_lut_LC_3_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19121\,
            lcout => \nx.n17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i880_3_lut_LC_3_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__21777\,
            in1 => \N__24053\,
            in2 => \_gnd_net_\,
            in3 => \N__21965\,
            lcout => \nx.n1309\,
            ltout => \nx.n1309_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i3_3_lut_LC_3_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25477\,
            in2 => \N__19098\,
            in3 => \N__20341\,
            lcout => \nx.n12_adj_669\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i6_4_lut_adj_158_LC_3_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011111010"
        )
    port map (
            in0 => \N__19302\,
            in1 => \N__22008\,
            in2 => \N__19284\,
            in3 => \N__19263\,
            lcout => n17_adj_816,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i879_3_lut_LC_3_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21761\,
            in2 => \N__21981\,
            in3 => \N__21741\,
            lcout => \nx.n1308\,
            ltout => \nx.n1308_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i8_4_lut_LC_3_23_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__19257\,
            in1 => \N__20290\,
            in2 => \N__19251\,
            in3 => \N__20496\,
            lcout => \nx.n1334\,
            ltout => \nx.n1334_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i941_3_lut_LC_3_23_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101000001010"
        )
    port map (
            in0 => \N__20291\,
            in1 => \_gnd_net_\,
            in2 => \N__19248\,
            in3 => \N__20274\,
            lcout => \nx.n1402\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i9149_3_lut_LC_3_24_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20313\,
            in2 => \N__20550\,
            in3 => \N__20475\,
            lcout => \nx.n1404\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i945_3_lut_LC_3_24_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20352\,
            in2 => \N__20480\,
            in3 => \N__20519\,
            lcout => \nx.n1406\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i942_3_lut_LC_3_24_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20573\,
            in2 => \N__20304\,
            in3 => \N__20474\,
            lcout => \nx.n1403\,
            ltout => \nx.n1403_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i3_3_lut_adj_72_LC_3_24_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24103\,
            in2 => \N__19245\,
            in3 => \N__19603\,
            lcout => \nx.n13_adj_729\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i6_4_lut_adj_71_LC_3_24_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__20252\,
            in1 => \N__19232\,
            in2 => \N__19387\,
            in3 => \N__20422\,
            lcout => OPEN,
            ltout => \nx.n16_adj_727_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i8_3_lut_LC_3_24_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19438\,
            in2 => \N__19461\,
            in3 => \N__19564\,
            lcout => \nx.n18_adj_728\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i947_3_lut_LC_3_24_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20210\,
            in2 => \N__20196\,
            in3 => \N__20470\,
            lcout => \nx.n1408\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1010_3_lut_LC_3_25_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19418\,
            in2 => \N__19458\,
            in3 => \N__19505\,
            lcout => \nx.n1503\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1012_3_lut_LC_3_25_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__19449\,
            in1 => \_gnd_net_\,
            in2 => \N__19520\,
            in3 => \N__19442\,
            lcout => \nx.n1505\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i9_4_lut_adj_73_LC_3_25_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__19318\,
            in1 => \N__19417\,
            in2 => \N__19404\,
            in3 => \N__19395\,
            lcout => \nx.n1433\,
            ltout => \nx.n1433_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1011_3_lut_LC_3_25_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19389\,
            in2 => \N__19365\,
            in3 => \N__19362\,
            lcout => \nx.n1504\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1009_3_lut_LC_3_25_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19356\,
            in2 => \N__19350\,
            in3 => \N__19509\,
            lcout => \nx.n1502\,
            ltout => \nx.n1502_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i5_2_lut_LC_3_25_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__19332\,
            in3 => \N__21007\,
            lcout => \nx.n16_adj_732\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1013_3_lut_LC_3_25_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19329\,
            in2 => \N__19323\,
            in3 => \N__19513\,
            lcout => \nx.n1506\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1015_3_lut_LC_3_25_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19614\,
            in2 => \N__19519\,
            in3 => \N__19607\,
            lcout => \nx.n1508\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1007_3_lut_LC_3_26_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20432\,
            in2 => \N__19587\,
            in3 => \N__19501\,
            lcout => \nx.n1500\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1014_3_lut_LC_3_26_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19578\,
            in2 => \N__19518\,
            in3 => \N__19572\,
            lcout => \nx.n1507\,
            ltout => \nx.n1507_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i7_4_lut_adj_75_LC_3_26_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__21028\,
            in1 => \N__20689\,
            in2 => \N__19548\,
            in3 => \N__19467\,
            lcout => OPEN,
            ltout => \nx.n18_adj_731_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i9_4_lut_adj_76_LC_3_26_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__20632\,
            in1 => \N__20957\,
            in2 => \N__19545\,
            in3 => \N__20941\,
            lcout => OPEN,
            ltout => \nx.n20_adj_733_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i10_4_lut_adj_77_LC_3_26_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__20909\,
            in1 => \N__20653\,
            in2 => \N__19542\,
            in3 => \N__19539\,
            lcout => \nx.n1532\,
            ltout => \nx.n1532_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i9208_1_lut_LC_3_26_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__19533\,
            in3 => \_gnd_net_\,
            lcout => \nx.n13604\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1016_3_lut_LC_3_26_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__19530\,
            in1 => \N__24104\,
            in2 => \_gnd_net_\,
            in3 => \N__19500\,
            lcout => \nx.n1509\,
            ltout => \nx.n1509_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i5936_2_lut_LC_3_26_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__19470\,
            in3 => \N__23826\,
            lcout => \nx.n9729\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i26_4_lut_adj_139_LC_3_27_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__20808\,
            in1 => \N__19647\,
            in2 => \N__24717\,
            in3 => \N__20823\,
            lcout => \nx.n54\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.start_103_LC_4_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23249\,
            in2 => \_gnd_net_\,
            in3 => \N__23492\,
            lcout => \nx.start\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46850\,
            ce => \N__19620\,
            sr => \_gnd_net_\
        );

    \nx.sub_14_inv_0_i31_1_lut_LC_4_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21089\,
            lcout => \nx.n3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i20_4_lut_adj_116_LC_4_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111011001111"
        )
    port map (
            in0 => \N__24945\,
            in1 => \N__23470\,
            in2 => \N__23259\,
            in3 => \N__21078\,
            lcout => OPEN,
            ltout => \nx.n7_adj_764_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i1_4_lut_adj_118_LC_4_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011010000"
        )
    port map (
            in0 => \N__21348\,
            in1 => \N__22872\,
            in2 => \N__19626\,
            in3 => \N__23479\,
            lcout => n11353,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i7535_3_lut_LC_4_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111010101010"
        )
    port map (
            in0 => \N__23248\,
            in1 => \N__24933\,
            in2 => \_gnd_net_\,
            in3 => \N__21347\,
            lcout => OPEN,
            ltout => \nx.n11864_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i15_4_lut_adj_150_LC_4_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111010000110000"
        )
    port map (
            in0 => \N__21390\,
            in1 => \N__23480\,
            in2 => \N__19623\,
            in3 => \N__21269\,
            lcout => \nx.n7_adj_667\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i7561_2_lut_LC_4_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__23243\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__23469\,
            lcout => \nx.n11892\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i9093_2_lut_3_lut_LC_4_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101110"
        )
    port map (
            in0 => \N__23244\,
            in1 => \N__21333\,
            in2 => \_gnd_net_\,
            in3 => \N__21384\,
            lcout => \nx.n13445\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i6_4_lut_adj_152_LC_4_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000100"
        )
    port map (
            in0 => \N__19989\,
            in1 => \N__19830\,
            in2 => \N__19824\,
            in3 => \N__20067\,
            lcout => \nx.n16_adj_785\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.sub_14_inv_0_i4_1_lut_LC_4_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19688\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \nx.n30_adj_712\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.sub_14_inv_0_i2_1_lut_LC_4_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19718\,
            lcout => \nx.n32\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.sub_14_inv_0_i6_1_lut_LC_4_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19751\,
            lcout => \nx.n28_adj_715\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.neo_pixel_transmitter_t0_i0_i5_LC_4_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__25117\,
            in1 => \_gnd_net_\,
            in2 => \N__19755\,
            in3 => \N__19773\,
            lcout => neo_pixel_transmitter_t0_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46851\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.neo_pixel_transmitter_t0_i0_i1_LC_4_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110001011100010"
        )
    port map (
            in0 => \N__19742\,
            in1 => \N__25116\,
            in2 => \N__19722\,
            in3 => \_gnd_net_\,
            lcout => neo_pixel_transmitter_t0_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46851\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i1_2_lut_adj_147_LC_4_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19670\,
            in2 => \_gnd_net_\,
            in3 => \N__20100\,
            lcout => \nx.n13211\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.neo_pixel_transmitter_t0_i0_i3_LC_4_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__25166\,
            in1 => \N__19709\,
            in2 => \_gnd_net_\,
            in3 => \N__19689\,
            lcout => neo_pixel_transmitter_t0_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46854\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i1_4_lut_adj_153_LC_4_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111011"
        )
    port map (
            in0 => \N__20049\,
            in1 => \N__19677\,
            in2 => \N__19671\,
            in3 => \N__19962\,
            lcout => OPEN,
            ltout => \nx.n6_adj_786_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i4_4_lut_adj_154_LC_4_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__20030\,
            in1 => \N__20009\,
            in2 => \N__20103\,
            in3 => \N__20099\,
            lcout => \nx.n13659\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i5953_4_lut_LC_4_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111100000"
        )
    port map (
            in0 => \N__20048\,
            in1 => \N__19988\,
            in2 => \N__20010\,
            in3 => \N__19961\,
            lcout => \nx.n9747\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i1_4_lut_adj_148_LC_4_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__20063\,
            in1 => \N__20047\,
            in2 => \N__20031\,
            in3 => \N__20016\,
            lcout => OPEN,
            ltout => \nx.n13217_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i1_4_lut_adj_149_LC_4_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__20005\,
            in1 => \N__19987\,
            in2 => \N__19965\,
            in3 => \N__19960\,
            lcout => \nx.n7564\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.sub_14_inv_0_i14_1_lut_LC_4_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19907\,
            lcout => \nx.n20_adj_726\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.neo_pixel_transmitter_t0_i0_i13_LC_4_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__19908\,
            in1 => \N__19928\,
            in2 => \_gnd_net_\,
            in3 => \N__25165\,
            lcout => neo_pixel_transmitter_t0_13,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46854\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.neo_pixel_transmitter_t0_i0_i25_LC_4_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__19899\,
            in1 => \N__20139\,
            in2 => \_gnd_net_\,
            in3 => \N__25217\,
            lcout => neo_pixel_transmitter_t0_25,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46860\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.neo_pixel_transmitter_t0_i0_i19_LC_4_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__19880\,
            in1 => \N__21414\,
            in2 => \_gnd_net_\,
            in3 => \N__25216\,
            lcout => neo_pixel_transmitter_t0_19,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46860\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i8987_3_lut_LC_4_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__19860\,
            in1 => \N__19842\,
            in2 => \_gnd_net_\,
            in3 => \N__46410\,
            lcout => n13382,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.neo_pixel_transmitter_t0_i0_i29_LC_4_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__20177\,
            in1 => \N__20153\,
            in2 => \_gnd_net_\,
            in3 => \N__25218\,
            lcout => neo_pixel_transmitter_t0_29,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46860\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i809_rep_49_3_lut_LC_4_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23628\,
            in2 => \N__21576\,
            in3 => \N__21816\,
            lcout => \nx.n1206\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.sub_14_inv_0_i26_1_lut_LC_4_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20138\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \nx.n8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i808_3_lut_LC_4_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21899\,
            in2 => \N__21827\,
            in3 => \N__21879\,
            lcout => \nx.n1205\,
            ltout => \nx.n1205_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i3_3_lut_adj_18_LC_4_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24054\,
            in2 => \N__20112\,
            in3 => \N__21760\,
            lcout => \nx.n11_adj_674\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i810_3_lut_LC_4_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21605\,
            in2 => \N__21826\,
            in3 => \N__21585\,
            lcout => \nx.n1207\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i811_3_lut_LC_4_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21632\,
            in2 => \N__21618\,
            in3 => \N__21809\,
            lcout => \nx.n1208\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i807_3_lut_LC_4_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23517\,
            in2 => \N__21825\,
            in3 => \N__21870\,
            lcout => \nx.n1204\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i7_4_lut_adj_20_LC_4_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__21670\,
            in1 => \N__21697\,
            in2 => \N__20235\,
            in3 => \N__20109\,
            lcout => \nx.n1235\,
            ltout => \nx.n1235_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i875_3_lut_LC_4_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22142\,
            in2 => \N__20241\,
            in3 => \N__22128\,
            lcout => \nx.n1304\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i812_3_lut_LC_4_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__21645\,
            in1 => \N__24000\,
            in2 => \_gnd_net_\,
            in3 => \N__21821\,
            lcout => \nx.n1209\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i806_3_lut_LC_4_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21861\,
            in2 => \N__21828\,
            in3 => \N__21837\,
            lcout => \nx.n1203\,
            ltout => \nx.n1203_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i5_4_lut_adj_19_LC_4_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__22073\,
            in1 => \N__21724\,
            in2 => \N__20238\,
            in3 => \N__22111\,
            lcout => \nx.n13_adj_675\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i878_3_lut_LC_4_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101000001010"
        )
    port map (
            in0 => \N__21725\,
            in1 => \_gnd_net_\,
            in2 => \N__21983\,
            in3 => \N__21708\,
            lcout => \nx.n1307\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i876_3_lut_LC_4_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010101010"
        )
    port map (
            in0 => \N__21671\,
            in1 => \_gnd_net_\,
            in2 => \N__22155\,
            in3 => \N__21973\,
            lcout => \nx.n1305\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i877_3_lut_LC_4_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101000001010"
        )
    port map (
            in0 => \N__21698\,
            in1 => \_gnd_net_\,
            in2 => \N__21984\,
            in3 => \N__21681\,
            lcout => \nx.n1306\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_937_2_lut_LC_4_23_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25476\,
            in2 => \_gnd_net_\,
            in3 => \N__20214\,
            lcout => \nx.n1377\,
            ltout => OPEN,
            carryin => \bfn_4_23_0_\,
            carryout => \nx.n10764\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_937_3_lut_LC_4_23_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__20211\,
            in3 => \N__20187\,
            lcout => \nx.n1376\,
            ltout => OPEN,
            carryin => \nx.n10764\,
            carryout => \nx.n10765\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_937_4_lut_LC_4_23_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41610\,
            in2 => \N__20382\,
            in3 => \N__20355\,
            lcout => \nx.n1375\,
            ltout => OPEN,
            carryin => \nx.n10765\,
            carryout => \nx.n10766\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_937_5_lut_LC_4_23_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41613\,
            in2 => \N__20520\,
            in3 => \N__20346\,
            lcout => \nx.n1374\,
            ltout => OPEN,
            carryin => \nx.n10766\,
            carryout => \nx.n10767\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_937_6_lut_LC_4_23_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41611\,
            in2 => \N__20343\,
            in3 => \N__20316\,
            lcout => \nx.n1373\,
            ltout => OPEN,
            carryin => \nx.n10767\,
            carryout => \nx.n10768\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_937_7_lut_LC_4_23_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41614\,
            in2 => \N__20549\,
            in3 => \N__20307\,
            lcout => \nx.n1372\,
            ltout => OPEN,
            carryin => \nx.n10768\,
            carryout => \nx.n10769\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_937_8_lut_LC_4_23_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41612\,
            in2 => \N__20574\,
            in3 => \N__20295\,
            lcout => \nx.n1371\,
            ltout => OPEN,
            carryin => \nx.n10769\,
            carryout => \nx.n10770\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_937_9_lut_LC_4_23_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41615\,
            in2 => \N__20292\,
            in3 => \N__20268\,
            lcout => \nx.n1370\,
            ltout => OPEN,
            carryin => \nx.n10770\,
            carryout => \nx.n10771\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_937_10_lut_LC_4_24_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42279\,
            in2 => \N__21930\,
            in3 => \N__20265\,
            lcout => \nx.n1369\,
            ltout => OPEN,
            carryin => \bfn_4_24_0_\,
            carryout => \nx.n10772\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_937_11_lut_LC_4_24_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000010001001000"
        )
    port map (
            in0 => \N__42280\,
            in1 => \N__20469\,
            in2 => \N__22059\,
            in3 => \N__20262\,
            lcout => \nx.n1400\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_2_lut_adj_156_LC_4_24_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20613\,
            in2 => \_gnd_net_\,
            in3 => \N__20598\,
            lcout => n6_adj_843,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i1_2_lut_LC_4_24_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__22058\,
            in3 => \N__21925\,
            lcout => OPEN,
            ltout => \nx.n10_adj_668_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i7_4_lut_LC_4_24_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__20572\,
            in1 => \N__20545\,
            in2 => \N__20523\,
            in3 => \N__20518\,
            lcout => \nx.n16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i940_3_lut_LC_4_24_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21929\,
            in2 => \N__20490\,
            in3 => \N__20468\,
            lcout => \nx.n1401\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_2_lut_3_lut_adj_185_LC_4_24_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101000000000"
        )
    port map (
            in0 => \N__47665\,
            in1 => \_gnd_net_\,
            in2 => \N__43940\,
            in3 => \N__26209\,
            lcout => n22_adj_795,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i11_4_lut_LC_4_25_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__22216\,
            in1 => \N__20799\,
            in2 => \N__22536\,
            in3 => \N__20388\,
            lcout => \nx.n1631\,
            ltout => \nx.n1631_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i9206_1_lut_LC_4_25_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__20394\,
            in3 => \_gnd_net_\,
            lcout => \nx.n13602\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i3_3_lut_adj_21_LC_4_25_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23866\,
            in2 => \N__22260\,
            in3 => \N__22174\,
            lcout => OPEN,
            ltout => \nx.n15_adj_676_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i10_4_lut_LC_4_25_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__22555\,
            in1 => \N__22416\,
            in2 => \N__20391\,
            in3 => \N__20817\,
            lcout => \nx.n22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i19_4_lut_adj_135_LC_4_25_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__30146\,
            in1 => \N__24052\,
            in2 => \N__25332\,
            in3 => \N__28213\,
            lcout => \nx.n47_adj_780\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i6_2_lut_LC_4_25_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__22512\,
            in3 => \N__22576\,
            lcout => \nx.n18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i8_4_lut_adj_159_LC_4_25_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__20793\,
            in1 => \N__20778\,
            in2 => \N__20763\,
            in3 => \N__20742\,
            lcout => n19_adj_814,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1071_2_lut_LC_4_26_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__23828\,
            in1 => \N__23827\,
            in2 => \N__20711\,
            in3 => \N__20727\,
            lcout => \nx.n1609\,
            ltout => OPEN,
            carryin => \bfn_4_26_0_\,
            carryout => \nx.n10783\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1071_3_lut_LC_4_26_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__20724\,
            in1 => \N__20723\,
            in2 => \N__20712\,
            in3 => \N__20694\,
            lcout => \nx.n1608\,
            ltout => OPEN,
            carryin => \nx.n10783\,
            carryout => \nx.n10784\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1071_4_lut_LC_4_26_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101000111010"
        )
    port map (
            in0 => \N__20691\,
            in1 => \N__20690\,
            in2 => \N__20889\,
            in3 => \N__20673\,
            lcout => \nx.n1607\,
            ltout => OPEN,
            carryin => \nx.n10784\,
            carryout => \nx.n10785\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1071_5_lut_LC_4_26_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101000111010"
        )
    port map (
            in0 => \N__20670\,
            in1 => \N__20669\,
            in2 => \N__20892\,
            in3 => \N__20658\,
            lcout => \nx.n1606\,
            ltout => OPEN,
            carryin => \nx.n10785\,
            carryout => \nx.n10786\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1071_6_lut_LC_4_26_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101000111010"
        )
    port map (
            in0 => \N__20655\,
            in1 => \N__20654\,
            in2 => \N__20890\,
            in3 => \N__20637\,
            lcout => \nx.n1605\,
            ltout => OPEN,
            carryin => \nx.n10786\,
            carryout => \nx.n10787\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1071_7_lut_LC_4_26_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101000111010"
        )
    port map (
            in0 => \N__20634\,
            in1 => \N__20633\,
            in2 => \N__20893\,
            in3 => \N__20616\,
            lcout => \nx.n1604\,
            ltout => OPEN,
            carryin => \nx.n10787\,
            carryout => \nx.n10788\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1071_8_lut_LC_4_26_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101000111010"
        )
    port map (
            in0 => \N__21030\,
            in1 => \N__21029\,
            in2 => \N__20891\,
            in3 => \N__21012\,
            lcout => \nx.n1603\,
            ltout => OPEN,
            carryin => \nx.n10788\,
            carryout => \nx.n10789\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1071_9_lut_LC_4_26_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101000111010"
        )
    port map (
            in0 => \N__21009\,
            in1 => \N__21008\,
            in2 => \N__20894\,
            in3 => \N__20991\,
            lcout => \nx.n1602\,
            ltout => OPEN,
            carryin => \nx.n10789\,
            carryout => \nx.n10790\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1071_10_lut_LC_4_27_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101000111010"
        )
    port map (
            in0 => \N__20988\,
            in1 => \N__20987\,
            in2 => \N__20895\,
            in3 => \N__20973\,
            lcout => \nx.n1601\,
            ltout => OPEN,
            carryin => \bfn_4_27_0_\,
            carryout => \nx.n10791\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1071_11_lut_LC_4_27_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101000111010"
        )
    port map (
            in0 => \N__20970\,
            in1 => \N__20969\,
            in2 => \N__20897\,
            in3 => \N__20946\,
            lcout => \nx.n1600\,
            ltout => OPEN,
            carryin => \nx.n10791\,
            carryout => \nx.n10792\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1071_12_lut_LC_4_27_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101000111010"
        )
    port map (
            in0 => \N__20942\,
            in1 => \N__20943\,
            in2 => \N__20896\,
            in3 => \N__20925\,
            lcout => \nx.n1599\,
            ltout => OPEN,
            carryin => \nx.n10792\,
            carryout => \nx.n10793\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1071_13_lut_LC_4_27_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101000111010"
        )
    port map (
            in0 => \N__20922\,
            in1 => \N__20921\,
            in2 => \N__20898\,
            in3 => \N__20826\,
            lcout => \nx.n1598\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i17_4_lut_adj_136_LC_4_27_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__28936\,
            in1 => \N__23952\,
            in2 => \N__26034\,
            in3 => \N__34340\,
            lcout => \nx.n45_adj_781\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i7_4_lut_adj_22_LC_4_27_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__22195\,
            in1 => \N__22483\,
            in2 => \N__22462\,
            in3 => \N__22435\,
            lcout => \nx.n19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_pin_0__bdd_4_lut_LC_5_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001110001000"
        )
    port map (
            in0 => \N__21234\,
            in1 => \N__46545\,
            in2 => \N__21216\,
            in3 => \N__46405\,
            lcout => n13649,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pin_output_enable__i6_LC_5_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101100011001100"
        )
    port map (
            in0 => \N__22893\,
            in1 => \N__21176\,
            in2 => \N__47675\,
            in3 => \N__47121\,
            lcout => pin_oe_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46861\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \n13649_bdd_4_lut_LC_5_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000110000"
        )
    port map (
            in0 => \N__21165\,
            in1 => \N__46566\,
            in2 => \N__21147\,
            in3 => \N__21126\,
            lcout => n13652,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.neo_pixel_transmitter_t0_i0_i30_LC_5_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__21120\,
            in1 => \N__21090\,
            in2 => \_gnd_net_\,
            in3 => \N__25157\,
            lcout => neo_pixel_transmitter_t0_30,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46855\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i7610_4_lut_LC_5_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001010"
        )
    port map (
            in0 => \N__23203\,
            in1 => \N__22855\,
            in2 => \N__26805\,
            in3 => \N__23183\,
            lcout => \nx.n11946\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i53_4_lut_LC_5_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011111010"
        )
    port map (
            in0 => \N__21072\,
            in1 => \N__21268\,
            in2 => \N__23187\,
            in3 => \N__23481\,
            lcout => OPEN,
            ltout => \nx.n11948_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i52_4_lut_LC_5_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000111101111"
        )
    port map (
            in0 => \N__24943\,
            in1 => \N__26795\,
            in2 => \N__21066\,
            in3 => \N__22887\,
            lcout => \nx.n11988\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i8984_3_lut_LC_5_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__21063\,
            in1 => \N__21048\,
            in2 => \_gnd_net_\,
            in3 => \N__46396\,
            lcout => OPEN,
            ltout => \n13379_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \n13613_bdd_4_lut_LC_5_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000100010"
        )
    port map (
            in0 => \N__21507\,
            in1 => \N__45645\,
            in2 => \N__21033\,
            in3 => \N__21447\,
            lcout => n13616,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i3_4_lut_4_lut_LC_5_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000100"
        )
    port map (
            in0 => \N__26796\,
            in1 => \N__23482\,
            in2 => \N__21276\,
            in3 => \N__24944\,
            lcout => \nx.n12451\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i9091_2_lut_LC_5_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__24942\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26794\,
            lcout => \nx.n13438\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \neopxl_color_i15_LC_5_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111011100010000"
        )
    port map (
            in0 => \N__47673\,
            in1 => \N__43939\,
            in2 => \N__43701\,
            in3 => \N__25757\,
            lcout => neopxl_color_15,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46856\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i1_2_lut_adj_145_LC_5_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21331\,
            in2 => \_gnd_net_\,
            in3 => \N__21383\,
            lcout => \nx.n11908\,
            ltout => \nx.n11908_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i7592_4_lut_LC_5_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111100100"
        )
    port map (
            in0 => \N__26802\,
            in1 => \N__22854\,
            in2 => \N__21351\,
            in3 => \N__23168\,
            lcout => \nx.n11926\,
            ltout => \nx.n11926_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i1_4_lut_adj_127_LC_5_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101000000000"
        )
    port map (
            in0 => \N__23472\,
            in1 => \N__22868\,
            in2 => \N__21339\,
            in3 => \N__21240\,
            lcout => n7671,
            ltout => \n7671_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.state_i1_LC_5_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101111111110000"
        )
    port map (
            in0 => \N__26803\,
            in1 => \N__26855\,
            in2 => \N__21336\,
            in3 => \N__23473\,
            lcout => state_1_adj_791,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46856\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i2_2_lut_adj_146_LC_5_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21332\,
            in2 => \_gnd_net_\,
            in3 => \N__21297\,
            lcout => \nx.n11113\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i1_3_lut_4_lut_LC_5_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011111110111011"
        )
    port map (
            in0 => \N__26801\,
            in1 => \N__23471\,
            in2 => \N__24957\,
            in3 => \N__21258\,
            lcout => \nx.n12381\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.neo_pixel_transmitter_t0_i0_i11_LC_5_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__21564\,
            in1 => \N__21438\,
            in2 => \_gnd_net_\,
            in3 => \N__25155\,
            lcout => neo_pixel_transmitter_t0_11,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46856\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i8983_3_lut_LC_5_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__21537\,
            in1 => \N__21522\,
            in2 => \_gnd_net_\,
            in3 => \N__46407\,
            lcout => n13378,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i8986_3_lut_LC_5_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__21498\,
            in1 => \N__21477\,
            in2 => \_gnd_net_\,
            in3 => \N__46406\,
            lcout => OPEN,
            ltout => \n13381_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_pin_1__bdd_4_lut_9226_LC_5_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110100000"
        )
    port map (
            in0 => \N__45644\,
            in1 => \N__21456\,
            in2 => \N__21450\,
            in3 => \N__46565\,
            lcout => n13613,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.sub_14_inv_0_i12_1_lut_LC_5_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21437\,
            lcout => \nx.n22_adj_749\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i739_3_lut_LC_5_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__23553\,
            in1 => \_gnd_net_\,
            in2 => \N__23604\,
            in3 => \N__23361\,
            lcout => \nx.n1104\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i743_3_lut_LC_5_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23582\,
            in2 => \N__23388\,
            in3 => \N__23552\,
            lcout => \nx.n1108\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.sub_14_inv_0_i20_1_lut_LC_5_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__21413\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \nx.n14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i741_3_lut_LC_5_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23548\,
            in2 => \N__23652\,
            in3 => \N__23373\,
            lcout => \nx.n1106\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i744_3_lut_LC_5_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23397\,
            in2 => \N__23558\,
            in3 => \N__23951\,
            lcout => \nx.n1109\,
            ltout => \nx.n1109_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i5944_2_lut_LC_5_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__21654\,
            in3 => \N__23998\,
            lcout => OPEN,
            ltout => \nx.n9737_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i5_4_lut_LC_5_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__21601\,
            in1 => \N__21895\,
            in2 => \N__21651\,
            in3 => \N__23509\,
            lcout => OPEN,
            ltout => \nx.n12_adj_673_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i6_4_lut_LC_5_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__23623\,
            in1 => \N__23348\,
            in2 => \N__21648\,
            in3 => \N__21853\,
            lcout => \nx.n1136\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_803_2_lut_LC_5_21_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23999\,
            in2 => \_gnd_net_\,
            in3 => \N__21636\,
            lcout => \nx.n1177\,
            ltout => OPEN,
            carryin => \bfn_5_21_0_\,
            carryout => \nx.n10749\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_803_3_lut_LC_5_21_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__21633\,
            in3 => \N__21609\,
            lcout => \nx.n1176\,
            ltout => OPEN,
            carryin => \nx.n10749\,
            carryout => \nx.n10750\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_803_4_lut_LC_5_21_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42219\,
            in2 => \N__21606\,
            in3 => \N__21579\,
            lcout => \nx.n1175\,
            ltout => OPEN,
            carryin => \nx.n10750\,
            carryout => \nx.n10751\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_803_5_lut_LC_5_21_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42193\,
            in2 => \N__23627\,
            in3 => \N__21567\,
            lcout => \nx.n1174\,
            ltout => OPEN,
            carryin => \nx.n10751\,
            carryout => \nx.n10752\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_803_6_lut_LC_5_21_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42220\,
            in2 => \N__21900\,
            in3 => \N__21873\,
            lcout => \nx.n1173\,
            ltout => OPEN,
            carryin => \nx.n10752\,
            carryout => \nx.n10753\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_803_7_lut_LC_5_21_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42194\,
            in2 => \N__23516\,
            in3 => \N__21864\,
            lcout => \nx.n1172\,
            ltout => OPEN,
            carryin => \nx.n10753\,
            carryout => \nx.n10754\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_803_8_lut_LC_5_21_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42221\,
            in2 => \N__21860\,
            in3 => \N__21831\,
            lcout => \nx.n1171\,
            ltout => OPEN,
            carryin => \nx.n10754\,
            carryout => \nx.n10755\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_803_9_lut_LC_5_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000010001001000"
        )
    port map (
            in0 => \N__42222\,
            in1 => \N__21820\,
            in2 => \N__23349\,
            in3 => \N__21780\,
            lcout => \nx.n1202\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_870_2_lut_LC_5_22_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24048\,
            in2 => \_gnd_net_\,
            in3 => \N__21765\,
            lcout => \nx.n1277\,
            ltout => OPEN,
            carryin => \bfn_5_22_0_\,
            carryout => \nx.n10756\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_870_3_lut_LC_5_22_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__21762\,
            in3 => \N__21729\,
            lcout => \nx.n1276\,
            ltout => OPEN,
            carryin => \nx.n10756\,
            carryout => \nx.n10757\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_870_4_lut_LC_5_22_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42096\,
            in2 => \N__21726\,
            in3 => \N__21702\,
            lcout => \nx.n1275\,
            ltout => OPEN,
            carryin => \nx.n10757\,
            carryout => \nx.n10758\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_870_5_lut_LC_5_22_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42195\,
            in2 => \N__21699\,
            in3 => \N__21675\,
            lcout => \nx.n1274\,
            ltout => OPEN,
            carryin => \nx.n10758\,
            carryout => \nx.n10759\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_870_6_lut_LC_5_22_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42097\,
            in2 => \N__21672\,
            in3 => \N__22146\,
            lcout => \nx.n1273\,
            ltout => OPEN,
            carryin => \nx.n10759\,
            carryout => \nx.n10760\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_870_7_lut_LC_5_22_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42196\,
            in2 => \N__22143\,
            in3 => \N__22122\,
            lcout => \nx.n1272\,
            ltout => OPEN,
            carryin => \nx.n10760\,
            carryout => \nx.n10761\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_870_8_lut_LC_5_22_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42098\,
            in2 => \N__22118\,
            in3 => \N__22086\,
            lcout => \nx.n1271\,
            ltout => OPEN,
            carryin => \nx.n10761\,
            carryout => \nx.n10762\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_870_9_lut_LC_5_22_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42197\,
            in2 => \N__21999\,
            in3 => \N__22083\,
            lcout => \nx.n1270\,
            ltout => OPEN,
            carryin => \nx.n10762\,
            carryout => \nx.n10763\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_870_10_lut_LC_5_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000010001001000"
        )
    port map (
            in0 => \N__42198\,
            in1 => \N__21972\,
            in2 => \N__22080\,
            in3 => \N__22062\,
            lcout => \nx.n1301\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_2_lut_adj_157_LC_5_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22044\,
            in2 => \_gnd_net_\,
            in3 => \N__22026\,
            lcout => n4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i873_3_lut_LC_5_23_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21998\,
            in2 => \N__21982\,
            in3 => \N__21936\,
            lcout => \nx.n1302\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i21_4_lut_adj_140_LC_5_24_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__31778\,
            in1 => \N__23864\,
            in2 => \N__26082\,
            in3 => \N__38912\,
            lcout => OPEN,
            ltout => \nx.n49_adj_784_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i27_4_lut_LC_5_24_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__25434\,
            in1 => \N__22269\,
            in2 => \N__21915\,
            in3 => \N__21912\,
            lcout => \state_3_N_448_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i9167_2_lut_3_lut_LC_5_24_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010000000000"
        )
    port map (
            in0 => \N__43652\,
            in1 => \N__43947\,
            in2 => \_gnd_net_\,
            in3 => \N__47664\,
            lcout => n7664,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i2_2_lut_adj_132_LC_5_24_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__26353\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__25899\,
            lcout => OPEN,
            ltout => \nx.n30_adj_777_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i15_4_lut_adj_138_LC_5_24_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111000"
        )
    port map (
            in0 => \N__30791\,
            in1 => \N__32391\,
            in2 => \N__22272\,
            in3 => \N__23997\,
            lcout => \nx.n43_adj_783\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1138_2_lut_LC_5_25_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__23868\,
            in1 => \N__23867\,
            in2 => \N__22238\,
            in3 => \N__22263\,
            lcout => \nx.n1709\,
            ltout => OPEN,
            carryin => \bfn_5_25_0_\,
            carryout => \nx.n10794\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1138_3_lut_LC_5_25_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__22259\,
            in1 => \N__22258\,
            in2 => \N__22239\,
            in3 => \N__22221\,
            lcout => \nx.n1708\,
            ltout => OPEN,
            carryin => \nx.n10794\,
            carryout => \nx.n10795\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1138_4_lut_LC_5_25_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101000111010"
        )
    port map (
            in0 => \N__22218\,
            in1 => \N__22217\,
            in2 => \N__22385\,
            in3 => \N__22200\,
            lcout => \nx.n1707\,
            ltout => OPEN,
            carryin => \nx.n10795\,
            carryout => \nx.n10796\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1138_5_lut_LC_5_25_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101000111010"
        )
    port map (
            in0 => \N__22197\,
            in1 => \N__22196\,
            in2 => \N__22388\,
            in3 => \N__22179\,
            lcout => \nx.n1706\,
            ltout => OPEN,
            carryin => \nx.n10796\,
            carryout => \nx.n10797\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1138_6_lut_LC_5_25_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101000111010"
        )
    port map (
            in0 => \N__22176\,
            in1 => \N__22175\,
            in2 => \N__22386\,
            in3 => \N__22158\,
            lcout => \nx.n1705\,
            ltout => OPEN,
            carryin => \nx.n10797\,
            carryout => \nx.n10798\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1138_7_lut_LC_5_25_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101000111010"
        )
    port map (
            in0 => \N__22578\,
            in1 => \N__22577\,
            in2 => \N__22389\,
            in3 => \N__22560\,
            lcout => \nx.n1704\,
            ltout => OPEN,
            carryin => \nx.n10798\,
            carryout => \nx.n10799\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1138_8_lut_LC_5_25_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101000111010"
        )
    port map (
            in0 => \N__22557\,
            in1 => \N__22556\,
            in2 => \N__22387\,
            in3 => \N__22539\,
            lcout => \nx.n1703\,
            ltout => OPEN,
            carryin => \nx.n10799\,
            carryout => \nx.n10800\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1138_9_lut_LC_5_25_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101000111010"
        )
    port map (
            in0 => \N__22535\,
            in1 => \N__22534\,
            in2 => \N__22390\,
            in3 => \N__22515\,
            lcout => \nx.n1702\,
            ltout => OPEN,
            carryin => \nx.n10800\,
            carryout => \nx.n10801\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1138_10_lut_LC_5_26_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101000111010"
        )
    port map (
            in0 => \N__22511\,
            in1 => \N__22510\,
            in2 => \N__22391\,
            in3 => \N__22491\,
            lcout => \nx.n1701\,
            ltout => OPEN,
            carryin => \bfn_5_26_0_\,
            carryout => \nx.n10802\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1138_11_lut_LC_5_26_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101000111010"
        )
    port map (
            in0 => \N__22487\,
            in1 => \N__22488\,
            in2 => \N__22394\,
            in3 => \N__22467\,
            lcout => \nx.n1700\,
            ltout => OPEN,
            carryin => \nx.n10802\,
            carryout => \nx.n10803\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1138_12_lut_LC_5_26_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101000111010"
        )
    port map (
            in0 => \N__22464\,
            in1 => \N__22463\,
            in2 => \N__22392\,
            in3 => \N__22440\,
            lcout => \nx.n1699\,
            ltout => OPEN,
            carryin => \nx.n10803\,
            carryout => \nx.n10804\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1138_13_lut_LC_5_26_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101000111010"
        )
    port map (
            in0 => \N__22437\,
            in1 => \N__22436\,
            in2 => \N__22395\,
            in3 => \N__22419\,
            lcout => \nx.n1698\,
            ltout => OPEN,
            carryin => \nx.n10804\,
            carryout => \nx.n10805\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1138_14_lut_LC_5_26_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101000111010"
        )
    port map (
            in0 => \N__22414\,
            in1 => \N__22415\,
            in2 => \N__22393\,
            in3 => \N__22317\,
            lcout => \nx.n1697\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i7_3_lut_adj_130_LC_5_26_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22654\,
            in2 => \N__22606\,
            in3 => \N__22822\,
            lcout => \nx.n20_adj_775\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i3_3_lut_adj_119_LC_5_26_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110100000"
        )
    port map (
            in0 => \N__24743\,
            in1 => \_gnd_net_\,
            in2 => \N__22690\,
            in3 => \N__22630\,
            lcout => \nx.n16_adj_766\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1205_2_lut_LC_5_27_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__24764\,
            in1 => \N__24763\,
            in2 => \N__22913\,
            in3 => \N__22695\,
            lcout => \nx.n1809\,
            ltout => OPEN,
            carryin => \bfn_5_27_0_\,
            carryout => \nx.n10806\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1205_3_lut_LC_5_27_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__22692\,
            in1 => \N__22691\,
            in2 => \N__22914\,
            in3 => \N__22668\,
            lcout => \nx.n1808\,
            ltout => OPEN,
            carryin => \nx.n10806\,
            carryout => \nx.n10807\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1205_4_lut_LC_5_27_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101000111010"
        )
    port map (
            in0 => \N__22665\,
            in1 => \N__22661\,
            in2 => \N__22999\,
            in3 => \N__22641\,
            lcout => \nx.n1807\,
            ltout => OPEN,
            carryin => \nx.n10807\,
            carryout => \nx.n10808\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1205_5_lut_LC_5_27_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101000111010"
        )
    port map (
            in0 => \N__22638\,
            in1 => \N__22637\,
            in2 => \N__23002\,
            in3 => \N__22617\,
            lcout => \nx.n1806\,
            ltout => OPEN,
            carryin => \nx.n10808\,
            carryout => \nx.n10809\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1205_6_lut_LC_5_27_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101000111010"
        )
    port map (
            in0 => \N__22764\,
            in1 => \N__22763\,
            in2 => \N__23000\,
            in3 => \N__22614\,
            lcout => \nx.n1805\,
            ltout => OPEN,
            carryin => \nx.n10809\,
            carryout => \nx.n10810\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1205_7_lut_LC_5_27_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101000111010"
        )
    port map (
            in0 => \N__22742\,
            in1 => \N__22741\,
            in2 => \N__23003\,
            in3 => \N__22611\,
            lcout => \nx.n1804\,
            ltout => OPEN,
            carryin => \nx.n10810\,
            carryout => \nx.n10811\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1205_8_lut_LC_5_27_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101000111010"
        )
    port map (
            in0 => \N__22608\,
            in1 => \N__22607\,
            in2 => \N__23001\,
            in3 => \N__22584\,
            lcout => \nx.n1803\,
            ltout => OPEN,
            carryin => \nx.n10811\,
            carryout => \nx.n10812\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1205_9_lut_LC_5_27_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101000111010"
        )
    port map (
            in0 => \N__22794\,
            in1 => \N__22787\,
            in2 => \N__23004\,
            in3 => \N__22581\,
            lcout => \nx.n1802\,
            ltout => OPEN,
            carryin => \nx.n10812\,
            carryout => \nx.n10813\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1205_10_lut_LC_5_28_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101000111010"
        )
    port map (
            in0 => \N__23112\,
            in1 => \N__23111\,
            in2 => \N__22993\,
            in3 => \N__22833\,
            lcout => \nx.n1801\,
            ltout => OPEN,
            carryin => \bfn_5_28_0_\,
            carryout => \nx.n10814\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1205_11_lut_LC_5_28_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101000111010"
        )
    port map (
            in0 => \N__22830\,
            in1 => \N__22829\,
            in2 => \N__22996\,
            in3 => \N__22809\,
            lcout => \nx.n1800\,
            ltout => OPEN,
            carryin => \nx.n10814\,
            carryout => \nx.n10815\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1205_12_lut_LC_5_28_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101000111010"
        )
    port map (
            in0 => \N__22716\,
            in1 => \N__22715\,
            in2 => \N__22994\,
            in3 => \N__22806\,
            lcout => \nx.n1799\,
            ltout => OPEN,
            carryin => \nx.n10815\,
            carryout => \nx.n10816\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1205_13_lut_LC_5_28_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101000111010"
        )
    port map (
            in0 => \N__23064\,
            in1 => \N__23063\,
            in2 => \N__22997\,
            in3 => \N__22803\,
            lcout => \nx.n1798\,
            ltout => OPEN,
            carryin => \nx.n10816\,
            carryout => \nx.n10817\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1205_14_lut_LC_5_28_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101000111010"
        )
    port map (
            in0 => \N__23088\,
            in1 => \N__23087\,
            in2 => \N__22995\,
            in3 => \N__22800\,
            lcout => \nx.n1797\,
            ltout => OPEN,
            carryin => \nx.n10817\,
            carryout => \nx.n10818\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1205_15_lut_LC_5_28_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101000111010"
        )
    port map (
            in0 => \N__23042\,
            in1 => \N__23043\,
            in2 => \N__22998\,
            in3 => \N__22797\,
            lcout => \nx.n1796\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i4_2_lut_LC_5_28_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__24138\,
            in3 => \N__24157\,
            lcout => \nx.n18_adj_716\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i9_4_lut_adj_129_LC_5_29_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__22786\,
            in1 => \N__22762\,
            in2 => \N__22743\,
            in3 => \N__22714\,
            lcout => OPEN,
            ltout => \nx.n22_adj_774_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i11_4_lut_adj_131_LC_5_29_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__23121\,
            in1 => \N__23110\,
            in2 => \N__23091\,
            in3 => \N__23086\,
            lcout => OPEN,
            ltout => \nx.n24_adj_776_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i12_4_lut_adj_143_LC_5_29_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__23062\,
            in1 => \N__23041\,
            in2 => \N__23016\,
            in3 => \N__23013\,
            lcout => \nx.n1730\,
            ltout => \nx.n1730_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i9205_1_lut_LC_5_29_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__22917\,
            in3 => \_gnd_net_\,
            lcout => \nx.n13601\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i10_4_lut_adj_67_LC_5_29_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__24372\,
            in1 => \N__24345\,
            in2 => \N__24321\,
            in3 => \N__24286\,
            lcout => \nx.n24_adj_717\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i7635_2_lut_3_lut_4_lut_4_lut_LC_6_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101100000000"
        )
    port map (
            in0 => \N__42628\,
            in1 => \N__45671\,
            in2 => \N__44439\,
            in3 => \N__47624\,
            lcout => n11972,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i9118_3_lut_4_lut_LC_6_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__23261\,
            in1 => \N__23478\,
            in2 => \N__22881\,
            in3 => \N__23182\,
            lcout => \nx.n13514\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i9133_4_lut_LC_6_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101111110000000"
        )
    port map (
            in0 => \N__24941\,
            in1 => \N__23205\,
            in2 => \N__26804\,
            in3 => \N__22856\,
            lcout => \nx.n13513\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.equal_372_i8_2_lut_LC_6_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23260\,
            in2 => \_gnd_net_\,
            in3 => \N__24940\,
            lcout => \nx.n7598\,
            ltout => \nx.n7598_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i9095_3_lut_LC_6_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22857\,
            in2 => \N__22836\,
            in3 => \N__23181\,
            lcout => \nx.n13435\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i4_4_lut_4_lut_LC_6_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__23476\,
            in1 => \N__23142\,
            in2 => \N__26797\,
            in3 => \N__26854\,
            lcout => \nx.n10_adj_760\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.neo_pixel_transmitter_t0_i0_i26_LC_6_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__23304\,
            in1 => \N__23331\,
            in2 => \_gnd_net_\,
            in3 => \N__25238\,
            lcout => neo_pixel_transmitter_t0_26,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46862\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i8969_3_lut_LC_6_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__26174\,
            in1 => \N__25756\,
            in2 => \_gnd_net_\,
            in3 => \N__24984\,
            lcout => \nx.n13364\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i4191_3_lut_LC_6_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011100000000"
        )
    port map (
            in0 => \N__23477\,
            in1 => \N__26777\,
            in2 => \_gnd_net_\,
            in3 => \N__26708\,
            lcout => \nx.n7983\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.sub_14_inv_0_i27_1_lut_LC_6_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__23303\,
            lcout => \nx.n7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i5_3_lut_adj_142_LC_6_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010001000"
        )
    port map (
            in0 => \N__26798\,
            in1 => \N__23283\,
            in2 => \_gnd_net_\,
            in3 => \N__23127\,
            lcout => \nx.n7994\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \update_color_126_LC_6_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__25053\,
            in1 => \N__25788\,
            in2 => \N__23277\,
            in3 => \N__24996\,
            lcout => update_color,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46866\,
            ce => 'H',
            sr => \N__25047\
        );

    \nx.i9076_3_lut_4_lut_LC_6_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111110111111"
        )
    port map (
            in0 => \N__23262\,
            in1 => \N__23204\,
            in2 => \N__24956\,
            in3 => \N__23169\,
            lcout => OPEN,
            ltout => \nx.n13436_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i822_4_lut_LC_6_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111001011111010"
        )
    port map (
            in0 => \N__23474\,
            in1 => \N__23141\,
            in2 => \N__23130\,
            in3 => \N__26853\,
            lcout => \nx.n3901\,
            ltout => \nx.n3901_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i9173_4_lut_4_lut_LC_6_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101000011011"
        )
    port map (
            in0 => \N__26799\,
            in1 => \N__23475\,
            in2 => \N__23409\,
            in3 => \N__23406\,
            lcout => \nx.n7657\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_736_2_lut_LC_6_20_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23940\,
            in2 => \_gnd_net_\,
            in3 => \N__23391\,
            lcout => \nx.n1077\,
            ltout => OPEN,
            carryin => \bfn_6_20_0_\,
            carryout => \nx.n10743\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_736_3_lut_LC_6_20_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__23583\,
            in3 => \N__23379\,
            lcout => \nx.n1076\,
            ltout => OPEN,
            carryin => \nx.n10743\,
            carryout => \nx.n10744\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_736_4_lut_LC_6_20_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42217\,
            in2 => \N__25415\,
            in3 => \N__23376\,
            lcout => \nx.n1075\,
            ltout => OPEN,
            carryin => \nx.n10744\,
            carryout => \nx.n10745\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_736_5_lut_LC_6_20_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42093\,
            in2 => \N__23651\,
            in3 => \N__23367\,
            lcout => \nx.n1074\,
            ltout => OPEN,
            carryin => \nx.n10745\,
            carryout => \nx.n10746\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_736_6_lut_LC_6_20_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42218\,
            in2 => \N__25395\,
            in3 => \N__23364\,
            lcout => \nx.n1073\,
            ltout => OPEN,
            carryin => \nx.n10746\,
            carryout => \nx.n10747\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_736_7_lut_LC_6_20_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42094\,
            in2 => \N__23603\,
            in3 => \N__23355\,
            lcout => \nx.n1072\,
            ltout => OPEN,
            carryin => \nx.n10747\,
            carryout => \nx.n10748\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_736_8_lut_LC_6_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001000001100000"
        )
    port map (
            in0 => \N__42095\,
            in1 => \N__25614\,
            in2 => \N__23559\,
            in3 => \N__23352\,
            lcout => \nx.n1103\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i676_3_lut_LC_6_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25328\,
            in2 => \N__25284\,
            in3 => \N__25357\,
            lcout => \nx.n1009\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.sub_14_inv_0_i29_1_lut_LC_6_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__25068\,
            lcout => \nx.n5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i9195_2_lut_LC_6_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__25695\,
            in3 => \N__25365\,
            lcout => \nx.n1007\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i742_3_lut_LC_6_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23634\,
            in2 => \N__25416\,
            in3 => \N__23554\,
            lcout => \nx.n1107\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i672_3_lut_LC_6_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25641\,
            in2 => \N__25665\,
            in3 => \N__25366\,
            lcout => \nx.n1005\,
            ltout => \nx.n1005_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i2_3_lut_LC_6_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23950\,
            in2 => \N__23586\,
            in3 => \N__23581\,
            lcout => OPEN,
            ltout => \nx.n7_adj_690_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i4_4_lut_LC_6_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111011"
        )
    port map (
            in0 => \N__25610\,
            in1 => \N__25422\,
            in2 => \N__23562\,
            in3 => \N__25411\,
            lcout => \nx.n1037\,
            ltout => \nx.n1037_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i740_3_lut_LC_6_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101000001010"
        )
    port map (
            in0 => \N__25394\,
            in1 => \_gnd_net_\,
            in2 => \N__23526\,
            in3 => \N__23523\,
            lcout => \nx.n1105\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i8903_4_lut_LC_6_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011110010010110"
        )
    port map (
            in0 => \N__25938\,
            in1 => \N__25898\,
            in2 => \N__23751\,
            in3 => \N__25559\,
            lcout => \nx.n7899\,
            ltout => \nx.n7899_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i1_3_lut_4_lut_adj_144_LC_6_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000011100001011"
        )
    port map (
            in0 => \N__25560\,
            in1 => \N__25326\,
            in2 => \N__23754\,
            in3 => \N__25940\,
            lcout => \nx.n12839\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i1_3_lut_LC_6_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__25856\,
            in3 => \N__25830\,
            lcout => \nx.n740\,
            ltout => \nx.n740_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i8902_4_lut_LC_6_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001001101101100"
        )
    port map (
            in0 => \N__25897\,
            in1 => \N__25947\,
            in2 => \N__23742\,
            in3 => \N__26081\,
            lcout => \nx.n11866\,
            ltout => \nx.n11866_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i1_4_lut_LC_6_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000001010"
        )
    port map (
            in0 => \N__26088\,
            in1 => \_gnd_net_\,
            in2 => \N__23739\,
            in3 => \N__25594\,
            lcout => \nx.n838\,
            ltout => \nx.n838_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i1_2_lut_adj_43_LC_6_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__23736\,
            in3 => \N__25939\,
            lcout => \nx.n7497\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i12_3_lut_LC_6_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26025\,
            in2 => \N__25984\,
            in3 => \N__26069\,
            lcout => \nx.n708\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i5701_4_lut_LC_6_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100110010"
        )
    port map (
            in0 => \N__23733\,
            in1 => \N__23718\,
            in2 => \N__23697\,
            in3 => \N__23682\,
            lcout => n1907,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.bit_ctr__i0_LC_6_23_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26155\,
            in2 => \_gnd_net_\,
            in3 => \N__23670\,
            lcout => \nx.bit_ctr_0\,
            ltout => OPEN,
            carryin => \bfn_6_23_0_\,
            carryout => \nx.n10613\,
            clk => \N__46875\,
            ce => \N__24240\,
            sr => \N__24208\
        );

    \nx.bit_ctr__i1_LC_6_23_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24842\,
            in2 => \_gnd_net_\,
            in3 => \N__23667\,
            lcout => \nx.bit_ctr_1\,
            ltout => OPEN,
            carryin => \nx.n10613\,
            carryout => \nx.n10614\,
            clk => \N__46875\,
            ce => \N__24240\,
            sr => \N__24208\
        );

    \nx.bit_ctr__i2_LC_6_23_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26870\,
            in2 => \_gnd_net_\,
            in3 => \N__23784\,
            lcout => \nx.bit_ctr_2\,
            ltout => OPEN,
            carryin => \nx.n10614\,
            carryout => \nx.n10615\,
            clk => \N__46875\,
            ce => \N__24240\,
            sr => \N__24208\
        );

    \nx.bit_ctr__i3_LC_6_23_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30792\,
            in2 => \_gnd_net_\,
            in3 => \N__23781\,
            lcout => \nx.bit_ctr_3\,
            ltout => OPEN,
            carryin => \nx.n10615\,
            carryout => \nx.n10616\,
            clk => \N__46875\,
            ce => \N__24240\,
            sr => \N__24208\
        );

    \nx.bit_ctr__i4_LC_6_23_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32392\,
            in2 => \_gnd_net_\,
            in3 => \N__23778\,
            lcout => \nx.bit_ctr_4\,
            ltout => OPEN,
            carryin => \nx.n10616\,
            carryout => \nx.n10617\,
            clk => \N__46875\,
            ce => \N__24240\,
            sr => \N__24208\
        );

    \nx.bit_ctr__i5_LC_6_23_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29329\,
            in2 => \_gnd_net_\,
            in3 => \N__23775\,
            lcout => \nx.bit_ctr_5\,
            ltout => OPEN,
            carryin => \nx.n10617\,
            carryout => \nx.n10618\,
            clk => \N__46875\,
            ce => \N__24240\,
            sr => \N__24208\
        );

    \nx.bit_ctr__i6_LC_6_23_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35233\,
            in2 => \_gnd_net_\,
            in3 => \N__23772\,
            lcout => \nx.bit_ctr_6\,
            ltout => OPEN,
            carryin => \nx.n10618\,
            carryout => \nx.n10619\,
            clk => \N__46875\,
            ce => \N__24240\,
            sr => \N__24208\
        );

    \nx.bit_ctr__i7_LC_6_23_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28205\,
            in2 => \_gnd_net_\,
            in3 => \N__23769\,
            lcout => \nx.bit_ctr_7\,
            ltout => OPEN,
            carryin => \nx.n10619\,
            carryout => \nx.n10620\,
            clk => \N__46875\,
            ce => \N__24240\,
            sr => \N__24208\
        );

    \nx.bit_ctr__i8_LC_6_24_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30123\,
            in2 => \_gnd_net_\,
            in3 => \N__23766\,
            lcout => \nx.bit_ctr_8\,
            ltout => OPEN,
            carryin => \bfn_6_24_0_\,
            carryout => \nx.n10621\,
            clk => \N__46876\,
            ce => \N__24250\,
            sr => \N__24212\
        );

    \nx.bit_ctr__i9_LC_6_24_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38913\,
            in2 => \_gnd_net_\,
            in3 => \N__23763\,
            lcout => \nx.bit_ctr_9\,
            ltout => OPEN,
            carryin => \nx.n10621\,
            carryout => \nx.n10622\,
            clk => \N__46876\,
            ce => \N__24250\,
            sr => \N__24212\
        );

    \nx.bit_ctr__i10_LC_6_24_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39899\,
            in2 => \_gnd_net_\,
            in3 => \N__23760\,
            lcout => \nx.bit_ctr_10\,
            ltout => OPEN,
            carryin => \nx.n10622\,
            carryout => \nx.n10623\,
            clk => \N__46876\,
            ce => \N__24250\,
            sr => \N__24212\
        );

    \nx.bit_ctr__i11_LC_6_24_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36045\,
            in2 => \_gnd_net_\,
            in3 => \N__23757\,
            lcout => \nx.bit_ctr_11\,
            ltout => OPEN,
            carryin => \nx.n10623\,
            carryout => \nx.n10624\,
            clk => \N__46876\,
            ce => \N__24250\,
            sr => \N__24212\
        );

    \nx.bit_ctr__i12_LC_6_24_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34328\,
            in2 => \_gnd_net_\,
            in3 => \N__23889\,
            lcout => \nx.bit_ctr_12\,
            ltout => OPEN,
            carryin => \nx.n10624\,
            carryout => \nx.n10625\,
            clk => \N__46876\,
            ce => \N__24250\,
            sr => \N__24212\
        );

    \nx.bit_ctr__i13_LC_6_24_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31779\,
            in2 => \_gnd_net_\,
            in3 => \N__23886\,
            lcout => \nx.bit_ctr_13\,
            ltout => OPEN,
            carryin => \nx.n10625\,
            carryout => \nx.n10626\,
            clk => \N__46876\,
            ce => \N__24250\,
            sr => \N__24212\
        );

    \nx.bit_ctr__i14_LC_6_24_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30510\,
            in2 => \_gnd_net_\,
            in3 => \N__23883\,
            lcout => \nx.bit_ctr_14\,
            ltout => OPEN,
            carryin => \nx.n10626\,
            carryout => \nx.n10627\,
            clk => \N__46876\,
            ce => \N__24250\,
            sr => \N__24212\
        );

    \nx.bit_ctr__i15_LC_6_24_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28917\,
            in2 => \_gnd_net_\,
            in3 => \N__23880\,
            lcout => \nx.bit_ctr_15\,
            ltout => OPEN,
            carryin => \nx.n10627\,
            carryout => \nx.n10628\,
            clk => \N__46876\,
            ce => \N__24250\,
            sr => \N__24212\
        );

    \nx.bit_ctr__i16_LC_6_25_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26354\,
            in2 => \_gnd_net_\,
            in3 => \N__23877\,
            lcout => \nx.bit_ctr_16\,
            ltout => OPEN,
            carryin => \bfn_6_25_0_\,
            carryout => \nx.n10629\,
            clk => \N__46878\,
            ce => \N__24255\,
            sr => \N__24213\
        );

    \nx.bit_ctr__i17_LC_6_25_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25514\,
            in2 => \_gnd_net_\,
            in3 => \N__23874\,
            lcout => \nx.bit_ctr_17\,
            ltout => OPEN,
            carryin => \nx.n10629\,
            carryout => \nx.n10630\,
            clk => \N__46878\,
            ce => \N__24255\,
            sr => \N__24213\
        );

    \nx.bit_ctr__i18_LC_6_25_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24753\,
            in2 => \_gnd_net_\,
            in3 => \N__23871\,
            lcout => \nx.bit_ctr_18\,
            ltout => OPEN,
            carryin => \nx.n10630\,
            carryout => \nx.n10631\,
            clk => \N__46878\,
            ce => \N__24255\,
            sr => \N__24213\
        );

    \nx.bit_ctr__i19_LC_6_25_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23865\,
            in2 => \_gnd_net_\,
            in3 => \N__23832\,
            lcout => \nx.bit_ctr_19\,
            ltout => OPEN,
            carryin => \nx.n10631\,
            carryout => \nx.n10632\,
            clk => \N__46878\,
            ce => \N__24255\,
            sr => \N__24213\
        );

    \nx.bit_ctr__i20_LC_6_25_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23813\,
            in2 => \_gnd_net_\,
            in3 => \N__24108\,
            lcout => \nx.bit_ctr_20\,
            ltout => OPEN,
            carryin => \nx.n10632\,
            carryout => \nx.n10633\,
            clk => \N__46878\,
            ce => \N__24255\,
            sr => \N__24213\
        );

    \nx.bit_ctr__i21_LC_6_25_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24092\,
            in2 => \_gnd_net_\,
            in3 => \N__24060\,
            lcout => \nx.bit_ctr_21\,
            ltout => OPEN,
            carryin => \nx.n10633\,
            carryout => \nx.n10634\,
            clk => \N__46878\,
            ce => \N__24255\,
            sr => \N__24213\
        );

    \nx.bit_ctr__i22_LC_6_25_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25463\,
            in2 => \_gnd_net_\,
            in3 => \N__24057\,
            lcout => \nx.bit_ctr_22\,
            ltout => OPEN,
            carryin => \nx.n10634\,
            carryout => \nx.n10635\,
            clk => \N__46878\,
            ce => \N__24255\,
            sr => \N__24213\
        );

    \nx.bit_ctr__i23_LC_6_25_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24044\,
            in2 => \_gnd_net_\,
            in3 => \N__24003\,
            lcout => \nx.bit_ctr_23\,
            ltout => OPEN,
            carryin => \nx.n10635\,
            carryout => \nx.n10636\,
            clk => \N__46878\,
            ce => \N__24255\,
            sr => \N__24213\
        );

    \nx.bit_ctr__i24_LC_6_26_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23987\,
            in2 => \_gnd_net_\,
            in3 => \N__23955\,
            lcout => \nx.bit_ctr_24\,
            ltout => OPEN,
            carryin => \bfn_6_26_0_\,
            carryout => \nx.n10637\,
            clk => \N__46882\,
            ce => \N__24254\,
            sr => \N__24204\
        );

    \nx.bit_ctr__i25_LC_6_26_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23939\,
            in2 => \_gnd_net_\,
            in3 => \N__23901\,
            lcout => \nx.bit_ctr_25\,
            ltout => OPEN,
            carryin => \nx.n10637\,
            carryout => \nx.n10638\,
            clk => \N__46882\,
            ce => \N__24254\,
            sr => \N__24204\
        );

    \nx.bit_ctr__i26_LC_6_26_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25313\,
            in2 => \_gnd_net_\,
            in3 => \N__23898\,
            lcout => \nx.bit_ctr_26\,
            ltout => OPEN,
            carryin => \nx.n10638\,
            carryout => \nx.n10639\,
            clk => \N__46882\,
            ce => \N__24254\,
            sr => \N__24204\
        );

    \nx.bit_ctr__i27_LC_6_26_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25925\,
            in2 => \_gnd_net_\,
            in3 => \N__23895\,
            lcout => \nx.bit_ctr_27\,
            ltout => OPEN,
            carryin => \nx.n10639\,
            carryout => \nx.n10640\,
            clk => \N__46882\,
            ce => \N__24254\,
            sr => \N__24204\
        );

    \nx.bit_ctr__i28_LC_6_26_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25893\,
            in2 => \_gnd_net_\,
            in3 => \N__23892\,
            lcout => \nx.bit_ctr_28\,
            ltout => OPEN,
            carryin => \nx.n10640\,
            carryout => \nx.n10641\,
            clk => \N__46882\,
            ce => \N__24254\,
            sr => \N__24204\
        );

    \nx.bit_ctr__i29_LC_6_26_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26068\,
            in2 => \_gnd_net_\,
            in3 => \N__24264\,
            lcout => \nx.bit_ctr_29\,
            ltout => OPEN,
            carryin => \nx.n10641\,
            carryout => \nx.n10642\,
            clk => \N__46882\,
            ce => \N__24254\,
            sr => \N__24204\
        );

    \nx.bit_ctr__i30_LC_6_26_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26016\,
            in2 => \_gnd_net_\,
            in3 => \N__24261\,
            lcout => \nx.bit_ctr_30\,
            ltout => OPEN,
            carryin => \nx.n10642\,
            carryout => \nx.n10643\,
            clk => \N__46882\,
            ce => \N__24254\,
            sr => \N__24204\
        );

    \nx.bit_ctr__i31_LC_6_26_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25974\,
            in2 => \_gnd_net_\,
            in3 => \N__24258\,
            lcout => \nx.bit_ctr_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46882\,
            ce => \N__24254\,
            sr => \N__24204\
        );

    \nx.mod_5_add_1272_2_lut_LC_6_27_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__25524\,
            in1 => \N__25523\,
            in2 => \N__24416\,
            in3 => \N__24168\,
            lcout => \nx.n1909\,
            ltout => OPEN,
            carryin => \bfn_6_27_0_\,
            carryout => \nx.n10819\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1272_3_lut_LC_6_27_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__24602\,
            in1 => \N__24601\,
            in2 => \N__24417\,
            in3 => \N__24165\,
            lcout => \nx.n1908\,
            ltout => OPEN,
            carryin => \nx.n10819\,
            carryout => \nx.n10820\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1272_4_lut_LC_6_27_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101000111010"
        )
    port map (
            in0 => \N__24626\,
            in1 => \N__24625\,
            in2 => \N__24511\,
            in3 => \N__24162\,
            lcout => \nx.n1907\,
            ltout => OPEN,
            carryin => \nx.n10820\,
            carryout => \nx.n10821\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1272_5_lut_LC_6_27_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101000111010"
        )
    port map (
            in0 => \N__24159\,
            in1 => \N__24158\,
            in2 => \N__24514\,
            in3 => \N__24141\,
            lcout => \nx.n1906\,
            ltout => OPEN,
            carryin => \nx.n10821\,
            carryout => \nx.n10822\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1272_6_lut_LC_6_27_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101000111010"
        )
    port map (
            in0 => \N__24134\,
            in1 => \N__24133\,
            in2 => \N__24512\,
            in3 => \N__24114\,
            lcout => \nx.n1905\,
            ltout => OPEN,
            carryin => \nx.n10822\,
            carryout => \nx.n10823\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1272_7_lut_LC_6_27_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101000111010"
        )
    port map (
            in0 => \N__24674\,
            in1 => \N__24673\,
            in2 => \N__24515\,
            in3 => \N__24111\,
            lcout => \nx.n1904\,
            ltout => OPEN,
            carryin => \nx.n10823\,
            carryout => \nx.n10824\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1272_8_lut_LC_6_27_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101000111010"
        )
    port map (
            in0 => \N__24371\,
            in1 => \N__24370\,
            in2 => \N__24513\,
            in3 => \N__24351\,
            lcout => \nx.n1903\,
            ltout => OPEN,
            carryin => \nx.n10824\,
            carryout => \nx.n10825\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1272_9_lut_LC_6_27_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101000111010"
        )
    port map (
            in0 => \N__24581\,
            in1 => \N__24580\,
            in2 => \N__24516\,
            in3 => \N__24348\,
            lcout => \nx.n1902\,
            ltout => OPEN,
            carryin => \nx.n10825\,
            carryout => \nx.n10826\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1272_10_lut_LC_6_28_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101000111010"
        )
    port map (
            in0 => \N__24344\,
            in1 => \N__24343\,
            in2 => \N__24504\,
            in3 => \N__24324\,
            lcout => \nx.n1901\,
            ltout => OPEN,
            carryin => \bfn_6_28_0_\,
            carryout => \nx.n10827\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1272_11_lut_LC_6_28_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101000111010"
        )
    port map (
            in0 => \N__24320\,
            in1 => \N__24319\,
            in2 => \N__24508\,
            in3 => \N__24300\,
            lcout => \nx.n1900\,
            ltout => OPEN,
            carryin => \nx.n10827\,
            carryout => \nx.n10828\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1272_12_lut_LC_6_28_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101000111010"
        )
    port map (
            in0 => \N__24561\,
            in1 => \N__24560\,
            in2 => \N__24505\,
            in3 => \N__24297\,
            lcout => \nx.n1899\,
            ltout => OPEN,
            carryin => \nx.n10828\,
            carryout => \nx.n10829\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1272_13_lut_LC_6_28_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101000111010"
        )
    port map (
            in0 => \N__24696\,
            in1 => \N__24695\,
            in2 => \N__24509\,
            in3 => \N__24294\,
            lcout => \nx.n1898\,
            ltout => OPEN,
            carryin => \nx.n10829\,
            carryout => \nx.n10830\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1272_14_lut_LC_6_28_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101000111010"
        )
    port map (
            in0 => \N__24648\,
            in1 => \N__24647\,
            in2 => \N__24506\,
            in3 => \N__24291\,
            lcout => \nx.n1897\,
            ltout => OPEN,
            carryin => \nx.n10830\,
            carryout => \nx.n10831\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1272_15_lut_LC_6_28_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101000111010"
        )
    port map (
            in0 => \N__24288\,
            in1 => \N__24287\,
            in2 => \N__24510\,
            in3 => \N__24270\,
            lcout => \nx.n1896\,
            ltout => OPEN,
            carryin => \nx.n10831\,
            carryout => \nx.n10832\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1272_16_lut_LC_6_28_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101000111010"
        )
    port map (
            in0 => \N__24539\,
            in1 => \N__24540\,
            in2 => \N__24507\,
            in3 => \N__24267\,
            lcout => \nx.n1895\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i20_4_lut_adj_133_LC_6_29_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__25941\,
            in1 => \N__25978\,
            in2 => \N__24765\,
            in3 => \N__39921\,
            lcout => \nx.n48_adj_778\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i12_4_lut_adj_69_LC_6_29_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__24702\,
            in1 => \N__24694\,
            in2 => \N__24678\,
            in3 => \N__24654\,
            lcout => OPEN,
            ltout => \nx.n26_adj_719_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i13_4_lut_adj_70_LC_6_29_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__24640\,
            in1 => \N__24627\,
            in2 => \N__24606\,
            in3 => \N__24522\,
            lcout => \nx.n1829\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i5924_2_lut_LC_6_29_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010001000"
        )
    port map (
            in0 => \N__25515\,
            in1 => \N__24603\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => \nx.n9717_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i8_4_lut_adj_68_LC_6_29_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__24582\,
            in1 => \N__24559\,
            in2 => \N__24543\,
            in3 => \N__24538\,
            lcout => \nx.n22_adj_718\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i9209_1_lut_LC_6_29_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__24450\,
            lcout => \nx.n13605\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i7629_2_lut_3_lut_4_lut_4_lut_LC_7_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011001000"
        )
    port map (
            in0 => \N__44435\,
            in1 => \N__47519\,
            in2 => \N__45682\,
            in3 => \N__42627\,
            lcout => n11966,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pin_output_enable__i7_LC_7_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011100010101010"
        )
    port map (
            in0 => \N__24383\,
            in1 => \N__32424\,
            in2 => \N__47610\,
            in3 => \N__47153\,
            lcout => pin_oe_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46867\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.one_wire_108_LC_7_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__24955\,
            lcout => \NEOPXL_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46857\,
            ce => \N__24864\,
            sr => \N__24855\
        );

    \nx.i8968_3_lut_LC_7_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__26170\,
            in1 => \N__25025\,
            in2 => \_gnd_net_\,
            in3 => \N__26605\,
            lcout => \nx.n13363\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i1_2_lut_adj_107_LC_7_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30811\,
            in2 => \_gnd_net_\,
            in3 => \N__26565\,
            lcout => \nx.n11156\,
            ltout => \nx.n11156_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.bit_ctr_1__bdd_4_lut_LC_7_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101101010001010"
        )
    port map (
            in0 => \N__24846\,
            in1 => \N__24828\,
            in2 => \N__24822\,
            in3 => \N__24819\,
            lcout => OPEN,
            ltout => \nx.n13619_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.n13619_bdd_4_lut_LC_7_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001010"
        )
    port map (
            in0 => \N__24771\,
            in1 => \N__26139\,
            in2 => \N__24813\,
            in3 => \N__24810\,
            lcout => \nx.n13622\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pin_output_enable__i2_LC_7_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101100011001100"
        )
    port map (
            in0 => \N__24804\,
            in1 => \N__24782\,
            in2 => \N__47674\,
            in3 => \N__47157\,
            lcout => pin_oe_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46868\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i8977_3_lut_LC_7_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101000001010"
        )
    port map (
            in0 => \N__32221\,
            in1 => \_gnd_net_\,
            in2 => \N__26175\,
            in3 => \N__27289\,
            lcout => \nx.n13372\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i17_4_lut_adj_84_LC_7_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__33164\,
            in1 => \N__33131\,
            in2 => \N__32767\,
            in3 => \N__33092\,
            lcout => \nx.n44_adj_741\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i9204_1_lut_LC_7_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__29669\,
            lcout => \nx.n13600\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.neo_pixel_transmitter_t0_i0_i28_LC_7_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__25269\,
            in1 => \N__25067\,
            in2 => \_gnd_net_\,
            in3 => \N__25219\,
            lcout => neo_pixel_transmitter_t0_28,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46872\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_LC_7_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110111111110110"
        )
    port map (
            in0 => \N__32222\,
            in1 => \N__24990\,
            in2 => \N__24983\,
            in3 => \N__25032\,
            lcout => n9_adj_847,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \neopxl_color_prev_i13_LC_7_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__25024\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => neopxl_color_prev_13,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46873\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \neopxl_color_i13_LC_7_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111011100010000"
        )
    port map (
            in0 => \N__47516\,
            in1 => \N__43894\,
            in2 => \N__43692\,
            in3 => \N__25023\,
            lcout => neopxl_color_13,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46873\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i9171_2_lut_3_lut_LC_7_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__43893\,
            in1 => \N__47515\,
            in2 => \_gnd_net_\,
            in3 => \N__43676\,
            lcout => \current_pin_7__N_153\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \neopxl_color_prev_i14_LC_7_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__24979\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => neopxl_color_prev_14,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46873\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i3_4_lut_LC_7_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110111111110110"
        )
    port map (
            in0 => \N__27027\,
            in1 => \N__27294\,
            in2 => \N__25026\,
            in3 => \N__25002\,
            lcout => n11_adj_845,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \neopxl_color_prev_i4_LC_7_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__32223\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => neopxl_color_prev_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46873\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \neopxl_color_i14_LC_7_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110101001100"
        )
    port map (
            in0 => \N__43895\,
            in1 => \N__24978\,
            in2 => \N__47631\,
            in3 => \N__43680\,
            lcout => neopxl_color_14,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46873\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i7605_3_lut_LC_7_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25694\,
            in2 => \N__25368\,
            in3 => \N__25677\,
            lcout => \nx.n11941\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i675_3_lut_LC_7_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25713\,
            in2 => \N__25731\,
            in3 => \N__25358\,
            lcout => \nx.n1008\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i9197_2_lut_LC_7_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__25367\,
            in3 => \N__25676\,
            lcout => \nx.n1006\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i1_2_lut_adj_25_LC_7_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110011111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25580\,
            in2 => \N__25599\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => \nx.n12837_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i604_4_lut_LC_7_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000101"
        )
    port map (
            in0 => \N__25563\,
            in1 => \_gnd_net_\,
            in2 => \N__25380\,
            in3 => \N__25807\,
            lcout => \nx.n905\,
            ltout => \nx.n905_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i1_4_lut_adj_44_LC_7_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000000"
        )
    port map (
            in0 => \N__25535\,
            in1 => \N__25657\,
            in2 => \N__25377\,
            in3 => \N__25374\,
            lcout => \nx.n11174\,
            ltout => \nx.n11174_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i9198_1_lut_LC_7_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__25335\,
            in3 => \_gnd_net_\,
            lcout => \nx.n13594\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i605_4_lut_LC_7_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010101001"
        )
    port map (
            in0 => \N__25595\,
            in1 => \N__25579\,
            in2 => \N__25809\,
            in3 => \N__25562\,
            lcout => \nx.n906\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_669_2_lut_LC_7_22_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25327\,
            in2 => \_gnd_net_\,
            in3 => \N__25272\,
            lcout => \nx.n977\,
            ltout => OPEN,
            carryin => \bfn_7_22_0_\,
            carryout => \nx.n10738\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_669_3_lut_LC_7_22_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__25730\,
            in3 => \N__25707\,
            lcout => \nx.n976\,
            ltout => OPEN,
            carryin => \nx.n10738\,
            carryout => \nx.n10739\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_669_4_lut_LC_7_22_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41616\,
            in2 => \N__25704\,
            in3 => \N__25680\,
            lcout => \nx.n975\,
            ltout => OPEN,
            carryin => \nx.n10739\,
            carryout => \nx.n10740\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_669_5_lut_LC_7_22_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41619\,
            in2 => \N__25539\,
            in3 => \N__25668\,
            lcout => \nx.n974\,
            ltout => OPEN,
            carryin => \nx.n10740\,
            carryout => \nx.n10741\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_669_6_lut_LC_7_22_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41617\,
            in2 => \N__25664\,
            in3 => \N__25635\,
            lcout => \nx.n973\,
            ltout => OPEN,
            carryin => \nx.n10741\,
            carryout => \nx.n10742\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_669_7_lut_LC_7_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000010001001000"
        )
    port map (
            in0 => \N__41618\,
            in1 => \N__25632\,
            in2 => \N__25626\,
            in3 => \N__25617\,
            lcout => \nx.n4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i538_3_lut_2_lut_LC_7_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__25855\,
            in3 => \N__25827\,
            lcout => \nx.n807\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i9153_3_lut_LC_7_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011000011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25808\,
            in2 => \N__25581\,
            in3 => \N__25561\,
            lcout => \nx.n11868\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i16_4_lut_adj_137_LC_7_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__35232\,
            in1 => \N__25522\,
            in2 => \N__25481\,
            in3 => \N__29328\,
            lcout => \nx.n44_adj_782\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i1665_3_lut_4_lut_LC_7_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000001000"
        )
    port map (
            in0 => \N__25894\,
            in1 => \N__26073\,
            in2 => \N__26033\,
            in3 => \N__25985\,
            lcout => \nx.n11912\,
            ltout => \nx.n11912_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i5757_2_lut_3_lut_4_lut_LC_7_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110111010111"
        )
    port map (
            in0 => \N__25926\,
            in1 => \N__25895\,
            in2 => \N__26091\,
            in3 => \N__25828\,
            lcout => \nx.n58\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i6008_2_lut_4_lut_3_lut_LC_7_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011100000111000"
        )
    port map (
            in0 => \N__26074\,
            in1 => \N__26029\,
            in2 => \N__25989\,
            in3 => \_gnd_net_\,
            lcout => \nx.n9803\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i20_4_lut_adj_87_LC_7_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__32975\,
            in1 => \N__33293\,
            in2 => \N__32847\,
            in3 => \N__32891\,
            lcout => \nx.n47\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i1940_2_lut_3_lut_4_lut_LC_7_23_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000101000"
        )
    port map (
            in0 => \N__25927\,
            in1 => \N__25896\,
            in2 => \N__25857\,
            in3 => \N__25829\,
            lcout => \nx.n5703\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i2_4_lut_adj_170_LC_7_24_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110111111110110"
        )
    port map (
            in0 => \N__25776\,
            in1 => \N__26127\,
            in2 => \N__25770\,
            in3 => \N__25737\,
            lcout => n10_adj_846,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \neopxl_color_prev_i7_LC_7_24_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__26129\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => neopxl_color_prev_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46879\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \neopxl_color_prev_i15_LC_7_24_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__25769\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => neopxl_color_prev_15,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46879\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_2_lut_3_lut_LC_7_24_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010001000"
        )
    port map (
            in0 => \N__26128\,
            in1 => \N__43897\,
            in2 => \_gnd_net_\,
            in3 => \N__47518\,
            lcout => n22_adj_793,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i8978_3_lut_LC_7_24_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__26126\,
            in1 => \N__26208\,
            in2 => \_gnd_net_\,
            in3 => \N__26161\,
            lcout => \nx.n13373\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_2_lut_3_lut_adj_191_LC_7_24_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010001000"
        )
    port map (
            in0 => \N__27293\,
            in1 => \N__43892\,
            in2 => \_gnd_net_\,
            in3 => \N__47514\,
            lcout => n22,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_2_lut_3_lut_adj_194_LC_7_24_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010001000"
        )
    port map (
            in0 => \N__32220\,
            in1 => \N__43896\,
            in2 => \_gnd_net_\,
            in3 => \N__47517\,
            lcout => n22_adj_787,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \neopxl_color_i7_LC_7_25_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0000111100001000"
        )
    port map (
            in0 => \N__47539\,
            in1 => \N__43898\,
            in2 => \N__43715\,
            in3 => \N__26130\,
            lcout => neopxl_color_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46883\,
            ce => 'H',
            sr => \N__26109\
        );

    \nx.i5_3_lut_LC_7_25_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26348\,
            in2 => \N__26313\,
            in3 => \N__26653\,
            lcout => \nx.n20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1356_3_lut_LC_7_25_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__26349\,
            in1 => \N__26325\,
            in2 => \_gnd_net_\,
            in3 => \N__27543\,
            lcout => \nx.n2009\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i1_2_lut_adj_27_LC_7_26_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__26505\,
            in3 => \N__26543\,
            lcout => \nx.n16_adj_678\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i11_4_lut_adj_26_LC_7_26_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__27127\,
            in1 => \N__26248\,
            in2 => \N__27089\,
            in3 => \N__26275\,
            lcout => OPEN,
            ltout => \nx.n26_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i13_4_lut_adj_28_LC_7_26_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__27601\,
            in1 => \N__27355\,
            in2 => \N__26100\,
            in3 => \N__26097\,
            lcout => OPEN,
            ltout => \nx.n28_adj_679_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i14_4_lut_adj_29_LC_7_26_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__26416\,
            in1 => \N__26523\,
            in2 => \N__26367\,
            in3 => \N__26364\,
            lcout => \nx.n1928\,
            ltout => \nx.n1928_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1354_3_lut_LC_7_26_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101000001010"
        )
    port map (
            in0 => \N__26276\,
            in1 => \_gnd_net_\,
            in2 => \N__26358\,
            in3 => \N__26259\,
            lcout => \nx.n2007\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1352_3_lut_LC_7_26_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101000001010"
        )
    port map (
            in0 => \N__26417\,
            in1 => \_gnd_net_\,
            in2 => \N__27545\,
            in3 => \N__26400\,
            lcout => \nx.n2005\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1353_3_lut_LC_7_26_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010101010"
        )
    port map (
            in0 => \N__26249\,
            in1 => \_gnd_net_\,
            in2 => \N__26232\,
            in3 => \N__27518\,
            lcout => \nx.n2006\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1355_3_lut_LC_7_26_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101011001010"
        )
    port map (
            in0 => \N__26308\,
            in1 => \N__26286\,
            in2 => \N__27544\,
            in3 => \_gnd_net_\,
            lcout => \nx.n2008\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1339_2_lut_LC_7_27_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26355\,
            in2 => \_gnd_net_\,
            in3 => \N__26316\,
            lcout => \nx.n1977\,
            ltout => OPEN,
            carryin => \bfn_7_27_0_\,
            carryout => \nx.n10833\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1339_3_lut_LC_7_27_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__26309\,
            in3 => \N__26280\,
            lcout => \nx.n1976\,
            ltout => OPEN,
            carryin => \nx.n10833\,
            carryout => \nx.n10834\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1339_4_lut_LC_7_27_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41627\,
            in2 => \N__26277\,
            in3 => \N__26253\,
            lcout => \nx.n1975\,
            ltout => OPEN,
            carryin => \nx.n10834\,
            carryout => \nx.n10835\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1339_5_lut_LC_7_27_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41630\,
            in2 => \N__26250\,
            in3 => \N__26223\,
            lcout => \nx.n1974\,
            ltout => OPEN,
            carryin => \nx.n10835\,
            carryout => \nx.n10836\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1339_6_lut_LC_7_27_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41628\,
            in2 => \N__26418\,
            in3 => \N__26394\,
            lcout => \nx.n1973\,
            ltout => OPEN,
            carryin => \nx.n10836\,
            carryout => \nx.n10837\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1339_7_lut_LC_7_27_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41631\,
            in2 => \N__27088\,
            in3 => \N__26391\,
            lcout => \nx.n1972\,
            ltout => OPEN,
            carryin => \nx.n10837\,
            carryout => \nx.n10838\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1339_8_lut_LC_7_27_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41629\,
            in2 => \N__26654\,
            in3 => \N__26388\,
            lcout => \nx.n1971\,
            ltout => OPEN,
            carryin => \nx.n10838\,
            carryout => \nx.n10839\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1339_9_lut_LC_7_27_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41632\,
            in2 => \N__27131\,
            in3 => \N__26385\,
            lcout => \nx.n1970\,
            ltout => OPEN,
            carryin => \nx.n10839\,
            carryout => \nx.n10840\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1339_10_lut_LC_7_28_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42201\,
            in2 => \N__27605\,
            in3 => \N__26382\,
            lcout => \nx.n1969\,
            ltout => OPEN,
            carryin => \bfn_7_28_0_\,
            carryout => \nx.n10841\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1339_11_lut_LC_7_28_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42205\,
            in2 => \N__27356\,
            in3 => \N__26379\,
            lcout => \nx.n1968\,
            ltout => OPEN,
            carryin => \nx.n10841\,
            carryout => \nx.n10842\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1339_12_lut_LC_7_28_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42202\,
            in2 => \N__27170\,
            in3 => \N__26376\,
            lcout => \nx.n1967\,
            ltout => OPEN,
            carryin => \nx.n10842\,
            carryout => \nx.n10843\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1339_13_lut_LC_7_28_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42206\,
            in2 => \N__27212\,
            in3 => \N__26373\,
            lcout => \nx.n1966\,
            ltout => OPEN,
            carryin => \nx.n10843\,
            carryout => \nx.n10844\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1339_14_lut_LC_7_28_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42203\,
            in2 => \N__26468\,
            in3 => \N__26370\,
            lcout => \nx.n1965\,
            ltout => OPEN,
            carryin => \nx.n10844\,
            carryout => \nx.n10845\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1339_15_lut_LC_7_28_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42207\,
            in2 => \N__26436\,
            in3 => \N__26550\,
            lcout => \nx.n1964\,
            ltout => OPEN,
            carryin => \nx.n10845\,
            carryout => \nx.n10846\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1339_16_lut_LC_7_28_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42204\,
            in2 => \N__26504\,
            in3 => \N__26547\,
            lcout => \nx.n1963\,
            ltout => OPEN,
            carryin => \nx.n10846\,
            carryout => \nx.n10847\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1339_17_lut_LC_7_28_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__27552\,
            in1 => \N__42208\,
            in2 => \N__26544\,
            in3 => \N__26526\,
            lcout => \nx.n1994\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i9_4_lut_LC_7_29_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__27163\,
            in1 => \N__27205\,
            in2 => \N__26467\,
            in3 => \N__26431\,
            lcout => \nx.n24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1342_3_lut_LC_7_29_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27551\,
            in2 => \N__26514\,
            in3 => \N__26500\,
            lcout => \nx.n1995\,
            ltout => \nx.n1995_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i9_4_lut_adj_33_LC_7_29_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__28964\,
            in1 => \N__29143\,
            in2 => \N__26478\,
            in3 => \N__27407\,
            lcout => \nx.n25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1344_3_lut_LC_7_29_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26475\,
            in2 => \N__26469\,
            in3 => \N__27546\,
            lcout => \nx.n1997\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1343_3_lut_LC_7_29_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110010101100"
        )
    port map (
            in0 => \N__26442\,
            in1 => \N__26432\,
            in2 => \N__27567\,
            in3 => \_gnd_net_\,
            lcout => \nx.n1996\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1350_3_lut_LC_7_29_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26667\,
            in2 => \N__26658\,
            in3 => \N__27550\,
            lcout => \nx.n2003\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i8965_4_lut_LC_7_31_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101000100010"
        )
    port map (
            in0 => \N__27884\,
            in1 => \N__27815\,
            in2 => \N__27843\,
            in3 => \N__27863\,
            lcout => n13360,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i8966_4_lut_LC_7_31_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011000100"
        )
    port map (
            in0 => \N__27864\,
            in1 => \N__27842\,
            in2 => \N__27819\,
            in3 => \N__27885\,
            lcout => OPEN,
            ltout => \n13361_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i8967_3_lut_LC_7_31_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111101010101"
        )
    port map (
            in0 => \N__26628\,
            in1 => \_gnd_net_\,
            in2 => \N__26622\,
            in3 => \N__27789\,
            lcout => \LED_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i1_4_lut_adj_103_LC_9_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101100"
        )
    port map (
            in0 => \N__33483\,
            in1 => \N__33516\,
            in2 => \N__34024\,
            in3 => \N__27924\,
            lcout => \nx.n12817\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \neopxl_color_i12_LC_9_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111011100010000"
        )
    port map (
            in0 => \N__47598\,
            in1 => \N__43932\,
            in2 => \N__43691\,
            in3 => \N__26596\,
            lcout => neopxl_color_12,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46869\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i2147_3_lut_LC_9_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34131\,
            in2 => \N__34025\,
            in3 => \N__34098\,
            lcout => \nx.n59\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i9112_3_lut_LC_9_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__30815\,
            in1 => \N__30747\,
            in2 => \_gnd_net_\,
            in3 => \N__26564\,
            lcout => \nx.color_bit_N_642_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i2146_3_lut_LC_9_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34047\,
            in2 => \N__34032\,
            in3 => \N__34080\,
            lcout => OPEN,
            ltout => \nx.n61_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i1_4_lut_adj_106_LC_9_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__26574\,
            in1 => \N__33861\,
            in2 => \N__26568\,
            in3 => \N__26676\,
            lcout => \nx.n11153\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.state_i0_LC_9_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0000001000000000"
        )
    port map (
            in0 => \N__26880\,
            in1 => \N__26859\,
            in2 => \N__26823\,
            in3 => \N__26814\,
            lcout => state_0_adj_792,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46874\,
            ce => \N__26715\,
            sr => \N__26697\
        );

    \nx.i1_4_lut_adj_104_LC_9_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101111111000"
        )
    port map (
            in0 => \N__33432\,
            in1 => \N__34027\,
            in2 => \N__26688\,
            in3 => \N__33468\,
            lcout => OPEN,
            ltout => \nx.n12819_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i1_4_lut_adj_105_LC_9_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110111111000"
        )
    port map (
            in0 => \N__34028\,
            in1 => \N__33387\,
            in2 => \N__26679\,
            in3 => \N__33417\,
            lcout => \nx.n12821\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i2036_3_lut_LC_9_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__35205\,
            in1 => \N__35259\,
            in2 => \_gnd_net_\,
            in3 => \N__37321\,
            lcout => \nx.n3009\,
            ltout => \nx.n3009_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i13_3_lut_LC_9_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29338\,
            in2 => \N__26670\,
            in3 => \N__29227\,
            lcout => \nx.n39_adj_671\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1967_3_lut_LC_9_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28233\,
            in2 => \N__26910\,
            in3 => \N__37517\,
            lcout => \nx.n2908\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1966_3_lut_LC_9_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26895\,
            in2 => \N__37564\,
            in3 => \N__28082\,
            lcout => \nx.n2907\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i14_4_lut_adj_66_LC_9_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__37766\,
            in1 => \N__27046\,
            in2 => \N__27974\,
            in3 => \N__26981\,
            lcout => \nx.n38_adj_713\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i17_4_lut_adj_117_LC_9_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__37339\,
            in1 => \N__35449\,
            in2 => \N__35517\,
            in3 => \N__35401\,
            lcout => \nx.n42_adj_765\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1899_3_lut_LC_9_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011110000"
        )
    port map (
            in0 => \N__28278\,
            in1 => \_gnd_net_\,
            in2 => \N__30009\,
            in3 => \N__31270\,
            lcout => \nx.n2808\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1950_3_lut_LC_9_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101011001010"
        )
    port map (
            in0 => \N__27047\,
            in1 => \N__27000\,
            in2 => \N__37595\,
            in3 => \_gnd_net_\,
            lcout => \nx.n2891\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1947_3_lut_LC_9_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26955\,
            in2 => \N__28344\,
            in3 => \N__37556\,
            lcout => \nx.n2888\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1882_3_lut_LC_9_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31574\,
            in2 => \N__31278\,
            in3 => \N__28458\,
            lcout => \nx.n2791\,
            ltout => \nx.n2791_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1949_3_lut_LC_9_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26970\,
            in2 => \N__26916\,
            in3 => \N__37560\,
            lcout => \nx.n2890\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1942_2_lut_LC_9_21_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28206\,
            in2 => \_gnd_net_\,
            in3 => \N__26913\,
            lcout => \nx.n2877\,
            ltout => OPEN,
            carryin => \bfn_9_21_0_\,
            carryout => \nx.n11004\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1942_3_lut_LC_9_21_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28229\,
            in2 => \_gnd_net_\,
            in3 => \N__26898\,
            lcout => \nx.n2876\,
            ltout => OPEN,
            carryin => \nx.n11004\,
            carryout => \nx.n11005\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1942_4_lut_LC_9_21_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41742\,
            in2 => \N__28083\,
            in3 => \N__26886\,
            lcout => \nx.n2875\,
            ltout => OPEN,
            carryin => \nx.n11005\,
            carryout => \nx.n11006\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1942_5_lut_LC_9_21_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41745\,
            in2 => \N__28031\,
            in3 => \N__26883\,
            lcout => \nx.n2874\,
            ltout => OPEN,
            carryin => \nx.n11006\,
            carryout => \nx.n11007\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1942_6_lut_LC_9_21_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41743\,
            in2 => \N__34817\,
            in3 => \N__26943\,
            lcout => \nx.n2873\,
            ltout => OPEN,
            carryin => \nx.n11007\,
            carryout => \nx.n11008\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1942_7_lut_LC_9_21_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41746\,
            in2 => \N__33844\,
            in3 => \N__26940\,
            lcout => \nx.n2872\,
            ltout => OPEN,
            carryin => \nx.n11008\,
            carryout => \nx.n11009\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1942_8_lut_LC_9_21_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41744\,
            in2 => \N__36845\,
            in3 => \N__26937\,
            lcout => \nx.n2871\,
            ltout => OPEN,
            carryin => \nx.n11009\,
            carryout => \nx.n11010\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1942_9_lut_LC_9_21_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41747\,
            in2 => \N__34172\,
            in3 => \N__26934\,
            lcout => \nx.n2870\,
            ltout => OPEN,
            carryin => \nx.n11010\,
            carryout => \nx.n11011\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1942_10_lut_LC_9_22_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41935\,
            in2 => \N__28161\,
            in3 => \N__26931\,
            lcout => \nx.n2869\,
            ltout => OPEN,
            carryin => \bfn_9_22_0_\,
            carryout => \nx.n11012\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1942_11_lut_LC_9_22_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41811\,
            in2 => \N__28108\,
            in3 => \N__26928\,
            lcout => \nx.n2868\,
            ltout => OPEN,
            carryin => \nx.n11012\,
            carryout => \nx.n11013\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1942_12_lut_LC_9_22_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41936\,
            in2 => \N__29774\,
            in3 => \N__26925\,
            lcout => \nx.n2867\,
            ltout => OPEN,
            carryin => \nx.n11013\,
            carryout => \nx.n11014\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1942_13_lut_LC_9_22_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41812\,
            in2 => \N__31440\,
            in3 => \N__26922\,
            lcout => \nx.n2866\,
            ltout => OPEN,
            carryin => \nx.n11014\,
            carryout => \nx.n11015\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1942_14_lut_LC_9_22_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41937\,
            in2 => \N__33804\,
            in3 => \N__26919\,
            lcout => \nx.n2865\,
            ltout => OPEN,
            carryin => \nx.n11015\,
            carryout => \nx.n11016\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1942_15_lut_LC_9_22_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41813\,
            in2 => \N__34882\,
            in3 => \N__27015\,
            lcout => \nx.n2864\,
            ltout => OPEN,
            carryin => \nx.n11016\,
            carryout => \nx.n11017\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1942_16_lut_LC_9_22_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41938\,
            in2 => \N__31143\,
            in3 => \N__27012\,
            lcout => \nx.n2863\,
            ltout => OPEN,
            carryin => \nx.n11017\,
            carryout => \nx.n11018\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1942_17_lut_LC_9_22_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41814\,
            in2 => \N__28136\,
            in3 => \N__27009\,
            lcout => \nx.n2862\,
            ltout => OPEN,
            carryin => \nx.n11018\,
            carryout => \nx.n11019\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1942_18_lut_LC_9_23_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41939\,
            in2 => \N__37654\,
            in3 => \N__27006\,
            lcout => \nx.n2861\,
            ltout => OPEN,
            carryin => \bfn_9_23_0_\,
            carryout => \nx.n11020\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1942_19_lut_LC_9_23_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37762\,
            in2 => \N__42187\,
            in3 => \N__27003\,
            lcout => \nx.n2860\,
            ltout => OPEN,
            carryin => \nx.n11020\,
            carryout => \nx.n11021\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1942_20_lut_LC_9_23_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41943\,
            in2 => \N__27048\,
            in3 => \N__26991\,
            lcout => \nx.n2859\,
            ltout => OPEN,
            carryin => \nx.n11021\,
            carryout => \nx.n11022\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1942_21_lut_LC_9_23_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41805\,
            in2 => \N__26988\,
            in3 => \N__26961\,
            lcout => \nx.n2858\,
            ltout => OPEN,
            carryin => \nx.n11022\,
            carryout => \nx.n11023\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1942_22_lut_LC_9_23_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41944\,
            in2 => \N__27970\,
            in3 => \N__26958\,
            lcout => \nx.n2857\,
            ltout => OPEN,
            carryin => \nx.n11023\,
            carryout => \nx.n11024\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1942_23_lut_LC_9_23_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41806\,
            in2 => \N__28340\,
            in3 => \N__26946\,
            lcout => \nx.n2856\,
            ltout => OPEN,
            carryin => \nx.n11024\,
            carryout => \nx.n11025\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1942_24_lut_LC_9_23_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31331\,
            in2 => \N__42071\,
            in3 => \N__27057\,
            lcout => \nx.n2855\,
            ltout => OPEN,
            carryin => \nx.n11025\,
            carryout => \nx.n11026\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1942_25_lut_LC_9_23_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41810\,
            in2 => \N__29946\,
            in3 => \N__27054\,
            lcout => \nx.n2854\,
            ltout => OPEN,
            carryin => \nx.n11026\,
            carryout => \nx.n11027\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1942_26_lut_LC_9_24_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000010001001000"
        )
    port map (
            in0 => \N__42060\,
            in1 => \N__37596\,
            in2 => \N__28608\,
            in3 => \N__27051\,
            lcout => \nx.n2885\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1885_3_lut_LC_9_24_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31667\,
            in2 => \N__28488\,
            in3 => \N__31269\,
            lcout => \nx.n2794\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1892_3_lut_LC_9_24_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28380\,
            in2 => \N__31277\,
            in3 => \N__34209\,
            lcout => \nx.n2801\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1880_3_lut_LC_9_24_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31268\,
            in2 => \N__31611\,
            in3 => \N__28434\,
            lcout => \nx.n2789\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1881_3_lut_LC_9_24_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31637\,
            in2 => \N__31276\,
            in3 => \N__28443\,
            lcout => \nx.n2790\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1883_3_lut_LC_9_24_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31261\,
            in2 => \N__30087\,
            in3 => \N__28467\,
            lcout => \nx.n2792\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \neopxl_color_prev_i5_LC_9_24_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__27271\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => neopxl_color_prev_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46886\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1884_3_lut_LC_9_24_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31260\,
            in2 => \N__30066\,
            in3 => \N__28476\,
            lcout => \nx.n2793\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \neopxl_color_i5_LC_9_25_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0011001100100000"
        )
    port map (
            in0 => \N__43951\,
            in1 => \N__43716\,
            in2 => \N__47696\,
            in3 => \N__27270\,
            lcout => neopxl_color_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46891\,
            ce => 'H',
            sr => \N__27243\
        );

    \nx.mod_5_i1345_3_lut_LC_9_25_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27228\,
            in2 => \N__27582\,
            in3 => \N__27216\,
            lcout => \nx.n1998\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1346_3_lut_LC_9_25_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27189\,
            in2 => \N__27177\,
            in3 => \N__27576\,
            lcout => \nx.n1999\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1349_3_lut_LC_9_25_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27147\,
            in2 => \N__27581\,
            in3 => \N__27135\,
            lcout => \nx.n2002\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1351_3_lut_LC_9_25_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27108\,
            in2 => \N__27096\,
            in3 => \N__27572\,
            lcout => \nx.n2004\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1547_3_lut_LC_9_25_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30213\,
            in2 => \N__32304\,
            in3 => \N__32579\,
            lcout => \nx.n2296\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1406_2_lut_LC_9_26_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28929\,
            in2 => \_gnd_net_\,
            in3 => \N__27063\,
            lcout => \nx.n2077\,
            ltout => OPEN,
            carryin => \bfn_9_26_0_\,
            carryout => \nx.n10848\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1406_3_lut_LC_9_26_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__29204\,
            in3 => \N__27060\,
            lcout => \nx.n2076\,
            ltout => OPEN,
            carryin => \nx.n10848\,
            carryout => \nx.n10849\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1406_4_lut_LC_9_26_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42086\,
            in2 => \N__29020\,
            in3 => \N__27321\,
            lcout => \nx.n2075\,
            ltout => OPEN,
            carryin => \nx.n10849\,
            carryout => \nx.n10850\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1406_5_lut_LC_9_26_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42061\,
            in2 => \N__28869\,
            in3 => \N__27318\,
            lcout => \nx.n2074\,
            ltout => OPEN,
            carryin => \nx.n10850\,
            carryout => \nx.n10851\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1406_6_lut_LC_9_26_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42087\,
            in2 => \N__28711\,
            in3 => \N__27315\,
            lcout => \nx.n2073\,
            ltout => OPEN,
            carryin => \nx.n10851\,
            carryout => \nx.n10852\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1406_7_lut_LC_9_26_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42062\,
            in2 => \N__28679\,
            in3 => \N__27312\,
            lcout => \nx.n2072\,
            ltout => OPEN,
            carryin => \nx.n10852\,
            carryout => \nx.n10853\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1406_8_lut_LC_9_26_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42088\,
            in2 => \N__28790\,
            in3 => \N__27309\,
            lcout => \nx.n2071\,
            ltout => OPEN,
            carryin => \nx.n10853\,
            carryout => \nx.n10854\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1406_9_lut_LC_9_26_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42063\,
            in2 => \N__28848\,
            in3 => \N__27306\,
            lcout => \nx.n2070\,
            ltout => OPEN,
            carryin => \nx.n10854\,
            carryout => \nx.n10855\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1406_10_lut_LC_9_27_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42089\,
            in2 => \N__28644\,
            in3 => \N__27303\,
            lcout => \nx.n2069\,
            ltout => OPEN,
            carryin => \bfn_9_27_0_\,
            carryout => \nx.n10856\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1406_11_lut_LC_9_27_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42064\,
            in2 => \N__28554\,
            in3 => \N__27300\,
            lcout => \nx.n2068\,
            ltout => OPEN,
            carryin => \nx.n10856\,
            carryout => \nx.n10857\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1406_12_lut_LC_9_27_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42090\,
            in2 => \N__28821\,
            in3 => \N__27297\,
            lcout => \nx.n2067\,
            ltout => OPEN,
            carryin => \nx.n10857\,
            carryout => \nx.n10858\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1406_13_lut_LC_9_27_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42065\,
            in2 => \N__28530\,
            in3 => \N__27426\,
            lcout => \nx.n2066\,
            ltout => OPEN,
            carryin => \nx.n10858\,
            carryout => \nx.n10859\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1406_14_lut_LC_9_27_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42091\,
            in2 => \N__28755\,
            in3 => \N__27423\,
            lcout => \nx.n2065\,
            ltout => OPEN,
            carryin => \nx.n10859\,
            carryout => \nx.n10860\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1406_15_lut_LC_9_27_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42066\,
            in2 => \N__28982\,
            in3 => \N__27420\,
            lcout => \nx.n2064\,
            ltout => OPEN,
            carryin => \nx.n10860\,
            carryout => \nx.n10861\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1406_16_lut_LC_9_27_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42092\,
            in2 => \N__29157\,
            in3 => \N__27417\,
            lcout => \nx.n2063\,
            ltout => OPEN,
            carryin => \nx.n10861\,
            carryout => \nx.n10862\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1406_17_lut_LC_9_27_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42067\,
            in2 => \N__27392\,
            in3 => \N__27414\,
            lcout => \nx.n2062\,
            ltout => OPEN,
            carryin => \nx.n10862\,
            carryout => \nx.n10863\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1406_18_lut_LC_9_28_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001000001100000"
        )
    port map (
            in0 => \N__42216\,
            in1 => \N__27411\,
            in2 => \N__29125\,
            in3 => \N__27396\,
            lcout => \nx.n2093\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1409_3_lut_LC_9_28_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29112\,
            in2 => \N__27393\,
            in3 => \N__27366\,
            lcout => \nx.n2094\,
            ltout => \nx.n2094_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i1_2_lut_adj_35_LC_9_28_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__27360\,
            in3 => \N__30854\,
            lcout => \nx.n18_adj_682\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1347_3_lut_LC_9_28_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27357\,
            in2 => \N__27580\,
            in3 => \N__27330\,
            lcout => \nx.n2000\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1348_3_lut_LC_9_28_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27621\,
            in2 => \N__27612\,
            in3 => \N__27568\,
            lcout => \nx.n2001\,
            ltout => \nx.n2001_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1415_3_lut_LC_9_28_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27489\,
            in2 => \N__27483\,
            in3 => \N__29111\,
            lcout => \nx.n2100\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1414_3_lut_LC_9_28_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28819\,
            in2 => \N__29126\,
            in3 => \N__27480\,
            lcout => \nx.n2099\,
            ltout => \nx.n2099_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i11_4_lut_adj_38_LC_9_28_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__30337\,
            in1 => \N__36580\,
            in2 => \N__27474\,
            in3 => \N__30712\,
            lcout => \nx.n28_adj_686\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_635__i0_LC_9_29_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27471\,
            in2 => \_gnd_net_\,
            in3 => \N__27465\,
            lcout => n26_adj_798,
            ltout => OPEN,
            carryin => \bfn_9_29_0_\,
            carryout => n10644,
            clk => \N__46913\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_635__i1_LC_9_29_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27462\,
            in2 => \_gnd_net_\,
            in3 => \N__27456\,
            lcout => n25,
            ltout => OPEN,
            carryin => n10644,
            carryout => n10645,
            clk => \N__46913\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_635__i2_LC_9_29_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27453\,
            in2 => \_gnd_net_\,
            in3 => \N__27447\,
            lcout => n24,
            ltout => OPEN,
            carryin => n10645,
            carryout => n10646,
            clk => \N__46913\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_635__i3_LC_9_29_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27444\,
            in2 => \_gnd_net_\,
            in3 => \N__27438\,
            lcout => n23,
            ltout => OPEN,
            carryin => n10646,
            carryout => n10647,
            clk => \N__46913\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_635__i4_LC_9_29_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27435\,
            in2 => \_gnd_net_\,
            in3 => \N__27429\,
            lcout => n22_adj_799,
            ltout => OPEN,
            carryin => n10647,
            carryout => n10648,
            clk => \N__46913\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_635__i5_LC_9_29_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27693\,
            in2 => \_gnd_net_\,
            in3 => \N__27687\,
            lcout => n21,
            ltout => OPEN,
            carryin => n10648,
            carryout => n10649,
            clk => \N__46913\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_635__i6_LC_9_29_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27684\,
            in2 => \_gnd_net_\,
            in3 => \N__27678\,
            lcout => n20,
            ltout => OPEN,
            carryin => n10649,
            carryout => n10650,
            clk => \N__46913\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_635__i7_LC_9_29_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27675\,
            in2 => \_gnd_net_\,
            in3 => \N__27669\,
            lcout => n19_adj_800,
            ltout => OPEN,
            carryin => n10650,
            carryout => n10651,
            clk => \N__46913\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_635__i8_LC_9_30_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27666\,
            in2 => \_gnd_net_\,
            in3 => \N__27660\,
            lcout => n18,
            ltout => OPEN,
            carryin => \bfn_9_30_0_\,
            carryout => n10652,
            clk => \N__46915\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_635__i9_LC_9_30_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27657\,
            in2 => \_gnd_net_\,
            in3 => \N__27651\,
            lcout => n17,
            ltout => OPEN,
            carryin => n10652,
            carryout => n10653,
            clk => \N__46915\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_635__i10_LC_9_30_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27648\,
            in2 => \_gnd_net_\,
            in3 => \N__27642\,
            lcout => n16,
            ltout => OPEN,
            carryin => n10653,
            carryout => n10654,
            clk => \N__46915\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_635__i11_LC_9_30_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27639\,
            in2 => \_gnd_net_\,
            in3 => \N__27633\,
            lcout => n15,
            ltout => OPEN,
            carryin => n10654,
            carryout => n10655,
            clk => \N__46915\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_635__i12_LC_9_30_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27630\,
            in2 => \_gnd_net_\,
            in3 => \N__27624\,
            lcout => n14_adj_802,
            ltout => OPEN,
            carryin => n10655,
            carryout => n10656,
            clk => \N__46915\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_635__i13_LC_9_30_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27765\,
            in2 => \_gnd_net_\,
            in3 => \N__27759\,
            lcout => n13,
            ltout => OPEN,
            carryin => n10656,
            carryout => n10657,
            clk => \N__46915\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_635__i14_LC_9_30_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27756\,
            in2 => \_gnd_net_\,
            in3 => \N__27750\,
            lcout => n12,
            ltout => OPEN,
            carryin => n10657,
            carryout => n10658,
            clk => \N__46915\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_635__i15_LC_9_30_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27747\,
            in2 => \_gnd_net_\,
            in3 => \N__27741\,
            lcout => n11,
            ltout => OPEN,
            carryin => n10658,
            carryout => n10659,
            clk => \N__46915\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_635__i16_LC_9_31_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27738\,
            in2 => \_gnd_net_\,
            in3 => \N__27732\,
            lcout => n10_adj_806,
            ltout => OPEN,
            carryin => \bfn_9_31_0_\,
            carryout => n10660,
            clk => \N__46921\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_635__i17_LC_9_31_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27729\,
            in2 => \_gnd_net_\,
            in3 => \N__27723\,
            lcout => n9_adj_807,
            ltout => OPEN,
            carryin => n10660,
            carryout => n10661,
            clk => \N__46921\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_635__i18_LC_9_31_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27720\,
            in2 => \_gnd_net_\,
            in3 => \N__27714\,
            lcout => n8,
            ltout => OPEN,
            carryin => n10661,
            carryout => n10662,
            clk => \N__46921\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_635__i19_LC_9_31_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27711\,
            in2 => \_gnd_net_\,
            in3 => \N__27705\,
            lcout => n7_adj_808,
            ltout => OPEN,
            carryin => n10662,
            carryout => n10663,
            clk => \N__46921\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_635__i20_LC_9_31_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27702\,
            in2 => \_gnd_net_\,
            in3 => \N__27696\,
            lcout => n6_adj_809,
            ltout => OPEN,
            carryin => n10663,
            carryout => n10664,
            clk => \N__46921\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_635__i21_LC_9_31_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27878\,
            in2 => \_gnd_net_\,
            in3 => \N__27867\,
            lcout => blink_counter_21,
            ltout => OPEN,
            carryin => n10664,
            carryout => n10665,
            clk => \N__46921\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_635__i22_LC_9_31_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27857\,
            in2 => \_gnd_net_\,
            in3 => \N__27846\,
            lcout => blink_counter_22,
            ltout => OPEN,
            carryin => n10665,
            carryout => n10666,
            clk => \N__46921\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_635__i23_LC_9_31_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27833\,
            in2 => \_gnd_net_\,
            in3 => \N__27822\,
            lcout => blink_counter_23,
            ltout => OPEN,
            carryin => n10666,
            carryout => n10667,
            clk => \N__46921\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_635__i24_LC_9_32_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27806\,
            in2 => \_gnd_net_\,
            in3 => \N__27795\,
            lcout => blink_counter_24,
            ltout => OPEN,
            carryin => \bfn_9_32_0_\,
            carryout => n10668,
            clk => \N__46923\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_635__i25_LC_9_32_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27782\,
            in2 => \_gnd_net_\,
            in3 => \N__27792\,
            lcout => blink_counter_25,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46923\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i1_4_lut_adj_96_LC_10_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101100"
        )
    port map (
            in0 => \N__32943\,
            in1 => \N__32962\,
            in2 => \N__34006\,
            in3 => \N__30945\,
            lcout => \nx.n12775\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i2154_3_lut_LC_10_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33663\,
            in2 => \N__33692\,
            in3 => \N__33984\,
            lcout => OPEN,
            ltout => \nx.n45_adj_754_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i1_4_lut_adj_99_LC_10_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__27918\,
            in1 => \N__30759\,
            in2 => \N__27771\,
            in3 => \N__27897\,
            lcout => OPEN,
            ltout => \nx.n12809_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i1_4_lut_adj_100_LC_10_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101011111100"
        )
    port map (
            in0 => \N__33618\,
            in1 => \N__33648\,
            in2 => \N__27768\,
            in3 => \N__33985\,
            lcout => OPEN,
            ltout => \nx.n12811_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i1_4_lut_adj_101_LC_10_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110111111000"
        )
    port map (
            in0 => \N__33986\,
            in1 => \N__33573\,
            in2 => \N__27930\,
            in3 => \N__33603\,
            lcout => OPEN,
            ltout => \nx.n12813_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i1_4_lut_adj_102_LC_10_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101011111100"
        )
    port map (
            in0 => \N__33531\,
            in1 => \N__33554\,
            in2 => \N__27927\,
            in3 => \N__33987\,
            lcout => \nx.n12815\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i2155_3_lut_LC_10_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33085\,
            in2 => \N__34007\,
            in3 => \N__33708\,
            lcout => \nx.n43_adj_753\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i19_4_lut_adj_80_LC_10_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__33238\,
            in1 => \N__33043\,
            in2 => \N__33205\,
            in3 => \N__32923\,
            lcout => OPEN,
            ltout => \nx.n46_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i23_4_lut_LC_10_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__32794\,
            in1 => \N__33361\,
            in2 => \N__27912\,
            in3 => \N__27891\,
            lcout => \nx.n50_adj_742\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i2170_3_lut_LC_10_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33027\,
            in2 => \N__33050\,
            in3 => \N__33988\,
            lcout => OPEN,
            ltout => \nx.n13_adj_743_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i1_4_lut_adj_94_LC_10_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110111111000"
        )
    port map (
            in0 => \N__33989\,
            in1 => \N__33264\,
            in2 => \N__27909\,
            in3 => \N__33286\,
            lcout => OPEN,
            ltout => \nx.n12787_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i1_4_lut_adj_98_LC_10_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__30933\,
            in1 => \N__27906\,
            in2 => \N__27900\,
            in3 => \N__30960\,
            lcout => \nx.n12803\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i8_3_lut_adj_81_LC_10_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110100000"
        )
    port map (
            in0 => \N__32399\,
            in1 => \_gnd_net_\,
            in2 => \N__32353\,
            in3 => \N__33004\,
            lcout => \nx.n35_adj_738\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i2035_3_lut_LC_10_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35186\,
            in2 => \N__37322\,
            in3 => \N__35166\,
            lcout => \nx.n3008\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i2014_3_lut_LC_10_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35611\,
            in2 => \N__35589\,
            in3 => \N__37311\,
            lcout => \nx.n2987\,
            ltout => \nx.n2987_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i15_4_lut_LC_10_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__29248\,
            in1 => \N__29476\,
            in2 => \N__28011\,
            in3 => \N__30919\,
            lcout => OPEN,
            ltout => \nx.n41_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i24_4_lut_LC_10_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__36933\,
            in1 => \N__34920\,
            in2 => \N__28008\,
            in3 => \N__31077\,
            lcout => OPEN,
            ltout => \nx.n50_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i25_4_lut_LC_10_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__28005\,
            in1 => \N__31383\,
            in2 => \N__27999\,
            in3 => \N__29514\,
            lcout => \nx.n3017\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i2034_3_lut_LC_10_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011110000"
        )
    port map (
            in0 => \N__35118\,
            in1 => \_gnd_net_\,
            in2 => \N__35150\,
            in3 => \N__37307\,
            lcout => \nx.n3007\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1968_3_lut_LC_10_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__27996\,
            in1 => \N__28215\,
            in2 => \_gnd_net_\,
            in3 => \N__37513\,
            lcout => \nx.n2909\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1948_3_lut_LC_10_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27987\,
            in2 => \N__37566\,
            in3 => \N__27975\,
            lcout => \nx.n2889\,
            ltout => \nx.n2889_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i5_3_lut_adj_112_LC_10_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35257\,
            in2 => \N__27942\,
            in3 => \N__35185\,
            lcout => \nx.n30_adj_759\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1959_3_lut_LC_10_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101000001010"
        )
    port map (
            in0 => \N__28110\,
            in1 => \_gnd_net_\,
            in2 => \N__37565\,
            in3 => \N__27939\,
            lcout => \nx.n2900\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i16_4_lut_adj_61_LC_10_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__28027\,
            in1 => \N__33845\,
            in2 => \N__34883\,
            in3 => \N__28109\,
            lcout => OPEN,
            ltout => \nx.n40_adj_705_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i20_4_lut_LC_10_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__37658\,
            in1 => \N__28081\,
            in2 => \N__28062\,
            in3 => \N__28167\,
            lcout => OPEN,
            ltout => \nx.n44_adj_721_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i23_4_lut_adj_90_LC_10_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__29484\,
            in1 => \N__28038\,
            in2 => \N__28059\,
            in3 => \N__28302\,
            lcout => \nx.n2819\,
            ltout => \nx.n2819_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1953_3_lut_LC_10_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28056\,
            in2 => \N__28047\,
            in3 => \N__28137\,
            lcout => \nx.n2894\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1965_3_lut_LC_10_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28044\,
            in2 => \N__28032\,
            in3 => \N__37521\,
            lcout => \nx.n2906\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i18_4_lut_adj_74_LC_10_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__28160\,
            in1 => \N__34804\,
            in2 => \N__29775\,
            in3 => \N__34168\,
            lcout => \nx.n42_adj_730\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1894_3_lut_LC_10_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__28407\,
            in1 => \_gnd_net_\,
            in2 => \N__31253\,
            in3 => \N__37817\,
            lcout => \nx.n2803\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i13_3_lut_adj_114_LC_10_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111010"
        )
    port map (
            in0 => \N__35528\,
            in1 => \_gnd_net_\,
            in2 => \N__35065\,
            in3 => \N__35861\,
            lcout => \nx.n38_adj_762\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1898_3_lut_LC_10_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28263\,
            in2 => \N__31252\,
            in3 => \N__35805\,
            lcout => \nx.n2807\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1900_3_lut_LC_10_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__28293\,
            in1 => \N__30147\,
            in2 => \_gnd_net_\,
            in3 => \N__31205\,
            lcout => \nx.n2809\,
            ltout => \nx.n2809_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i6_3_lut_LC_10_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28129\,
            in2 => \N__28218\,
            in3 => \N__28214\,
            lcout => \nx.n30_adj_704\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1893_3_lut_LC_10_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35771\,
            in2 => \N__28395\,
            in3 => \N__31212\,
            lcout => \nx.n2802\,
            ltout => \nx.n2802_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1960_3_lut_LC_10_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28146\,
            in2 => \N__28140\,
            in3 => \N__37555\,
            lcout => \nx.n2901\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1886_3_lut_LC_10_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30035\,
            in2 => \N__31255\,
            in3 => \N__28500\,
            lcout => \nx.n2795\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i9135_3_lut_LC_10_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28371\,
            in2 => \N__29898\,
            in3 => \N__31216\,
            lcout => \nx.n2800\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1895_3_lut_LC_10_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28239\,
            in2 => \N__31254\,
            in3 => \N__37856\,
            lcout => \nx.n2804\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i22_4_lut_LC_10_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__29961\,
            in1 => \N__29832\,
            in2 => \N__29874\,
            in3 => \N__35745\,
            lcout => \nx.n2720\,
            ltout => \nx.n2720_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i9137_3_lut_LC_10_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28248\,
            in2 => \N__28113\,
            in3 => \N__29741\,
            lcout => \nx.n2805\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1879_3_lut_LC_10_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31220\,
            in2 => \N__31479\,
            in3 => \N__28425\,
            lcout => \nx.n2788\,
            ltout => \nx.n2788_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i2_2_lut_LC_10_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__28347\,
            in3 => \N__28336\,
            lcout => OPEN,
            ltout => \nx.n26_adj_706_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i19_4_lut_adj_78_LC_10_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__28607\,
            in1 => \N__29938\,
            in2 => \N__28314\,
            in3 => \N__28311\,
            lcout => \nx.n43_adj_735\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1875_2_lut_LC_10_23_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30142\,
            in2 => \_gnd_net_\,
            in3 => \N__28281\,
            lcout => \nx.n2777\,
            ltout => OPEN,
            carryin => \bfn_10_23_0_\,
            carryout => \nx.n10981\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1875_3_lut_LC_10_23_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__29999\,
            in3 => \N__28266\,
            lcout => \nx.n2776\,
            ltout => OPEN,
            carryin => \nx.n10981\,
            carryout => \nx.n10982\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1875_4_lut_LC_10_23_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41748\,
            in2 => \N__35803\,
            in3 => \N__28254\,
            lcout => \nx.n2775\,
            ltout => OPEN,
            carryin => \nx.n10982\,
            carryout => \nx.n10983\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1875_5_lut_LC_10_23_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41751\,
            in2 => \N__31818\,
            in3 => \N__28251\,
            lcout => \nx.n2774\,
            ltout => OPEN,
            carryin => \nx.n10983\,
            carryout => \nx.n10984\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1875_6_lut_LC_10_23_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41749\,
            in2 => \N__29742\,
            in3 => \N__28242\,
            lcout => \nx.n2773\,
            ltout => OPEN,
            carryin => \nx.n10984\,
            carryout => \nx.n10985\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1875_7_lut_LC_10_23_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41752\,
            in2 => \N__37857\,
            in3 => \N__28410\,
            lcout => \nx.n2772\,
            ltout => OPEN,
            carryin => \nx.n10985\,
            carryout => \nx.n10986\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1875_8_lut_LC_10_23_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41750\,
            in2 => \N__37821\,
            in3 => \N__28398\,
            lcout => \nx.n2771\,
            ltout => OPEN,
            carryin => \nx.n10986\,
            carryout => \nx.n10987\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1875_9_lut_LC_10_23_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41753\,
            in2 => \N__35775\,
            in3 => \N__28383\,
            lcout => \nx.n2770\,
            ltout => OPEN,
            carryin => \nx.n10987\,
            carryout => \nx.n10988\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1875_10_lut_LC_10_24_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42047\,
            in2 => \N__34208\,
            in3 => \N__28374\,
            lcout => \nx.n2769\,
            ltout => OPEN,
            carryin => \bfn_10_24_0_\,
            carryout => \nx.n10989\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1875_11_lut_LC_10_24_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42051\,
            in2 => \N__29894\,
            in3 => \N__28362\,
            lcout => \nx.n2768\,
            ltout => OPEN,
            carryin => \nx.n10989\,
            carryout => \nx.n10990\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1875_12_lut_LC_10_24_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42048\,
            in2 => \N__31536\,
            in3 => \N__28359\,
            lcout => \nx.n2767\,
            ltout => OPEN,
            carryin => \nx.n10990\,
            carryout => \nx.n10991\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1875_13_lut_LC_10_24_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42052\,
            in2 => \N__29922\,
            in3 => \N__28356\,
            lcout => \nx.n2766\,
            ltout => OPEN,
            carryin => \nx.n10991\,
            carryout => \nx.n10992\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1875_14_lut_LC_10_24_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42049\,
            in2 => \N__29858\,
            in3 => \N__28353\,
            lcout => \nx.n2765\,
            ltout => OPEN,
            carryin => \nx.n10992\,
            carryout => \nx.n10993\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1875_15_lut_LC_10_24_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42053\,
            in2 => \N__31301\,
            in3 => \N__28350\,
            lcout => \nx.n2764\,
            ltout => OPEN,
            carryin => \nx.n10993\,
            carryout => \nx.n10994\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1875_16_lut_LC_10_24_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42050\,
            in2 => \N__30036\,
            in3 => \N__28491\,
            lcout => \nx.n2763\,
            ltout => OPEN,
            carryin => \nx.n10994\,
            carryout => \nx.n10995\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1875_17_lut_LC_10_24_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42054\,
            in2 => \N__31668\,
            in3 => \N__28479\,
            lcout => \nx.n2762\,
            ltout => OPEN,
            carryin => \nx.n10995\,
            carryout => \nx.n10996\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1875_18_lut_LC_10_25_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42055\,
            in2 => \N__30062\,
            in3 => \N__28470\,
            lcout => \nx.n2761\,
            ltout => OPEN,
            carryin => \bfn_10_25_0_\,
            carryout => \nx.n10997\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1875_19_lut_LC_10_25_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41966\,
            in2 => \N__30083\,
            in3 => \N__28461\,
            lcout => \nx.n2760\,
            ltout => OPEN,
            carryin => \nx.n10997\,
            carryout => \nx.n10998\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1875_20_lut_LC_10_25_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42056\,
            in2 => \N__31575\,
            in3 => \N__28446\,
            lcout => \nx.n2759\,
            ltout => OPEN,
            carryin => \nx.n10998\,
            carryout => \nx.n10999\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1875_21_lut_LC_10_25_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41967\,
            in2 => \N__31638\,
            in3 => \N__28437\,
            lcout => \nx.n2758\,
            ltout => OPEN,
            carryin => \nx.n10999\,
            carryout => \nx.n11000\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1875_22_lut_LC_10_25_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42057\,
            in2 => \N__31607\,
            in3 => \N__28428\,
            lcout => \nx.n2757\,
            ltout => OPEN,
            carryin => \nx.n11000\,
            carryout => \nx.n11001\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1875_23_lut_LC_10_25_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41968\,
            in2 => \N__31478\,
            in3 => \N__28416\,
            lcout => \nx.n2756\,
            ltout => OPEN,
            carryin => \nx.n11001\,
            carryout => \nx.n11002\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1875_24_lut_LC_10_25_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42058\,
            in2 => \N__31509\,
            in3 => \N__28413\,
            lcout => \nx.n2755\,
            ltout => OPEN,
            carryin => \nx.n11002\,
            carryout => \nx.n11003\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1875_25_lut_LC_10_25_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001000001100000"
        )
    port map (
            in0 => \N__42059\,
            in1 => \N__39983\,
            in2 => \N__31275\,
            in3 => \N__28611\,
            lcout => \nx.n2786\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1417_3_lut_LC_10_26_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28843\,
            in2 => \N__28590\,
            in3 => \N__29120\,
            lcout => \nx.n2102\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i5916_2_lut_LC_10_26_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28937\,
            in2 => \_gnd_net_\,
            in3 => \N__29200\,
            lcout => OPEN,
            ltout => \nx.n9709_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i10_4_lut_adj_31_LC_10_26_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__28522\,
            in1 => \N__28744\,
            in2 => \N__28581\,
            in3 => \N__28636\,
            lcout => OPEN,
            ltout => \nx.n26_adj_681_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i15_4_lut_adj_34_LC_10_26_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__28797\,
            in1 => \N__28578\,
            in2 => \N__28566\,
            in3 => \N__28536\,
            lcout => \nx.n2027\,
            ltout => \nx.n2027_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1421_3_lut_LC_10_26_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101000001010"
        )
    port map (
            in0 => \N__28868\,
            in1 => \_gnd_net_\,
            in2 => \N__28563\,
            in3 => \N__28560\,
            lcout => \nx.n2106\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i12_4_lut_adj_30_LC_10_26_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__28672\,
            in1 => \N__28712\,
            in2 => \N__28789\,
            in3 => \N__28553\,
            lcout => \nx.n28_adj_680\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1413_3_lut_LC_10_26_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010101010"
        )
    port map (
            in0 => \N__28523\,
            in1 => \_gnd_net_\,
            in2 => \N__28509\,
            in3 => \N__29121\,
            lcout => \nx.n2098\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i11_4_lut_adj_32_LC_10_26_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__29021\,
            in1 => \N__28867\,
            in2 => \N__28847\,
            in3 => \N__28820\,
            lcout => \nx.n27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1418_3_lut_LC_10_27_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101000001010"
        )
    port map (
            in0 => \N__28791\,
            in1 => \_gnd_net_\,
            in2 => \N__29122\,
            in3 => \N__28764\,
            lcout => \nx.n2103\,
            ltout => \nx.n2103_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i7_2_lut_LC_10_27_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__28758\,
            in3 => \N__30365\,
            lcout => \nx.n24_adj_684\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1412_3_lut_LC_10_27_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28754\,
            in2 => \N__29124\,
            in3 => \N__28728\,
            lcout => \nx.n2097\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1420_3_lut_LC_10_27_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28722\,
            in2 => \N__28716\,
            in3 => \N__29094\,
            lcout => \nx.n2105\,
            ltout => \nx.n2105_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1487_3_lut_LC_10_27_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101100011011000"
        )
    port map (
            in0 => \N__36533\,
            in1 => \N__30354\,
            in2 => \N__28683\,
            in3 => \_gnd_net_\,
            lcout => \nx.n2204\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1419_3_lut_LC_10_27_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28680\,
            in2 => \N__28653\,
            in3 => \N__29095\,
            lcout => \nx.n2104\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1416_3_lut_LC_10_27_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28643\,
            in2 => \N__29123\,
            in3 => \N__28617\,
            lcout => \nx.n2101\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1492_3_lut_LC_10_27_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30528\,
            in2 => \N__30486\,
            in3 => \N__36532\,
            lcout => \nx.n2209\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1422_3_lut_LC_10_28_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29034\,
            in2 => \N__29025\,
            in3 => \N__29106\,
            lcout => \nx.n2107\,
            ltout => \nx.n2107_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i12_4_lut_adj_39_LC_10_28_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111000"
        )
    port map (
            in0 => \N__30470\,
            in1 => \N__30533\,
            in2 => \N__28992\,
            in3 => \N__28989\,
            lcout => \nx.n29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1411_3_lut_LC_10_28_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28983\,
            in2 => \N__28953\,
            in3 => \N__29107\,
            lcout => \nx.n2096\,
            ltout => \nx.n2096_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i10_4_lut_adj_45_LC_10_28_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__30671\,
            in1 => \N__30628\,
            in2 => \N__28944\,
            in3 => \N__30562\,
            lcout => \nx.n27_adj_691\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1424_3_lut_LC_10_28_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__28941\,
            in1 => \N__28893\,
            in2 => \_gnd_net_\,
            in3 => \N__29105\,
            lcout => \nx.n2109\,
            ltout => \nx.n2109_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1491_3_lut_LC_10_28_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011110000"
        )
    port map (
            in0 => \N__30456\,
            in1 => \_gnd_net_\,
            in2 => \N__28881\,
            in3 => \N__36534\,
            lcout => \nx.n2208\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1485_3_lut_LC_10_28_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30291\,
            in2 => \N__36559\,
            in3 => \N__30305\,
            lcout => \nx.n2202\,
            ltout => \nx.n2202_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i4_3_lut_LC_10_28_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101011110000"
        )
    port map (
            in0 => \N__31696\,
            in1 => \_gnd_net_\,
            in2 => \N__28878\,
            in3 => \N__31789\,
            lcout => \nx.n22_adj_693\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i13_4_lut_adj_37_LC_10_29_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__30446\,
            in1 => \N__30398\,
            in2 => \N__32707\,
            in3 => \N__28875\,
            lcout => \nx.n30_adj_685\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1478_3_lut_LC_10_29_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010101010"
        )
    port map (
            in0 => \N__30596\,
            in1 => \_gnd_net_\,
            in2 => \N__30582\,
            in3 => \N__36525\,
            lcout => \nx.n2195\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1476_3_lut_LC_10_29_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30887\,
            in2 => \N__36558\,
            in3 => \N__30873\,
            lcout => \nx.n2193\,
            ltout => \nx.n2193_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i10_4_lut_adj_47_LC_10_29_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__32596\,
            in1 => \N__32638\,
            in2 => \N__29208\,
            in3 => \N__30833\,
            lcout => \nx.n28_adj_692\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1423_3_lut_LC_10_29_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29205\,
            in2 => \N__29175\,
            in3 => \N__29116\,
            lcout => \nx.n2108\,
            ltout => \nx.n2108_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1490_3_lut_LC_10_29_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30432\,
            in2 => \N__29160\,
            in3 => \N__36524\,
            lcout => \nx.n2207\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1488_3_lut_LC_10_29_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__30381\,
            in1 => \_gnd_net_\,
            in2 => \N__36557\,
            in3 => \N__30399\,
            lcout => \nx.n2205\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1410_3_lut_LC_10_29_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29153\,
            in2 => \N__29127\,
            in3 => \N__29043\,
            lcout => \nx.n2095\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONSTANT_ONE_LUT4_LC_11_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \CONSTANT_ONE_NET\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i15_4_lut_adj_82_LC_11_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__33508\,
            in1 => \N__33412\,
            in2 => \N__33466\,
            in3 => \N__34126\,
            lcout => OPEN,
            ltout => \nx.n42_adj_739_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i21_4_lut_adj_85_LC_11_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__33328\,
            in1 => \N__34078\,
            in2 => \N__29397\,
            in3 => \N__33887\,
            lcout => \nx.n48\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i5_2_lut_adj_83_LC_11_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33685\,
            in2 => \_gnd_net_\,
            in3 => \N__33640\,
            lcout => OPEN,
            ltout => \nx.n32_adj_740_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i22_4_lut_adj_86_LC_11_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__33595\,
            in1 => \N__33553\,
            in2 => \N__29394\,
            in3 => \N__29391\,
            lcout => OPEN,
            ltout => \nx.n49_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i26_4_lut_LC_11_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__29379\,
            in1 => \N__29373\,
            in2 => \N__29358\,
            in3 => \N__29355\,
            lcout => \nx.n3116\,
            ltout => \nx.n3116_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i2167_3_lut_LC_11_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32924\,
            in2 => \N__29349\,
            in3 => \N__32904\,
            lcout => \nx.n19_adj_745\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_2076_2_lut_LC_11_18_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__29346\,
            in1 => \N__29345\,
            in2 => \N__29276\,
            in3 => \N__29301\,
            lcout => \nx.n3109\,
            ltout => OPEN,
            carryin => \bfn_11_18_0_\,
            carryout => \nx.n11053\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_2076_3_lut_LC_11_18_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__29298\,
            in1 => \N__29297\,
            in2 => \N__29277\,
            in3 => \N__29253\,
            lcout => \nx.n3108\,
            ltout => OPEN,
            carryin => \nx.n11053\,
            carryout => \nx.n11054\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_2076_4_lut_LC_11_18_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101000111010"
        )
    port map (
            in0 => \N__29250\,
            in1 => \N__29249\,
            in2 => \N__29670\,
            in3 => \N__29232\,
            lcout => \nx.n3107\,
            ltout => OPEN,
            carryin => \nx.n11054\,
            carryout => \nx.n11055\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_2076_5_lut_LC_11_18_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101000111010"
        )
    port map (
            in0 => \N__29229\,
            in1 => \N__29228\,
            in2 => \N__29673\,
            in3 => \N__29211\,
            lcout => \nx.n3106\,
            ltout => OPEN,
            carryin => \nx.n11055\,
            carryout => \nx.n11056\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_2076_6_lut_LC_11_18_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101000111010"
        )
    port map (
            in0 => \N__34959\,
            in1 => \N__34958\,
            in2 => \N__29671\,
            in3 => \N__29424\,
            lcout => \nx.n3105\,
            ltout => OPEN,
            carryin => \nx.n11056\,
            carryout => \nx.n11057\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_2076_7_lut_LC_11_18_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101000111010"
        )
    port map (
            in0 => \N__31050\,
            in1 => \N__31049\,
            in2 => \N__29674\,
            in3 => \N__29421\,
            lcout => \nx.n3104\,
            ltout => OPEN,
            carryin => \nx.n11057\,
            carryout => \nx.n11058\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_2076_8_lut_LC_11_18_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101000111010"
        )
    port map (
            in0 => \N__34944\,
            in1 => \N__34943\,
            in2 => \N__29672\,
            in3 => \N__29418\,
            lcout => \nx.n3103\,
            ltout => OPEN,
            carryin => \nx.n11058\,
            carryout => \nx.n11059\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_2076_9_lut_LC_11_18_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101000111010"
        )
    port map (
            in0 => \N__31068\,
            in1 => \N__31067\,
            in2 => \N__29675\,
            in3 => \N__29415\,
            lcout => \nx.n3102\,
            ltout => OPEN,
            carryin => \nx.n11059\,
            carryout => \nx.n11060\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_2076_10_lut_LC_11_19_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101000111010"
        )
    port map (
            in0 => \N__36978\,
            in1 => \N__36977\,
            in2 => \N__29676\,
            in3 => \N__29412\,
            lcout => \nx.n3101\,
            ltout => OPEN,
            carryin => \bfn_11_19_0_\,
            carryout => \nx.n11061\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_2076_11_lut_LC_11_19_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101000111010"
        )
    port map (
            in0 => \N__31092\,
            in1 => \N__31091\,
            in2 => \N__29680\,
            in3 => \N__29409\,
            lcout => \nx.n3100\,
            ltout => OPEN,
            carryin => \nx.n11061\,
            carryout => \nx.n11062\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_2076_12_lut_LC_11_19_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101000111010"
        )
    port map (
            in0 => \N__31112\,
            in1 => \N__31111\,
            in2 => \N__29677\,
            in3 => \N__29406\,
            lcout => \nx.n3099\,
            ltout => OPEN,
            carryin => \nx.n11062\,
            carryout => \nx.n11063\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_2076_13_lut_LC_11_19_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101000111010"
        )
    port map (
            in0 => \N__34908\,
            in1 => \N__34907\,
            in2 => \N__29681\,
            in3 => \N__29403\,
            lcout => \nx.n3098\,
            ltout => OPEN,
            carryin => \nx.n11063\,
            carryout => \nx.n11064\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_2076_14_lut_LC_11_19_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101000111010"
        )
    port map (
            in0 => \N__29478\,
            in1 => \N__29477\,
            in2 => \N__29678\,
            in3 => \N__29400\,
            lcout => \nx.n3097\,
            ltout => OPEN,
            carryin => \nx.n11064\,
            carryout => \nx.n11065\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_2076_15_lut_LC_11_19_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101000111010"
        )
    port map (
            in0 => \N__31398\,
            in1 => \N__31397\,
            in2 => \N__29682\,
            in3 => \N__29451\,
            lcout => \nx.n3096\,
            ltout => OPEN,
            carryin => \nx.n11065\,
            carryout => \nx.n11066\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_2076_16_lut_LC_11_19_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101000111010"
        )
    port map (
            in0 => \N__29505\,
            in1 => \N__29504\,
            in2 => \N__29679\,
            in3 => \N__29448\,
            lcout => \nx.n3095\,
            ltout => OPEN,
            carryin => \nx.n11066\,
            carryout => \nx.n11067\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_2076_17_lut_LC_11_19_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101000111010"
        )
    port map (
            in0 => \N__36960\,
            in1 => \N__36959\,
            in2 => \N__29683\,
            in3 => \N__29445\,
            lcout => \nx.n3094\,
            ltout => OPEN,
            carryin => \nx.n11067\,
            carryout => \nx.n11068\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_2076_18_lut_LC_11_20_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101000111010"
        )
    port map (
            in0 => \N__31013\,
            in1 => \N__31012\,
            in2 => \N__29684\,
            in3 => \N__29442\,
            lcout => \nx.n3093\,
            ltout => OPEN,
            carryin => \bfn_11_20_0_\,
            carryout => \nx.n11069\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_2076_19_lut_LC_11_20_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101000111010"
        )
    port map (
            in0 => \N__37167\,
            in1 => \N__37166\,
            in2 => \N__29688\,
            in3 => \N__29439\,
            lcout => \nx.n3092\,
            ltout => OPEN,
            carryin => \nx.n11069\,
            carryout => \nx.n11070\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_2076_20_lut_LC_11_20_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101000111010"
        )
    port map (
            in0 => \N__37686\,
            in1 => \N__37685\,
            in2 => \N__29685\,
            in3 => \N__29436\,
            lcout => \nx.n3091\,
            ltout => OPEN,
            carryin => \nx.n11070\,
            carryout => \nx.n11071\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_2076_21_lut_LC_11_20_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101000111010"
        )
    port map (
            in0 => \N__33732\,
            in1 => \N__33731\,
            in2 => \N__29689\,
            in3 => \N__29433\,
            lcout => \nx.n3090\,
            ltout => OPEN,
            carryin => \nx.n11071\,
            carryout => \nx.n11072\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_2076_22_lut_LC_11_20_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101000111010"
        )
    port map (
            in0 => \N__36873\,
            in1 => \N__36872\,
            in2 => \N__29686\,
            in3 => \N__29430\,
            lcout => \nx.n3089\,
            ltout => OPEN,
            carryin => \nx.n11072\,
            carryout => \nx.n11073\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_2076_23_lut_LC_11_20_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101000111010"
        )
    port map (
            in0 => \N__30924\,
            in1 => \N__30920\,
            in2 => \N__29690\,
            in3 => \N__29427\,
            lcout => \nx.n3088\,
            ltout => OPEN,
            carryin => \nx.n11073\,
            carryout => \nx.n11074\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_2076_24_lut_LC_11_20_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101000111010"
        )
    port map (
            in0 => \N__31371\,
            in1 => \N__31370\,
            in2 => \N__29687\,
            in3 => \N__29727\,
            lcout => \nx.n3087\,
            ltout => OPEN,
            carryin => \nx.n11074\,
            carryout => \nx.n11075\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_2076_25_lut_LC_11_20_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101000111010"
        )
    port map (
            in0 => \N__29724\,
            in1 => \N__29723\,
            in2 => \N__29691\,
            in3 => \N__29712\,
            lcout => \nx.n3086\,
            ltout => OPEN,
            carryin => \nx.n11075\,
            carryout => \nx.n11076\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_2076_26_lut_LC_11_21_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101000111010"
        )
    port map (
            in0 => \N__33753\,
            in1 => \N__33752\,
            in2 => \N__29701\,
            in3 => \N__29709\,
            lcout => \nx.n3085\,
            ltout => OPEN,
            carryin => \bfn_11_21_0_\,
            carryout => \nx.n11077\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_2076_27_lut_LC_11_21_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101000111010"
        )
    port map (
            in0 => \N__29799\,
            in1 => \N__29798\,
            in2 => \N__29703\,
            in3 => \N__29706\,
            lcout => \nx.n3084\,
            ltout => OPEN,
            carryin => \nx.n11077\,
            carryout => \nx.n11078\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_2076_28_lut_LC_11_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101000111010"
        )
    port map (
            in0 => \N__35844\,
            in1 => \N__35843\,
            in2 => \N__29702\,
            in3 => \N__29517\,
            lcout => \nx.n3083\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i14_4_lut_LC_11_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__29497\,
            in1 => \N__31113\,
            in2 => \N__31014\,
            in3 => \N__29797\,
            lcout => \nx.n40_adj_670\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i2023_3_lut_LC_11_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35307\,
            in2 => \N__37392\,
            in3 => \N__37313\,
            lcout => \nx.n2996\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i17_4_lut_adj_79_LC_11_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__31432\,
            in1 => \N__36841\,
            in2 => \N__31139\,
            in3 => \N__33796\,
            lcout => \nx.n41_adj_736\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i2025_3_lut_LC_11_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35334\,
            in2 => \N__37323\,
            in3 => \N__35356\,
            lcout => \nx.n2998\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1888_3_lut_LC_11_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29841\,
            in2 => \N__29862\,
            in3 => \N__31230\,
            lcout => \nx.n2797\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i18_4_lut_adj_41_LC_11_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__31495\,
            in1 => \N__34201\,
            in2 => \N__39984\,
            in3 => \N__31542\,
            lcout => \nx.n41_adj_688\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1890_3_lut_LC_11_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110010101100"
        )
    port map (
            in0 => \N__29826\,
            in1 => \N__31529\,
            in2 => \N__31259\,
            in3 => \_gnd_net_\,
            lcout => \nx.n2799\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1945_3_lut_LC_11_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29942\,
            in2 => \N__29817\,
            in3 => \N__37575\,
            lcout => \nx.n2886\,
            ltout => \nx.n2886_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i2012_3_lut_LC_11_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__37317\,
            in1 => \_gnd_net_\,
            in2 => \N__29802\,
            in3 => \N__35883\,
            lcout => \nx.n2985\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1897_3_lut_LC_11_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31814\,
            in2 => \N__29784\,
            in3 => \N__31226\,
            lcout => \nx.n2806\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1958_3_lut_LC_11_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29773\,
            in2 => \N__37602\,
            in3 => \N__29751\,
            lcout => \nx.n2899\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1813_3_lut_LC_11_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101100011011000"
        )
    port map (
            in0 => \N__40098\,
            in1 => \N__39384\,
            in2 => \N__39410\,
            in3 => \_gnd_net_\,
            lcout => \nx.n2690\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1829_3_lut_LC_11_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38784\,
            in2 => \N__38757\,
            in3 => \N__40097\,
            lcout => \nx.n2706\,
            ltout => \nx.n2706_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i17_4_lut_adj_40_LC_11_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__29921\,
            in1 => \N__31813\,
            in2 => \N__29964\,
            in3 => \N__31528\,
            lcout => \nx.n40_adj_687\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1819_3_lut_LC_11_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39683\,
            in2 => \N__39669\,
            in3 => \N__40096\,
            lcout => \nx.n2696\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1820_3_lut_LC_11_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101100011011000"
        )
    port map (
            in0 => \N__40099\,
            in1 => \N__39705\,
            in2 => \N__39735\,
            in3 => \_gnd_net_\,
            lcout => \nx.n2697\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1878_3_lut_LC_11_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31222\,
            in2 => \N__31505\,
            in3 => \N__29955\,
            lcout => \nx.n2787\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1822_3_lut_LC_11_23_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__40100\,
            in1 => \_gnd_net_\,
            in2 => \N__39108\,
            in3 => \N__39138\,
            lcout => \nx.n2699\,
            ltout => \nx.n2699_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1889_3_lut_LC_11_23_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011110000"
        )
    port map (
            in0 => \N__29907\,
            in1 => \_gnd_net_\,
            in2 => \N__29901\,
            in3 => \N__31221\,
            lcout => \nx.n2798\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i9134_3_lut_LC_11_24_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101000001010"
        )
    port map (
            in0 => \N__39221\,
            in1 => \_gnd_net_\,
            in2 => \N__40094\,
            in3 => \N__39195\,
            lcout => \nx.n2701\,
            ltout => \nx.n2701_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i19_4_lut_adj_36_LC_11_24_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__30093\,
            in1 => \N__31294\,
            in2 => \N__29877\,
            in3 => \N__30015\,
            lcout => \nx.n42_adj_683\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1821_3_lut_LC_11_24_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39086\,
            in2 => \N__40093\,
            in3 => \N__39057\,
            lcout => \nx.n2698\,
            ltout => \nx.n2698_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i7_3_lut_LC_11_24_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30132\,
            in2 => \N__30096\,
            in3 => \N__29995\,
            lcout => \nx.n30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1817_3_lut_LC_11_24_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39567\,
            in2 => \N__40092\,
            in3 => \N__39600\,
            lcout => \nx.n2694\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1816_3_lut_LC_11_24_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39549\,
            in2 => \N__39522\,
            in3 => \N__40058\,
            lcout => \nx.n2693\,
            ltout => \nx.n2693_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i14_4_lut_adj_23_LC_11_24_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__30055\,
            in1 => \N__31657\,
            in2 => \N__30039\,
            in3 => \N__30031\,
            lcout => \nx.n37_adj_677\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1832_3_lut_LC_11_24_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__38920\,
            in1 => \N__38883\,
            in2 => \_gnd_net_\,
            in3 => \N__40051\,
            lcout => \nx.n2709\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1540_2_lut_LC_11_25_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31794\,
            in2 => \_gnd_net_\,
            in3 => \N__29976\,
            lcout => \nx.n2277\,
            ltout => OPEN,
            carryin => \bfn_11_25_0_\,
            carryout => \nx.n10881\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1540_3_lut_LC_11_25_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__31703\,
            in3 => \N__29973\,
            lcout => \nx.n2276\,
            ltout => OPEN,
            carryin => \nx.n10881\,
            carryout => \nx.n10882\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1540_4_lut_LC_11_25_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41559\,
            in2 => \N__32072\,
            in3 => \N__29970\,
            lcout => \nx.n2275\,
            ltout => OPEN,
            carryin => \nx.n10882\,
            carryout => \nx.n10883\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1540_5_lut_LC_11_25_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41561\,
            in2 => \N__32106\,
            in3 => \N__29967\,
            lcout => \nx.n2274\,
            ltout => OPEN,
            carryin => \nx.n10883\,
            carryout => \nx.n10884\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1540_6_lut_LC_11_25_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31724\,
            in2 => \N__41963\,
            in3 => \N__30174\,
            lcout => \nx.n2273\,
            ltout => OPEN,
            carryin => \nx.n10884\,
            carryout => \nx.n10885\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1540_7_lut_LC_11_25_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41565\,
            in2 => \N__32025\,
            in3 => \N__30171\,
            lcout => \nx.n2272\,
            ltout => OPEN,
            carryin => \nx.n10885\,
            carryout => \nx.n10886\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1540_8_lut_LC_11_25_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41560\,
            in2 => \N__31955\,
            in3 => \N__30168\,
            lcout => \nx.n2271\,
            ltout => OPEN,
            carryin => \nx.n10886\,
            carryout => \nx.n10887\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1540_9_lut_LC_11_25_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41566\,
            in2 => \N__31883\,
            in3 => \N__30165\,
            lcout => \nx.n2270\,
            ltout => OPEN,
            carryin => \nx.n10887\,
            carryout => \nx.n10888\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1540_10_lut_LC_11_26_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41567\,
            in2 => \N__31904\,
            in3 => \N__30162\,
            lcout => \nx.n2269\,
            ltout => OPEN,
            carryin => \bfn_11_26_0_\,
            carryout => \nx.n10889\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1540_11_lut_LC_11_26_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41573\,
            in2 => \N__32673\,
            in3 => \N__30159\,
            lcout => \nx.n2268\,
            ltout => OPEN,
            carryin => \nx.n10889\,
            carryout => \nx.n10890\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1540_12_lut_LC_11_26_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41568\,
            in2 => \N__36459\,
            in3 => \N__30156\,
            lcout => \nx.n2267\,
            ltout => OPEN,
            carryin => \nx.n10890\,
            carryout => \nx.n10891\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1540_13_lut_LC_11_26_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31979\,
            in2 => \N__41964\,
            in3 => \N__30153\,
            lcout => \nx.n2266\,
            ltout => OPEN,
            carryin => \nx.n10891\,
            carryout => \nx.n10892\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1540_14_lut_LC_11_26_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32133\,
            in2 => \N__41965\,
            in3 => \N__30150\,
            lcout => \nx.n2265\,
            ltout => OPEN,
            carryin => \nx.n10892\,
            carryout => \nx.n10893\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1540_15_lut_LC_11_26_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41577\,
            in2 => \N__32297\,
            in3 => \N__30201\,
            lcout => \nx.n2264\,
            ltout => OPEN,
            carryin => \nx.n10893\,
            carryout => \nx.n10894\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1540_16_lut_LC_11_26_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41572\,
            in2 => \N__32274\,
            in3 => \N__30198\,
            lcout => \nx.n2263\,
            ltout => OPEN,
            carryin => \nx.n10894\,
            carryout => \nx.n10895\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1540_17_lut_LC_11_26_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41578\,
            in2 => \N__32609\,
            in3 => \N__30195\,
            lcout => \nx.n2262\,
            ltout => OPEN,
            carryin => \nx.n10895\,
            carryout => \nx.n10896\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1540_18_lut_LC_11_27_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41589\,
            in2 => \N__32643\,
            in3 => \N__30192\,
            lcout => \nx.n2261\,
            ltout => OPEN,
            carryin => \bfn_11_27_0_\,
            carryout => \nx.n10897\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1540_19_lut_LC_11_27_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41590\,
            in2 => \N__30281\,
            in3 => \N__30189\,
            lcout => \nx.n2260\,
            ltout => OPEN,
            carryin => \nx.n10897\,
            carryout => \nx.n10898\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1540_20_lut_LC_11_27_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000010001001000"
        )
    port map (
            in0 => \N__41591\,
            in1 => \N__32560\,
            in2 => \N__30840\,
            in3 => \N__30186\,
            lcout => \nx.n2291\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1479_3_lut_LC_11_27_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30612\,
            in2 => \N__30636\,
            in3 => \N__36538\,
            lcout => \nx.n2196\,
            ltout => \nx.n2196_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1546_3_lut_LC_11_27_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30183\,
            in2 => \N__30177\,
            in3 => \N__32558\,
            lcout => \nx.n2295\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i12_4_lut_adj_49_LC_11_27_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__32128\,
            in1 => \N__32062\,
            in2 => \N__31951\,
            in3 => \N__32665\,
            lcout => \nx.n30_adj_694\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1480_3_lut_LC_11_27_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101000001010"
        )
    port map (
            in0 => \N__30670\,
            in1 => \_gnd_net_\,
            in2 => \N__36560\,
            in3 => \N__30648\,
            lcout => \nx.n2197\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1543_3_lut_LC_11_27_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__32559\,
            in1 => \_gnd_net_\,
            in2 => \N__30282\,
            in3 => \N__30264\,
            lcout => \nx.n2292\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1477_3_lut_LC_11_28_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36548\,
            in2 => \N__30570\,
            in3 => \N__30546\,
            lcout => \nx.n2194\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i16_4_lut_adj_46_LC_11_28_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__30258\,
            in1 => \N__30252\,
            in2 => \N__30243\,
            in3 => \N__30234\,
            lcout => \nx.n2126\,
            ltout => \nx.n2126_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1489_3_lut_LC_11_28_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__30408\,
            in1 => \_gnd_net_\,
            in2 => \N__30228\,
            in3 => \N__30422\,
            lcout => \nx.n2206\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1482_3_lut_LC_11_28_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__36552\,
            in1 => \_gnd_net_\,
            in2 => \N__30696\,
            in3 => \N__30722\,
            lcout => \nx.n2199\,
            ltout => \nx.n2199_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i13_4_lut_adj_48_LC_11_28_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__31723\,
            in1 => \N__32092\,
            in2 => \N__30225\,
            in3 => \N__32011\,
            lcout => OPEN,
            ltout => \nx.n31_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i16_4_lut_adj_50_LC_11_28_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__36455\,
            in1 => \N__31873\,
            in2 => \N__30222\,
            in3 => \N__30219\,
            lcout => \nx.n34_adj_695\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1486_3_lut_LC_11_28_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30318\,
            in2 => \N__36563\,
            in3 => \N__30338\,
            lcout => \nx.n2203\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1473_2_lut_LC_11_29_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30532\,
            in2 => \_gnd_net_\,
            in3 => \N__30474\,
            lcout => \nx.n2177\,
            ltout => OPEN,
            carryin => \bfn_11_29_0_\,
            carryout => \nx.n10864\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1473_3_lut_LC_11_29_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__30471\,
            in3 => \N__30450\,
            lcout => \nx.n2176\,
            ltout => OPEN,
            carryin => \nx.n10864\,
            carryout => \nx.n10865\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1473_4_lut_LC_11_29_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42199\,
            in2 => \N__30447\,
            in3 => \N__30426\,
            lcout => \nx.n2175\,
            ltout => OPEN,
            carryin => \nx.n10865\,
            carryout => \nx.n10866\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1473_5_lut_LC_11_29_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41592\,
            in2 => \N__30423\,
            in3 => \N__30402\,
            lcout => \nx.n2174\,
            ltout => OPEN,
            carryin => \nx.n10866\,
            carryout => \nx.n10867\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1473_6_lut_LC_11_29_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30397\,
            in2 => \N__41974\,
            in3 => \N__30375\,
            lcout => \nx.n2173\,
            ltout => OPEN,
            carryin => \nx.n10867\,
            carryout => \nx.n10868\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1473_7_lut_LC_11_29_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41596\,
            in2 => \N__30372\,
            in3 => \N__30345\,
            lcout => \nx.n2172\,
            ltout => OPEN,
            carryin => \nx.n10868\,
            carryout => \nx.n10869\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1473_8_lut_LC_11_29_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42200\,
            in2 => \N__30342\,
            in3 => \N__30312\,
            lcout => \nx.n2171\,
            ltout => OPEN,
            carryin => \nx.n10869\,
            carryout => \nx.n10870\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1473_9_lut_LC_11_29_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41597\,
            in2 => \N__30309\,
            in3 => \N__30285\,
            lcout => \nx.n2170\,
            ltout => OPEN,
            carryin => \nx.n10870\,
            carryout => \nx.n10871\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1473_10_lut_LC_11_30_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41598\,
            in2 => \N__32708\,
            in3 => \N__30732\,
            lcout => \nx.n2169\,
            ltout => OPEN,
            carryin => \bfn_11_30_0_\,
            carryout => \nx.n10872\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1473_11_lut_LC_11_30_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41605\,
            in2 => \N__36593\,
            in3 => \N__30729\,
            lcout => \nx.n2168\,
            ltout => OPEN,
            carryin => \nx.n10872\,
            carryout => \nx.n10873\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1473_12_lut_LC_11_30_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41599\,
            in2 => \N__30726\,
            in3 => \N__30684\,
            lcout => \nx.n2167\,
            ltout => OPEN,
            carryin => \nx.n10873\,
            carryout => \nx.n10874\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1473_13_lut_LC_11_30_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41606\,
            in2 => \N__32166\,
            in3 => \N__30681\,
            lcout => \nx.n2166\,
            ltout => OPEN,
            carryin => \nx.n10874\,
            carryout => \nx.n10875\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1473_14_lut_LC_11_30_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41600\,
            in2 => \N__30678\,
            in3 => \N__30639\,
            lcout => \nx.n2165\,
            ltout => OPEN,
            carryin => \nx.n10875\,
            carryout => \nx.n10876\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1473_15_lut_LC_11_30_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30635\,
            in2 => \N__41975\,
            in3 => \N__30603\,
            lcout => \nx.n2164\,
            ltout => OPEN,
            carryin => \nx.n10876\,
            carryout => \nx.n10877\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1473_16_lut_LC_11_30_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41604\,
            in2 => \N__30600\,
            in3 => \N__30573\,
            lcout => \nx.n2163\,
            ltout => OPEN,
            carryin => \nx.n10877\,
            carryout => \nx.n10878\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1473_17_lut_LC_11_30_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41607\,
            in2 => \N__30569\,
            in3 => \N__30537\,
            lcout => \nx.n2162\,
            ltout => OPEN,
            carryin => \nx.n10878\,
            carryout => \nx.n10879\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1473_18_lut_LC_11_31_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41608\,
            in2 => \N__30894\,
            in3 => \N__30864\,
            lcout => \nx.n2161\,
            ltout => OPEN,
            carryin => \bfn_11_31_0_\,
            carryout => \nx.n10880\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1473_19_lut_LC_11_31_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001000001100000"
        )
    port map (
            in0 => \N__41609\,
            in1 => \N__30861\,
            in2 => \N__36561\,
            in3 => \N__30843\,
            lcout => \nx.n2192\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i2166_3_lut_LC_12_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__32856\,
            in1 => \_gnd_net_\,
            in2 => \N__34005\,
            in3 => \N__32884\,
            lcout => OPEN,
            ltout => \nx.n21_adj_750_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i1_4_lut_adj_93_LC_12_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110011111010"
        )
    port map (
            in0 => \N__33248\,
            in1 => \N__33222\,
            in2 => \N__30819\,
            in3 => \N__33977\,
            lcout => OPEN,
            ltout => \nx.n12781_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i1_4_lut_adj_97_LC_12_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111000"
        )
    port map (
            in0 => \N__30816\,
            in1 => \N__30743\,
            in2 => \N__30762\,
            in3 => \N__30990\,
            lcout => \nx.n12801\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i2163_3_lut_LC_12_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32727\,
            in2 => \N__32769\,
            in3 => \N__33967\,
            lcout => OPEN,
            ltout => \nx.n27_adj_744_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i1_4_lut_adj_89_LC_12_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110111111000"
        )
    port map (
            in0 => \N__33968\,
            in1 => \N__33306\,
            in2 => \N__30750\,
            in3 => \N__33329\,
            lcout => \nx.n12779\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i2172_3_lut_LC_12_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__32370\,
            in1 => \N__32412\,
            in2 => \_gnd_net_\,
            in3 => \N__33972\,
            lcout => \nx.n3209\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i2164_3_lut_LC_12_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32798\,
            in2 => \N__34004\,
            in3 => \N__32778\,
            lcout => OPEN,
            ltout => \nx.n25_adj_748_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i1_4_lut_adj_92_LC_12_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101011111100"
        )
    port map (
            in0 => \N__33180\,
            in1 => \N__33209\,
            in2 => \N__30993\,
            in3 => \N__33973\,
            lcout => \nx.n12785\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i1_4_lut_adj_88_LC_12_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101100"
        )
    port map (
            in0 => \N__32811\,
            in1 => \N__32833\,
            in2 => \N__34001\,
            in3 => \N__30984\,
            lcout => OPEN,
            ltout => \nx.n12777_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i1_4_lut_adj_91_LC_12_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101011111100"
        )
    port map (
            in0 => \N__32985\,
            in1 => \N__33005\,
            in2 => \N__30978\,
            in3 => \N__33962\,
            lcout => \nx.n12789\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i2157_3_lut_LC_12_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33141\,
            in2 => \N__34003\,
            in3 => \N__33163\,
            lcout => OPEN,
            ltout => \nx.n39_adj_747_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i1_4_lut_adj_95_LC_12_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__30951\,
            in1 => \N__30975\,
            in2 => \N__30969\,
            in3 => \N__30966\,
            lcout => \nx.n12799\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i2162_3_lut_LC_12_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33345\,
            in2 => \N__34002\,
            in3 => \N__33365\,
            lcout => \nx.n29_adj_746\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i2171_3_lut_LC_12_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32325\,
            in2 => \N__32354\,
            in3 => \N__33955\,
            lcout => \nx.n11_adj_751\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i2156_3_lut_LC_12_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33124\,
            in2 => \N__33105\,
            in3 => \N__33966\,
            lcout => \nx.n41_adj_752\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i2016_3_lut_LC_12_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35673\,
            in2 => \N__37103\,
            in3 => \N__37298\,
            lcout => \nx.n2989\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i2027_3_lut_LC_12_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35462\,
            in2 => \N__35430\,
            in3 => \N__37294\,
            lcout => \nx.n3000\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i2028_3_lut_LC_12_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35515\,
            in2 => \N__35481\,
            in3 => \N__37299\,
            lcout => \nx.n3001\,
            ltout => \nx.n3001_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i18_4_lut_adj_125_LC_12_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__31066\,
            in1 => \N__31048\,
            in2 => \N__31080\,
            in3 => \N__35836\,
            lcout => \nx.n44\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i2030_3_lut_LC_12_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37417\,
            in2 => \N__35001\,
            in3 => \N__37293\,
            lcout => \nx.n3003\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i2032_3_lut_LC_12_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101011001010"
        )
    port map (
            in0 => \N__35069\,
            in1 => \N__35040\,
            in2 => \N__37320\,
            in3 => \_gnd_net_\,
            lcout => \nx.n3005\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i14_4_lut_adj_113_LC_12_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__35560\,
            in1 => \N__35612\,
            in2 => \N__36904\,
            in3 => \N__35282\,
            lcout => \nx.n39_adj_761\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1954_3_lut_LC_12_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31138\,
            in2 => \N__31032\,
            in3 => \N__37588\,
            lcout => \nx.n2895\,
            ltout => \nx.n2895_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i2021_3_lut_LC_12_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35271\,
            in2 => \N__31017\,
            in3 => \N__37318\,
            lcout => \nx.n2994\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_2_lut_3_lut_adj_196_LC_12_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100000000"
        )
    port map (
            in0 => \N__43925\,
            in1 => \N__47594\,
            in2 => \_gnd_net_\,
            in3 => \N__43681\,
            lcout => n7992,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1957_3_lut_LC_12_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101000001010"
        )
    port map (
            in0 => \N__31439\,
            in1 => \_gnd_net_\,
            in2 => \N__37606\,
            in3 => \N__31413\,
            lcout => \nx.n2898\,
            ltout => \nx.n2898_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i2024_3_lut_LC_12_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__37319\,
            in1 => \_gnd_net_\,
            in2 => \N__31401\,
            in3 => \N__35319\,
            lcout => \nx.n2997\,
            ltout => \nx.n2997_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i19_4_lut_LC_12_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__33719\,
            in1 => \N__33745\,
            in2 => \N__31386\,
            in3 => \N__31369\,
            lcout => \nx.n45\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i2015_3_lut_LC_12_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35657\,
            in2 => \N__35637\,
            in3 => \N__37312\,
            lcout => \nx.n2988\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1946_3_lut_LC_12_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011110000"
        )
    port map (
            in0 => \N__31353\,
            in1 => \_gnd_net_\,
            in2 => \N__31341\,
            in3 => \N__37607\,
            lcout => \nx.n2887\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1815_3_lut_LC_12_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39471\,
            in2 => \N__39501\,
            in3 => \N__40106\,
            lcout => \nx.n2692\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1887_3_lut_LC_12_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31320\,
            in2 => \N__31308\,
            in3 => \N__31274\,
            lcout => \nx.n2796\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i16_4_lut_adj_16_LC_12_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__39251\,
            in1 => \N__39169\,
            in2 => \N__39306\,
            in3 => \N__39124\,
            lcout => \nx.n38\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1757_rep_22_3_lut_LC_12_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40374\,
            in2 => \N__40347\,
            in3 => \N__40914\,
            lcout => \nx.n2602\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1752_3_lut_LC_12_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40729\,
            in2 => \N__40927\,
            in3 => \N__40707\,
            lcout => \nx.n2597\,
            ltout => \nx.n2597_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i15_4_lut_adj_17_LC_12_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__39214\,
            in1 => \N__39727\,
            in2 => \N__31641\,
            in3 => \N__39079\,
            lcout => \nx.n37\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1814_3_lut_LC_12_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39453\,
            in2 => \N__39435\,
            in3 => \N__40079\,
            lcout => \nx.n2691\,
            ltout => \nx.n2691_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i13_4_lut_adj_24_LC_12_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__31459\,
            in1 => \N__31594\,
            in2 => \N__31578\,
            in3 => \N__31558\,
            lcout => \nx.n36\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i9151_3_lut_LC_12_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39173\,
            in2 => \N__39153\,
            in3 => \N__40078\,
            lcout => \nx.n2700\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1811_3_lut_LC_12_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101000001010"
        )
    port map (
            in0 => \N__39951\,
            in1 => \_gnd_net_\,
            in2 => \N__40091\,
            in3 => \N__40119\,
            lcout => \nx.n2688\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1812_3_lut_LC_12_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010101010"
        )
    port map (
            in0 => \N__40159\,
            in1 => \_gnd_net_\,
            in2 => \N__40134\,
            in3 => \N__40047\,
            lcout => \nx.n2689\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i12_4_lut_LC_12_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__40802\,
            in1 => \N__39400\,
            in2 => \N__40163\,
            in3 => \N__39950\,
            lcout => OPEN,
            ltout => \nx.n34_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i17_3_lut_LC_12_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39342\,
            in2 => \N__31443\,
            in3 => \N__39372\,
            lcout => OPEN,
            ltout => \nx.n39_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i21_4_lut_LC_12_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__31839\,
            in1 => \N__31830\,
            in2 => \N__31824\,
            in3 => \N__37146\,
            lcout => \nx.n2621\,
            ltout => \nx.n2621_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1831_rep_15_3_lut_LC_12_23_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__38844\,
            in1 => \_gnd_net_\,
            in2 => \N__31821\,
            in3 => \N__38865\,
            lcout => \nx.n2708\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1830_3_lut_LC_12_23_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38829\,
            in2 => \N__38802\,
            in3 => \N__40046\,
            lcout => \nx.n2707\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1560_3_lut_LC_12_24_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__31790\,
            in1 => \N__31746\,
            in2 => \_gnd_net_\,
            in3 => \N__32561\,
            lcout => \nx.n2309\,
            ltout => \nx.n2309_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i5904_2_lut_LC_12_24_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__31740\,
            in3 => \N__34329\,
            lcout => OPEN,
            ltout => \nx.n9697_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i13_4_lut_adj_54_LC_12_24_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__34528\,
            in1 => \N__37898\,
            in2 => \N__31737\,
            in3 => \N__34249\,
            lcout => \nx.n32_adj_698\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1556_3_lut_LC_12_24_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31734\,
            in2 => \N__32578\,
            in3 => \N__31728\,
            lcout => \nx.n2305\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1559_3_lut_LC_12_24_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31704\,
            in2 => \N__31677\,
            in3 => \N__32562\,
            lcout => \nx.n2308\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1818_3_lut_LC_12_24_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39648\,
            in2 => \N__39618\,
            in3 => \N__40076\,
            lcout => \nx.n2695\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1746_3_lut_LC_12_24_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40527\,
            in2 => \N__40500\,
            in3 => \N__40928\,
            lcout => \nx.n2591\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i14_4_lut_adj_55_LC_12_25_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__36415\,
            in1 => \N__34469\,
            in2 => \N__34572\,
            in3 => \N__34442\,
            lcout => \nx.n33_adj_699\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1554_3_lut_LC_12_25_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31956\,
            in2 => \N__31923\,
            in3 => \N__32572\,
            lcout => \nx.n2303\,
            ltout => \nx.n2303_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1621_3_lut_LC_12_25_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011110000"
        )
    port map (
            in0 => \N__34455\,
            in1 => \_gnd_net_\,
            in2 => \N__31914\,
            in3 => \N__37987\,
            lcout => \nx.n2402\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1552_3_lut_LC_12_25_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31911\,
            in2 => \N__32580\,
            in3 => \N__31905\,
            lcout => \nx.n2301\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1553_3_lut_LC_12_25_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31884\,
            in2 => \N__31854\,
            in3 => \N__32571\,
            lcout => \nx.n2302\,
            ltout => \nx.n2302_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1620_3_lut_LC_12_25_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011110000"
        )
    port map (
            in0 => \N__34428\,
            in1 => \_gnd_net_\,
            in2 => \N__31845\,
            in3 => \N__37988\,
            lcout => \nx.n2401\,
            ltout => \nx.n2401_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i14_4_lut_adj_58_LC_12_25_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__35936\,
            in1 => \N__36274\,
            in2 => \N__31842\,
            in3 => \N__36202\,
            lcout => \nx.n34_adj_701\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1612_3_lut_LC_12_26_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101000001010"
        )
    port map (
            in0 => \N__34678\,
            in1 => \_gnd_net_\,
            in2 => \N__38015\,
            in3 => \N__34656\,
            lcout => \nx.n2393\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1557_3_lut_LC_12_26_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__32112\,
            in1 => \_gnd_net_\,
            in2 => \N__32569\,
            in3 => \N__32105\,
            lcout => \nx.n2306\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1558_3_lut_LC_12_26_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010101010"
        )
    port map (
            in0 => \N__32073\,
            in1 => \_gnd_net_\,
            in2 => \N__32043\,
            in3 => \N__32538\,
            lcout => \nx.n2307\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1555_3_lut_LC_12_26_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__32031\,
            in1 => \_gnd_net_\,
            in2 => \N__32570\,
            in3 => \N__32024\,
            lcout => \nx.n2304\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1610_3_lut_LC_12_26_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34601\,
            in2 => \N__38016\,
            in3 => \N__34587\,
            lcout => \nx.n2391\,
            ltout => \nx.n2391_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i11_4_lut_adj_62_LC_12_26_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__36359\,
            in1 => \N__38573\,
            in2 => \N__31992\,
            in3 => \N__38518\,
            lcout => \nx.n31_adj_707\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i11_4_lut_adj_52_LC_12_26_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__36307\,
            in1 => \N__34643\,
            in2 => \N__34680\,
            in3 => \N__34717\,
            lcout => OPEN,
            ltout => \nx.n30_adj_696_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i15_4_lut_adj_53_LC_12_26_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__34600\,
            in1 => \N__34498\,
            in2 => \N__31989\,
            in3 => \N__34973\,
            lcout => \nx.n34_adj_697\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1549_3_lut_LC_12_27_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31986\,
            in2 => \N__31980\,
            in3 => \N__32554\,
            lcout => \nx.n2298\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1550_3_lut_LC_12_27_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31962\,
            in2 => \N__32577\,
            in3 => \N__36454\,
            lcout => \nx.n2299\,
            ltout => \nx.n2299_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i12_4_lut_adj_56_LC_12_27_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__34405\,
            in1 => \N__36664\,
            in2 => \N__32316\,
            in3 => \N__36631\,
            lcout => \nx.n31_adj_700\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1611_3_lut_LC_12_27_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101000001010"
        )
    port map (
            in0 => \N__34642\,
            in1 => \_gnd_net_\,
            in2 => \N__38021\,
            in3 => \N__34620\,
            lcout => \nx.n2392\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1548_3_lut_LC_12_27_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32132\,
            in2 => \N__32313\,
            in3 => \N__32553\,
            lcout => \nx.n2297\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i3_2_lut_LC_12_27_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32290\,
            in2 => \_gnd_net_\,
            in3 => \N__32270\,
            lcout => OPEN,
            ltout => \nx.n21_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i17_4_lut_adj_51_LC_12_27_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__32259\,
            in1 => \N__32253\,
            in2 => \N__32241\,
            in3 => \N__32238\,
            lcout => \nx.n2225\,
            ltout => \nx.n2225_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1551_3_lut_LC_12_27_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__32232\,
            in1 => \_gnd_net_\,
            in2 => \N__32226\,
            in3 => \N__32669\,
            lcout => \nx.n2300\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \neopxl_color_i4_LC_12_28_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0000000011101010"
        )
    port map (
            in0 => \N__32203\,
            in1 => \N__47693\,
            in2 => \N__43956\,
            in3 => \N__43711\,
            lcout => neopxl_color_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46916\,
            ce => 'H',
            sr => \N__32181\
        );

    \nx.mod_5_i1481_3_lut_LC_12_28_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32162\,
            in2 => \N__36564\,
            in3 => \N__32142\,
            lcout => \nx.n2198\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1484_3_lut_LC_12_28_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32718\,
            in2 => \N__32709\,
            in3 => \N__36553\,
            lcout => \nx.n2201\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1544_3_lut_LC_12_28_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32649\,
            in2 => \N__32576\,
            in3 => \N__32642\,
            lcout => \nx.n2293\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1545_3_lut_LC_12_28_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32622\,
            in2 => \N__32613\,
            in3 => \N__32552\,
            lcout => \nx.n2294\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pin_output_enable__i4_LC_13_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101100011001100"
        )
    port map (
            in0 => \N__37119\,
            in1 => \N__32462\,
            in2 => \N__47657\,
            in3 => \N__47072\,
            lcout => pin_oe_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46881\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i7633_2_lut_3_lut_4_lut_4_lut_LC_13_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111000000000"
        )
    port map (
            in0 => \N__42614\,
            in1 => \N__44106\,
            in2 => \N__45649\,
            in3 => \N__47549\,
            lcout => OPEN,
            ltout => \n11970_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pin_output_enable__i0_LC_13_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010110010101010"
        )
    port map (
            in0 => \N__32435\,
            in1 => \N__47581\,
            in2 => \N__32451\,
            in3 => \N__47146\,
            lcout => pin_oe_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46877\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i7631_3_lut_4_lut_4_lut_LC_13_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000001110000"
        )
    port map (
            in0 => \N__43429\,
            in1 => \N__45592\,
            in2 => \N__47635\,
            in3 => \N__42613\,
            lcout => n11968,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_2143_2_lut_LC_13_17_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32411\,
            in2 => \_gnd_net_\,
            in3 => \N__32361\,
            lcout => \nx.n3177\,
            ltout => OPEN,
            carryin => \bfn_13_17_0_\,
            carryout => \nx.n11079\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_2143_3_lut_LC_13_17_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__32358\,
            in3 => \N__32319\,
            lcout => \nx.n3176\,
            ltout => OPEN,
            carryin => \nx.n11079\,
            carryout => \nx.n11080\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_2143_4_lut_LC_13_17_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41308\,
            in2 => \N__33054\,
            in3 => \N__33015\,
            lcout => \nx.n3175\,
            ltout => OPEN,
            carryin => \nx.n11080\,
            carryout => \nx.n11081\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_2143_5_lut_LC_13_17_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41314\,
            in2 => \N__33012\,
            in3 => \N__32979\,
            lcout => \nx.n3174\,
            ltout => OPEN,
            carryin => \nx.n11081\,
            carryout => \nx.n11082\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_2143_6_lut_LC_13_17_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41309\,
            in2 => \N__32976\,
            in3 => \N__32934\,
            lcout => \nx.n3173\,
            ltout => OPEN,
            carryin => \nx.n11082\,
            carryout => \nx.n11083\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_2143_7_lut_LC_13_17_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41315\,
            in2 => \N__32931\,
            in3 => \N__32895\,
            lcout => \nx.n3172\,
            ltout => OPEN,
            carryin => \nx.n11083\,
            carryout => \nx.n11084\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_2143_8_lut_LC_13_17_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41310\,
            in2 => \N__32892\,
            in3 => \N__32850\,
            lcout => \nx.n3171\,
            ltout => OPEN,
            carryin => \nx.n11084\,
            carryout => \nx.n11085\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_2143_9_lut_LC_13_17_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32843\,
            in2 => \N__41638\,
            in3 => \N__32805\,
            lcout => \nx.n3170\,
            ltout => OPEN,
            carryin => \nx.n11085\,
            carryout => \nx.n11086\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_2143_10_lut_LC_13_18_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41472\,
            in2 => \N__32802\,
            in3 => \N__32772\,
            lcout => \nx.n3169\,
            ltout => OPEN,
            carryin => \bfn_13_18_0_\,
            carryout => \nx.n11087\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_2143_11_lut_LC_13_18_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41476\,
            in2 => \N__32768\,
            in3 => \N__32721\,
            lcout => \nx.n3168\,
            ltout => OPEN,
            carryin => \nx.n11087\,
            carryout => \nx.n11088\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_2143_12_lut_LC_13_18_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41473\,
            in2 => \N__33372\,
            in3 => \N__33339\,
            lcout => \nx.n3167\,
            ltout => OPEN,
            carryin => \nx.n11088\,
            carryout => \nx.n11089\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_2143_13_lut_LC_13_18_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41477\,
            in2 => \N__33336\,
            in3 => \N__33300\,
            lcout => \nx.n3166\,
            ltout => OPEN,
            carryin => \nx.n11089\,
            carryout => \nx.n11090\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_2143_14_lut_LC_13_18_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41474\,
            in2 => \N__33297\,
            in3 => \N__33255\,
            lcout => \nx.n3165\,
            ltout => OPEN,
            carryin => \nx.n11090\,
            carryout => \nx.n11091\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_2143_15_lut_LC_13_18_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41478\,
            in2 => \N__33252\,
            in3 => \N__33216\,
            lcout => \nx.n3164\,
            ltout => OPEN,
            carryin => \nx.n11091\,
            carryout => \nx.n11092\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_2143_16_lut_LC_13_18_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41475\,
            in2 => \N__33213\,
            in3 => \N__33174\,
            lcout => \nx.n3163\,
            ltout => OPEN,
            carryin => \nx.n11092\,
            carryout => \nx.n11093\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_2143_17_lut_LC_13_18_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41479\,
            in2 => \N__33171\,
            in3 => \N__33135\,
            lcout => \nx.n3162\,
            ltout => OPEN,
            carryin => \nx.n11093\,
            carryout => \nx.n11094\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_2143_18_lut_LC_13_19_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33132\,
            in2 => \N__41862\,
            in3 => \N__33096\,
            lcout => \nx.n3161\,
            ltout => OPEN,
            carryin => \bfn_13_19_0_\,
            carryout => \nx.n11095\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_2143_19_lut_LC_13_19_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41483\,
            in2 => \N__33093\,
            in3 => \N__33696\,
            lcout => \nx.n3160\,
            ltout => OPEN,
            carryin => \nx.n11095\,
            carryout => \nx.n11096\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_2143_20_lut_LC_13_19_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33693\,
            in2 => \N__41863\,
            in3 => \N__33651\,
            lcout => \nx.n3159\,
            ltout => OPEN,
            carryin => \nx.n11096\,
            carryout => \nx.n11097\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_2143_21_lut_LC_13_19_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33647\,
            in2 => \N__41866\,
            in3 => \N__33606\,
            lcout => \nx.n3158\,
            ltout => OPEN,
            carryin => \nx.n11097\,
            carryout => \nx.n11098\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_2143_22_lut_LC_13_19_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33602\,
            in2 => \N__41864\,
            in3 => \N__33561\,
            lcout => \nx.n3157\,
            ltout => OPEN,
            carryin => \nx.n11098\,
            carryout => \nx.n11099\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_2143_23_lut_LC_13_19_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33558\,
            in2 => \N__41867\,
            in3 => \N__33519\,
            lcout => \nx.n3156\,
            ltout => OPEN,
            carryin => \nx.n11099\,
            carryout => \nx.n11100\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_2143_24_lut_LC_13_19_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33515\,
            in2 => \N__41865\,
            in3 => \N__33471\,
            lcout => \nx.n3155\,
            ltout => OPEN,
            carryin => \nx.n11100\,
            carryout => \nx.n11101\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_2143_25_lut_LC_13_19_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33467\,
            in2 => \N__41868\,
            in3 => \N__33420\,
            lcout => \nx.n3154\,
            ltout => OPEN,
            carryin => \nx.n11101\,
            carryout => \nx.n11102\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_2143_26_lut_LC_13_20_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33413\,
            in2 => \N__42120\,
            in3 => \N__33375\,
            lcout => \nx.n3153\,
            ltout => OPEN,
            carryin => \bfn_13_20_0_\,
            carryout => \nx.n11103\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_2143_27_lut_LC_13_20_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34127\,
            in2 => \N__42122\,
            in3 => \N__34083\,
            lcout => \nx.n3152\,
            ltout => OPEN,
            carryin => \nx.n11103\,
            carryout => \nx.n11104\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_2143_28_lut_LC_13_20_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34079\,
            in2 => \N__42121\,
            in3 => \N__34035\,
            lcout => \nx.n3151\,
            ltout => OPEN,
            carryin => \nx.n11104\,
            carryout => \nx.n11105\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_2143_29_lut_LC_13_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__34026\,
            in1 => \N__41875\,
            in2 => \N__33891\,
            in3 => \N__33864\,
            lcout => \nx.n13280\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1963_3_lut_LC_13_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33849\,
            in2 => \N__33819\,
            in3 => \N__37579\,
            lcout => \nx.n2904\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1956_3_lut_LC_13_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33803\,
            in2 => \N__33771\,
            in3 => \N__37580\,
            lcout => \nx.n2897\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i2013_3_lut_LC_13_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35570\,
            in2 => \N__35547\,
            in3 => \N__37306\,
            lcout => \nx.n2986\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1826_rep_14_3_lut_LC_13_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39304\,
            in2 => \N__39273\,
            in3 => \N__40105\,
            lcout => \nx.n2703\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i2018_3_lut_LC_13_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35685\,
            in2 => \N__37725\,
            in3 => \N__37305\,
            lcout => \nx.n2991\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1755_3_lut_LC_13_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40263\,
            in2 => \N__40283\,
            in3 => \N__40907\,
            lcout => \nx.n2600\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1756_3_lut_LC_13_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40302\,
            in2 => \N__40922\,
            in3 => \N__40322\,
            lcout => \nx.n2601\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1758_3_lut_LC_13_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40389\,
            in2 => \N__40415\,
            in3 => \N__40903\,
            lcout => \nx.n2603\,
            ltout => \nx.n2603_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1825_3_lut_LC_13_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39237\,
            in2 => \N__34212\,
            in3 => \N__40077\,
            lcout => \nx.n2702\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1961_3_lut_LC_13_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34176\,
            in2 => \N__34149\,
            in3 => \N__37597\,
            lcout => \nx.n2902\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1685_3_lut_LC_13_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36099\,
            in2 => \N__36132\,
            in3 => \N__38478\,
            lcout => \nx.n2498\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1687_3_lut_LC_13_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36147\,
            in2 => \N__36174\,
            in3 => \N__38461\,
            lcout => \nx.n2500\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1688_3_lut_LC_13_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36186\,
            in2 => \N__38497\,
            in3 => \N__36212\,
            lcout => \nx.n2501\,
            ltout => \nx.n2501_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i6_3_lut_adj_110_LC_13_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101011110000"
        )
    port map (
            in0 => \N__39923\,
            in1 => \_gnd_net_\,
            in2 => \N__34134\,
            in3 => \N__39838\,
            lcout => \nx.n27_adj_757\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1694_3_lut_LC_13_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35979\,
            in2 => \N__36003\,
            in3 => \N__38456\,
            lcout => \nx.n2507\,
            ltout => \nx.n2507_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i15_4_lut_adj_109_LC_13_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__40321\,
            in1 => \N__40237\,
            in2 => \N__34215\,
            in3 => \N__40408\,
            lcout => \nx.n36_adj_756\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1689_rep_26_3_lut_LC_13_23_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36222\,
            in2 => \N__36249\,
            in3 => \N__38460\,
            lcout => \nx.n2502\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1691_3_lut_LC_13_23_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__35889\,
            in1 => \_gnd_net_\,
            in2 => \N__38496\,
            in3 => \N__35913\,
            lcout => \nx.n2504\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1690_3_lut_LC_13_24_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36258\,
            in2 => \N__36282\,
            in3 => \N__38474\,
            lcout => \nx.n2503\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1626_3_lut_LC_13_24_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34250\,
            in2 => \N__34230\,
            in3 => \N__37999\,
            lcout => \nx.n2407\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1614_3_lut_LC_13_24_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34695\,
            in2 => \N__34731\,
            in3 => \N__38000\,
            lcout => \nx.n2395\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1627_3_lut_LC_13_24_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34266\,
            in2 => \N__38017\,
            in3 => \N__34280\,
            lcout => \nx.n2408\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1628_3_lut_LC_13_24_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__34296\,
            in1 => \N__34333\,
            in2 => \_gnd_net_\,
            in3 => \N__37995\,
            lcout => \nx.n2409\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1623_3_lut_LC_13_25_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34509\,
            in2 => \N__34535\,
            in3 => \N__37967\,
            lcout => \nx.n2404\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1618_3_lut_LC_13_25_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34413\,
            in2 => \N__38008\,
            in3 => \N__34389\,
            lcout => \nx.n2399\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1624_3_lut_LC_13_25_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34570\,
            in2 => \N__34548\,
            in3 => \N__37968\,
            lcout => \nx.n2405\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1617_3_lut_LC_13_25_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101000001010"
        )
    port map (
            in0 => \N__34767\,
            in1 => \_gnd_net_\,
            in2 => \N__38010\,
            in3 => \N__34749\,
            lcout => \nx.n2398\,
            ltout => \nx.n2398_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i15_4_lut_adj_63_LC_13_25_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__35905\,
            in1 => \N__35995\,
            in2 => \N__34377\,
            in3 => \N__36238\,
            lcout => \nx.n35_adj_708\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1622_3_lut_LC_13_25_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101011001010"
        )
    port map (
            in0 => \N__34499\,
            in1 => \N__34479\,
            in2 => \N__38009\,
            in3 => \_gnd_net_\,
            lcout => \nx.n2403\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i18_4_lut_adj_57_LC_13_25_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__34374\,
            in1 => \N__34365\,
            in2 => \N__34359\,
            in3 => \N__34350\,
            lcout => \nx.n2324\,
            ltout => \nx.n2324_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1625_3_lut_LC_13_25_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36071\,
            in2 => \N__34344\,
            in3 => \N__37896\,
            lcout => \nx.n2406\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1607_2_lut_LC_13_26_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34341\,
            in2 => \_gnd_net_\,
            in3 => \N__34287\,
            lcout => \nx.n2377\,
            ltout => OPEN,
            carryin => \bfn_13_26_0_\,
            carryout => \nx.n10899\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1607_3_lut_LC_13_26_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__34284\,
            in3 => \N__34257\,
            lcout => \nx.n2376\,
            ltout => OPEN,
            carryin => \nx.n10899\,
            carryout => \nx.n10900\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1607_4_lut_LC_13_26_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41998\,
            in2 => \N__34254\,
            in3 => \N__34218\,
            lcout => \nx.n2375\,
            ltout => OPEN,
            carryin => \nx.n10900\,
            carryout => \nx.n10901\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1607_5_lut_LC_13_26_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42015\,
            in2 => \N__37897\,
            in3 => \N__34575\,
            lcout => \nx.n2374\,
            ltout => OPEN,
            carryin => \nx.n10901\,
            carryout => \nx.n10902\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1607_6_lut_LC_13_26_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34571\,
            in2 => \N__42210\,
            in3 => \N__34539\,
            lcout => \nx.n2373\,
            ltout => OPEN,
            carryin => \nx.n10902\,
            carryout => \nx.n10903\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1607_7_lut_LC_13_26_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42019\,
            in2 => \N__34536\,
            in3 => \N__34503\,
            lcout => \nx.n2372\,
            ltout => OPEN,
            carryin => \nx.n10903\,
            carryout => \nx.n10904\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1607_8_lut_LC_13_26_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41999\,
            in2 => \N__34500\,
            in3 => \N__34473\,
            lcout => \nx.n2371\,
            ltout => OPEN,
            carryin => \nx.n10904\,
            carryout => \nx.n10905\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1607_9_lut_LC_13_26_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42020\,
            in2 => \N__34470\,
            in3 => \N__34449\,
            lcout => \nx.n2370\,
            ltout => OPEN,
            carryin => \nx.n10905\,
            carryout => \nx.n10906\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1607_10_lut_LC_13_27_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42025\,
            in2 => \N__34446\,
            in3 => \N__34419\,
            lcout => \nx.n2369\,
            ltout => OPEN,
            carryin => \bfn_13_27_0_\,
            carryout => \nx.n10907\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1607_11_lut_LC_13_27_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41976\,
            in2 => \N__36422\,
            in3 => \N__34416\,
            lcout => \nx.n2368\,
            ltout => OPEN,
            carryin => \nx.n10907\,
            carryout => \nx.n10908\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1607_12_lut_LC_13_27_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42026\,
            in2 => \N__34412\,
            in3 => \N__34380\,
            lcout => \nx.n2367\,
            ltout => OPEN,
            carryin => \nx.n10908\,
            carryout => \nx.n10909\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1607_13_lut_LC_13_27_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34760\,
            in2 => \N__42211\,
            in3 => \N__34740\,
            lcout => \nx.n2366\,
            ltout => OPEN,
            carryin => \nx.n10909\,
            carryout => \nx.n10910\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1607_14_lut_LC_13_27_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42030\,
            in2 => \N__36638\,
            in3 => \N__34737\,
            lcout => \nx.n2365\,
            ltout => OPEN,
            carryin => \nx.n10910\,
            carryout => \nx.n10911\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1607_15_lut_LC_13_27_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41977\,
            in2 => \N__36671\,
            in3 => \N__34734\,
            lcout => \nx.n2364\,
            ltout => OPEN,
            carryin => \nx.n10911\,
            carryout => \nx.n10912\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1607_16_lut_LC_13_27_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42031\,
            in2 => \N__34730\,
            in3 => \N__34686\,
            lcout => \nx.n2363\,
            ltout => OPEN,
            carryin => \nx.n10912\,
            carryout => \nx.n10913\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1607_17_lut_LC_13_27_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41978\,
            in2 => \N__36318\,
            in3 => \N__34683\,
            lcout => \nx.n2362\,
            ltout => OPEN,
            carryin => \nx.n10913\,
            carryout => \nx.n10914\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1607_18_lut_LC_13_28_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42212\,
            in2 => \N__34679\,
            in3 => \N__34647\,
            lcout => \nx.n2361\,
            ltout => OPEN,
            carryin => \bfn_13_28_0_\,
            carryout => \nx.n10915\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1607_19_lut_LC_13_28_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42215\,
            in2 => \N__34644\,
            in3 => \N__34614\,
            lcout => \nx.n2360\,
            ltout => OPEN,
            carryin => \nx.n10915\,
            carryout => \nx.n10916\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1607_20_lut_LC_13_28_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42213\,
            in2 => \N__34611\,
            in3 => \N__34578\,
            lcout => \nx.n2359\,
            ltout => OPEN,
            carryin => \nx.n10916\,
            carryout => \nx.n10917\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1607_21_lut_LC_13_28_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000010001001000"
        )
    port map (
            in0 => \N__42214\,
            in1 => \N__38004\,
            in2 => \N__34983\,
            in3 => \N__34962\,
            lcout => \nx.n2390\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i2031_3_lut_LC_14_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35028\,
            in2 => \N__35013\,
            in3 => \N__37255\,
            lcout => \nx.n3004\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i2033_3_lut_LC_14_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35079\,
            in2 => \N__37304\,
            in3 => \N__35106\,
            lcout => \nx.n3006\,
            ltout => \nx.n3006_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i17_4_lut_LC_14_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__34936\,
            in1 => \N__34895\,
            in2 => \N__34923\,
            in3 => \N__36871\,
            lcout => \nx.n43\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i2026_3_lut_LC_14_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35412\,
            in2 => \N__37303\,
            in3 => \N__35382\,
            lcout => \nx.n2999\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1955_3_lut_LC_14_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34884\,
            in2 => \N__37608\,
            in3 => \N__34851\,
            lcout => \nx.n2896\,
            ltout => \nx.n2896_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i18_4_lut_adj_115_LC_14_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__35151\,
            in1 => \N__35369\,
            in2 => \N__34836\,
            in3 => \N__35105\,
            lcout => OPEN,
            ltout => \nx.n43_adj_763_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i22_4_lut_adj_123_LC_14_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__36803\,
            in1 => \N__35027\,
            in2 => \N__34833\,
            in3 => \N__34830\,
            lcout => \nx.n47_adj_770\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1964_3_lut_LC_14_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34818\,
            in2 => \N__34785\,
            in3 => \N__37598\,
            lcout => \nx.n2905\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_2009_2_lut_LC_14_19_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35258\,
            in2 => \_gnd_net_\,
            in3 => \N__35193\,
            lcout => \nx.n2977\,
            ltout => OPEN,
            carryin => \bfn_14_19_0_\,
            carryout => \nx.n11028\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_2009_3_lut_LC_14_19_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__35190\,
            in3 => \N__35154\,
            lcout => \nx.n2976\,
            ltout => OPEN,
            carryin => \nx.n11028\,
            carryout => \nx.n11029\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_2009_4_lut_LC_14_19_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41316\,
            in2 => \N__35146\,
            in3 => \N__35109\,
            lcout => \nx.n2975\,
            ltout => OPEN,
            carryin => \nx.n11029\,
            carryout => \nx.n11030\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_2009_5_lut_LC_14_19_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41322\,
            in2 => \N__35099\,
            in3 => \N__35073\,
            lcout => \nx.n2974\,
            ltout => OPEN,
            carryin => \nx.n11030\,
            carryout => \nx.n11031\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_2009_6_lut_LC_14_19_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41317\,
            in2 => \N__35070\,
            in3 => \N__35031\,
            lcout => \nx.n2973\,
            ltout => OPEN,
            carryin => \nx.n11031\,
            carryout => \nx.n11032\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_2009_7_lut_LC_14_19_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35026\,
            in2 => \N__41639\,
            in3 => \N__35004\,
            lcout => \nx.n2972\,
            ltout => OPEN,
            carryin => \nx.n11032\,
            carryout => \nx.n11033\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_2009_8_lut_LC_14_19_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41321\,
            in2 => \N__37418\,
            in3 => \N__34989\,
            lcout => \nx.n2971\,
            ltout => OPEN,
            carryin => \nx.n11033\,
            carryout => \nx.n11034\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_2009_9_lut_LC_14_19_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41323\,
            in2 => \N__36802\,
            in3 => \N__34986\,
            lcout => \nx.n2970\,
            ltout => OPEN,
            carryin => \nx.n11034\,
            carryout => \nx.n11035\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_2009_10_lut_LC_14_20_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41640\,
            in2 => \N__35516\,
            in3 => \N__35466\,
            lcout => \nx.n2969\,
            ltout => OPEN,
            carryin => \bfn_14_20_0_\,
            carryout => \nx.n11036\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_2009_11_lut_LC_14_20_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41644\,
            in2 => \N__35463\,
            in3 => \N__35415\,
            lcout => \nx.n2968\,
            ltout => OPEN,
            carryin => \nx.n11036\,
            carryout => \nx.n11037\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_2009_12_lut_LC_14_20_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41641\,
            in2 => \N__35411\,
            in3 => \N__35373\,
            lcout => \nx.n2967\,
            ltout => OPEN,
            carryin => \nx.n11037\,
            carryout => \nx.n11038\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_2009_13_lut_LC_14_20_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41645\,
            in2 => \N__35370\,
            in3 => \N__35322\,
            lcout => \nx.n2966\,
            ltout => OPEN,
            carryin => \nx.n11038\,
            carryout => \nx.n11039\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_2009_14_lut_LC_14_20_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41642\,
            in2 => \N__37437\,
            in3 => \N__35310\,
            lcout => \nx.n2965\,
            ltout => OPEN,
            carryin => \nx.n11039\,
            carryout => \nx.n11040\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_2009_15_lut_LC_14_20_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41646\,
            in2 => \N__37381\,
            in3 => \N__35295\,
            lcout => \nx.n2964\,
            ltout => OPEN,
            carryin => \nx.n11040\,
            carryout => \nx.n11041\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_2009_16_lut_LC_14_20_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41643\,
            in2 => \N__37011\,
            in3 => \N__35292\,
            lcout => \nx.n2963\,
            ltout => OPEN,
            carryin => \nx.n11041\,
            carryout => \nx.n11042\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_2009_17_lut_LC_14_20_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41647\,
            in2 => \N__35289\,
            in3 => \N__35262\,
            lcout => \nx.n2962\,
            ltout => OPEN,
            carryin => \nx.n11042\,
            carryout => \nx.n11043\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_2009_18_lut_LC_14_21_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41648\,
            in2 => \N__37353\,
            in3 => \N__35691\,
            lcout => \nx.n2961\,
            ltout => OPEN,
            carryin => \bfn_14_21_0_\,
            carryout => \nx.n11044\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_2009_19_lut_LC_14_21_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37448\,
            in2 => \N__41997\,
            in3 => \N__35688\,
            lcout => \nx.n2960\,
            ltout => OPEN,
            carryin => \nx.n11044\,
            carryout => \nx.n11045\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_2009_20_lut_LC_14_21_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41652\,
            in2 => \N__37718\,
            in3 => \N__35679\,
            lcout => \nx.n2959\,
            ltout => OPEN,
            carryin => \nx.n11045\,
            carryout => \nx.n11046\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_2009_21_lut_LC_14_21_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41655\,
            in2 => \N__36915\,
            in3 => \N__35676\,
            lcout => \nx.n2958\,
            ltout => OPEN,
            carryin => \nx.n11046\,
            carryout => \nx.n11047\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_2009_22_lut_LC_14_21_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41653\,
            in2 => \N__37107\,
            in3 => \N__35661\,
            lcout => \nx.n2957\,
            ltout => OPEN,
            carryin => \nx.n11047\,
            carryout => \nx.n11048\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_2009_23_lut_LC_14_21_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41656\,
            in2 => \N__35658\,
            in3 => \N__35625\,
            lcout => \nx.n2956\,
            ltout => OPEN,
            carryin => \nx.n11048\,
            carryout => \nx.n11049\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_2009_24_lut_LC_14_21_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41654\,
            in2 => \N__35622\,
            in3 => \N__35574\,
            lcout => \nx.n2955\,
            ltout => OPEN,
            carryin => \nx.n11049\,
            carryout => \nx.n11050\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_2009_25_lut_LC_14_21_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41657\,
            in2 => \N__35571\,
            in3 => \N__35538\,
            lcout => \nx.n2954\,
            ltout => OPEN,
            carryin => \nx.n11050\,
            carryout => \nx.n11051\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_2009_26_lut_LC_14_22_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41679\,
            in2 => \N__35535\,
            in3 => \N__35874\,
            lcout => \nx.n2953\,
            ltout => OPEN,
            carryin => \bfn_14_22_0_\,
            carryout => \nx.n11052\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_2009_27_lut_LC_14_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000010001001000"
        )
    port map (
            in0 => \N__41680\,
            in1 => \N__37263\,
            in2 => \N__35871\,
            in3 => \N__35847\,
            lcout => \nx.n2984\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i18_4_lut_adj_128_LC_14_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__35817\,
            in1 => \N__35811\,
            in2 => \N__40203\,
            in3 => \N__40373\,
            lcout => \nx.n39_adj_773\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i16_4_lut_adj_42_LC_14_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__35804\,
            in1 => \N__35764\,
            in2 => \N__37846\,
            in3 => \N__37804\,
            lcout => \nx.n39_adj_689\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1754_rep_17_3_lut_LC_14_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40241\,
            in2 => \N__40221\,
            in3 => \N__40902\,
            lcout => \nx.n2599\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i12_4_lut_adj_60_LC_14_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__38104\,
            in1 => \N__38254\,
            in2 => \N__36131\,
            in3 => \N__38173\,
            lcout => \nx.n32_adj_703\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i5_3_lut_adj_59_LC_14_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101011110000"
        )
    port map (
            in0 => \N__36058\,
            in1 => \_gnd_net_\,
            in2 => \N__35970\,
            in3 => \N__38317\,
            lcout => OPEN,
            ltout => \nx.n25_adj_702_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i17_4_lut_adj_64_LC_14_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__38290\,
            in1 => \N__38143\,
            in2 => \N__35736\,
            in3 => \N__35733\,
            lcout => OPEN,
            ltout => \nx.n37_adj_709_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i19_4_lut_adj_65_LC_14_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__35721\,
            in1 => \N__35712\,
            in2 => \N__35706\,
            in3 => \N__35703\,
            lcout => \nx.n2423\,
            ltout => \nx.n2423_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1696_3_lut_LC_14_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36059\,
            in2 => \N__36078\,
            in3 => \N__36015\,
            lcout => \nx.n2509\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1693_3_lut_LC_14_23_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35949\,
            in2 => \N__38498\,
            in3 => \N__35968\,
            lcout => \nx.n2506\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1625_rep_29_3_lut_LC_14_23_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36075\,
            in2 => \N__35925\,
            in3 => \N__38465\,
            lcout => \nx.n13321\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1674_2_lut_LC_14_24_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36057\,
            in2 => \_gnd_net_\,
            in3 => \N__36009\,
            lcout => \nx.n2477\,
            ltout => OPEN,
            carryin => \bfn_14_24_0_\,
            carryout => \nx.n10918\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1674_3_lut_LC_14_24_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__38321\,
            in3 => \N__36006\,
            lcout => \nx.n2476\,
            ltout => OPEN,
            carryin => \nx.n10918\,
            carryout => \nx.n10919\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1674_4_lut_LC_14_24_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42009\,
            in2 => \N__36002\,
            in3 => \N__35973\,
            lcout => \nx.n2475\,
            ltout => OPEN,
            carryin => \nx.n10919\,
            carryout => \nx.n10920\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1674_5_lut_LC_14_24_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42012\,
            in2 => \N__35969\,
            in3 => \N__35943\,
            lcout => \nx.n2474\,
            ltout => OPEN,
            carryin => \nx.n10920\,
            carryout => \nx.n10921\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1674_6_lut_LC_14_24_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42010\,
            in2 => \N__35940\,
            in3 => \N__35916\,
            lcout => \nx.n2473\,
            ltout => OPEN,
            carryin => \nx.n10921\,
            carryout => \nx.n10922\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1674_7_lut_LC_14_24_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42013\,
            in2 => \N__35912\,
            in3 => \N__36285\,
            lcout => \nx.n2472\,
            ltout => OPEN,
            carryin => \nx.n10922\,
            carryout => \nx.n10923\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1674_8_lut_LC_14_24_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42011\,
            in2 => \N__36281\,
            in3 => \N__36252\,
            lcout => \nx.n2471\,
            ltout => OPEN,
            carryin => \nx.n10923\,
            carryout => \nx.n10924\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1674_9_lut_LC_14_24_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42014\,
            in2 => \N__36245\,
            in3 => \N__36216\,
            lcout => \nx.n2470\,
            ltout => OPEN,
            carryin => \nx.n10924\,
            carryout => \nx.n10925\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1674_10_lut_LC_14_25_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42000\,
            in2 => \N__36213\,
            in3 => \N__36177\,
            lcout => \nx.n2469\,
            ltout => OPEN,
            carryin => \bfn_14_25_0_\,
            carryout => \nx.n10926\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1674_11_lut_LC_14_25_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42021\,
            in2 => \N__36170\,
            in3 => \N__36138\,
            lcout => \nx.n2468\,
            ltout => OPEN,
            carryin => \nx.n10926\,
            carryout => \nx.n10927\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1674_12_lut_LC_14_25_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42001\,
            in2 => \N__38297\,
            in3 => \N__36135\,
            lcout => \nx.n2467\,
            ltout => OPEN,
            carryin => \nx.n10927\,
            carryout => \nx.n10928\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1674_13_lut_LC_14_25_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42022\,
            in2 => \N__36127\,
            in3 => \N__36087\,
            lcout => \nx.n2466\,
            ltout => OPEN,
            carryin => \nx.n10928\,
            carryout => \nx.n10929\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1674_14_lut_LC_14_25_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42002\,
            in2 => \N__38204\,
            in3 => \N__36084\,
            lcout => \nx.n2465\,
            ltout => OPEN,
            carryin => \nx.n10929\,
            carryout => \nx.n10930\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1674_15_lut_LC_14_25_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42023\,
            in2 => \N__38148\,
            in3 => \N__36081\,
            lcout => \nx.n2464\,
            ltout => OPEN,
            carryin => \nx.n10930\,
            carryout => \nx.n10931\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1674_16_lut_LC_14_25_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42003\,
            in2 => \N__38259\,
            in3 => \N__36381\,
            lcout => \nx.n2463\,
            ltout => OPEN,
            carryin => \nx.n10931\,
            carryout => \nx.n10932\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1674_17_lut_LC_14_25_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42024\,
            in2 => \N__38180\,
            in3 => \N__36378\,
            lcout => \nx.n2462\,
            ltout => OPEN,
            carryin => \nx.n10932\,
            carryout => \nx.n10933\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1674_18_lut_LC_14_26_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42004\,
            in2 => \N__38105\,
            in3 => \N__36375\,
            lcout => \nx.n2461\,
            ltout => OPEN,
            carryin => \bfn_14_26_0_\,
            carryout => \nx.n10934\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1674_19_lut_LC_14_26_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42032\,
            in2 => \N__38531\,
            in3 => \N__36372\,
            lcout => \nx.n2460\,
            ltout => OPEN,
            carryin => \nx.n10934\,
            carryout => \nx.n10935\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1674_20_lut_LC_14_26_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42005\,
            in2 => \N__38591\,
            in3 => \N__36369\,
            lcout => \nx.n2459\,
            ltout => OPEN,
            carryin => \nx.n10935\,
            carryout => \nx.n10936\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1674_21_lut_LC_14_26_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38054\,
            in2 => \N__42209\,
            in3 => \N__36366\,
            lcout => \nx.n2458\,
            ltout => OPEN,
            carryin => \nx.n10936\,
            carryout => \nx.n10937\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1674_22_lut_LC_14_26_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000010001001000"
        )
    port map (
            in0 => \N__42033\,
            in1 => \N__38500\,
            in2 => \N__36363\,
            in3 => \N__36342\,
            lcout => \nx.n2489\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pin_output_enable__i18_LC_14_26_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101100011001100"
        )
    port map (
            in0 => \N__38964\,
            in1 => \N__36329\,
            in2 => \N__47694\,
            in3 => \N__47154\,
            lcout => pin_oe_18,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46917\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1613_3_lut_LC_14_27_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36317\,
            in2 => \N__36294\,
            in3 => \N__38011\,
            lcout => \nx.n2394\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1615_3_lut_LC_14_27_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36672\,
            in2 => \N__36648\,
            in3 => \N__38012\,
            lcout => \nx.n2396\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1616_3_lut_LC_14_27_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010011100100"
        )
    port map (
            in0 => \N__38014\,
            in1 => \N__36639\,
            in2 => \N__36615\,
            in3 => \_gnd_net_\,
            lcout => \nx.n2397\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1483_3_lut_LC_14_27_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36606\,
            in2 => \N__36594\,
            in3 => \N__36562\,
            lcout => \nx.n2200\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1619_3_lut_LC_14_27_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010011100100"
        )
    port map (
            in0 => \N__38013\,
            in1 => \N__36423\,
            in2 => \N__36396\,
            in3 => \_gnd_net_\,
            lcout => \nx.n2400\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \state__i0_LC_15_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47325\,
            in2 => \N__43191\,
            in3 => \N__43822\,
            lcout => state_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46893\,
            ce => \N__42399\,
            sr => \N__38390\
        );

    \state__i2_LC_15_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000100000000"
        )
    port map (
            in0 => \N__47324\,
            in1 => \N__43186\,
            in2 => \_gnd_net_\,
            in3 => \N__43823\,
            lcout => state_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46893\,
            ce => \N__42399\,
            sr => \N__38390\
        );

    \i1_2_lut_LC_15_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101010101"
        )
    port map (
            in0 => \N__43817\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__43584\,
            lcout => n7602,
            ltout => \n7602_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_3_lut_4_lut_adj_195_LC_15_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011000100"
        )
    port map (
            in0 => \N__36729\,
            in1 => \N__45902\,
            in2 => \N__36387\,
            in3 => \N__47299\,
            lcout => n7730,
            ltout => \n7730_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pin_output_enable__i9_LC_15_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101100"
        )
    port map (
            in0 => \N__47301\,
            in1 => \N__36767\,
            in2 => \N__36384\,
            in3 => \N__42381\,
            lcout => pin_oe_9,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46888\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pin_output_enable__i10_LC_15_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011100010101010"
        )
    port map (
            in0 => \N__36746\,
            in1 => \N__36735\,
            in2 => \N__47431\,
            in3 => \N__47039\,
            lcout => pin_oe_10,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46888\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i7623_2_lut_3_lut_4_lut_4_lut_LC_15_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011001000"
        )
    port map (
            in0 => \N__44430\,
            in1 => \N__47300\,
            in2 => \N__45681\,
            in3 => \N__44532\,
            lcout => n11960,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i308_2_lut_LC_15_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38627\,
            in2 => \_gnd_net_\,
            in3 => \N__43184\,
            lcout => n2618,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pin_output_enable__i3_LC_15_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010001011100010"
        )
    port map (
            in0 => \N__36713\,
            in1 => \N__47038\,
            in2 => \N__47577\,
            in3 => \N__38646\,
            lcout => pin_oe_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46885\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_2_lut_3_lut_4_lut_adj_164_LC_15_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011001101"
        )
    port map (
            in0 => \N__44968\,
            in1 => \N__44831\,
            in2 => \N__45664\,
            in3 => \N__44503\,
            lcout => OPEN,
            ltout => \n8_adj_825_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pin_output_i0_i9_LC_15_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111100100000"
        )
    port map (
            in0 => \N__45898\,
            in1 => \N__46147\,
            in2 => \N__36702\,
            in3 => \N__36689\,
            lcout => pin_out_9,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46880\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i9176_2_lut_3_lut_4_lut_3_lut_LC_15_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001100110"
        )
    port map (
            in0 => \N__43836\,
            in1 => \N__47367\,
            in2 => \_gnd_net_\,
            in3 => \N__43596\,
            lcout => n11789,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i8974_3_lut_LC_15_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__46385\,
            in1 => \N__36688\,
            in2 => \_gnd_net_\,
            in3 => \N__43340\,
            lcout => n13369,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \equal_240_i6_2_lut_LC_15_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46564\,
            in2 => \_gnd_net_\,
            in3 => \N__46386\,
            lcout => n6_adj_813,
            ltout => \n6_adj_813_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i7637_2_lut_3_lut_4_lut_4_lut_LC_15_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100100011001100"
        )
    port map (
            in0 => \N__42578\,
            in1 => \N__47590\,
            in2 => \N__37122\,
            in3 => \N__45627\,
            lcout => n11974,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i20_4_lut_adj_122_LC_15_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__37714\,
            in1 => \N__37102\,
            in2 => \N__37065\,
            in3 => \N__37047\,
            lcout => OPEN,
            ltout => \nx.n45_adj_769_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i24_4_lut_adj_124_LC_15_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__37359\,
            in1 => \N__37035\,
            in2 => \N__37020\,
            in3 => \N__37017\,
            lcout => \nx.n2918\,
            ltout => \nx.n2918_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i2022_3_lut_LC_15_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37007\,
            in2 => \N__36993\,
            in3 => \N__36990\,
            lcout => \nx.n2995\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i2029_3_lut_LC_15_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36984\,
            in2 => \N__36804\,
            in3 => \N__37262\,
            lcout => \nx.n3002\,
            ltout => \nx.n3002_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i16_4_lut_LC_15_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__36947\,
            in1 => \N__37159\,
            in2 => \N__36936\,
            in3 => \N__37673\,
            lcout => \nx.n42\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i2017_3_lut_LC_15_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36921\,
            in2 => \N__36911\,
            in3 => \N__37227\,
            lcout => \nx.n2990\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1962_3_lut_LC_15_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36849\,
            in2 => \N__36822\,
            in3 => \N__37603\,
            lcout => \nx.n2903\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1951_3_lut_LC_15_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37773\,
            in2 => \N__37743\,
            in3 => \N__37605\,
            lcout => \nx.n2892\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i2019_3_lut_LC_15_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37449\,
            in2 => \N__37695\,
            in3 => \N__37231\,
            lcout => \nx.n2992\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1952_3_lut_LC_15_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37662\,
            in2 => \N__37626\,
            in3 => \N__37604\,
            lcout => \nx.n2893\,
            ltout => \nx.n2893_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i16_4_lut_adj_121_LC_15_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__37436\,
            in1 => \N__37419\,
            in2 => \N__37395\,
            in3 => \N__37382\,
            lcout => \nx.n41_adj_768\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i2020_3_lut_LC_15_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37349\,
            in2 => \N__37276\,
            in3 => \N__37173\,
            lcout => \nx.n2993\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i18_4_lut_LC_15_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__38821\,
            in1 => \N__39592\,
            in2 => \N__37131\,
            in3 => \N__38067\,
            lcout => \nx.n40\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1764_3_lut_LC_15_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__39927\,
            in1 => \N__39864\,
            in2 => \_gnd_net_\,
            in3 => \N__40894\,
            lcout => \nx.n2609\,
            ltout => \nx.n2609_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i6_3_lut_adj_155_LC_15_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110100000"
        )
    port map (
            in0 => \N__38927\,
            in1 => \_gnd_net_\,
            in2 => \N__37134\,
            in3 => \N__39643\,
            lcout => \nx.n28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1761_3_lut_LC_15_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39747\,
            in2 => \N__39774\,
            in3 => \N__40898\,
            lcout => \nx.n2606\,
            ltout => \nx.n2606_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1828_3_lut_LC_15_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39351\,
            in2 => \N__37860\,
            in3 => \N__40101\,
            lcout => \nx.n2705\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1763_3_lut_LC_15_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39819\,
            in2 => \N__40921\,
            in3 => \N__39848\,
            lcout => \nx.n2608\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1827_3_lut_LC_15_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39337\,
            in2 => \N__40107\,
            in3 => \N__39315\,
            lcout => \nx.n2704\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1762_3_lut_LC_15_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39806\,
            in2 => \N__39789\,
            in3 => \N__40863\,
            lcout => \nx.n2607\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i16_4_lut_adj_126_LC_15_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__39805\,
            in1 => \N__40474\,
            in2 => \N__40446\,
            in3 => \N__38028\,
            lcout => OPEN,
            ltout => \nx.n37_adj_772_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i20_4_lut_adj_141_LC_15_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__38217\,
            in1 => \N__38550\,
            in2 => \N__37785\,
            in3 => \N__37782\,
            lcout => \nx.n2522\,
            ltout => \nx.n2522_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1760_3_lut_LC_15_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40458\,
            in2 => \N__37776\,
            in3 => \N__40475\,
            lcout => \nx.n2605\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1753_3_lut_LC_15_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101000001010"
        )
    port map (
            in0 => \N__40201\,
            in1 => \_gnd_net_\,
            in2 => \N__40900\,
            in3 => \N__40176\,
            lcout => \nx.n2598\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1747_3_lut_LC_15_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40864\,
            in2 => \N__40569\,
            in3 => \N__40542\,
            lcout => \nx.n2592\,
            ltout => \nx.n2592_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i13_4_lut_LC_15_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__38773\,
            in1 => \N__39538\,
            in2 => \N__38070\,
            in3 => \N__39487\,
            lcout => \nx.n35\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1677_3_lut_LC_15_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38061\,
            in2 => \N__38499\,
            in3 => \N__38040\,
            lcout => \nx.n2490\,
            ltout => \nx.n2490_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i1_2_lut_adj_108_LC_15_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__38031\,
            in3 => \N__40946\,
            lcout => \nx.n22_adj_755\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1749_3_lut_LC_15_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40637\,
            in2 => \N__40623\,
            in3 => \N__40861\,
            lcout => \nx.n2594\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1748_3_lut_LC_15_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__40860\,
            in1 => \_gnd_net_\,
            in2 => \N__40584\,
            in3 => \N__40604\,
            lcout => \nx.n2593\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1751_3_lut_LC_15_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40692\,
            in2 => \N__40674\,
            in3 => \N__40859\,
            lcout => \nx.n2596\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i9121_3_lut_4_lut_LC_15_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111000010000"
        )
    port map (
            in0 => \N__38022\,
            in1 => \N__38470\,
            in2 => \N__37905\,
            in3 => \N__37869\,
            lcout => \nx.n2505\,
            ltout => \nx.n2505_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1759_3_lut_LC_15_23_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011110000"
        )
    port map (
            in0 => \N__40428\,
            in1 => \_gnd_net_\,
            in2 => \N__37863\,
            in3 => \N__40862\,
            lcout => \nx.n2604\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1695_3_lut_LC_15_23_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011110000"
        )
    port map (
            in0 => \N__38334\,
            in1 => \_gnd_net_\,
            in2 => \N__38328\,
            in3 => \N__38469\,
            lcout => \nx.n2508\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1686_3_lut_LC_15_24_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38298\,
            in2 => \N__38268\,
            in3 => \N__38492\,
            lcout => \nx.n2499\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1682_3_lut_LC_15_24_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101000001010"
        )
    port map (
            in0 => \N__38258\,
            in1 => \_gnd_net_\,
            in2 => \N__38505\,
            in3 => \N__38229\,
            lcout => \nx.n2495\,
            ltout => \nx.n2495_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i13_4_lut_adj_111_LC_15_24_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__40658\,
            in1 => \N__40690\,
            in2 => \N__38220\,
            in3 => \N__40736\,
            lcout => \nx.n34_adj_758\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1684_3_lut_LC_15_24_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38208\,
            in2 => \N__38504\,
            in3 => \N__38187\,
            lcout => \nx.n2497\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1681_3_lut_LC_15_24_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38181\,
            in2 => \N__38157\,
            in3 => \N__38487\,
            lcout => \nx.n2494\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1683_3_lut_LC_15_24_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010101010"
        )
    port map (
            in0 => \N__38147\,
            in1 => \_gnd_net_\,
            in2 => \N__38118\,
            in3 => \N__38488\,
            lcout => \nx.n2496\,
            ltout => \nx.n2496_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1750_3_lut_LC_15_24_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011110000"
        )
    port map (
            in0 => \N__40647\,
            in1 => \_gnd_net_\,
            in2 => \N__38109\,
            in3 => \N__40901\,
            lcout => \nx.n2595\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1680_3_lut_LC_15_25_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38106\,
            in2 => \N__38079\,
            in3 => \N__38502\,
            lcout => \nx.n2493\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pin_output_enable__i22_LC_15_25_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101000011001100"
        )
    port map (
            in0 => \N__42663\,
            in1 => \N__38603\,
            in2 => \N__47695\,
            in3 => \N__47155\,
            lcout => pin_oe_22,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46918\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1678_3_lut_LC_15_25_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38592\,
            in2 => \N__38562\,
            in3 => \N__38503\,
            lcout => \nx.n2491\,
            ltout => \nx.n2491_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i12_4_lut_adj_120_LC_15_25_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__40516\,
            in1 => \N__40600\,
            in2 => \N__38553\,
            in3 => \N__40558\,
            lcout => \nx.n33_adj_767\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1679_3_lut_LC_15_26_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38541\,
            in2 => \N__38535\,
            in3 => \N__38501\,
            lcout => \nx.n2492\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1745_3_lut_LC_15_26_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40926\,
            in2 => \N__42363\,
            in3 => \N__42345\,
            lcout => \nx.n2590\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \state__i1_LC_16_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100101000001010"
        )
    port map (
            in0 => \N__47323\,
            in1 => \N__38631\,
            in2 => \N__43875\,
            in3 => \N__43190\,
            lcout => state_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46897\,
            ce => \N__42398\,
            sr => \N__38391\
        );

    \counter_633__i0_LC_16_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000000100"
        )
    port map (
            in0 => \N__38370\,
            in1 => \N__40758\,
            in2 => \N__47459\,
            in3 => \N__42888\,
            lcout => counter_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46894\,
            ce => \N__45961\,
            sr => \_gnd_net_\
        );

    \pin_output_enable__i11_LC_16_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100010011100100"
        )
    port map (
            in0 => \N__47037\,
            in1 => \N__38345\,
            in2 => \N__47489\,
            in3 => \N__44219\,
            lcout => pin_oe_11,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46889\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \equal_243_i6_2_lut_LC_16_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46509\,
            in2 => \_gnd_net_\,
            in3 => \N__46321\,
            lcout => n6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_2_lut_3_lut_4_lut_adj_197_LC_16_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011101111"
        )
    port map (
            in0 => \N__43600\,
            in1 => \N__47368\,
            in2 => \N__43890\,
            in3 => \N__42887\,
            lcout => n6_adj_819,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \equal_244_i7_2_lut_LC_16_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43240\,
            in2 => \_gnd_net_\,
            in3 => \N__45263\,
            lcout => n7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \equal_241_i9_2_lut_3_lut_4_lut_LC_16_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111011"
        )
    port map (
            in0 => \N__43241\,
            in1 => \N__43398\,
            in2 => \N__45270\,
            in3 => \N__45481\,
            lcout => n9,
            ltout => \n9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_2_lut_adj_193_LC_16_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__38640\,
            in3 => \N__44830\,
            lcout => OPEN,
            ltout => \n8_adj_820_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pin_output_i0_i3_LC_16_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111100100000"
        )
    port map (
            in0 => \N__45899\,
            in1 => \N__46145\,
            in2 => \N__38637\,
            in3 => \N__38707\,
            lcout => pin_out_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46884\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i2_2_lut_adj_180_LC_16_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42494\,
            in2 => \_gnd_net_\,
            in3 => \N__42509\,
            lcout => OPEN,
            ltout => \n6_adj_805_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i3_4_lut_adj_181_LC_16_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011111010"
        )
    port map (
            in0 => \N__42476\,
            in1 => \N__43239\,
            in2 => \N__38634\,
            in3 => \N__45262\,
            lcout => n1788,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pin_output_i0_i4_LC_16_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111100100000"
        )
    port map (
            in0 => \N__45900\,
            in1 => \N__46146\,
            in2 => \N__38730\,
            in3 => \N__42694\,
            lcout => pin_out_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46884\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i5698_2_lut_LC_16_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46322\,
            in2 => \_gnd_net_\,
            in3 => \N__46508\,
            lcout => n9488,
            ltout => \n9488_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \equal_233_i9_2_lut_3_lut_4_lut_LC_16_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111011111"
        )
    port map (
            in0 => \N__45254\,
            in1 => \N__43242\,
            in2 => \N__38736\,
            in3 => \N__45454\,
            lcout => n9_adj_812,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \equal_234_i7_2_lut_LC_16_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011111111"
        )
    port map (
            in0 => \N__43243\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__45253\,
            lcout => n7_adj_811,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_2_lut_3_lut_4_lut_adj_172_LC_16_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000001"
        )
    port map (
            in0 => \N__42583\,
            in1 => \N__44389\,
            in2 => \N__45568\,
            in3 => \N__44873\,
            lcout => OPEN,
            ltout => \n7_adj_818_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pin_output_i0_i2_LC_16_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111100100000"
        )
    port map (
            in0 => \N__45901\,
            in1 => \N__46142\,
            in2 => \N__38733\,
            in3 => \N__38672\,
            lcout => pin_out_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46890\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_2_lut_3_lut_4_lut_adj_166_LC_16_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100010000"
        )
    port map (
            in0 => \N__42582\,
            in1 => \N__44063\,
            in2 => \N__45567\,
            in3 => \N__44872\,
            lcout => n7_adj_821,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_2_lut_3_lut_4_lut_adj_173_LC_16_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000001"
        )
    port map (
            in0 => \N__42603\,
            in1 => \N__44990\,
            in2 => \N__45588\,
            in3 => \N__44874\,
            lcout => n8_adj_817,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i8960_3_lut_LC_16_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__38711\,
            in1 => \N__38671\,
            in2 => \_gnd_net_\,
            in3 => \N__46384\,
            lcout => OPEN,
            ltout => \n13355_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \n13625_bdd_4_lut_LC_16_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101001000100"
        )
    port map (
            in0 => \N__45493\,
            in1 => \N__38652\,
            in2 => \N__38655\,
            in3 => \N__42672\,
            lcout => n13628,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i8959_3_lut_LC_16_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__38977\,
            in1 => \N__39019\,
            in2 => \_gnd_net_\,
            in3 => \N__46383\,
            lcout => n13354,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_2_lut_3_lut_4_lut_adj_174_LC_16_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011110001"
        )
    port map (
            in0 => \N__44091\,
            in1 => \N__45498\,
            in2 => \N__44913\,
            in3 => \N__42604\,
            lcout => OPEN,
            ltout => \n7_adj_840_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pin_output_i0_i0_LC_16_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011101010101010"
        )
    port map (
            in0 => \N__39020\,
            in1 => \N__46143\,
            in2 => \N__39039\,
            in3 => \N__45973\,
            lcout => pin_out_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46898\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pin_output_i0_i1_LC_16_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010111010101010"
        )
    port map (
            in0 => \N__38978\,
            in1 => \N__39003\,
            in2 => \N__46152\,
            in3 => \N__45972\,
            lcout => pin_out_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46898\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i7615_2_lut_3_lut_4_lut_4_lut_LC_16_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011100000"
        )
    port map (
            in0 => \N__45497\,
            in1 => \N__44387\,
            in2 => \N__47599\,
            in3 => \N__45107\,
            lcout => n11952,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pin_output_enable__i8_LC_16_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010110010101010"
        )
    port map (
            in0 => \N__38942\,
            in1 => \N__47502\,
            in2 => \N__42648\,
            in3 => \N__47156\,
            lcout => pin_oe_8,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46898\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1808_2_lut_LC_16_21_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38931\,
            in2 => \_gnd_net_\,
            in3 => \N__38868\,
            lcout => \nx.n2677\,
            ltout => OPEN,
            carryin => \bfn_16_21_0_\,
            carryout => \nx.n10959\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1808_3_lut_LC_16_21_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__38861\,
            in3 => \N__38832\,
            lcout => \nx.n2676\,
            ltout => OPEN,
            carryin => \nx.n10959\,
            carryout => \nx.n10960\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1808_4_lut_LC_16_21_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42123\,
            in2 => \N__38825\,
            in3 => \N__38787\,
            lcout => \nx.n2675\,
            ltout => OPEN,
            carryin => \nx.n10960\,
            carryout => \nx.n10961\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1808_5_lut_LC_16_21_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42126\,
            in2 => \N__38780\,
            in3 => \N__38739\,
            lcout => \nx.n2674\,
            ltout => OPEN,
            carryin => \nx.n10961\,
            carryout => \nx.n10962\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1808_6_lut_LC_16_21_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42124\,
            in2 => \N__39368\,
            in3 => \N__39345\,
            lcout => \nx.n2673\,
            ltout => OPEN,
            carryin => \nx.n10962\,
            carryout => \nx.n10963\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1808_7_lut_LC_16_21_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42127\,
            in2 => \N__39338\,
            in3 => \N__39309\,
            lcout => \nx.n2672\,
            ltout => OPEN,
            carryin => \nx.n10963\,
            carryout => \nx.n10964\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1808_8_lut_LC_16_21_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42125\,
            in2 => \N__39305\,
            in3 => \N__39261\,
            lcout => \nx.n2671\,
            ltout => OPEN,
            carryin => \nx.n10964\,
            carryout => \nx.n10965\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1808_9_lut_LC_16_21_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42128\,
            in2 => \N__39258\,
            in3 => \N__39225\,
            lcout => \nx.n2670\,
            ltout => OPEN,
            carryin => \nx.n10965\,
            carryout => \nx.n10966\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1808_10_lut_LC_16_22_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42138\,
            in2 => \N__39222\,
            in3 => \N__39180\,
            lcout => \nx.n2669\,
            ltout => OPEN,
            carryin => \bfn_16_22_0_\,
            carryout => \nx.n10967\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1808_11_lut_LC_16_22_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42168\,
            in2 => \N__39177\,
            in3 => \N__39141\,
            lcout => \nx.n2668\,
            ltout => OPEN,
            carryin => \nx.n10967\,
            carryout => \nx.n10968\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1808_12_lut_LC_16_22_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42139\,
            in2 => \N__39137\,
            in3 => \N__39090\,
            lcout => \nx.n2667\,
            ltout => OPEN,
            carryin => \nx.n10968\,
            carryout => \nx.n10969\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1808_13_lut_LC_16_22_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42169\,
            in2 => \N__39087\,
            in3 => \N__39042\,
            lcout => \nx.n2666\,
            ltout => OPEN,
            carryin => \nx.n10969\,
            carryout => \nx.n10970\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1808_14_lut_LC_16_22_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42140\,
            in2 => \N__39731\,
            in3 => \N__39690\,
            lcout => \nx.n2665\,
            ltout => OPEN,
            carryin => \nx.n10970\,
            carryout => \nx.n10971\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1808_15_lut_LC_16_22_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42170\,
            in2 => \N__39687\,
            in3 => \N__39651\,
            lcout => \nx.n2664\,
            ltout => OPEN,
            carryin => \nx.n10971\,
            carryout => \nx.n10972\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1808_16_lut_LC_16_22_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42141\,
            in2 => \N__39644\,
            in3 => \N__39603\,
            lcout => \nx.n2663\,
            ltout => OPEN,
            carryin => \nx.n10972\,
            carryout => \nx.n10973\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1808_17_lut_LC_16_22_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42171\,
            in2 => \N__39599\,
            in3 => \N__39552\,
            lcout => \nx.n2662\,
            ltout => OPEN,
            carryin => \nx.n10973\,
            carryout => \nx.n10974\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1808_18_lut_LC_16_23_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42041\,
            in2 => \N__39545\,
            in3 => \N__39504\,
            lcout => \nx.n2661\,
            ltout => OPEN,
            carryin => \bfn_16_23_0_\,
            carryout => \nx.n10975\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1808_19_lut_LC_16_23_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42172\,
            in2 => \N__39494\,
            in3 => \N__39456\,
            lcout => \nx.n2660\,
            ltout => OPEN,
            carryin => \nx.n10975\,
            carryout => \nx.n10976\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1808_20_lut_LC_16_23_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42042\,
            in2 => \N__39452\,
            in3 => \N__39417\,
            lcout => \nx.n2659\,
            ltout => OPEN,
            carryin => \nx.n10976\,
            carryout => \nx.n10977\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1808_21_lut_LC_16_23_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42173\,
            in2 => \N__39414\,
            in3 => \N__39375\,
            lcout => \nx.n2658\,
            ltout => OPEN,
            carryin => \nx.n10977\,
            carryout => \nx.n10978\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1808_22_lut_LC_16_23_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42043\,
            in2 => \N__40164\,
            in3 => \N__40122\,
            lcout => \nx.n2657\,
            ltout => OPEN,
            carryin => \nx.n10978\,
            carryout => \nx.n10979\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1808_23_lut_LC_16_23_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42174\,
            in2 => \N__39949\,
            in3 => \N__40110\,
            lcout => \nx.n2656\,
            ltout => OPEN,
            carryin => \nx.n10979\,
            carryout => \nx.n10980\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1808_24_lut_LC_16_23_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000010001001000"
        )
    port map (
            in0 => \N__42175\,
            in1 => \N__40095\,
            in2 => \N__40803\,
            in3 => \N__39987\,
            lcout => \nx.n2687\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1744_3_lut_LC_16_23_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40899\,
            in2 => \N__42332\,
            in3 => \N__42312\,
            lcout => \nx.n2589\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1741_2_lut_LC_16_24_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39922\,
            in2 => \_gnd_net_\,
            in3 => \N__39852\,
            lcout => \nx.n2577\,
            ltout => OPEN,
            carryin => \bfn_16_24_0_\,
            carryout => \nx.n10938\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1741_3_lut_LC_16_24_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__39849\,
            in3 => \N__39810\,
            lcout => \nx.n2576\,
            ltout => OPEN,
            carryin => \nx.n10938\,
            carryout => \nx.n10939\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1741_4_lut_LC_16_24_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42270\,
            in2 => \N__39807\,
            in3 => \N__39777\,
            lcout => \nx.n2575\,
            ltout => OPEN,
            carryin => \nx.n10939\,
            carryout => \nx.n10940\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1741_5_lut_LC_16_24_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39770\,
            in2 => \N__42297\,
            in3 => \N__39738\,
            lcout => \nx.n2574\,
            ltout => OPEN,
            carryin => \nx.n10940\,
            carryout => \nx.n10941\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1741_6_lut_LC_16_24_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42274\,
            in2 => \N__40482\,
            in3 => \N__40449\,
            lcout => \nx.n2573\,
            ltout => OPEN,
            carryin => \nx.n10941\,
            carryout => \nx.n10942\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1741_7_lut_LC_16_24_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42255\,
            in2 => \N__40445\,
            in3 => \N__40422\,
            lcout => \nx.n2572\,
            ltout => OPEN,
            carryin => \nx.n10942\,
            carryout => \nx.n10943\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1741_8_lut_LC_16_24_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42275\,
            in2 => \N__40419\,
            in3 => \N__40377\,
            lcout => \nx.n2571\,
            ltout => OPEN,
            carryin => \nx.n10943\,
            carryout => \nx.n10944\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1741_9_lut_LC_16_24_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40372\,
            in2 => \N__42298\,
            in3 => \N__40332\,
            lcout => \nx.n2570\,
            ltout => OPEN,
            carryin => \nx.n10944\,
            carryout => \nx.n10945\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1741_10_lut_LC_16_25_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42256\,
            in2 => \N__40329\,
            in3 => \N__40290\,
            lcout => \nx.n2569\,
            ltout => OPEN,
            carryin => \bfn_16_25_0_\,
            carryout => \nx.n10946\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1741_11_lut_LC_16_25_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42262\,
            in2 => \N__40287\,
            in3 => \N__40251\,
            lcout => \nx.n2568\,
            ltout => OPEN,
            carryin => \nx.n10946\,
            carryout => \nx.n10947\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1741_12_lut_LC_16_25_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42257\,
            in2 => \N__40248\,
            in3 => \N__40206\,
            lcout => \nx.n2567\,
            ltout => OPEN,
            carryin => \nx.n10947\,
            carryout => \nx.n10948\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1741_13_lut_LC_16_25_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42263\,
            in2 => \N__40202\,
            in3 => \N__40167\,
            lcout => \nx.n2566\,
            ltout => OPEN,
            carryin => \nx.n10948\,
            carryout => \nx.n10949\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1741_14_lut_LC_16_25_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42258\,
            in2 => \N__40740\,
            in3 => \N__40695\,
            lcout => \nx.n2565\,
            ltout => OPEN,
            carryin => \nx.n10949\,
            carryout => \nx.n10950\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1741_15_lut_LC_16_25_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40691\,
            in2 => \N__42295\,
            in3 => \N__40662\,
            lcout => \nx.n2564\,
            ltout => OPEN,
            carryin => \nx.n10950\,
            carryout => \nx.n10951\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1741_16_lut_LC_16_25_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40659\,
            in2 => \N__42296\,
            in3 => \N__40641\,
            lcout => \nx.n2563\,
            ltout => OPEN,
            carryin => \nx.n10951\,
            carryout => \nx.n10952\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1741_17_lut_LC_16_25_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42267\,
            in2 => \N__40638\,
            in3 => \N__40611\,
            lcout => \nx.n2562\,
            ltout => OPEN,
            carryin => \nx.n10952\,
            carryout => \nx.n10953\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1741_18_lut_LC_16_26_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42251\,
            in2 => \N__40608\,
            in3 => \N__40572\,
            lcout => \nx.n2561\,
            ltout => OPEN,
            carryin => \bfn_16_26_0_\,
            carryout => \nx.n10954\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1741_19_lut_LC_16_26_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42268\,
            in2 => \N__40565\,
            in3 => \N__40530\,
            lcout => \nx.n2560\,
            ltout => OPEN,
            carryin => \nx.n10954\,
            carryout => \nx.n10955\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1741_20_lut_LC_16_26_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42252\,
            in2 => \N__40523\,
            in3 => \N__40485\,
            lcout => \nx.n2559\,
            ltout => OPEN,
            carryin => \nx.n10955\,
            carryout => \nx.n10956\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1741_21_lut_LC_16_26_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42269\,
            in2 => \N__42362\,
            in3 => \N__42339\,
            lcout => \nx.n2558\,
            ltout => OPEN,
            carryin => \nx.n10956\,
            carryout => \nx.n10957\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1741_22_lut_LC_16_26_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42253\,
            in2 => \N__42336\,
            in3 => \N__42303\,
            lcout => \nx.n2557\,
            ltout => OPEN,
            carryin => \nx.n10957\,
            carryout => \nx.n10958\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1741_23_lut_LC_16_26_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001000001100000"
        )
    port map (
            in0 => \N__42254\,
            in1 => \N__40947\,
            in2 => \N__40929\,
            in3 => \N__40806\,
            lcout => \nx.n2588\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i9207_1_lut_2_lut_3_lut_LC_17_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__43818\,
            in1 => \N__47363\,
            in2 => \_gnd_net_\,
            in3 => \N__43592\,
            lcout => n13603,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pin_output_enable__i12_LC_17_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011100010101010"
        )
    port map (
            in0 => \N__40769\,
            in1 => \N__42807\,
            in2 => \N__47488\,
            in3 => \N__47120\,
            lcout => pin_oe_12,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46902\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \counter_633_add_4_2_lut_LC_17_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42785\,
            in2 => \N__43183\,
            in3 => \N__40752\,
            lcout => n45,
            ltout => OPEN,
            carryin => \bfn_17_15_0_\,
            carryout => n10700,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \counter_633__i1_LC_17_15_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100101000111010"
        )
    port map (
            in0 => \N__42878\,
            in1 => \N__42756\,
            in2 => \N__42433\,
            in3 => \N__40749\,
            lcout => counter_1,
            ltout => OPEN,
            carryin => n10700,
            carryout => n10701,
            clk => \N__46899\,
            ce => \N__45981\,
            sr => \_gnd_net_\
        );

    \counter_633__i2_LC_17_15_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1110001000101110"
        )
    port map (
            in0 => \N__42874\,
            in1 => \N__42423\,
            in2 => \N__43092\,
            in3 => \N__40746\,
            lcout => counter_2,
            ltout => OPEN,
            carryin => n10701,
            carryout => n10702,
            clk => \N__46899\,
            ce => \N__45981\,
            sr => \_gnd_net_\
        );

    \counter_633__i3_LC_17_15_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100101000111010"
        )
    port map (
            in0 => \N__42879\,
            in1 => \N__43074\,
            in2 => \N__42434\,
            in3 => \N__40743\,
            lcout => counter_3,
            ltout => OPEN,
            carryin => n10702,
            carryout => n10703,
            clk => \N__46899\,
            ce => \N__45981\,
            sr => \_gnd_net_\
        );

    \counter_633__i4_LC_17_15_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1110001000101110"
        )
    port map (
            in0 => \N__42875\,
            in1 => \N__42427\,
            in2 => \N__43119\,
            in3 => \N__42444\,
            lcout => counter_4,
            ltout => OPEN,
            carryin => n10703,
            carryout => n10704,
            clk => \N__46899\,
            ce => \N__45981\,
            sr => \_gnd_net_\
        );

    \counter_633__i5_LC_17_15_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100101000111010"
        )
    port map (
            in0 => \N__42880\,
            in1 => \N__43104\,
            in2 => \N__42435\,
            in3 => \N__42441\,
            lcout => counter_5,
            ltout => OPEN,
            carryin => n10704,
            carryout => n10705,
            clk => \N__46899\,
            ce => \N__45981\,
            sr => \_gnd_net_\
        );

    \counter_633__i6_LC_17_15_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1110001000101110"
        )
    port map (
            in0 => \N__42876\,
            in1 => \N__42431\,
            in2 => \N__42771\,
            in3 => \N__42438\,
            lcout => counter_6,
            ltout => OPEN,
            carryin => n10705,
            carryout => n10706,
            clk => \N__46899\,
            ce => \N__45981\,
            sr => \_gnd_net_\
        );

    \counter_633__i7_LC_17_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110010001001110"
        )
    port map (
            in0 => \N__42432\,
            in1 => \N__42877\,
            in2 => \N__42801\,
            in3 => \N__42402\,
            lcout => counter_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46899\,
            ce => \N__45981\,
            sr => \_gnd_net_\
        );

    \i9193_4_lut_4_lut_LC_17_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001101110111"
        )
    port map (
            in0 => \N__43128\,
            in1 => \N__43874\,
            in2 => \N__47677\,
            in3 => \N__43641\,
            lcout => n7681,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_2_lut_3_lut_4_lut_4_lut_adj_190_LC_17_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011001000"
        )
    port map (
            in0 => \N__44964\,
            in1 => \N__47646\,
            in2 => \N__45569\,
            in3 => \N__44529\,
            lcout => n11824,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i7627_2_lut_3_lut_4_lut_4_lut_LC_17_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010101000"
        )
    port map (
            in0 => \N__47647\,
            in1 => \N__45106\,
            in2 => \N__44113\,
            in3 => \N__45466\,
            lcout => n11964,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_pin_i0_i0_LC_17_17_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46323\,
            in2 => \_gnd_net_\,
            in3 => \N__42369\,
            lcout => current_pin_0,
            ltout => OPEN,
            carryin => \bfn_17_17_0_\,
            carryout => n10575,
            clk => \N__46887\,
            ce => \N__42456\,
            sr => \N__42465\
        );

    \current_pin_i0_i1_LC_17_17_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46510\,
            in2 => \_gnd_net_\,
            in3 => \N__42366\,
            lcout => current_pin_1,
            ltout => OPEN,
            carryin => n10575,
            carryout => n10576,
            clk => \N__46887\,
            ce => \N__42456\,
            sr => \N__42465\
        );

    \current_pin_i0_i2_LC_17_17_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45560\,
            in2 => \_gnd_net_\,
            in3 => \N__42519\,
            lcout => current_pin_2,
            ltout => OPEN,
            carryin => n10576,
            carryout => n10577,
            clk => \N__46887\,
            ce => \N__42456\,
            sr => \N__42465\
        );

    \current_pin_i0_i3_LC_17_17_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45267\,
            in2 => \_gnd_net_\,
            in3 => \N__42516\,
            lcout => current_pin_3,
            ltout => OPEN,
            carryin => n10577,
            carryout => n10578,
            clk => \N__46887\,
            ce => \N__42456\,
            sr => \N__42465\
        );

    \current_pin_i0_i4_LC_17_17_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43244\,
            in2 => \_gnd_net_\,
            in3 => \N__42513\,
            lcout => current_pin_4,
            ltout => OPEN,
            carryin => n10578,
            carryout => n10579,
            clk => \N__46887\,
            ce => \N__42456\,
            sr => \N__42465\
        );

    \current_pin_i0_i5_LC_17_17_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42510\,
            in2 => \_gnd_net_\,
            in3 => \N__42498\,
            lcout => current_pin_5,
            ltout => OPEN,
            carryin => n10579,
            carryout => n10580,
            clk => \N__46887\,
            ce => \N__42456\,
            sr => \N__42465\
        );

    \current_pin_i0_i6_LC_17_17_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42495\,
            in2 => \_gnd_net_\,
            in3 => \N__42483\,
            lcout => current_pin_6,
            ltout => OPEN,
            carryin => n10580,
            carryout => n10581,
            clk => \N__46887\,
            ce => \N__42456\,
            sr => \N__42465\
        );

    \current_pin_i0_i7_LC_17_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42477\,
            in2 => \_gnd_net_\,
            in3 => \N__42480\,
            lcout => current_pin_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46887\,
            ce => \N__42456\,
            sr => \N__42465\
        );

    \i4198_2_lut_3_lut_4_lut_LC_17_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110100000000"
        )
    port map (
            in0 => \N__43911\,
            in1 => \N__43640\,
            in2 => \N__47658\,
            in3 => \N__42455\,
            lcout => n7985,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i9181_2_lut_4_lut_LC_17_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001000000011"
        )
    port map (
            in0 => \N__43174\,
            in1 => \N__47586\,
            in2 => \N__43668\,
            in3 => \N__43910\,
            lcout => n7635,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_3_lut_4_lut_LC_17_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011101100"
        )
    port map (
            in0 => \N__43414\,
            in1 => \N__44891\,
            in2 => \N__45597\,
            in3 => \N__42588\,
            lcout => OPEN,
            ltout => \n9_adj_824_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pin_output_i0_i7_LC_17_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111100100000"
        )
    port map (
            in0 => \N__45971\,
            in1 => \N__46098\,
            in2 => \N__42741\,
            in3 => \N__42946\,
            lcout => pin_out_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46895\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_2_lut_3_lut_4_lut_adj_167_LC_17_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011011100"
        )
    port map (
            in0 => \N__44995\,
            in1 => \N__44890\,
            in2 => \N__45596\,
            in3 => \N__42587\,
            lcout => OPEN,
            ltout => \n8_adj_822_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pin_output_i0_i5_LC_17_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111100100000"
        )
    port map (
            in0 => \N__45970\,
            in1 => \N__46097\,
            in2 => \N__42738\,
            in3 => \N__42724\,
            lcout => pin_out_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46895\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i8962_3_lut_LC_17_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__46344\,
            in1 => \N__42728\,
            in2 => \_gnd_net_\,
            in3 => \N__42698\,
            lcout => OPEN,
            ltout => \n13357_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_pin_1__bdd_4_lut_9236_LC_17_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110110001100100"
        )
    port map (
            in0 => \N__45487\,
            in1 => \N__46511\,
            in2 => \N__42675\,
            in3 => \N__42894\,
            lcout => n13625,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \equal_234_i6_2_lut_LC_17_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46512\,
            in2 => \_gnd_net_\,
            in3 => \N__46345\,
            lcout => n6_adj_810,
            ltout => \n6_adj_810_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i7543_2_lut_3_lut_4_lut_LC_17_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110111111111"
        )
    port map (
            in0 => \N__43248\,
            in1 => \N__45268\,
            in2 => \N__42666\,
            in3 => \N__45488\,
            lcout => n11874,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_2_lut_3_lut_4_lut_4_lut_adj_188_LC_17_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011001000"
        )
    port map (
            in0 => \N__44530\,
            in1 => \N__47636\,
            in2 => \N__44114\,
            in3 => \N__45507\,
            lcout => n11823,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_2_lut_3_lut_4_lut_adj_168_LC_17_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011110100"
        )
    port map (
            in0 => \N__44388\,
            in1 => \N__45508\,
            in2 => \N__44909\,
            in3 => \N__42615\,
            lcout => OPEN,
            ltout => \n7_adj_823_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pin_output_i0_i6_LC_17_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010101011101010"
        )
    port map (
            in0 => \N__42908\,
            in1 => \N__45974\,
            in2 => \N__42993\,
            in3 => \N__46144\,
            lcout => pin_out_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46903\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pin_output_enable__i19_LC_17_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110010001100"
        )
    port map (
            in0 => \N__43365\,
            in1 => \N__42977\,
            in2 => \N__47149\,
            in3 => \N__47637\,
            lcout => pin_oe_19,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46903\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i8963_3_lut_LC_17_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__46343\,
            in1 => \N__42950\,
            in2 => \_gnd_net_\,
            in3 => \N__42907\,
            lcout => n13358,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_2_lut_3_lut_4_lut_adj_165_LC_17_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011001101"
        )
    port map (
            in0 => \N__44107\,
            in1 => \N__44907\,
            in2 => \N__45587\,
            in3 => \N__44531\,
            lcout => n8_adj_826,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i2_3_lut_LC_18_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__43824\,
            in1 => \N__47329\,
            in2 => \_gnd_net_\,
            in3 => \N__43588\,
            lcout => n3762,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pin_output_enable__i16_LC_18_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011100010101010"
        )
    port map (
            in0 => \N__42818\,
            in1 => \N__42843\,
            in2 => \N__47460\,
            in3 => \N__47122\,
            lcout => pin_oe_16,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46908\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_2_lut_3_lut_4_lut_4_lut_adj_202_LC_18_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010001010"
        )
    port map (
            in0 => \N__47479\,
            in1 => \N__44112\,
            in2 => \N__45642\,
            in3 => \N__44537\,
            lcout => n11820,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i2_2_lut_LC_18_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42797\,
            in2 => \_gnd_net_\,
            in3 => \N__42786\,
            lcout => OPEN,
            ltout => \n10_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i9165_4_lut_LC_18_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__42767\,
            in1 => \N__42755\,
            in2 => \N__42744\,
            in3 => \N__43062\,
            lcout => \state_7_N_167_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i6_4_lut_adj_179_LC_18_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__43115\,
            in1 => \N__43103\,
            in2 => \N__43091\,
            in3 => \N__43073\,
            lcout => n14,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i8975_3_lut_LC_18_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__43042\,
            in1 => \N__43009\,
            in2 => \_gnd_net_\,
            in3 => \N__46320\,
            lcout => n13370,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pin_output_i0_i11_LC_18_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101110011001100"
        )
    port map (
            in0 => \N__46094\,
            in1 => \N__43043\,
            in2 => \N__44199\,
            in3 => \N__45994\,
            lcout => pin_out_11,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46900\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_2_lut_3_lut_4_lut_adj_163_LC_18_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010101011"
        )
    port map (
            in0 => \N__44854\,
            in1 => \N__44426\,
            in2 => \N__45643\,
            in3 => \N__44534\,
            lcout => OPEN,
            ltout => \n7_adj_827_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pin_output_i0_i10_LC_18_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111100100000"
        )
    port map (
            in0 => \N__45993\,
            in1 => \N__46095\,
            in2 => \N__43029\,
            in3 => \N__43010\,
            lcout => pin_out_10,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46900\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_2_lut_3_lut_4_lut_adj_160_LC_18_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010101110"
        )
    port map (
            in0 => \N__44853\,
            in1 => \N__45461\,
            in2 => \N__44996\,
            in3 => \N__44533\,
            lcout => n7_adj_830,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_2_lut_3_lut_4_lut_adj_161_LC_18_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011001110"
        )
    port map (
            in0 => \N__45556\,
            in1 => \N__44878\,
            in2 => \N__44111\,
            in3 => \N__44535\,
            lcout => n8_adj_829,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i5882_2_lut_3_lut_4_lut_LC_18_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111011"
        )
    port map (
            in0 => \N__47478\,
            in1 => \N__43891\,
            in2 => \N__43651\,
            in3 => \N__43302\,
            lcout => n9675,
            ltout => \n9675_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pin_output_i0_i15_LC_18_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111100001000"
        )
    port map (
            in0 => \N__45979\,
            in1 => \N__43308\,
            in2 => \N__42996\,
            in3 => \N__45787\,
            lcout => pin_out_15,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46892\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_2_lut_3_lut_4_lut_adj_162_LC_18_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011101100"
        )
    port map (
            in0 => \N__43431\,
            in1 => \N__44879\,
            in2 => \N__45634\,
            in3 => \N__44536\,
            lcout => n8_adj_832,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_2_lut_3_lut_4_lut_4_lut_LC_18_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011100000"
        )
    port map (
            in0 => \N__45462\,
            in1 => \N__44991\,
            in2 => \N__47600\,
            in3 => \N__45062\,
            lcout => n11822,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i9145_4_lut_LC_18_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000010111000"
        )
    port map (
            in0 => \N__44676\,
            in1 => \N__43236\,
            in2 => \N__43257\,
            in3 => \N__45251\,
            lcout => \pin_out_22__N_216\,
            ltout => \pin_out_22__N_216_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i9155_4_lut_LC_18_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010110101111000"
        )
    port map (
            in0 => \N__43237\,
            in1 => \N__45201\,
            in2 => \N__43296\,
            in3 => \N__44124\,
            lcout => n13551,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \n13637_bdd_4_lut_LC_18_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001010000"
        )
    port map (
            in0 => \N__45452\,
            in1 => \N__43293\,
            in2 => \N__43284\,
            in3 => \N__46206\,
            lcout => OPEN,
            ltout => \n13640_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i9144_3_lut_LC_18_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__45250\,
            in1 => \_gnd_net_\,
            in2 => \N__43272\,
            in3 => \N__43269\,
            lcout => n13540,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \equal_224_i7_2_lut_LC_18_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43238\,
            in2 => \_gnd_net_\,
            in3 => \N__45252\,
            lcout => n7_adj_797,
            ltout => \n7_adj_797_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_2_lut_4_lut_adj_199_LC_18_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010101110"
        )
    port map (
            in0 => \N__44886\,
            in1 => \N__43424\,
            in2 => \N__43200\,
            in3 => \N__45453\,
            lcout => n8_adj_836,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i41_4_lut_LC_18_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000110101011"
        )
    port map (
            in0 => \N__47583\,
            in1 => \N__43197\,
            in2 => \N__43185\,
            in3 => \N__43976\,
            lcout => n26,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_2_lut_3_lut_4_lut_4_lut_adj_189_LC_18_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100010011001100"
        )
    port map (
            in0 => \N__43430\,
            in1 => \N__47584\,
            in2 => \N__44544\,
            in3 => \N__45574\,
            lcout => OPEN,
            ltout => \n11825_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pin_output_enable__i15_LC_18_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100101011001100"
        )
    port map (
            in0 => \N__47585\,
            in1 => \N__43988\,
            in2 => \N__44007\,
            in3 => \N__47123\,
            lcout => pin_oe_15,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46904\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i4262_2_lut_3_lut_4_lut_LC_18_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__43977\,
            in1 => \N__47582\,
            in2 => \N__43912\,
            in3 => \N__43625\,
            lcout => n8025,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i7617_2_lut_3_lut_4_lut_4_lut_LC_18_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111100000000"
        )
    port map (
            in0 => \N__44105\,
            in1 => \N__45101\,
            in2 => \N__45641\,
            in3 => \N__47641\,
            lcout => OPEN,
            ltout => \n11954_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pin_output_enable__i20_LC_18_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010110010101010"
        )
    port map (
            in0 => \N__43442\,
            in1 => \N__47642\,
            in2 => \N__43458\,
            in3 => \N__47130\,
            lcout => pin_oe_20,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46909\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_2_lut_4_lut_4_lut_LC_18_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011010000"
        )
    port map (
            in0 => \N__43428\,
            in1 => \N__45570\,
            in2 => \N__47676\,
            in3 => \N__45091\,
            lcout => n11821,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_2_lut_3_lut_4_lut_adj_177_LC_18_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110111001100"
        )
    port map (
            in0 => \N__45100\,
            in1 => \N__44908\,
            in2 => \N__44115\,
            in3 => \N__45668\,
            lcout => n7_adj_837,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pin_output_i0_i8_LC_18_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111001011110000"
        )
    port map (
            in0 => \N__43359\,
            in1 => \N__46141\,
            in2 => \N__43336\,
            in3 => \N__45980\,
            lcout => pin_out_8,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46919\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i7625_2_lut_3_lut_4_lut_4_lut_LC_19_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010001100"
        )
    port map (
            in0 => \N__44431\,
            in1 => \N__47481\,
            in2 => \N__45669\,
            in3 => \N__44539\,
            lcout => OPEN,
            ltout => \n11962_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pin_output_enable__i14_LC_19_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100101011001100"
        )
    port map (
            in0 => \N__47482\,
            in1 => \N__44231\,
            in2 => \N__44250\,
            in3 => \N__47119\,
            lcout => pin_oe_14,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46910\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_2_lut_adj_198_LC_19_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44220\,
            in2 => \_gnd_net_\,
            in3 => \N__44871\,
            lcout => n8_adj_828,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i7621_2_lut_3_lut_4_lut_4_lut_LC_19_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010001100"
        )
    port map (
            in0 => \N__44981\,
            in1 => \N__47483\,
            in2 => \N__45670\,
            in3 => \N__45105\,
            lcout => OPEN,
            ltout => \n11958_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pin_output_enable__i21_LC_19_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100101011001100"
        )
    port map (
            in0 => \N__47484\,
            in1 => \N__44168\,
            in2 => \N__44190\,
            in3 => \N__47124\,
            lcout => pin_oe_21,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46905\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i9140_3_lut_LC_19_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__45534\,
            in1 => \N__45117\,
            in2 => \_gnd_net_\,
            in3 => \N__44157\,
            lcout => OPEN,
            ltout => \n13536_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i9146_3_lut_LC_19_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45261\,
            in2 => \N__44139\,
            in3 => \N__44136\,
            lcout => n13542,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_2_lut_3_lut_4_lut_LC_19_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100010000"
        )
    port map (
            in0 => \N__44538\,
            in1 => \N__44422\,
            in2 => \N__45615\,
            in3 => \N__44902\,
            lcout => OPEN,
            ltout => \n7_adj_831_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pin_output_i0_i14_LC_19_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111100100000"
        )
    port map (
            in0 => \N__45995\,
            in1 => \N__46137\,
            in2 => \N__44118\,
            in3 => \N__45752\,
            lcout => pin_out_14,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46896\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_2_lut_3_lut_4_lut_adj_201_LC_19_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011110001"
        )
    port map (
            in0 => \N__45090\,
            in1 => \N__44095\,
            in2 => \N__44912\,
            in3 => \N__45538\,
            lcout => OPEN,
            ltout => \n7_adj_833_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pin_output_i0_i16_LC_19_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111101000000"
        )
    port map (
            in0 => \N__46136\,
            in1 => \N__45996\,
            in2 => \N__44553\,
            in3 => \N__44698\,
            lcout => pin_out_16,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46896\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pin_output_i0_i19_LC_19_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111001011110000"
        )
    port map (
            in0 => \N__44550\,
            in1 => \N__46096\,
            in2 => \N__44278\,
            in3 => \N__45959\,
            lcout => pin_out_19,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46906\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i7619_2_lut_3_lut_4_lut_4_lut_LC_19_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111100000000"
        )
    port map (
            in0 => \N__44540\,
            in1 => \N__45010\,
            in2 => \N__45652\,
            in3 => \N__47480\,
            lcout => n11956,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_2_lut_3_lut_4_lut_adj_178_LC_19_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010101011"
        )
    port map (
            in0 => \N__44903\,
            in1 => \N__44405\,
            in2 => \N__45654\,
            in3 => \N__45089\,
            lcout => OPEN,
            ltout => \n7_adj_835_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pin_output_i0_i18_LC_19_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011101010101010"
        )
    port map (
            in0 => \N__44309\,
            in1 => \N__46110\,
            in2 => \N__44442\,
            in3 => \N__45960\,
            lcout => pin_out_18,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46911\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_2_lut_4_lut_LC_19_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000111110000"
        )
    port map (
            in0 => \N__44421\,
            in1 => \N__45099\,
            in2 => \N__44910\,
            in3 => \N__45611\,
            lcout => OPEN,
            ltout => \n7_adj_839_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pin_output_i0_i22_LC_19_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111100100000"
        )
    port map (
            in0 => \N__45956\,
            in1 => \N__46111\,
            in2 => \N__44328\,
            in3 => \N__44581\,
            lcout => pin_out_22,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46914\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_pin_0__bdd_4_lut_9241_LC_19_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001110001000"
        )
    port map (
            in0 => \N__44308\,
            in1 => \N__46559\,
            in2 => \N__44282\,
            in3 => \N__46392\,
            lcout => n13631,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_2_lut_3_lut_4_lut_adj_176_LC_19_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100010000"
        )
    port map (
            in0 => \N__45098\,
            in1 => \N__45006\,
            in2 => \N__45653\,
            in3 => \N__44892\,
            lcout => n7_adj_838,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_2_lut_3_lut_4_lut_adj_200_LC_19_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000001"
        )
    port map (
            in0 => \N__45108\,
            in1 => \N__45019\,
            in2 => \N__45650\,
            in3 => \N__44911\,
            lcout => OPEN,
            ltout => \n8_adj_834_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pin_output_i0_i17_LC_19_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100110011101100"
        )
    port map (
            in0 => \N__45957\,
            in1 => \N__44738\,
            in2 => \N__44754\,
            in3 => \N__46139\,
            lcout => pin_out_17,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46920\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \n13631_bdd_4_lut_LC_19_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010111000"
        )
    port map (
            in0 => \N__44737\,
            in1 => \N__44724\,
            in2 => \N__44708\,
            in3 => \N__46563\,
            lcout => OPEN,
            ltout => \n13634_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i8994_3_lut_LC_19_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45598\,
            in2 => \N__44679\,
            in3 => \N__44559\,
            lcout => n13389,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pin_output_i0_i21_LC_19_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111010011110000"
        )
    port map (
            in0 => \N__46138\,
            in1 => \N__44667\,
            in2 => \N__44642\,
            in3 => \N__45958\,
            lcout => pin_out_21,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46920\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pin_output_i0_i20_LC_19_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111000011111000"
        )
    port map (
            in0 => \N__45952\,
            in1 => \N__44661\,
            in2 => \N__44615\,
            in3 => \N__46140\,
            lcout => pin_out_20,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46922\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_pin_4__I_0_i19_3_lut_LC_19_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__44635\,
            in1 => \N__44608\,
            in2 => \_gnd_net_\,
            in3 => \N__46408\,
            lcout => OPEN,
            ltout => \n19_adj_790_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i8993_4_lut_LC_19_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010011110000"
        )
    port map (
            in0 => \N__46409\,
            in1 => \N__44585\,
            in2 => \N__44562\,
            in3 => \N__46571\,
            lcout => n13388,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i8980_3_lut_LC_20_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__45811\,
            in1 => \N__46165\,
            in2 => \_gnd_net_\,
            in3 => \N__46336\,
            lcout => OPEN,
            ltout => \n13375_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_pin_1__bdd_4_lut_LC_20_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110110001100100"
        )
    port map (
            in0 => \N__45492\,
            in1 => \N__46513\,
            in2 => \N__46209\,
            in3 => \N__45735\,
            lcout => n13637,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pin_output_i0_i12_LC_20_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100111011001100"
        )
    port map (
            in0 => \N__46194\,
            in1 => \N__46166\,
            in2 => \N__46151\,
            in3 => \N__45978\,
            lcout => pin_out_12,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46901\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pin_output_i0_i13_LC_20_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111101000000"
        )
    port map (
            in0 => \N__46132\,
            in1 => \N__46008\,
            in2 => \N__45992\,
            in3 => \N__45812\,
            lcout => pin_out_13,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46901\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i8981_3_lut_LC_20_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__45788\,
            in1 => \N__45751\,
            in2 => \_gnd_net_\,
            in3 => \N__46335\,
            lcout => n13376,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pin_output_enable__i13_LC_20_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101100011001100"
        )
    port map (
            in0 => \N__45729\,
            in1 => \N__45707\,
            in2 => \N__47659\,
            in3 => \N__47147\,
            lcout => pin_oe_13,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46912\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i9075_4_lut_LC_20_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010101100"
        )
    port map (
            in0 => \N__46656\,
            in1 => \N__46605\,
            in2 => \N__45651\,
            in3 => \N__45269\,
            lcout => n13465,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_pin_0__bdd_4_lut_9246_LC_21_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011100011001100"
        )
    port map (
            in0 => \N__45189\,
            in1 => \N__46337\,
            in2 => \N__45174\,
            in3 => \N__46522\,
            lcout => OPEN,
            ltout => \n13643_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \n13643_bdd_4_lut_LC_21_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010111100000"
        )
    port map (
            in0 => \N__46523\,
            in1 => \N__45150\,
            in2 => \N__45138\,
            in3 => \N__45135\,
            lcout => n13646,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pin_output_enable__i17_LC_21_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101100011001100"
        )
    port map (
            in0 => \N__47706\,
            in1 => \N__46934\,
            in2 => \N__47663\,
            in3 => \N__47148\,
            lcout => pin_oe_17,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46907\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i8957_4_lut_LC_23_32_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010111000100010"
        )
    port map (
            in0 => \N__46215\,
            in1 => \N__46572\,
            in2 => \N__46419\,
            in3 => \N__46662\,
            lcout => n13352,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \n13607_bdd_4_lut_LC_24_27_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010111000"
        )
    port map (
            in0 => \N__46644\,
            in1 => \N__46428\,
            in2 => \N__46632\,
            in3 => \N__46555\,
            lcout => n13610,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_pin_0__bdd_4_lut_9231_LC_24_32_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101100010101010"
        )
    port map (
            in0 => \N__46411\,
            in1 => \N__46593\,
            in2 => \N__46587\,
            in3 => \N__46567\,
            lcout => n13607,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Mux_82_i19_3_lut_LC_24_32_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__46412\,
            in1 => \N__46233\,
            in2 => \_gnd_net_\,
            in3 => \N__46227\,
            lcout => n19_adj_789,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );
end \INTERFACE\;
