// Verilog netlist produced by program LSE :  version Diamond Version 0.0.0
// Netlist written on Fri Jan 31 00:25:13 2020
//
// Verilog Description of module TinyFPGA_B
//

module TinyFPGA_B (CLK, LED, USBPU, ENCODER0_A, ENCODER0_B, ENCODER1_A, 
            ENCODER1_B, HALL1, HALL2, HALL3, FAULT_N, NEOPXL, DE, 
            TX, RX, CS_CLK, CS, CS_MISO, SCL, SDA, INLC, INHC, 
            INLB, INHB, INLA, INHA) /* synthesis syn_module_defined=1 */ ;   // verilog/TinyFPGA_B.v(2[8:18])
    input CLK;   // verilog/TinyFPGA_B.v(3[9:12])
    output LED;   // verilog/TinyFPGA_B.v(4[10:13])
    output USBPU;   // verilog/TinyFPGA_B.v(5[10:15])
    input ENCODER0_A;   // verilog/TinyFPGA_B.v(6[9:19])
    input ENCODER0_B;   // verilog/TinyFPGA_B.v(7[9:19])
    input ENCODER1_A;   // verilog/TinyFPGA_B.v(8[9:19])
    input ENCODER1_B;   // verilog/TinyFPGA_B.v(9[9:19])
    input HALL1 /* synthesis black_box_pad_pin=1 */ ;   // verilog/TinyFPGA_B.v(10[9:14])
    input HALL2 /* synthesis black_box_pad_pin=1 */ ;   // verilog/TinyFPGA_B.v(11[9:14])
    input HALL3 /* synthesis black_box_pad_pin=1 */ ;   // verilog/TinyFPGA_B.v(12[9:14])
    input FAULT_N;   // verilog/TinyFPGA_B.v(13[9:16])
    output NEOPXL;   // verilog/TinyFPGA_B.v(14[10:16])
    output DE;   // verilog/TinyFPGA_B.v(15[10:12])
    output TX /* synthesis black_box_pad_pin=1 */ ;   // verilog/TinyFPGA_B.v(16[10:12])
    input RX;   // verilog/TinyFPGA_B.v(17[9:11])
    output CS_CLK;   // verilog/TinyFPGA_B.v(18[10:16])
    output CS;   // verilog/TinyFPGA_B.v(19[10:12])
    input CS_MISO;   // verilog/TinyFPGA_B.v(20[9:16])
    inout SCL /* synthesis black_box_pad_pin=1 */ ;   // verilog/TinyFPGA_B.v(21[9:12])
    inout SDA /* synthesis black_box_pad_pin=1 */ ;   // verilog/TinyFPGA_B.v(22[9:12])
    output INLC;   // verilog/TinyFPGA_B.v(23[10:14])
    output INHC;   // verilog/TinyFPGA_B.v(24[10:14])
    output INLB;   // verilog/TinyFPGA_B.v(25[10:14])
    output INHB;   // verilog/TinyFPGA_B.v(26[10:14])
    output INLA;   // verilog/TinyFPGA_B.v(27[10:14])
    output INHA;   // verilog/TinyFPGA_B.v(28[10:14])
    
    wire CLK_c /* synthesis SET_AS_NETWORK=CLK_c, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(3[9:12])
    wire clk32MHz /* synthesis SET_AS_NETWORK=clk32MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(33[6:14])
    
    wire GND_net, VCC_net, LED_c, ENCODER0_A_c_1, ENCODER0_B_c_0, 
        ENCODER1_A_c_1, ENCODER1_B_c_0, NEOPXL_c, DE_c, RX_c, INHC_c, 
        INLB_c, INHB_c, INLA_c, INHA_c;
    wire [7:0]ID;   // verilog/TinyFPGA_B.v(39[11:13])
    wire [23:0]neopxl_color;   // verilog/TinyFPGA_B.v(41[13:25])
    
    wire hall1, hall2, hall3;
    wire [22:0]pwm_setpoint;   // verilog/TinyFPGA_B.v(87[13:25])
    wire [23:0]duty;   // verilog/TinyFPGA_B.v(88[21:25])
    
    wire tx_o, tx_enable;
    wire [23:0]encoder0_position;   // verilog/TinyFPGA_B.v(122[22:39])
    wire [23:0]encoder0_position_scaled;   // verilog/TinyFPGA_B.v(123[21:45])
    wire [23:0]encoder1_position;   // verilog/TinyFPGA_B.v(124[22:39])
    wire [23:0]displacement;   // verilog/TinyFPGA_B.v(125[21:33])
    wire [23:0]setpoint;   // verilog/TinyFPGA_B.v(126[22:30])
    
    wire n33471;
    wire [23:0]Kp;   // verilog/TinyFPGA_B.v(127[22:24])
    
    wire n28352, n32323;
    wire [23:0]Ki;   // verilog/TinyFPGA_B.v(128[22:24])
    
    wire n28351, n28164, n28163;
    wire [7:0]control_mode;   // verilog/TinyFPGA_B.v(130[14:26])
    wire [23:0]PWMLimit;   // verilog/TinyFPGA_B.v(131[22:30])
    wire [23:0]IntegralLimit;   // verilog/TinyFPGA_B.v(132[22:35])
    
    wire n28162;
    wire [23:0]motor_state;   // verilog/TinyFPGA_B.v(162[22:33])
    
    wire n28350, n28349;
    wire [7:0]data;   // verilog/TinyFPGA_B.v(206[14:18])
    
    wire data_ready, sda_out, n17360, sda_enable, scl, scl_enable;
    wire [31:0]delay_counter;   // verilog/TinyFPGA_B.v(230[11:24])
    
    wire read;
    wire [2:0]\ID_READOUT_FSM.state ;   // verilog/TinyFPGA_B.v(238[15:20])
    wire [22:0]pwm_setpoint_22__N_11;
    
    wire RX_N_10;
    wire [31:0]timer;   // verilog/neopixel.v(9[12:17])
    wire [31:0]motor_state_23__N_82;
    wire [25:0]encoder0_position_scaled_23__N_34;
    wire [23:0]displacement_23__N_58;
    
    wire n573, n574, n575, n576, n577, n578, n579, n580, n581, 
        n582, n583, n584, n585, n586, n587, n588, n589, n590, 
        n591, n592, n593, n594, n595, n596, n597, n598, n599, 
        n600, n601, n602, n603, n604, read_N_295, n691, n6028, 
        n7, n425;
    wire [3:0]state;   // verilog/neopixel.v(16[20:25])
    
    wire start, \neo_pixel_transmitter.done ;
    wire [31:0]\neo_pixel_transmitter.t0 ;   // verilog/neopixel.v(28[14:16])
    
    wire n28161, n32009, n24759;
    wire [3:0]state_3__N_402;
    
    wire n4, n2970, n28348, n28347, n28160, n28346, n10, n28345, 
        n28344, n28343, n28342, n28159, n6, n17513, n28158, n28341, 
        n36960, n33535, n36943;
    wire [31:0]pwm_counter;   // verilog/pwm.v(11[9:20])
    
    wire n28340, n28157, n28339, n3, n4_adj_4884, n5, n6_adj_4885, 
        n7_adj_4886, n8, n9, n10_adj_4887, n11, n12, n13, n14, 
        n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, 
        n25, n28338, rx_data_ready;
    wire [7:0]rx_data;   // verilog/coms.v(91[13:20])
    wire [7:0]\data_in[3] ;   // verilog/coms.v(95[12:19])
    wire [7:0]\data_in[2] ;   // verilog/coms.v(95[12:19])
    wire [7:0]\data_in[1] ;   // verilog/coms.v(95[12:19])
    wire [7:0]\data_in[0] ;   // verilog/coms.v(95[12:19])
    
    wire n28156, n10524, n28337, n33425;
    wire [7:0]\data_in_frame[21] ;   // verilog/coms.v(96[12:25])
    wire [7:0]\data_in_frame[13] ;   // verilog/coms.v(96[12:25])
    wire [7:0]\data_in_frame[12] ;   // verilog/coms.v(96[12:25])
    wire [7:0]\data_in_frame[11] ;   // verilog/coms.v(96[12:25])
    wire [7:0]\data_in_frame[10] ;   // verilog/coms.v(96[12:25])
    wire [7:0]\data_in_frame[9] ;   // verilog/coms.v(96[12:25])
    wire [7:0]\data_in_frame[8] ;   // verilog/coms.v(96[12:25])
    wire [7:0]\data_in_frame[6] ;   // verilog/coms.v(96[12:25])
    wire [7:0]\data_in_frame[5] ;   // verilog/coms.v(96[12:25])
    wire [7:0]\data_in_frame[4] ;   // verilog/coms.v(96[12:25])
    wire [7:0]\data_in_frame[3] ;   // verilog/coms.v(96[12:25])
    wire [7:0]\data_in_frame[2] ;   // verilog/coms.v(96[12:25])
    wire [7:0]\data_in_frame[1] ;   // verilog/coms.v(96[12:25])
    wire [7:0]\data_out_frame[25] ;   // verilog/coms.v(97[12:26])
    wire [7:0]\data_out_frame[24] ;   // verilog/coms.v(97[12:26])
    wire [7:0]\data_out_frame[23] ;   // verilog/coms.v(97[12:26])
    wire [7:0]\data_out_frame[20] ;   // verilog/coms.v(97[12:26])
    wire [7:0]\data_out_frame[19] ;   // verilog/coms.v(97[12:26])
    wire [7:0]\data_out_frame[18] ;   // verilog/coms.v(97[12:26])
    wire [7:0]\data_out_frame[17] ;   // verilog/coms.v(97[12:26])
    wire [7:0]\data_out_frame[16] ;   // verilog/coms.v(97[12:26])
    wire [7:0]\data_out_frame[15] ;   // verilog/coms.v(97[12:26])
    wire [7:0]\data_out_frame[14] ;   // verilog/coms.v(97[12:26])
    wire [7:0]\data_out_frame[13] ;   // verilog/coms.v(97[12:26])
    wire [7:0]\data_out_frame[12] ;   // verilog/coms.v(97[12:26])
    wire [7:0]\data_out_frame[11] ;   // verilog/coms.v(97[12:26])
    wire [7:0]\data_out_frame[10] ;   // verilog/coms.v(97[12:26])
    wire [7:0]\data_out_frame[9] ;   // verilog/coms.v(97[12:26])
    wire [7:0]\data_out_frame[8] ;   // verilog/coms.v(97[12:26])
    wire [7:0]\data_out_frame[7] ;   // verilog/coms.v(97[12:26])
    wire [7:0]\data_out_frame[6] ;   // verilog/coms.v(97[12:26])
    wire [7:0]\data_out_frame[5] ;   // verilog/coms.v(97[12:26])
    wire [7:0]\data_out_frame[4] ;   // verilog/coms.v(97[12:26])
    
    wire n28155, tx_active;
    wire [31:0]\FRAME_MATCHER.state ;   // verilog/coms.v(112[11:16])
    
    wire n28336, n33401, n33399, n33397, n123, n4_adj_4888, n7_adj_4889, 
        n28154, n24721, n24_adj_4890, n10417, n24717, n21_adj_4891, 
        n20_adj_4892, n17_adj_4893, n25_adj_4894, n17_adj_4895, n31783, 
        n771, n28335, n28334, n28333, n28153, n28152, n34265, 
        n27756, n28332, n28331, n28330, n27755, n28329, n28151, 
        n28150, n28328, n24685, n28327, n24683, n28149, n28148, 
        n24833, n28326, n28325, n28147, n28324, n24747, n27754, 
        n24673, n28146, n28323, n27753, n28322, n28321, n24829, 
        n23879, n27752, n24707, n28145, n23736, n28320, n28319, 
        n28318, n28144, n28143, n28317, n28142, n28316, n28003, 
        n28315, n28141, n28314, n28313, n28140, n28139, n28138, 
        n28312, n28137, n28002, n28001, n28136, n28311, n28000, 
        n28310, n28309, n27751, n28135, n28308, n28307, n28134, 
        n28133, n27999, n27740, n28306, n28305, n28304, n28303, 
        n27847, n27739, n28302, n28301, n27846, n28132, n28131, 
        n28300, n27845, n28299, n28298, n28130, n28129, n28128, 
        n28297, n28127, n28126, n28125, n28124, n28123, n28122, 
        n28121, n27844, n28120, n28296, n28295, n28119, n27843, 
        n28294, n28293, n27842, n28118, n28292, n28291, n27841, 
        n27738, n28117, n28290, n28116, n28115, n28289, n28288, 
        n28287, n14_adj_4896, n28286, n27840, n28114, n28113, n28285, 
        n28284, n27750, n28283, n28282, n28281, n28280, n28279, 
        n28278, n28277, n28276, n31453, n28275, n28274, n27839, 
        n28273, n28272, n28271, n28270, n28269, n28268, n27838, 
        n28267, n27837, n28266, n27836, n28265, n27749, n28264, 
        n28263, n28262, n28261, n28260, n27835, n28259, n28258, 
        n28257, n24577, n28256, n28255, n5_adj_4897, n28254, n28096, 
        n37323, n28253, n28095, n3303;
    wire [31:0]\FRAME_MATCHER.state_31__N_2662 ;
    
    wire n28252, n28251, n28094, n28250, n28249, n28248, n28093, 
        n28247, n28246, n28245, n28092, n28091, n28090, n28244, 
        n28089, n28243, n28088, n28087, n28086, n28085, n28242, 
        n28084, n27834, n28241, n28240, n28239, n28238, n28237, 
        n28083, n28082, n28236, n28081, n27833, n4452, n28235, 
        n28234, n28233, n27832, n28080, n28079, n27831, n6_adj_4898, 
        n33923, n28078, n28077, n28076, n28232, n28231, n27830, 
        n28230, n27829, n28229, n28228, n28075, n28227, n28226, 
        n27828, n20830, n27748, n24244, n28225, n28074, n39, n17552, 
        n30, n29, n28, n27, n18_adj_4899, n8_adj_4900, n12_adj_4901, 
        n1247, n28224, n35293, n34503, n35117, n24835, n24729, 
        n34039, n19600, n19599, n19598, n19597, n19596, n19595, 
        n19594, n19593, n19592, n19588, n27747, n28223, n25_adj_4902, 
        n24_adj_4903, n23_adj_4904, n22_adj_4905, n21_adj_4906, n20_adj_4907, 
        n19_adj_4908, n18_adj_4909, n17_adj_4910, n16_adj_4911, n15_adj_4912, 
        n14_adj_4913, n13_adj_4914, n12_adj_4915, n19584, n19583, 
        n19582, n19581, n19580, n19579, n19578, n19577, n19576, 
        n19575, n19574, n19573, n19572, n19571, n19570, n19569, 
        n19568, n19567, n19566, n19565, n19564, n19563, n19562, 
        n19561, n19560, n19559, n19558, n19557, n19556, n19555, 
        n19554, n19553, n19552, n19551, n19550, n19549, n19548, 
        n19547, n19546, n19545, n19544, n19543, n19542, n19541, 
        n19540, n11_adj_4916, n10_adj_4917, n9_adj_4918, n8_adj_4919, 
        n7_adj_4920, n6_adj_4921, n5_adj_4922, n4_adj_4923, n3_adj_4924, 
        n2, n19539, n3647, n17358, n19538, n19537, n19536, n19535, 
        n19534, n19533, n19529, n19528, n19527, n19526, n19525, 
        n19524, n19521, n19520, n19519, n19518, n19517, n19516, 
        n19515, n19514, n19513, n19512, n19511, n19510, n19509, 
        n19508, n19507, n19101, n19100, n19099, n19098, n19097, 
        n19096, n19095, n19094, n19093, n19092, n19091, n19090, 
        n19089, n19088, n19087, n19086, n19085, n19084, n19083, 
        n19082, n19081, n19080, n19079, n19078, n19077, n19076, 
        n19075, n19074, n19073, n19506, n19505, n19504, n19503, 
        n19502, n19501, n19500, n19499, n19498, n19497, n19496, 
        n19495, n19494, n19493, n19492, n19491, n19490, n19489, 
        n19488, n19487, n19486, n19485, n6024, n19484, n19483, 
        n19482, n19481, n19480, n19479, n19478, n19477, n19476, 
        n19475, n19474, n19473, n19472, n19471, n19470, n19469, 
        n19468, n19467, n19466, n19465, n19464, n19463, n19462, 
        n19461, n4_adj_4925, n19460, n5523, n38214, n27827, n27826, 
        n28222, n28221, n28220, n32331, n27746, n28219, n19452, 
        n28218, n27745, n19072, n19071, n19070, n19451, n19450, 
        n19449, n19448, n34263, n28217, n19447, n28216, n19446, 
        n19445, quadA_debounced, quadB_debounced, n19444, n19443, 
        n19442, n19441, n24036, n19440, n19439, n19438, quadA_debounced_adj_4926, 
        quadB_debounced_adj_4927, n28215, n19437, n19436, n19435, 
        n4_adj_4928, n28214, n19434, n19069, n19068, n28213, n27737, 
        n28212, n28211, n19433, rw;
    wire [7:0]state_adj_5128;   // verilog/eeprom.v(23[11:16])
    
    wire n19432, n19431, n19430, n19429, n4_adj_4931, n19428, n19427, 
        n19426, n19425, n19424, n19423, n19422, n19421, n19420, 
        n19419, n6_adj_4932, n19418, n19417, n19416, n19415, n19414, 
        n19413, n19412, n19411, n19410, n19409, n19408, n19407, 
        n19406, r_Rx_Data;
    wire [2:0]r_Bit_Index;   // verilog/uart_rx.v(33[17:28])
    
    wire n28210, n19405, n19404, n19403, n19402, n19401, n19400, 
        n19399, n19398, n19397, n19396, n19395, n33367, n8_adj_4933, 
        n19067, n19394, n19393, n19392, n19066, n19391, n19390, 
        n38206, n15_adj_4934, n19389, n19388, n19387, n19386, n19385, 
        n19384, n19383, n19382, n19381, n19380, n19379, n19378, 
        n19377, n19376, n19375;
    wire [2:0]r_SM_Main_adj_5135;   // verilog/uart_tx.v(31[16:25])
    wire [2:0]r_Bit_Index_adj_5137;   // verilog/uart_tx.v(33[16:27])
    
    wire n37126, n6_adj_4936;
    wire [2:0]r_SM_Main_2__N_3487;
    
    wire n19374, n19373, n38205, n19372, n19371, n19370, n19369, 
        n19368, n19367, n19366, n19365, n19364, n63, n19363, n19362, 
        n19361, n19360, n19359, n19358, n19357, n19356, n19355, 
        n19354, n19353, n19352, n19351, n19350, n19349, n19348, 
        n19347, n19346, n19345;
    wire [1:0]reg_B;   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(142[19:24])
    
    wire n19344, n6027, n37058, n5690;
    wire [1:0]reg_B_adj_5146;   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(142[19:24])
    
    wire n37057, n19343, n19342, n19065;
    wire [7:0]state_adj_5158;   // verilog/i2c_controller.v(33[12:17])
    wire [7:0]saved_addr;   // verilog/i2c_controller.v(34[12:22])
    
    wire n19341, n19064, enable_slow_N_4001, n6026, n37130, n19340, 
        n31031, n15_adj_4940, n19339;
    wire [7:0]state_7__N_3898;
    
    wire n19338, n19337, n4_adj_4941, n19336, n37077, n5212, n19335, 
        n19334, n19333;
    wire [7:0]state_7__N_3914;
    
    wire n19332, n5410, n19331, n19330, n19329, n19328, n19327, 
        n19326, n19325, n19324, n19323, n5592, n19322, n19061, 
        n19060, n19057, n19056, n19321, n19320, n19319, n19318, 
        n19317, n19316, n19315, n19314, n19313, n19312, n19311, 
        n19310, n19309, n19308, n19307, n19306, n19305, n19304, 
        n19303, n19302, n19301, n19300, n19299, n19298, n19297, 
        n19296, n19295, n19294, n19293, n4_adj_4942, n19292, n19291, 
        n19290, n19289, n3_adj_4943, n19288, n19287, n19286, n19285, 
        n19284, n19283, n19282, n19281, n19280, n19279, n19278, 
        n19277, n19276, n19275, n19274, n19273, n19272, n19271, 
        n19270, n19269, n36967, n36965, n3_adj_4944, n5_adj_4945, 
        n6_adj_4946, n7_adj_4947, n8_adj_4948, n9_adj_4949, n10_adj_4950, 
        n11_adj_4951, n12_adj_4952, n13_adj_4953, n14_adj_4954, n15_adj_4955, 
        n16_adj_4956, n17_adj_4957, n18_adj_4958, n19_adj_4959, n20_adj_4960, 
        n21_adj_4961, n22_adj_4962, n23_adj_4963, n24_adj_4964, n25_adj_4965, 
        n5_adj_4966, n32660, n509, n510, n511, n36951, n513, n515, 
        n516, n517, n518, n519, n521, n523, n526, n36945, n598_adj_4967, 
        n619, n28209, n674, n675, n676, n677, n678, n679, n700, 
        n728, n729, n730, n731, n732, n733, n24827, n752, n753, 
        n754, n755, n756, n757, n758, n763, n765, n767, n768, 
        n770, n771_adj_4968, n772, n773, n774, n775, n778, n806, 
        n807, n808, n809, n810, n811, n812, n830, n831, n832, 
        n833, n834, n835, n836, n837, n856, n883, n884, n885, 
        n886, n887, n888, n889, n890, n891, n908, n909, n910, 
        n911, n912, n913, n914, n915, n916, n934, n961, n962, 
        n963, n964, n965, n966, n967, n968, n969, n970, n986, 
        n987, n988, n989, n990, n991, n992, n993, n994, n995, 
        n1012, n1039, n1040, n1041, n1042, n1043, n1044, n1045, 
        n1046, n1047, n1048, n1049, n28208, n1064, n1065, n1066, 
        n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, 
        n1090, n1117, n1118, n1119, n1120, n1121, n1122, n1123, 
        n1124, n1125, n1126, n1127, n1128, n1142, n1143, n1144, 
        n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, 
        n1153, n1168, n1195, n1196, n1197, n1198, n1199, n1200, 
        n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1220, 
        n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, 
        n1229, n1230, n1231, n1232, n1246, n1273, n1274, n1275, 
        n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, 
        n1284, n1285, n1286, n1298, n1299, n1300, n1301, n1302, 
        n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, 
        n1311, n1324, n1351, n1352, n1353, n1354, n1355, n1356, 
        n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364, 
        n1365, n1376, n1377, n1378, n1379, n1380, n1381, n1382, 
        n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, 
        n1402, n1429, n1430, n1431, n1432, n1433, n1434, n1435, 
        n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443, 
        n1444, n1454, n1455, n1456, n1457, n1458, n1459, n1460, 
        n1461, n1462, n1463, n1464, n1465, n1466, n1467, n1468, 
        n1469, n1480, n1507, n1508, n1509, n1510, n1511, n1512, 
        n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, 
        n1521, n1522, n1523, n1532, n1533, n1534, n1535, n1536, 
        n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544, 
        n1545, n1546, n1547, n1548, n1558, n32667, n1585, n1586, 
        n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594, 
        n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602, 
        n1610, n1611, n1612, n1613, n1614, n1615, n1616, n1617, 
        n1618, n1619, n1620, n1621, n1622, n1623, n1624, n1625, 
        n1626, n1627, n1636, n1663, n1664, n1665, n1666, n1667, 
        n1668, n1669, n1670, n1671, n1672, n1673, n1674, n1675, 
        n1676, n1677, n1678, n1679, n1680, n1681, n1688, n1689, 
        n1690, n1691, n1692, n1693, n1694, n1695, n1696, n1697, 
        n1698, n1699, n1700, n1701, n1702, n1703, n1704, n1705, 
        n1706, n1714, n1741, n1742, n1743, n1744, n1745, n1746, 
        n1747, n1748, n1749, n1750, n1751, n1752, n1753, n1754, 
        n1755, n1756, n1757, n1758, n1759, n1760, n1766, n1767, 
        n1768, n1769, n1770, n1771, n1772, n1773, n1774, n1775, 
        n1776, n1777, n1778, n1779, n1780, n1781, n1782, n1783, 
        n1784, n1785, n1792, n18956, n1819, n1820, n1821, n1822, 
        n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, 
        n1831, n1832, n1833, n1834, n1835, n1836, n1837, n1838, 
        n1839, n1844, n1845, n1846, n1847, n1848, n1849, n1850, 
        n1851, n1852, n1853, n1854, n1855, n1856, n1857, n1858, 
        n1859, n1860, n1861, n1862, n1863, n1864, n1870, n1897, 
        n1898, n1899, n1900, n1901, n1902, n1903, n1904, n1905, 
        n1906, n1907, n1908, n1909, n1910, n1911, n1912, n1913, 
        n1914, n1915, n1916, n1917, n1918, n1922, n1923, n1924, 
        n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932, 
        n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, 
        n1941, n1942, n1943, n1948, n1975, n1976, n1977, n1978, 
        n1979, n1980, n1981, n1982, n1983, n1984, n1985, n1986, 
        n1987, n1988, n1989, n1990, n1991, n1992, n1993, n1994, 
        n1995, n1996, n1997, n2000, n2001, n2002, n2003, n2004, 
        n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012, 
        n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020, 
        n2021, n2022, n2026, n2053, n2054, n2055, n2056, n2057, 
        n2058, n2059, n2060, n2061, n2062, n2063, n2064, n2065, 
        n2066, n2067, n2068, n2069, n2070, n2071, n2073, n2076, 
        n6223, n6222, n6221, n6220, n6219, n6218, n6217, n6216, 
        n6215, n6214, n6213, n6212, n6211, n6210, n6209, n6208, 
        n6207, n6206, n6205, n6203, n6202, n24_adj_4969, n18738, 
        n62, n18732, n17379, n17382, n32173, n17362, n18685, n4_adj_4970, 
        n18963, n35256, n32425, n19229, n18954, n19228, n19227, 
        n19226, n63_adj_4971, n19055, n19225, n34006, n7_adj_4972, 
        n19054, n19053, n17376, n17474, n19052, n19051, n19049, 
        n19047, n28207, n36878, n4_adj_4973, n6_adj_4974, n7_adj_4975, 
        n8_adj_4976, n9_adj_4977, n10_adj_4978, n11_adj_4979, n12_adj_4980, 
        n13_adj_4981, n15_adj_4982, n17_adj_4983, n19_adj_4984, n21_adj_4985, 
        n36966, n23_adj_4986, n25_adj_4987, n27_adj_4988, n36964, 
        n29_adj_4989, n30_adj_4990, n31, n33, n35, n36900, n28206, 
        n5_adj_4991, n16_adj_4992, n13_adj_4993, n12_adj_4994, n36814, 
        n36816, n28403, n36644, n6029, n28402, n33926, n36634, 
        n19224, n19223, n19222, n20_adj_4995, n18_adj_4996, n16_adj_4997, 
        n19046, n19044, n19043, n19042, n19041, n19040, n19035, 
        n19034, n19033, n19032, n19031, n19030, n8_adj_4998, n7_adj_4999, 
        n19165, n19164, n19163, n19162, n19161, n19160, n19159, 
        n19158, n12_adj_5000, n34, n31_adj_5001, n30_adj_5002, n28_adj_5003, 
        n2_adj_5004, n3_adj_5005, n4_adj_5006, n5_adj_5007, n6_adj_5008, 
        n7_adj_5009, n8_adj_5010, n9_adj_5011, n10_adj_5012, n11_adj_5013, 
        n12_adj_5014, n13_adj_5015, n14_adj_5016, n15_adj_5017, n16_adj_5018, 
        n17_adj_5019, n18_adj_5020, n19_adj_5021, n20_adj_5022, n21_adj_5023, 
        n22_adj_5024, n23_adj_5025, n24_adj_5026, n25_adj_5027, n22_adj_5028, 
        n21_adj_5029, n6_adj_5030, n38579, n35305, n12_adj_5031, n34_adj_5032, 
        n33_adj_5033, n32, n31_adj_5034, n30_adj_5035, n37, n36, 
        n30_adj_5036, n29_adj_5037, n32679, n28_adj_5038, n27_adj_5039, 
        n26, n25_adj_5040, n24_adj_5041, n35348, n23_adj_5042, n22_adj_5043, 
        n21_adj_5044, n32688, n7_adj_5045, n28401, n28400, n28205, 
        n28204, n13_adj_5046, n15_adj_5047, n17_adj_5048, n28399, 
        n28203, n33_adj_5049, n28398, n35_adj_5050, n28202, n37_adj_5051, 
        n39_adj_5052, n41, n43, n22_adj_5053, n20_adj_5054, n18_adj_5055, 
        n13_adj_5056, n15_adj_5057, n14_adj_5058, n36289, n14_adj_5059, 
        n10_adj_5060, n14_adj_5061, n9_adj_5062, n17_adj_5063, n16_adj_5064, 
        n28397, n7_adj_5065, n37131, n28396, n36277, n36276, n36275, 
        n10_adj_5066, n7_adj_5067, n14_adj_5068, n10_adj_5069, n32_adj_5070, 
        n48, n5_adj_5071, n19029, n34901, n36263, n14711, n28_adj_5072, 
        n17504, n27_adj_5073, n26_adj_5074, n25_adj_5075, n17534, 
        n17476, n28395, n10_adj_5076, n28201, n28200, n28199, n37129, 
        n28394, n36363, n36357, n36355, n36351, n36349, n28716, 
        n28715, n28714, n28713, n28712, n34410, n28711, n28710, 
        n28393, n28709, n28708, n28392, n28707, n35211, n35209, 
        n28706, n28705, n28704, n28703, n28391, n28702, n19023, 
        n28701, n19022, n28700, n28699, n28698, n28697, n28696, 
        n28695, n28694, n28_adj_5077, n28693, n26_adj_5078, n24_adj_5079, 
        n34029, n19_adj_5080, n28390, n28198, n28389, n28388, n34028, 
        n28387, n16_adj_5081, n35190, n28386, n27744, n28197, n34021, 
        n28385, n28384, n27743, n27742, n36224, n28383, n24819, 
        n24817, n17355, n17539, n28382, n24807, n23836, n34429, 
        n37281, n28381, n28380, n28379, n17506, n17518, n28188, 
        n28378, n24797, n28377, n28187, n28186, n28185, n28376, 
        n28184, n28183, n28182, n28375, n28374, n28181, n28180, 
        n28373, n27763, n37633, n28179, n28178, n28372, n28371, 
        n28177, n28370, n4_adj_5082, n24787, n28369, n28176, n28175, 
        n28368, n26_adj_5083, n24_adj_5084, n22_adj_5085, n14867, 
        n28367, n28366, n18_adj_5086, n28174, n27762, n28173, n28365, 
        n28172, n28171, n28364, n28363, n27761, n28362, n28361, 
        n28170, n27760, n36211, n8_adj_5087, n28169, n28360, n7_adj_5088, 
        n28168, n33567, n28359, n28167, n36208, n27759, n28166, 
        n27736, n27758, n36206, n17359, n28358, n28357, n28165, 
        n27735, n27734, n28356, n28355, n27757, n27733, n28354, 
        n27741, n28353;
    
    VCC i2 (.Y(VCC_net));
    \quad(DEBOUNCE_TICKS=100)_U1  quad_counter0 (.encoder0_position({encoder0_position}), 
            .GND_net(GND_net), .data_o({quadA_debounced, quadB_debounced}), 
            .clk32MHz(clk32MHz), .reg_B({reg_B}), .VCC_net(VCC_net), .n35256(n35256), 
            .n19049(n19049), .ENCODER0_B_c_0(ENCODER0_B_c_0), .n19588(n19588), 
            .ENCODER0_A_c_1(ENCODER0_A_c_1)) /* synthesis syn_module_defined=1 */ ;   // verilog/TinyFPGA_B.v(185[15] 190[4])
    SB_IO hall2_input (.PACKAGE_PIN(HALL2), .LATCH_INPUT_VALUE(GND_net), 
          .INPUT_CLK(GND_net), .OUTPUT_CLK(GND_net), .OUTPUT_ENABLE(GND_net), 
          .D_OUT_1(GND_net), .D_OUT_0(GND_net), .D_IN_0(hall2)) /* synthesis syn_instantiated=1, IO_FF_IN=TRUE */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam hall2_input.PIN_TYPE = 6'b000001;
    defparam hall2_input.PULLUP = 1'b1;
    defparam hall2_input.NEG_TRIGGER = 1'b0;
    defparam hall2_input.IO_STANDARD = "SB_LVCMOS";
    SB_IO hall3_input (.PACKAGE_PIN(HALL3), .LATCH_INPUT_VALUE(GND_net), 
          .INPUT_CLK(GND_net), .OUTPUT_CLK(GND_net), .OUTPUT_ENABLE(GND_net), 
          .D_OUT_1(GND_net), .D_OUT_0(GND_net), .D_IN_0(hall3)) /* synthesis syn_instantiated=1, IO_FF_IN=TRUE */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam hall3_input.PIN_TYPE = 6'b000001;
    defparam hall3_input.PULLUP = 1'b1;
    defparam hall3_input.NEG_TRIGGER = 1'b0;
    defparam hall3_input.IO_STANDARD = "SB_LVCMOS";
    SB_IO tx_output (.PACKAGE_PIN(TX), .LATCH_INPUT_VALUE(GND_net), .INPUT_CLK(GND_net), 
          .OUTPUT_CLK(GND_net), .OUTPUT_ENABLE(tx_enable), .D_OUT_1(GND_net), 
          .D_OUT_0(tx_o)) /* synthesis syn_instantiated=1 */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam tx_output.PIN_TYPE = 6'b101001;
    defparam tx_output.PULLUP = 1'b1;
    defparam tx_output.NEG_TRIGGER = 1'b0;
    defparam tx_output.IO_STANDARD = "SB_LVCMOS";
    SB_DFF h3_54 (.Q(INLB_c), .C(clk32MHz), .D(hall3));   // verilog/TinyFPGA_B.v(96[10] 109[6])
    SB_DFF displacement_i0 (.Q(displacement[0]), .C(clk32MHz), .D(displacement_23__N_58[0]));   // verilog/TinyFPGA_B.v(200[10] 203[6])
    SB_DFF h2_53 (.Q(INHB_c), .C(clk32MHz), .D(hall2));   // verilog/TinyFPGA_B.v(96[10] 109[6])
    SB_IO sda_output (.PACKAGE_PIN(SDA), .LATCH_INPUT_VALUE(GND_net), .INPUT_CLK(GND_net), 
          .OUTPUT_CLK(GND_net), .OUTPUT_ENABLE(sda_enable), .D_OUT_1(GND_net), 
          .D_OUT_0(sda_out), .D_IN_0(state_7__N_3914[3])) /* synthesis syn_instantiated=1 */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam sda_output.PIN_TYPE = 6'b101001;
    defparam sda_output.PULLUP = 1'b1;
    defparam sda_output.NEG_TRIGGER = 1'b0;
    defparam sda_output.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 i1_4_lut (.I0(n32_adj_5070), .I1(n2970), .I2(n17552), .I3(n4452), 
            .O(n32688));   // verilog/coms.v(127[12] 300[6])
    defparam i1_4_lut.LUT_INIT = 16'heeef;
    SB_IO CS_pad (.PACKAGE_PIN(CS), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(GND_net));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam CS_pad.PIN_TYPE = 6'b011001;
    defparam CS_pad.PULLUP = 1'b0;
    defparam CS_pad.NEG_TRIGGER = 1'b0;
    defparam CS_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO scl_output (.PACKAGE_PIN(SCL), .LATCH_INPUT_VALUE(GND_net), .INPUT_CLK(GND_net), 
          .OUTPUT_CLK(GND_net), .OUTPUT_ENABLE(scl_enable), .D_OUT_1(GND_net), 
          .D_OUT_0(scl)) /* synthesis syn_instantiated=1 */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam scl_output.PIN_TYPE = 6'b101001;
    defparam scl_output.PULLUP = 1'b1;
    defparam scl_output.NEG_TRIGGER = 1'b0;
    defparam scl_output.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 encoder0_position_23__I_0_unary_minus_2_add_3_25_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n3_adj_5005), .I3(n28715), .O(n3_adj_4924)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_unary_minus_2_add_3_25_lut.LUT_INIT = 16'hC33C;
    SB_IO hall1_input (.PACKAGE_PIN(HALL1), .LATCH_INPUT_VALUE(GND_net), 
          .INPUT_CLK(GND_net), .OUTPUT_CLK(GND_net), .OUTPUT_ENABLE(GND_net), 
          .D_OUT_1(GND_net), .D_OUT_0(GND_net), .D_IN_0(hall1)) /* synthesis syn_instantiated=1, IO_FF_IN=TRUE */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam hall1_input.PIN_TYPE = 6'b000001;
    defparam hall1_input.PULLUP = 1'b1;
    defparam hall1_input.NEG_TRIGGER = 1'b0;
    defparam hall1_input.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 i1_3_lut (.I0(n123), .I1(n32688), .I2(n63_adj_4971), .I3(GND_net), 
            .O(n7_adj_5067));   // verilog/coms.v(127[12] 300[6])
    defparam i1_3_lut.LUT_INIT = 16'h8c8c;
    SB_CARRY encoder0_position_23__I_0_unary_minus_2_add_3_25 (.CI(n28715), 
            .I0(GND_net), .I1(n3_adj_5005), .CO(n28716));
    neopixel nx (.\neo_pixel_transmitter.done (\neo_pixel_transmitter.done ), 
            .clk32MHz(clk32MHz), .\neo_pixel_transmitter.t0 ({\neo_pixel_transmitter.t0 }), 
            .GND_net(GND_net), .VCC_net(VCC_net), .timer({timer}), .start(start), 
            .n14(n14_adj_4896), .n24759(n24759), .\state[0] (state[0]), 
            .\state[1] (state[1]), .\state_3__N_402[1] (state_3__N_402[1]), 
            .LED_c(LED_c), .neopxl_color({neopxl_color}), .n18685(n18685), 
            .n33425(n33425), .n19040(n19040), .n19557(n19557), .n19556(n19556), 
            .n19555(n19555), .n19554(n19554), .n19553(n19553), .n19552(n19552), 
            .n19551(n19551), .n19550(n19550), .n19549(n19549), .n19548(n19548), 
            .n19547(n19547), .n19546(n19546), .n19545(n19545), .n19544(n19544), 
            .n19543(n19543), .n19542(n19542), .n19541(n19541), .n19540(n19540), 
            .n19539(n19539), .n19538(n19538), .n19537(n19537), .n19536(n19536), 
            .n19535(n19535), .n19534(n19534), .n19533(n19533), .n19529(n19529), 
            .n19528(n19528), .n19527(n19527), .n19526(n19526), .n19525(n19525), 
            .n19521(n19521), .NEOPXL_c(NEOPXL_c), .n33926(n33926), .n31453(n31453), 
            .n19022(n19022), .n34265(n34265)) /* synthesis syn_module_defined=1 */ ;   // verilog/TinyFPGA_B.v(43[10] 49[2])
    SB_LUT4 encoder0_position_23__I_0_unary_minus_2_add_3_24_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n4_adj_5006), .I3(n28714), .O(n4_adj_4923)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_unary_minus_2_add_3_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_unary_minus_2_add_3_24 (.CI(n28714), 
            .I0(GND_net), .I1(n4_adj_5006), .CO(n28715));
    SB_LUT4 encoder0_position_23__I_0_unary_minus_2_add_3_23_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n5_adj_5007), .I3(n28713), .O(n5_adj_4922)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_unary_minus_2_add_3_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i2_4_lut (.I0(n7_adj_5067), .I1(n123), .I2(n17476), .I3(n10417), 
            .O(n6_adj_4936));   // verilog/coms.v(127[12] 300[6])
    defparam i2_4_lut.LUT_INIT = 16'haeaf;
    SB_CARRY encoder0_position_23__I_0_unary_minus_2_add_3_23 (.CI(n28713), 
            .I0(GND_net), .I1(n5_adj_5007), .CO(n28714));
    SB_LUT4 i3_4_lut (.I0(n63), .I1(n6_adj_4936), .I2(n39), .I3(\FRAME_MATCHER.state_31__N_2662 [1]), 
            .O(n38205));   // verilog/coms.v(127[12] 300[6])
    defparam i3_4_lut.LUT_INIT = 16'hdfdd;
    SB_LUT4 encoder0_position_23__I_0_add_566_7_lut (.I0(GND_net), .I1(n833), 
            .I2(GND_net), .I3(n28130), .O(n886)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_566_7_lut.LUT_INIT = 16'hC33C;
    SB_DFFESR delay_counter_i0_i11 (.Q(delay_counter[11]), .C(CLK_c), .E(n5410), 
            .D(n593), .R(n18963));   // verilog/TinyFPGA_B.v(237[10] 265[6])
    SB_LUT4 encoder0_position_23__I_0_unary_minus_2_add_3_22_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n6_adj_5008), .I3(n28712), .O(n6_adj_4921)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_unary_minus_2_add_3_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_unary_minus_2_add_3_22 (.CI(n28712), 
            .I0(GND_net), .I1(n6_adj_5008), .CO(n28713));
    SB_LUT4 i13922_3_lut (.I0(PWMLimit[23]), .I1(\data_in_frame[8] [7]), 
            .I2(n33567), .I3(GND_net), .O(n19064));   // verilog/coms.v(127[12] 300[6])
    defparam i13922_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_23__I_0_add_566_7 (.CI(n28130), .I0(n833), 
            .I1(GND_net), .CO(n28131));
    SB_LUT4 i13923_3_lut (.I0(PWMLimit[22]), .I1(\data_in_frame[8] [6]), 
            .I2(n33567), .I3(GND_net), .O(n19065));   // verilog/coms.v(127[12] 300[6])
    defparam i13923_3_lut.LUT_INIT = 16'hacac;
    SB_DFF dir_58 (.Q(INHC_c), .C(clk32MHz), .D(duty[23]));   // verilog/TinyFPGA_B.v(96[10] 109[6])
    SB_LUT4 encoder0_position_23__I_0_unary_minus_2_add_3_21_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n7_adj_5009), .I3(n28711), .O(n7_adj_4920)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_unary_minus_2_add_3_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_unary_minus_2_add_3_21 (.CI(n28711), 
            .I0(GND_net), .I1(n7_adj_5009), .CO(n28712));
    SB_LUT4 encoder0_position_23__I_0_unary_minus_2_add_3_20_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n8_adj_5010), .I3(n28710), .O(n8_adj_4919)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_unary_minus_2_add_3_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i13924_3_lut (.I0(PWMLimit[21]), .I1(\data_in_frame[8] [5]), 
            .I2(n33567), .I3(GND_net), .O(n19066));   // verilog/coms.v(127[12] 300[6])
    defparam i13924_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_add_566_6_lut (.I0(GND_net), .I1(n834), 
            .I2(GND_net), .I3(n28129), .O(n887)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_566_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_566_6 (.CI(n28129), .I0(n834), 
            .I1(GND_net), .CO(n28130));
    SB_LUT4 encoder0_position_23__I_0_add_566_5_lut (.I0(GND_net), .I1(n835), 
            .I2(VCC_net), .I3(n28128), .O(n888)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_566_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_unary_minus_2_add_3_20 (.CI(n28710), 
            .I0(GND_net), .I1(n8_adj_5010), .CO(n28711));
    SB_LUT4 i13925_3_lut (.I0(PWMLimit[20]), .I1(\data_in_frame[8] [4]), 
            .I2(n33567), .I3(GND_net), .O(n19067));   // verilog/coms.v(127[12] 300[6])
    defparam i13925_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13926_3_lut (.I0(PWMLimit[19]), .I1(\data_in_frame[8] [3]), 
            .I2(n33567), .I3(GND_net), .O(n19068));   // verilog/coms.v(127[12] 300[6])
    defparam i13926_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_unary_minus_2_add_3_19_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n9_adj_5011), .I3(n28709), .O(n9_adj_4918)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_unary_minus_2_add_3_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i13927_3_lut (.I0(PWMLimit[18]), .I1(\data_in_frame[8] [2]), 
            .I2(n33567), .I3(GND_net), .O(n19069));   // verilog/coms.v(127[12] 300[6])
    defparam i13927_3_lut.LUT_INIT = 16'hacac;
    SB_DFFESR delay_counter_i0_i8 (.Q(delay_counter[8]), .C(CLK_c), .E(n5410), 
            .D(n596), .R(n18963));   // verilog/TinyFPGA_B.v(237[10] 265[6])
    SB_LUT4 i13928_3_lut (.I0(PWMLimit[17]), .I1(\data_in_frame[8] [1]), 
            .I2(n33567), .I3(GND_net), .O(n19070));   // verilog/coms.v(127[12] 300[6])
    defparam i13928_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13929_3_lut (.I0(PWMLimit[16]), .I1(\data_in_frame[8] [0]), 
            .I2(n33567), .I3(GND_net), .O(n19071));   // verilog/coms.v(127[12] 300[6])
    defparam i13929_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13930_3_lut (.I0(PWMLimit[15]), .I1(\data_in_frame[9] [7]), 
            .I2(n33567), .I3(GND_net), .O(n19072));   // verilog/coms.v(127[12] 300[6])
    defparam i13930_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13931_3_lut (.I0(PWMLimit[14]), .I1(\data_in_frame[9] [6]), 
            .I2(n33567), .I3(GND_net), .O(n19073));   // verilog/coms.v(127[12] 300[6])
    defparam i13931_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13932_3_lut (.I0(PWMLimit[13]), .I1(\data_in_frame[9] [5]), 
            .I2(n33567), .I3(GND_net), .O(n19074));   // verilog/coms.v(127[12] 300[6])
    defparam i13932_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13933_3_lut (.I0(PWMLimit[12]), .I1(\data_in_frame[9] [4]), 
            .I2(n33567), .I3(GND_net), .O(n19075));   // verilog/coms.v(127[12] 300[6])
    defparam i13933_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 unary_minus_4_inv_0_i8_1_lut (.I0(duty[7]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n18));   // verilog/TinyFPGA_B.v(106[23:28])
    defparam unary_minus_4_inv_0_i8_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_4_inv_0_i9_1_lut (.I0(duty[8]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n17));   // verilog/TinyFPGA_B.v(106[23:28])
    defparam unary_minus_4_inv_0_i9_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i13934_3_lut (.I0(PWMLimit[11]), .I1(\data_in_frame[9] [3]), 
            .I2(n33567), .I3(GND_net), .O(n19076));   // verilog/coms.v(127[12] 300[6])
    defparam i13934_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13935_3_lut (.I0(PWMLimit[10]), .I1(\data_in_frame[9] [2]), 
            .I2(n33567), .I3(GND_net), .O(n19077));   // verilog/coms.v(127[12] 300[6])
    defparam i13935_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13936_3_lut (.I0(PWMLimit[9]), .I1(\data_in_frame[9] [1]), 
            .I2(n33567), .I3(GND_net), .O(n19078));   // verilog/coms.v(127[12] 300[6])
    defparam i13936_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13937_3_lut (.I0(PWMLimit[8]), .I1(\data_in_frame[9] [0]), 
            .I2(n33567), .I3(GND_net), .O(n19079));   // verilog/coms.v(127[12] 300[6])
    defparam i13937_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13938_3_lut (.I0(PWMLimit[7]), .I1(\data_in_frame[10] [7]), 
            .I2(n33567), .I3(GND_net), .O(n19080));   // verilog/coms.v(127[12] 300[6])
    defparam i13938_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13939_3_lut (.I0(PWMLimit[6]), .I1(\data_in_frame[10] [6]), 
            .I2(n33567), .I3(GND_net), .O(n19081));   // verilog/coms.v(127[12] 300[6])
    defparam i13939_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13940_3_lut (.I0(PWMLimit[5]), .I1(\data_in_frame[10] [5]), 
            .I2(n33567), .I3(GND_net), .O(n19082));   // verilog/coms.v(127[12] 300[6])
    defparam i13940_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_23__I_0_add_566_5 (.CI(n28128), .I0(n835), 
            .I1(VCC_net), .CO(n28129));
    SB_LUT4 i13941_3_lut (.I0(PWMLimit[4]), .I1(\data_in_frame[10] [4]), 
            .I2(n33567), .I3(GND_net), .O(n19083));   // verilog/coms.v(127[12] 300[6])
    defparam i13941_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_add_566_4_lut (.I0(GND_net), .I1(n836), 
            .I2(GND_net), .I3(n28127), .O(n889)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_566_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_566_4 (.CI(n28127), .I0(n836), 
            .I1(GND_net), .CO(n28128));
    SB_DFFESR delay_counter_i0_i7 (.Q(delay_counter[7]), .C(CLK_c), .E(n5410), 
            .D(n597), .R(n18963));   // verilog/TinyFPGA_B.v(237[10] 265[6])
    SB_LUT4 i13942_3_lut (.I0(PWMLimit[3]), .I1(\data_in_frame[10] [3]), 
            .I2(n33567), .I3(GND_net), .O(n19084));   // verilog/coms.v(127[12] 300[6])
    defparam i13942_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_23__I_0_unary_minus_2_add_3_19 (.CI(n28709), 
            .I0(GND_net), .I1(n9_adj_5011), .CO(n28710));
    SB_DFFESR delay_counter_i0_i6 (.Q(delay_counter[6]), .C(CLK_c), .E(n5410), 
            .D(n598), .R(n18963));   // verilog/TinyFPGA_B.v(237[10] 265[6])
    SB_LUT4 encoder0_position_23__I_0_unary_minus_2_add_3_18_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n10_adj_5012), .I3(n28708), .O(n10_adj_4917)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_unary_minus_2_add_3_18_lut.LUT_INIT = 16'hC33C;
    SB_DFFESR delay_counter_i0_i5 (.Q(delay_counter[5]), .C(CLK_c), .E(n5410), 
            .D(n599), .R(n18963));   // verilog/TinyFPGA_B.v(237[10] 265[6])
    SB_LUT4 i13943_3_lut (.I0(PWMLimit[2]), .I1(\data_in_frame[10] [2]), 
            .I2(n33567), .I3(GND_net), .O(n19085));   // verilog/coms.v(127[12] 300[6])
    defparam i13943_3_lut.LUT_INIT = 16'hacac;
    SB_DFFESR delay_counter_i0_i4 (.Q(delay_counter[4]), .C(CLK_c), .E(n5410), 
            .D(n600), .R(n18963));   // verilog/TinyFPGA_B.v(237[10] 265[6])
    SB_DFFESR delay_counter_i0_i3 (.Q(delay_counter[3]), .C(CLK_c), .E(n5410), 
            .D(n601), .R(n18963));   // verilog/TinyFPGA_B.v(237[10] 265[6])
    SB_LUT4 mux_3363_i20_3_lut (.I0(encoder0_position[19]), .I1(n6_adj_4921), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n513));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam mux_3363_i20_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13944_3_lut (.I0(PWMLimit[1]), .I1(\data_in_frame[10] [1]), 
            .I2(n33567), .I3(GND_net), .O(n19086));   // verilog/coms.v(127[12] 300[6])
    defparam i13944_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mux_3363_i21_3_lut (.I0(encoder0_position[20]), .I1(n5_adj_4922), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n425));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam mux_3363_i21_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_3363_i22_3_lut (.I0(encoder0_position[21]), .I1(n4_adj_4923), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n511));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam mux_3363_i22_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_23__I_0_unary_minus_2_add_3_18 (.CI(n28708), 
            .I0(GND_net), .I1(n10_adj_5012), .CO(n28709));
    SB_LUT4 i13945_3_lut (.I0(control_mode[7]), .I1(\data_in_frame[1] [7]), 
            .I2(n33567), .I3(GND_net), .O(n19087));   // verilog/coms.v(127[12] 300[6])
    defparam i13945_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13946_3_lut (.I0(control_mode[6]), .I1(\data_in_frame[1] [6]), 
            .I2(n33567), .I3(GND_net), .O(n19088));   // verilog/coms.v(127[12] 300[6])
    defparam i13946_3_lut.LUT_INIT = 16'hacac;
    SB_DFFESR delay_counter_i0_i2 (.Q(delay_counter[2]), .C(CLK_c), .E(n5410), 
            .D(n602), .R(n18963));   // verilog/TinyFPGA_B.v(237[10] 265[6])
    SB_DFFESR delay_counter_i0_i1 (.Q(delay_counter[1]), .C(CLK_c), .E(n5410), 
            .D(n603), .R(n18963));   // verilog/TinyFPGA_B.v(237[10] 265[6])
    SB_LUT4 i13947_3_lut (.I0(control_mode[5]), .I1(\data_in_frame[1] [5]), 
            .I2(n33567), .I3(GND_net), .O(n19089));   // verilog/coms.v(127[12] 300[6])
    defparam i13947_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13948_3_lut (.I0(control_mode[4]), .I1(\data_in_frame[1] [4]), 
            .I2(n33567), .I3(GND_net), .O(n19090));   // verilog/coms.v(127[12] 300[6])
    defparam i13948_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13949_3_lut (.I0(control_mode[3]), .I1(\data_in_frame[1] [3]), 
            .I2(n33567), .I3(GND_net), .O(n19091));   // verilog/coms.v(127[12] 300[6])
    defparam i13949_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13950_3_lut (.I0(control_mode[2]), .I1(\data_in_frame[1] [2]), 
            .I2(n33567), .I3(GND_net), .O(n19092));   // verilog/coms.v(127[12] 300[6])
    defparam i13950_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13951_3_lut (.I0(control_mode[1]), .I1(\data_in_frame[1] [1]), 
            .I2(n33567), .I3(GND_net), .O(n19093));   // verilog/coms.v(127[12] 300[6])
    defparam i13951_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13952_3_lut (.I0(\data_in_frame[21] [7]), .I1(rx_data[7]), 
            .I2(n32679), .I3(GND_net), .O(n19094));   // verilog/coms.v(127[12] 300[6])
    defparam i13952_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13953_3_lut (.I0(\data_in_frame[21] [6]), .I1(rx_data[6]), 
            .I2(n32679), .I3(GND_net), .O(n19095));   // verilog/coms.v(127[12] 300[6])
    defparam i13953_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13954_3_lut (.I0(\data_in_frame[21] [5]), .I1(rx_data[5]), 
            .I2(n32679), .I3(GND_net), .O(n19096));   // verilog/coms.v(127[12] 300[6])
    defparam i13954_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13955_3_lut (.I0(\data_in_frame[21] [4]), .I1(rx_data[4]), 
            .I2(n32679), .I3(GND_net), .O(n19097));   // verilog/coms.v(127[12] 300[6])
    defparam i13955_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13956_3_lut (.I0(\data_in_frame[21] [3]), .I1(rx_data[3]), 
            .I2(n32679), .I3(GND_net), .O(n19098));   // verilog/coms.v(127[12] 300[6])
    defparam i13956_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13957_3_lut (.I0(\data_in_frame[21] [2]), .I1(rx_data[2]), 
            .I2(n32679), .I3(GND_net), .O(n19099));   // verilog/coms.v(127[12] 300[6])
    defparam i13957_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13958_3_lut (.I0(\data_in_frame[21] [1]), .I1(rx_data[1]), 
            .I2(n32679), .I3(GND_net), .O(n19100));   // verilog/coms.v(127[12] 300[6])
    defparam i13958_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13959_3_lut (.I0(\data_in_frame[21] [0]), .I1(rx_data[0]), 
            .I2(n32679), .I3(GND_net), .O(n19101));   // verilog/coms.v(127[12] 300[6])
    defparam i13959_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_unary_minus_2_add_3_17_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n11_adj_5013), .I3(n28707), .O(n11_adj_4916)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_unary_minus_2_add_3_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_unary_minus_2_add_3_17 (.CI(n28707), 
            .I0(GND_net), .I1(n11_adj_5013), .CO(n28708));
    SB_LUT4 encoder0_position_23__I_0_add_566_3_lut (.I0(GND_net), .I1(n837), 
            .I2(VCC_net), .I3(n28126), .O(n890)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_566_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_23__I_0_unary_minus_2_add_3_16_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n12_adj_5014), .I3(n28706), .O(n12_adj_4915)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_unary_minus_2_add_3_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_unary_minus_2_add_3_16 (.CI(n28706), 
            .I0(GND_net), .I1(n12_adj_5014), .CO(n28707));
    SB_LUT4 encoder0_position_23__I_0_unary_minus_2_add_3_15_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n13_adj_5015), .I3(n28705), .O(n13_adj_4914)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_unary_minus_2_add_3_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_unary_minus_2_add_3_15 (.CI(n28705), 
            .I0(GND_net), .I1(n13_adj_5015), .CO(n28706));
    SB_LUT4 encoder0_position_23__I_0_unary_minus_2_add_3_14_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n14_adj_5016), .I3(n28704), .O(n14_adj_4913)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_unary_minus_2_add_3_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_4_inv_0_i10_1_lut (.I0(duty[9]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n16));   // verilog/TinyFPGA_B.v(106[23:28])
    defparam unary_minus_4_inv_0_i10_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_4_inv_0_i11_1_lut (.I0(duty[10]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n15));   // verilog/TinyFPGA_B.v(106[23:28])
    defparam unary_minus_4_inv_0_i11_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY encoder0_position_23__I_0_unary_minus_2_add_3_14 (.CI(n28704), 
            .I0(GND_net), .I1(n14_adj_5016), .CO(n28705));
    SB_LUT4 encoder0_position_23__I_0_unary_minus_2_add_3_13_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n15_adj_5017), .I3(n28703), .O(n15_adj_4912)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_unary_minus_2_add_3_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_4_inv_0_i12_1_lut (.I0(duty[11]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n14));   // verilog/TinyFPGA_B.v(106[23:28])
    defparam unary_minus_4_inv_0_i12_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i26654_3_lut (.I0(encoder0_position[20]), .I1(n33397), .I2(encoder0_position[23]), 
            .I3(GND_net), .O(n677));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam i26654_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_23__I_0_unary_minus_2_add_3_13 (.CI(n28703), 
            .I0(GND_net), .I1(n15_adj_5017), .CO(n28704));
    SB_LUT4 encoder0_position_23__I_0_unary_minus_2_add_3_12_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n16_adj_5018), .I3(n28702), .O(n16_adj_4911)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_unary_minus_2_add_3_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_566_3 (.CI(n28126), .I0(n837), 
            .I1(VCC_net), .CO(n28127));
    SB_CARRY encoder0_position_23__I_0_unary_minus_2_add_3_12 (.CI(n28702), 
            .I0(GND_net), .I1(n16_adj_5018), .CO(n28703));
    SB_LUT4 encoder0_position_23__I_0_unary_minus_2_add_3_11_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n17_adj_5019), .I3(n28701), .O(n17_adj_4910)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_unary_minus_2_add_3_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_23__I_0_add_566_2_lut (.I0(GND_net), .I1(n517), 
            .I2(GND_net), .I3(VCC_net), .O(n891)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_566_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_unary_minus_2_add_3_11 (.CI(n28701), 
            .I0(GND_net), .I1(n17_adj_5019), .CO(n28702));
    SB_LUT4 encoder0_position_23__I_0_unary_minus_2_add_3_10_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n18_adj_5020), .I3(n28700), .O(n18_adj_4909)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_unary_minus_2_add_3_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i28543_1_lut (.I0(n4_adj_4970), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n35293));
    defparam i28543_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mux_3363_i23_3_lut (.I0(encoder0_position[22]), .I1(n3_adj_4924), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n510));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam mux_3363_i23_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_23__I_0_unary_minus_2_add_3_10 (.CI(n28700), 
            .I0(GND_net), .I1(n18_adj_5020), .CO(n28701));
    SB_LUT4 encoder0_position_23__I_0_unary_minus_2_add_3_9_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n19_adj_5021), .I3(n28699), .O(n19_adj_4908)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_unary_minus_2_add_3_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_unary_minus_2_add_3_9 (.CI(n28699), 
            .I0(GND_net), .I1(n19_adj_5021), .CO(n28700));
    SB_LUT4 encoder0_position_23__I_0_unary_minus_2_add_3_8_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n20_adj_5022), .I3(n28698), .O(n20_adj_4907)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_unary_minus_2_add_3_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_unary_minus_2_add_3_8 (.CI(n28698), 
            .I0(GND_net), .I1(n20_adj_5022), .CO(n28699));
    SB_LUT4 encoder0_position_23__I_0_unary_minus_2_add_3_7_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n21_adj_5023), .I3(n28697), .O(n21_adj_4906)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_unary_minus_2_add_3_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_unary_minus_2_add_3_7 (.CI(n28697), 
            .I0(GND_net), .I1(n21_adj_5023), .CO(n28698));
    SB_LUT4 encoder0_position_23__I_0_unary_minus_2_add_3_6_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n22_adj_5024), .I3(n28696), .O(n22_adj_4905)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_unary_minus_2_add_3_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_unary_minus_2_add_3_6 (.CI(n28696), 
            .I0(GND_net), .I1(n22_adj_5024), .CO(n28697));
    SB_LUT4 encoder0_position_23__I_0_unary_minus_2_add_3_5_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n23_adj_5025), .I3(n28695), .O(n23_adj_4904)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_unary_minus_2_add_3_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_unary_minus_2_add_3_5 (.CI(n28695), 
            .I0(GND_net), .I1(n23_adj_5025), .CO(n28696));
    SB_LUT4 encoder0_position_23__I_0_unary_minus_2_add_3_4_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n24_adj_5026), .I3(n28694), .O(n24_adj_4903)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_unary_minus_2_add_3_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_unary_minus_2_add_3_4 (.CI(n28694), 
            .I0(GND_net), .I1(n24_adj_5026), .CO(n28695));
    SB_LUT4 encoder0_position_23__I_0_unary_minus_2_add_3_3_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n25_adj_5027), .I3(n28693), .O(n25_adj_4902)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_unary_minus_2_add_3_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_unary_minus_2_add_3_3 (.CI(n28693), 
            .I0(GND_net), .I1(n25_adj_5027), .CO(n28694));
    SB_CARRY encoder0_position_23__I_0_unary_minus_2_add_3_2 (.CI(VCC_net), 
            .I0(GND_net), .I1(VCC_net), .CO(n28693));
    SB_LUT4 unary_minus_4_inv_0_i13_1_lut (.I0(duty[12]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n13));   // verilog/TinyFPGA_B.v(106[23:28])
    defparam unary_minus_4_inv_0_i13_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mux_3363_i18_3_lut (.I0(encoder0_position[17]), .I1(n8_adj_4919), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n515));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam mux_3363_i18_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i30526_1_lut (.I0(n700), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n37281));
    defparam i30526_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i30568_1_lut (.I0(n778), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n37323));
    defparam i30568_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 LessThan_744_i9_2_lut (.I0(pwm_counter[4]), .I1(pwm_setpoint[4]), 
            .I2(GND_net), .I3(GND_net), .O(n9_adj_4977));   // verilog/pwm.v(21[8:24])
    defparam LessThan_744_i9_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_744_i11_2_lut (.I0(pwm_counter[5]), .I1(pwm_setpoint[5]), 
            .I2(GND_net), .I3(GND_net), .O(n11_adj_4979));   // verilog/pwm.v(21[8:24])
    defparam LessThan_744_i11_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_744_i17_2_lut (.I0(pwm_counter[8]), .I1(pwm_setpoint[8]), 
            .I2(GND_net), .I3(GND_net), .O(n17_adj_4983));   // verilog/pwm.v(21[8:24])
    defparam LessThan_744_i17_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_744_i27_2_lut (.I0(pwm_counter[13]), .I1(pwm_setpoint[13]), 
            .I2(GND_net), .I3(GND_net), .O(n27_adj_4988));   // verilog/pwm.v(21[8:24])
    defparam LessThan_744_i27_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_744_i15_2_lut (.I0(pwm_counter[7]), .I1(pwm_setpoint[7]), 
            .I2(GND_net), .I3(GND_net), .O(n15_adj_4982));   // verilog/pwm.v(21[8:24])
    defparam LessThan_744_i15_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_744_i13_2_lut (.I0(pwm_counter[6]), .I1(pwm_setpoint[6]), 
            .I2(GND_net), .I3(GND_net), .O(n13_adj_4981));   // verilog/pwm.v(21[8:24])
    defparam LessThan_744_i13_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_744_i7_2_lut (.I0(pwm_counter[3]), .I1(pwm_setpoint[3]), 
            .I2(GND_net), .I3(GND_net), .O(n7_adj_4975));   // verilog/pwm.v(21[8:24])
    defparam LessThan_744_i7_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_744_i21_2_lut (.I0(pwm_counter[10]), .I1(pwm_setpoint[10]), 
            .I2(GND_net), .I3(GND_net), .O(n21_adj_4985));   // verilog/pwm.v(21[8:24])
    defparam LessThan_744_i21_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_744_i23_2_lut (.I0(pwm_counter[11]), .I1(pwm_setpoint[11]), 
            .I2(GND_net), .I3(GND_net), .O(n23_adj_4986));   // verilog/pwm.v(21[8:24])
    defparam LessThan_744_i23_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_744_i19_2_lut (.I0(pwm_counter[9]), .I1(pwm_setpoint[9]), 
            .I2(GND_net), .I3(GND_net), .O(n19_adj_4984));   // verilog/pwm.v(21[8:24])
    defparam LessThan_744_i19_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_744_i29_2_lut (.I0(pwm_counter[14]), .I1(pwm_setpoint[14]), 
            .I2(GND_net), .I3(GND_net), .O(n29_adj_4989));   // verilog/pwm.v(21[8:24])
    defparam LessThan_744_i29_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_744_i31_2_lut (.I0(pwm_counter[15]), .I1(pwm_setpoint[15]), 
            .I2(GND_net), .I3(GND_net), .O(n31));   // verilog/pwm.v(21[8:24])
    defparam LessThan_744_i31_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_744_i33_2_lut (.I0(pwm_counter[16]), .I1(pwm_setpoint[16]), 
            .I2(GND_net), .I3(GND_net), .O(n33));   // verilog/pwm.v(21[8:24])
    defparam LessThan_744_i33_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_744_i25_2_lut (.I0(pwm_counter[12]), .I1(pwm_setpoint[12]), 
            .I2(GND_net), .I3(GND_net), .O(n25_adj_4987));   // verilog/pwm.v(21[8:24])
    defparam LessThan_744_i25_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 unary_minus_4_inv_0_i14_1_lut (.I0(duty[13]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n12));   // verilog/TinyFPGA_B.v(106[23:28])
    defparam unary_minus_4_inv_0_i14_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY encoder0_position_23__I_0_add_566_2 (.CI(VCC_net), .I0(n517), 
            .I1(GND_net), .CO(n28126));
    SB_DFFESR delay_counter_i0_i10 (.Q(delay_counter[10]), .C(CLK_c), .E(n5410), 
            .D(n594), .R(n18963));   // verilog/TinyFPGA_B.v(237[10] 265[6])
    SB_LUT4 encoder0_position_23__I_0_i1371_3_lut (.I0(n2008), .I1(n2061), 
            .I2(n2026), .I3(GND_net), .O(n33_adj_5049));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1371_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1380_3_lut (.I0(n2017), .I1(n2070), 
            .I2(n2026), .I3(GND_net), .O(n15_adj_5047));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1380_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1367_3_lut (.I0(n2004), .I1(n2057), 
            .I2(n2026), .I3(GND_net), .O(n41));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1367_3_lut.LUT_INIT = 16'hacac;
    SB_DFFESR delay_counter_i0_i18 (.Q(delay_counter[18]), .C(CLK_c), .E(n5410), 
            .D(n586), .R(n18963));   // verilog/TinyFPGA_B.v(237[10] 265[6])
    SB_LUT4 encoder0_position_23__I_0_i1370_3_lut (.I0(n2007), .I1(n2060), 
            .I2(n2026), .I3(GND_net), .O(n35_adj_5050));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1370_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1368_3_lut (.I0(n2005), .I1(n2058), 
            .I2(n2026), .I3(GND_net), .O(n39_adj_5052));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1368_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1381_3_lut (.I0(n2018), .I1(n2071), 
            .I2(n2026), .I3(GND_net), .O(n13_adj_5046));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1381_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1379_3_lut (.I0(n2016), .I1(n2069), 
            .I2(n2026), .I3(GND_net), .O(n17_adj_5048));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1379_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1366_3_lut (.I0(n2003), .I1(n2056), 
            .I2(n2026), .I3(GND_net), .O(n43));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1366_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i4_4_lut (.I0(n2010), .I1(n33_adj_5049), .I2(n2063), .I3(n2026), 
            .O(n24_adj_5041));
    defparam i4_4_lut.LUT_INIT = 16'heefc;
    SB_LUT4 i2_4_lut_adj_1630 (.I0(n2001), .I1(n17_adj_5048), .I2(n2054), 
            .I3(n2026), .O(n22_adj_5043));
    defparam i2_4_lut_adj_1630.LUT_INIT = 16'heefc;
    SB_LUT4 i3_4_lut_adj_1631 (.I0(n2012), .I1(n13_adj_5046), .I2(n2065), 
            .I3(n2026), .O(n23_adj_5042));
    defparam i3_4_lut_adj_1631.LUT_INIT = 16'heefc;
    SB_LUT4 i1_4_lut_adj_1632 (.I0(n2014), .I1(n43), .I2(n2067), .I3(n2026), 
            .O(n21_adj_5044));
    defparam i1_4_lut_adj_1632.LUT_INIT = 16'heefc;
    SB_LUT4 encoder0_position_23__I_0_i1369_3_lut (.I0(n2006), .I1(n2059), 
            .I2(n2026), .I3(GND_net), .O(n37_adj_5051));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1369_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16_4_lut (.I0(n2020), .I1(n36224), .I2(n2026), .I3(n2019), 
            .O(n5_adj_4897));
    defparam i16_4_lut.LUT_INIT = 16'hac0c;
    SB_DFFESR delay_counter_i0_i17 (.Q(delay_counter[17]), .C(CLK_c), .E(n5410), 
            .D(n587), .R(n18963));   // verilog/TinyFPGA_B.v(237[10] 265[6])
    SB_LUT4 i29636_3_lut (.I0(n775), .I1(n2021), .I2(n2022), .I3(GND_net), 
            .O(n36276));
    defparam i29636_3_lut.LUT_INIT = 16'hecec;
    SB_LUT4 i19604_4_lut (.I0(n515), .I1(n677), .I2(n678), .I3(n679), 
            .O(n24747));
    defparam i19604_4_lut.LUT_INIT = 16'hfcec;
    SB_LUT4 i1_4_lut_adj_1633 (.I0(n36276), .I1(n5_adj_4897), .I2(n36277), 
            .I3(n2026), .O(n31031));
    defparam i1_4_lut_adj_1633.LUT_INIT = 16'h88c0;
    SB_LUT4 i14016_3_lut (.I0(\data_in_frame[13] [7]), .I1(rx_data[7]), 
            .I2(n32667), .I3(GND_net), .O(n19158));   // verilog/coms.v(127[12] 300[6])
    defparam i14016_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14017_3_lut (.I0(\data_in_frame[13] [6]), .I1(rx_data[6]), 
            .I2(n32667), .I3(GND_net), .O(n19159));   // verilog/coms.v(127[12] 300[6])
    defparam i14017_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i8_4_lut (.I0(n2013), .I1(n15_adj_5047), .I2(n2066), .I3(n2026), 
            .O(n28_adj_5038));
    defparam i8_4_lut.LUT_INIT = 16'heefc;
    SB_DFF pwm_setpoint_i0 (.Q(pwm_setpoint[0]), .C(clk32MHz), .D(pwm_setpoint_22__N_11[0]));   // verilog/TinyFPGA_B.v(96[10] 109[6])
    SB_LUT4 i6_4_lut (.I0(n2000), .I1(n41), .I2(n2053), .I3(n2026), 
            .O(n26));
    defparam i6_4_lut.LUT_INIT = 16'heefc;
    SB_LUT4 i7_4_lut (.I0(n2002), .I1(n35_adj_5050), .I2(n2055), .I3(n2026), 
            .O(n27_adj_5039));
    defparam i7_4_lut.LUT_INIT = 16'heefc;
    SB_LUT4 i5_4_lut (.I0(n2011), .I1(n31031), .I2(n2064), .I3(n2026), 
            .O(n25_adj_5040));
    defparam i5_4_lut.LUT_INIT = 16'heefc;
    SB_LUT4 i10_4_lut (.I0(n2009), .I1(n39_adj_5052), .I2(n2062), .I3(n2026), 
            .O(n30_adj_5036));
    defparam i10_4_lut.LUT_INIT = 16'heefc;
    SB_LUT4 i16_4_lut_adj_1634 (.I0(n21_adj_5044), .I1(n23_adj_5042), .I2(n22_adj_5043), 
            .I3(n24_adj_5041), .O(n36));
    defparam i16_4_lut_adj_1634.LUT_INIT = 16'hfffe;
    SB_LUT4 i14018_3_lut (.I0(\data_in_frame[13] [5]), .I1(rx_data[5]), 
            .I2(n32667), .I3(GND_net), .O(n19160));   // verilog/coms.v(127[12] 300[6])
    defparam i14018_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i9_4_lut (.I0(n2015), .I1(n37_adj_5051), .I2(n2068), .I3(n2026), 
            .O(n29_adj_5037));
    defparam i9_4_lut.LUT_INIT = 16'heefc;
    SB_LUT4 i17_4_lut (.I0(n25_adj_5040), .I1(n27_adj_5039), .I2(n26), 
            .I3(n28_adj_5038), .O(n37));
    defparam i17_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i14019_3_lut (.I0(\data_in_frame[13] [4]), .I1(rx_data[4]), 
            .I2(n32667), .I3(GND_net), .O(n19161));   // verilog/coms.v(127[12] 300[6])
    defparam i14019_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i30837_4_lut (.I0(n37), .I1(n29_adj_5037), .I2(n36), .I3(n30_adj_5036), 
            .O(n24787));
    defparam i30837_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 i14020_3_lut (.I0(\data_in_frame[13] [3]), .I1(rx_data[3]), 
            .I2(n32667), .I3(GND_net), .O(n19162));   // verilog/coms.v(127[12] 300[6])
    defparam i14020_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14021_3_lut (.I0(\data_in_frame[13] [2]), .I1(rx_data[2]), 
            .I2(n32667), .I3(GND_net), .O(n19163));   // verilog/coms.v(127[12] 300[6])
    defparam i14021_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14022_3_lut (.I0(\data_in_frame[13] [1]), .I1(rx_data[1]), 
            .I2(n32667), .I3(GND_net), .O(n19164));   // verilog/coms.v(127[12] 300[6])
    defparam i14022_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 unary_minus_4_inv_0_i15_1_lut (.I0(duty[14]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n11));   // verilog/TinyFPGA_B.v(106[23:28])
    defparam unary_minus_4_inv_0_i15_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i14023_3_lut (.I0(\data_in_frame[13] [0]), .I1(rx_data[0]), 
            .I2(n32667), .I3(GND_net), .O(n19165));   // verilog/coms.v(127[12] 300[6])
    defparam i14023_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_add_513_9_lut (.I0(n37323), .I1(n752), 
            .I2(VCC_net), .I3(n28125), .O(n830)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_513_9_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i30536_4_lut (.I0(n676), .I1(n674), .I2(n675), .I3(n24747), 
            .O(n700));
    defparam i30536_4_lut.LUT_INIT = 16'h1333;
    SB_LUT4 i26658_3_lut (.I0(encoder0_position[18]), .I1(n33401), .I2(encoder0_position[23]), 
            .I3(GND_net), .O(n679));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam i26658_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_23__I_0_i467_3_lut (.I0(n679), .I1(n732), 
            .I2(n700), .I3(GND_net), .O(n757));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i467_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i466_3_lut (.I0(n678), .I1(n731), 
            .I2(n700), .I3(GND_net), .O(n756));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i466_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_add_513_8_lut (.I0(GND_net), .I1(n753), 
            .I2(VCC_net), .I3(n28124), .O(n806)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_513_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_513_8 (.CI(n28124), .I0(n753), 
            .I1(VCC_net), .CO(n28125));
    SB_LUT4 i30861_2_lut_3_lut (.I0(n3_adj_4924), .I1(n4_adj_4970), .I2(encoder0_position[23]), 
            .I3(GND_net), .O(n619));
    defparam i30861_2_lut_3_lut.LUT_INIT = 16'h7f7f;
    SB_DFF h1_52 (.Q(INLA_c), .C(clk32MHz), .D(hall1));   // verilog/TinyFPGA_B.v(96[10] 109[6])
    SB_LUT4 i26626_3_lut_4_lut (.I0(n3_adj_4924), .I1(n4_adj_4970), .I2(n6026), 
            .I3(n4_adj_4923), .O(n33367));
    defparam i26626_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_IO INLC_pad (.PACKAGE_PIN(INLC), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(VCC_net));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam INLC_pad.PIN_TYPE = 6'b011001;
    defparam INLC_pad.PULLUP = 1'b0;
    defparam INLC_pad.NEG_TRIGGER = 1'b0;
    defparam INLC_pad.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 encoder0_position_23__I_0_i464_3_lut (.I0(n676), .I1(n729), 
            .I2(n700), .I3(GND_net), .O(n754));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i464_3_lut.LUT_INIT = 16'hacac;
    SB_DFFESR delay_counter_i0_i9 (.Q(delay_counter[9]), .C(CLK_c), .E(n5410), 
            .D(n595), .R(n18963));   // verilog/TinyFPGA_B.v(237[10] 265[6])
    SB_LUT4 encoder0_position_23__I_0_i468_3_lut (.I0(n515), .I1(n733), 
            .I2(n700), .I3(GND_net), .O(n758));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i468_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mux_3363_i17_3_lut (.I0(encoder0_position[16]), .I1(n9_adj_4918), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n516));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam mux_3363_i17_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 unary_minus_4_inv_0_i1_1_lut (.I0(duty[0]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n25));   // verilog/TinyFPGA_B.v(106[23:28])
    defparam unary_minus_4_inv_0_i1_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_23__I_0_add_513_7_lut (.I0(GND_net), .I1(n754), 
            .I2(GND_net), .I3(n28123), .O(n807)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_513_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i26655_3_lut_4_lut (.I0(n3_adj_4924), .I1(n4_adj_4970), .I2(n6028), 
            .I3(n6_adj_4921), .O(n33399));
    defparam i26655_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i26653_3_lut_4_lut (.I0(n3_adj_4924), .I1(n4_adj_4970), .I2(n6027), 
            .I3(n5_adj_4922), .O(n33397));
    defparam i26653_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i26657_3_lut_4_lut (.I0(n3_adj_4924), .I1(n4_adj_4970), .I2(n6029), 
            .I3(n7_adj_4920), .O(n33401));
    defparam i26657_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 encoder1_position_23__I_0_inv_0_i1_1_lut (.I0(encoder0_position_scaled[0]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n25_adj_4965));   // verilog/TinyFPGA_B.v(202[21:65])
    defparam encoder1_position_23__I_0_inv_0_i1_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_4_inv_0_i16_1_lut (.I0(duty[15]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n10_adj_4887));   // verilog/TinyFPGA_B.v(106[23:28])
    defparam unary_minus_4_inv_0_i16_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder1_position_23__I_0_inv_0_i2_1_lut (.I0(encoder0_position_scaled[1]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n24_adj_4964));   // verilog/TinyFPGA_B.v(202[21:65])
    defparam encoder1_position_23__I_0_inv_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder1_position_23__I_0_inv_0_i3_1_lut (.I0(encoder0_position_scaled[2]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n23_adj_4963));   // verilog/TinyFPGA_B.v(202[21:65])
    defparam encoder1_position_23__I_0_inv_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder1_position_23__I_0_inv_0_i4_1_lut (.I0(encoder0_position_scaled[3]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n22_adj_4962));   // verilog/TinyFPGA_B.v(202[21:65])
    defparam encoder1_position_23__I_0_inv_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY encoder0_position_23__I_0_add_513_7 (.CI(n28123), .I0(n754), 
            .I1(GND_net), .CO(n28124));
    SB_LUT4 encoder1_position_23__I_0_inv_0_i5_1_lut (.I0(encoder0_position_scaled[4]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n21_adj_4961));   // verilog/TinyFPGA_B.v(202[21:65])
    defparam encoder1_position_23__I_0_inv_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_4_inv_0_i17_1_lut (.I0(duty[16]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n9));   // verilog/TinyFPGA_B.v(106[23:28])
    defparam unary_minus_4_inv_0_i17_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder1_position_23__I_0_inv_0_i6_1_lut (.I0(encoder0_position_scaled[5]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n20_adj_4960));   // verilog/TinyFPGA_B.v(202[21:65])
    defparam encoder1_position_23__I_0_inv_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i19111_2_lut (.I0(n516), .I1(n758), .I2(GND_net), .I3(GND_net), 
            .O(n24244));
    defparam i19111_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 encoder0_position_23__I_0_add_513_6_lut (.I0(GND_net), .I1(n755), 
            .I2(GND_net), .I3(n28122), .O(n808)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_513_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_513_6 (.CI(n28122), .I0(n755), 
            .I1(GND_net), .CO(n28123));
    SB_LUT4 encoder0_position_23__I_0_add_513_5_lut (.I0(GND_net), .I1(n756), 
            .I2(VCC_net), .I3(n28121), .O(n809)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_513_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_4_inv_0_i18_1_lut (.I0(duty[17]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n8));   // verilog/TinyFPGA_B.v(106[23:28])
    defparam unary_minus_4_inv_0_i18_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder1_position_23__I_0_inv_0_i7_1_lut (.I0(encoder0_position_scaled[6]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n19_adj_4959));   // verilog/TinyFPGA_B.v(202[21:65])
    defparam encoder1_position_23__I_0_inv_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_4_inv_0_i19_1_lut (.I0(duty[18]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n7_adj_4886));   // verilog/TinyFPGA_B.v(106[23:28])
    defparam unary_minus_4_inv_0_i19_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder1_position_23__I_0_inv_0_i8_1_lut (.I0(encoder0_position_scaled[7]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n18_adj_4958));   // verilog/TinyFPGA_B.v(202[21:65])
    defparam encoder1_position_23__I_0_inv_0_i8_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY encoder0_position_23__I_0_add_513_5 (.CI(n28121), .I0(n756), 
            .I1(VCC_net), .CO(n28122));
    SB_LUT4 add_25_13_lut (.I0(GND_net), .I1(delay_counter[11]), .I2(GND_net), 
            .I3(n27743), .O(n593)) /* synthesis syn_instantiated=1 */ ;
    defparam add_25_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_23__I_0_add_513_4_lut (.I0(GND_net), .I1(n757), 
            .I2(GND_net), .I3(n28120), .O(n810)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_513_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_513_4 (.CI(n28120), .I0(n757), 
            .I1(GND_net), .CO(n28121));
    SB_LUT4 encoder0_position_23__I_0_add_513_3_lut (.I0(GND_net), .I1(n758), 
            .I2(VCC_net), .I3(n28119), .O(n811)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_513_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_513_3 (.CI(n28119), .I0(n758), 
            .I1(VCC_net), .CO(n28120));
    SB_LUT4 encoder0_position_23__I_0_add_513_2_lut (.I0(GND_net), .I1(n516), 
            .I2(GND_net), .I3(VCC_net), .O(n812)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_513_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_513_2 (.CI(VCC_net), .I0(n516), 
            .I1(GND_net), .CO(n28119));
    SB_LUT4 add_25_5_lut (.I0(GND_net), .I1(delay_counter[3]), .I2(GND_net), 
            .I3(n27735), .O(n601)) /* synthesis syn_instantiated=1 */ ;
    defparam add_25_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_23__I_0_add_460_8_lut (.I0(n37281), .I1(n674), 
            .I2(VCC_net), .I3(n28118), .O(n752)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_460_8_lut.LUT_INIT = 16'h8228;
    SB_LUT4 encoder0_position_23__I_0_add_460_7_lut (.I0(GND_net), .I1(n675), 
            .I2(GND_net), .I3(n28117), .O(n728)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_460_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_25_13 (.CI(n27743), .I0(delay_counter[11]), .I1(GND_net), 
            .CO(n27744));
    SB_CARRY encoder0_position_23__I_0_add_460_7 (.CI(n28117), .I0(n675), 
            .I1(GND_net), .CO(n28118));
    SB_LUT4 add_25_12_lut (.I0(GND_net), .I1(delay_counter[10]), .I2(GND_net), 
            .I3(n27742), .O(n594)) /* synthesis syn_instantiated=1 */ ;
    defparam add_25_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_23__I_0_add_460_6_lut (.I0(GND_net), .I1(n676), 
            .I2(GND_net), .I3(n28116), .O(n729)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_460_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_460_6 (.CI(n28116), .I0(n676), 
            .I1(GND_net), .CO(n28117));
    SB_LUT4 encoder0_position_23__I_0_add_460_5_lut (.I0(GND_net), .I1(n677), 
            .I2(VCC_net), .I3(n28115), .O(n730)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_460_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_460_5 (.CI(n28115), .I0(n677), 
            .I1(VCC_net), .CO(n28116));
    SB_CARRY add_25_12 (.CI(n27742), .I0(delay_counter[10]), .I1(GND_net), 
            .CO(n27743));
    SB_IO RX_pad (.PACKAGE_PIN(RX), .OUTPUT_ENABLE(VCC_net), .D_IN_0(RX_c));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam RX_pad.PIN_TYPE = 6'b000001;
    defparam RX_pad.PULLUP = 1'b0;
    defparam RX_pad.NEG_TRIGGER = 1'b0;
    defparam RX_pad.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 encoder0_position_23__I_0_add_460_4_lut (.I0(GND_net), .I1(n678), 
            .I2(GND_net), .I3(n28114), .O(n731)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_460_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_4_lut_adj_1635 (.I0(n754), .I1(n24244), .I2(n756), .I3(n757), 
            .O(n4_adj_4925));
    defparam i1_4_lut_adj_1635.LUT_INIT = 16'ha8a0;
    SB_CARRY add_25_5 (.CI(n27735), .I0(delay_counter[3]), .I1(GND_net), 
            .CO(n27736));
    SB_CARRY encoder0_position_23__I_0_add_460_4 (.CI(n28114), .I0(n678), 
            .I1(GND_net), .CO(n28115));
    SB_LUT4 encoder0_position_23__I_0_add_460_3_lut (.I0(GND_net), .I1(n679), 
            .I2(VCC_net), .I3(n28113), .O(n732)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_460_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_25_11_lut (.I0(GND_net), .I1(delay_counter[9]), .I2(GND_net), 
            .I3(n27741), .O(n595)) /* synthesis syn_instantiated=1 */ ;
    defparam add_25_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_460_3 (.CI(n28113), .I0(n679), 
            .I1(VCC_net), .CO(n28114));
    SB_LUT4 encoder0_position_23__I_0_add_460_2_lut (.I0(GND_net), .I1(n515), 
            .I2(GND_net), .I3(VCC_net), .O(n733)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_460_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_460_2 (.CI(VCC_net), .I0(n515), 
            .I1(GND_net), .CO(n28113));
    SB_LUT4 add_1872_7_lut (.I0(GND_net), .I1(n509), .I2(GND_net), .I3(n28003), 
            .O(n6024)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1872_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_1872_6_lut (.I0(n35293), .I1(n510), .I2(GND_net), .I3(n28002), 
            .O(n36211)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1872_6_lut.LUT_INIT = 16'hebbe;
    SB_CARRY add_1872_6 (.CI(n28002), .I0(n510), .I1(GND_net), .CO(n28003));
    SB_LUT4 add_1872_5_lut (.I0(GND_net), .I1(n511), .I2(VCC_net), .I3(n28001), 
            .O(n6026)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1872_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1872_5 (.CI(n28001), .I0(n511), .I1(VCC_net), .CO(n28002));
    SB_LUT4 add_1872_4_lut (.I0(GND_net), .I1(n425), .I2(GND_net), .I3(n28000), 
            .O(n6027)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1872_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1872_4 (.CI(n28000), .I0(n425), .I1(GND_net), .CO(n28001));
    SB_LUT4 add_1872_3_lut (.I0(GND_net), .I1(n513), .I2(VCC_net), .I3(n27999), 
            .O(n6028)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1872_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1872_3 (.CI(n27999), .I0(n513), .I1(VCC_net), .CO(n28000));
    SB_LUT4 add_1872_2_lut (.I0(GND_net), .I1(n598_adj_4967), .I2(GND_net), 
            .I3(VCC_net), .O(n6029)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1872_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder1_position_23__I_0_inv_0_i9_1_lut (.I0(encoder0_position_scaled[8]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n17_adj_4957));   // verilog/TinyFPGA_B.v(202[21:65])
    defparam encoder1_position_23__I_0_inv_0_i9_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_1872_2 (.CI(VCC_net), .I0(n598_adj_4967), .I1(GND_net), 
            .CO(n27999));
    SB_LUT4 unary_minus_4_inv_0_i20_1_lut (.I0(duty[19]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_4885));   // verilog/TinyFPGA_B.v(106[23:28])
    defparam unary_minus_4_inv_0_i20_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mux_77_i1_4_lut (.I0(encoder1_position[0]), .I1(displacement[0]), 
            .I2(n15_adj_4934), .I3(n15_adj_4940), .O(motor_state_23__N_82[0]));   // verilog/TinyFPGA_B.v(166[5] 168[10])
    defparam mux_77_i1_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i14080_3_lut (.I0(\data_in_frame[5] [7]), .I1(rx_data[7]), .I2(n32660), 
            .I3(GND_net), .O(n19222));   // verilog/coms.v(127[12] 300[6])
    defparam i14080_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14081_3_lut (.I0(\data_in_frame[5] [6]), .I1(rx_data[6]), .I2(n32660), 
            .I3(GND_net), .O(n19223));   // verilog/coms.v(127[12] 300[6])
    defparam i14081_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14082_3_lut (.I0(\data_in_frame[5] [5]), .I1(rx_data[5]), .I2(n32660), 
            .I3(GND_net), .O(n19224));   // verilog/coms.v(127[12] 300[6])
    defparam i14082_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14083_3_lut (.I0(\data_in_frame[5] [4]), .I1(rx_data[4]), .I2(n32660), 
            .I3(GND_net), .O(n19225));   // verilog/coms.v(127[12] 300[6])
    defparam i14083_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14084_3_lut (.I0(\data_in_frame[5] [3]), .I1(rx_data[3]), .I2(n32660), 
            .I3(GND_net), .O(n19226));   // verilog/coms.v(127[12] 300[6])
    defparam i14084_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14085_3_lut (.I0(\data_in_frame[5] [2]), .I1(rx_data[2]), .I2(n32660), 
            .I3(GND_net), .O(n19227));   // verilog/coms.v(127[12] 300[6])
    defparam i14085_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14086_3_lut (.I0(\data_in_frame[5] [1]), .I1(rx_data[1]), .I2(n32660), 
            .I3(GND_net), .O(n19228));   // verilog/coms.v(127[12] 300[6])
    defparam i14086_3_lut.LUT_INIT = 16'hacac;
    SB_DFFESR delay_counter_i0_i0 (.Q(delay_counter[0]), .C(CLK_c), .E(n5410), 
            .D(n604), .R(n18963));   // verilog/TinyFPGA_B.v(237[10] 265[6])
    SB_LUT4 i14087_3_lut (.I0(\data_in_frame[5] [0]), .I1(rx_data[0]), .I2(n32660), 
            .I3(GND_net), .O(n19229));   // verilog/coms.v(127[12] 300[6])
    defparam i14087_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder1_position_23__I_0_inv_0_i10_1_lut (.I0(encoder0_position_scaled[9]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n16_adj_4956));   // verilog/TinyFPGA_B.v(202[21:65])
    defparam encoder1_position_23__I_0_inv_0_i10_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_4_inv_0_i21_1_lut (.I0(duty[20]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n5));   // verilog/TinyFPGA_B.v(106[23:28])
    defparam unary_minus_4_inv_0_i21_1_lut.LUT_INIT = 16'h5555;
    SB_IO ENCODER1_B_pad (.PACKAGE_PIN(ENCODER1_B), .OUTPUT_ENABLE(VCC_net), 
          .D_IN_0(ENCODER1_B_c_0)) /* synthesis IO_FF_IN=TRUE */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam ENCODER1_B_pad.PIN_TYPE = 6'b000001;
    defparam ENCODER1_B_pad.PULLUP = 1'b0;
    defparam ENCODER1_B_pad.NEG_TRIGGER = 1'b0;
    defparam ENCODER1_B_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO ENCODER1_A_pad (.PACKAGE_PIN(ENCODER1_A), .OUTPUT_ENABLE(VCC_net), 
          .D_IN_0(ENCODER1_A_c_1)) /* synthesis IO_FF_IN=TRUE */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam ENCODER1_A_pad.PIN_TYPE = 6'b000001;
    defparam ENCODER1_A_pad.PULLUP = 1'b0;
    defparam ENCODER1_A_pad.NEG_TRIGGER = 1'b0;
    defparam ENCODER1_A_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO ENCODER0_B_pad (.PACKAGE_PIN(ENCODER0_B), .OUTPUT_ENABLE(VCC_net), 
          .D_IN_0(ENCODER0_B_c_0)) /* synthesis IO_FF_IN=TRUE */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam ENCODER0_B_pad.PIN_TYPE = 6'b000001;
    defparam ENCODER0_B_pad.PULLUP = 1'b0;
    defparam ENCODER0_B_pad.NEG_TRIGGER = 1'b0;
    defparam ENCODER0_B_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO ENCODER0_A_pad (.PACKAGE_PIN(ENCODER0_A), .OUTPUT_ENABLE(VCC_net), 
          .D_IN_0(ENCODER0_A_c_1)) /* synthesis IO_FF_IN=TRUE */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam ENCODER0_A_pad.PIN_TYPE = 6'b000001;
    defparam ENCODER0_A_pad.PULLUP = 1'b0;
    defparam ENCODER0_A_pad.NEG_TRIGGER = 1'b0;
    defparam ENCODER0_A_pad.IO_STANDARD = "SB_LVCMOS";
    SB_GB_IO CLK_pad (.PACKAGE_PIN(CLK), .OUTPUT_ENABLE(VCC_net), .GLOBAL_BUFFER_OUTPUT(CLK_c));   // verilog/TinyFPGA_B.v(3[9:12])
    defparam CLK_pad.PIN_TYPE = 6'b000001;
    defparam CLK_pad.PULLUP = 1'b0;
    defparam CLK_pad.NEG_TRIGGER = 1'b0;
    defparam CLK_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO INHA_pad (.PACKAGE_PIN(INHA), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(INHA_c));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam INHA_pad.PIN_TYPE = 6'b011001;
    defparam INHA_pad.PULLUP = 1'b0;
    defparam INHA_pad.NEG_TRIGGER = 1'b0;
    defparam INHA_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO INLA_pad (.PACKAGE_PIN(INLA), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(INLA_c));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam INLA_pad.PIN_TYPE = 6'b011001;
    defparam INLA_pad.PULLUP = 1'b0;
    defparam INLA_pad.NEG_TRIGGER = 1'b0;
    defparam INLA_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO INHB_pad (.PACKAGE_PIN(INHB), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(INHB_c));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam INHB_pad.PIN_TYPE = 6'b011001;
    defparam INHB_pad.PULLUP = 1'b0;
    defparam INHB_pad.NEG_TRIGGER = 1'b0;
    defparam INHB_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO INLB_pad (.PACKAGE_PIN(INLB), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(INLB_c));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam INLB_pad.PIN_TYPE = 6'b011001;
    defparam INLB_pad.PULLUP = 1'b0;
    defparam INLB_pad.NEG_TRIGGER = 1'b0;
    defparam INLB_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO INHC_pad (.PACKAGE_PIN(INHC), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(INHC_c)) /* synthesis IO_FF_OUT=TRUE */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam INHC_pad.PIN_TYPE = 6'b011001;
    defparam INHC_pad.PULLUP = 1'b0;
    defparam INHC_pad.NEG_TRIGGER = 1'b0;
    defparam INHC_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO CS_CLK_pad (.PACKAGE_PIN(CS_CLK), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(GND_net));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam CS_CLK_pad.PIN_TYPE = 6'b011001;
    defparam CS_CLK_pad.PULLUP = 1'b0;
    defparam CS_CLK_pad.NEG_TRIGGER = 1'b0;
    defparam CS_CLK_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO DE_pad (.PACKAGE_PIN(DE), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(DE_c));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DE_pad.PIN_TYPE = 6'b011001;
    defparam DE_pad.PULLUP = 1'b0;
    defparam DE_pad.NEG_TRIGGER = 1'b0;
    defparam DE_pad.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 add_25_4_lut (.I0(GND_net), .I1(delay_counter[2]), .I2(GND_net), 
            .I3(n27734), .O(n602)) /* synthesis syn_instantiated=1 */ ;
    defparam add_25_4_lut.LUT_INIT = 16'hC33C;
    SB_DFF displacement_i23 (.Q(displacement[23]), .C(clk32MHz), .D(displacement_23__N_58[23]));   // verilog/TinyFPGA_B.v(200[10] 203[6])
    SB_LUT4 i2_2_lut (.I0(pwm_counter[27]), .I1(pwm_counter[28]), .I2(GND_net), 
            .I3(GND_net), .O(n10_adj_5060));
    defparam i2_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i6_4_lut_adj_1636 (.I0(pwm_counter[23]), .I1(pwm_counter[29]), 
            .I2(pwm_counter[25]), .I3(pwm_counter[26]), .O(n14_adj_5059));
    defparam i6_4_lut_adj_1636.LUT_INIT = 16'hfffe;
    SB_LUT4 i7_4_lut_adj_1637 (.I0(pwm_counter[30]), .I1(n14_adj_5059), 
            .I2(n10_adj_5060), .I3(pwm_counter[24]), .O(n17360));
    defparam i7_4_lut_adj_1637.LUT_INIT = 16'hfffe;
    SB_LUT4 encoder0_position_23__I_0_i1322_3_lut (.I0(n1934), .I1(n1987), 
            .I2(n1948), .I3(GND_net), .O(n2012));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1322_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1315_3_lut (.I0(n1927), .I1(n1980), 
            .I2(n1948), .I3(GND_net), .O(n2005));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1315_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1327_3_lut (.I0(n1939), .I1(n1992), 
            .I2(n1948), .I3(GND_net), .O(n2017));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1327_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1324_3_lut (.I0(n1936), .I1(n1989), 
            .I2(n1948), .I3(GND_net), .O(n2014));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1324_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1325_3_lut (.I0(n1937), .I1(n1990), 
            .I2(n1948), .I3(GND_net), .O(n2015));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1325_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1313_3_lut (.I0(n1925), .I1(n1978), 
            .I2(n1948), .I3(GND_net), .O(n2003));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1313_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1332_3_lut (.I0(n774), .I1(n1997), 
            .I2(n1948), .I3(GND_net), .O(n2022));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1332_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1331_3_lut (.I0(n1943), .I1(n1996), 
            .I2(n1948), .I3(GND_net), .O(n2021));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1331_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mux_3363_i1_3_lut (.I0(encoder0_position[0]), .I1(n25_adj_4902), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n775));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam mux_3363_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_23__I_0_i1317_3_lut (.I0(n1929), .I1(n1982), 
            .I2(n1948), .I3(GND_net), .O(n2007));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1317_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1323_3_lut (.I0(n1935), .I1(n1988), 
            .I2(n1948), .I3(GND_net), .O(n2013));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1323_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1314_3_lut (.I0(n1926), .I1(n1979), 
            .I2(n1948), .I3(GND_net), .O(n2004));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1314_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1319_3_lut (.I0(n1931), .I1(n1984), 
            .I2(n1948), .I3(GND_net), .O(n2009));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1319_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1316_3_lut (.I0(n1928), .I1(n1981), 
            .I2(n1948), .I3(GND_net), .O(n2006));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1316_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1320_3_lut (.I0(n1932), .I1(n1985), 
            .I2(n1948), .I3(GND_net), .O(n2010));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1320_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder1_position_23__I_0_add_2_25_lut (.I0(GND_net), .I1(encoder1_position[23]), 
            .I2(n3_adj_4944), .I3(n28096), .O(displacement_23__N_58[23])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder1_position_23__I_0_add_2_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_23__I_0_i1326_3_lut (.I0(n1938), .I1(n1991), 
            .I2(n1948), .I3(GND_net), .O(n2016));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1326_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder1_position_23__I_0_add_2_24_lut (.I0(GND_net), .I1(encoder1_position[22]), 
            .I2(n3_adj_4944), .I3(n28095), .O(displacement_23__N_58[22])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder1_position_23__I_0_add_2_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder1_position_23__I_0_add_2_24 (.CI(n28095), .I0(encoder1_position[22]), 
            .I1(n3_adj_4944), .CO(n28096));
    SB_LUT4 encoder1_position_23__I_0_add_2_23_lut (.I0(GND_net), .I1(encoder1_position[21]), 
            .I2(n3_adj_4944), .I3(n28094), .O(displacement_23__N_58[21])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder1_position_23__I_0_add_2_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_23__I_0_i1310_3_lut (.I0(n1922), .I1(n1975), 
            .I2(n1948), .I3(GND_net), .O(n2000));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1310_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1330_3_lut (.I0(n1942), .I1(n1995), 
            .I2(n1948), .I3(GND_net), .O(n2020));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1330_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1328_3_lut (.I0(n1940), .I1(n1993), 
            .I2(n1948), .I3(GND_net), .O(n2018));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1328_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder1_position_23__I_0_add_2_23 (.CI(n28094), .I0(encoder1_position[21]), 
            .I1(n3_adj_4944), .CO(n28095));
    SB_LUT4 encoder0_position_23__I_0_i1329_3_lut (.I0(n1941), .I1(n1994), 
            .I2(n1948), .I3(GND_net), .O(n2019));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1329_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1311_3_lut (.I0(n1923), .I1(n1976), 
            .I2(n1948), .I3(GND_net), .O(n2001));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1311_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1318_3_lut (.I0(n1930), .I1(n1983), 
            .I2(n1948), .I3(GND_net), .O(n2008));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1318_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1321_3_lut (.I0(n1933), .I1(n1986), 
            .I2(n1948), .I3(GND_net), .O(n2011));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1321_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1312_3_lut (.I0(n1924), .I1(n1977), 
            .I2(n1948), .I3(GND_net), .O(n2002));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1312_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i11_4_lut (.I0(n2002), .I1(n2011), .I2(n2008), .I3(n2001), 
            .O(n30_adj_5035));
    defparam i11_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i19530_3_lut (.I0(n775), .I1(n2021), .I2(n2022), .I3(GND_net), 
            .O(n24673));
    defparam i19530_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i2_4_lut_adj_1638 (.I0(n2019), .I1(n2018), .I2(n24673), .I3(n2020), 
            .O(n35117));
    defparam i2_4_lut_adj_1638.LUT_INIT = 16'h8880;
    SB_LUT4 i15_4_lut (.I0(n2003), .I1(n30_adj_5035), .I2(n2015), .I3(n2014), 
            .O(n34_adj_5032));
    defparam i15_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i13_4_lut (.I0(n2000), .I1(n2016), .I2(n2010), .I3(n2006), 
            .O(n32));
    defparam i13_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i14_4_lut (.I0(n2009), .I1(n2004), .I2(n2013), .I3(n2007), 
            .O(n33_adj_5033));
    defparam i14_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i12_4_lut (.I0(n2017), .I1(n2005), .I2(n2012), .I3(n35117), 
            .O(n31_adj_5034));
    defparam i12_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i30830_4_lut (.I0(n31_adj_5034), .I1(n33_adj_5033), .I2(n32), 
            .I3(n34_adj_5032), .O(n2026));
    defparam i30830_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 encoder0_position_23__I_0_i1494_3_lut (.I0(n2026), .I1(n6222), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(encoder0_position_scaled_23__N_34[1]));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1494_3_lut.LUT_INIT = 16'hc5c5;
    SB_LUT4 encoder0_position_23__I_0_i1274_3_lut (.I0(n1861), .I1(n1914), 
            .I2(n1870), .I3(GND_net), .O(n1939));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1274_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1269_3_lut (.I0(n1856), .I1(n1909), 
            .I2(n1870), .I3(GND_net), .O(n1934));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1269_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1275_3_lut (.I0(n1862), .I1(n1915), 
            .I2(n1870), .I3(GND_net), .O(n1940));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1275_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder1_position_23__I_0_add_2_22_lut (.I0(GND_net), .I1(encoder1_position[20]), 
            .I2(n5_adj_4945), .I3(n28093), .O(displacement_23__N_58[20])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder1_position_23__I_0_add_2_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder1_position_23__I_0_add_2_22 (.CI(n28093), .I0(encoder1_position[20]), 
            .I1(n5_adj_4945), .CO(n28094));
    SB_LUT4 encoder1_position_23__I_0_add_2_21_lut (.I0(GND_net), .I1(encoder1_position[19]), 
            .I2(n6_adj_4946), .I3(n28092), .O(displacement_23__N_58[19])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder1_position_23__I_0_add_2_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder1_position_23__I_0_add_2_21 (.CI(n28092), .I0(encoder1_position[19]), 
            .I1(n6_adj_4946), .CO(n28093));
    SB_LUT4 encoder1_position_23__I_0_add_2_20_lut (.I0(GND_net), .I1(encoder1_position[18]), 
            .I2(n7_adj_4947), .I3(n28091), .O(displacement_23__N_58[18])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder1_position_23__I_0_add_2_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_23__I_0_i1278_3_lut (.I0(n773), .I1(n1918), 
            .I2(n1870), .I3(GND_net), .O(n1943));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1278_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder1_position_23__I_0_add_2_20 (.CI(n28091), .I0(encoder1_position[18]), 
            .I1(n7_adj_4947), .CO(n28092));
    SB_LUT4 encoder0_position_23__I_0_i1277_3_lut (.I0(n1864), .I1(n1917), 
            .I2(n1870), .I3(GND_net), .O(n1942));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1277_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1276_3_lut (.I0(n1863), .I1(n1916), 
            .I2(n1870), .I3(GND_net), .O(n1941));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1276_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mux_3363_i2_3_lut (.I0(encoder0_position[1]), .I1(n24_adj_4903), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n774));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam mux_3363_i2_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_23__I_0_i1259_3_lut (.I0(n1846), .I1(n1899), 
            .I2(n1870), .I3(GND_net), .O(n1924));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1259_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1264_3_lut (.I0(n1851), .I1(n1904), 
            .I2(n1870), .I3(GND_net), .O(n1929));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1264_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1268_3_lut (.I0(n1855), .I1(n1908), 
            .I2(n1870), .I3(GND_net), .O(n1933));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1268_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1261_3_lut (.I0(n1848), .I1(n1901), 
            .I2(n1870), .I3(GND_net), .O(n1926));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1261_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1258_3_lut (.I0(n1845), .I1(n1898), 
            .I2(n1870), .I3(GND_net), .O(n1923));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1258_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1262_3_lut (.I0(n1849), .I1(n1902), 
            .I2(n1870), .I3(GND_net), .O(n1927));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1262_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1271_3_lut (.I0(n1858), .I1(n1911), 
            .I2(n1870), .I3(GND_net), .O(n1936));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1271_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY add_25_11 (.CI(n27741), .I0(delay_counter[9]), .I1(GND_net), 
            .CO(n27742));
    SB_LUT4 encoder0_position_23__I_0_i1257_3_lut (.I0(n1844), .I1(n1897), 
            .I2(n1870), .I3(GND_net), .O(n1922));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1257_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1265_3_lut (.I0(n1852), .I1(n1905), 
            .I2(n1870), .I3(GND_net), .O(n1930));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1265_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1266_3_lut (.I0(n1853), .I1(n1906), 
            .I2(n1870), .I3(GND_net), .O(n1931));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1266_3_lut.LUT_INIT = 16'hacac;
    SB_DFF displacement_i22 (.Q(displacement[22]), .C(clk32MHz), .D(displacement_23__N_58[22]));   // verilog/TinyFPGA_B.v(200[10] 203[6])
    SB_LUT4 encoder0_position_23__I_0_i1270_3_lut (.I0(n1857), .I1(n1910), 
            .I2(n1870), .I3(GND_net), .O(n1935));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1270_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1263_3_lut (.I0(n1850), .I1(n1903), 
            .I2(n1870), .I3(GND_net), .O(n1928));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1263_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1267_3_lut (.I0(n1854), .I1(n1907), 
            .I2(n1870), .I3(GND_net), .O(n1932));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1267_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1272_3_lut (.I0(n1859), .I1(n1912), 
            .I2(n1870), .I3(GND_net), .O(n1937));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1272_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1273_3_lut (.I0(n1860), .I1(n1913), 
            .I2(n1870), .I3(GND_net), .O(n1938));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1273_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1260_3_lut (.I0(n1847), .I1(n1900), 
            .I2(n1870), .I3(GND_net), .O(n1925));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1260_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i10_4_lut_adj_1639 (.I0(n1925), .I1(n1938), .I2(n1937), .I3(n1932), 
            .O(n28_adj_5003));
    defparam i10_4_lut_adj_1639.LUT_INIT = 16'hfffe;
    SB_LUT4 i13_4_lut_adj_1640 (.I0(n1926), .I1(n1933), .I2(n1929), .I3(n1924), 
            .O(n31_adj_5001));
    defparam i13_4_lut_adj_1640.LUT_INIT = 16'hfffe;
    SB_LUT4 i19653_4_lut (.I0(n774), .I1(n1941), .I2(n1942), .I3(n1943), 
            .O(n24797));
    defparam i19653_4_lut.LUT_INIT = 16'hfcec;
    SB_LUT4 i4_2_lut (.I0(n1928), .I1(n1935), .I2(GND_net), .I3(GND_net), 
            .O(n22_adj_5028));
    defparam i4_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i12_4_lut_adj_1641 (.I0(n1931), .I1(n1930), .I2(n1922), .I3(n1936), 
            .O(n30_adj_5002));
    defparam i12_4_lut_adj_1641.LUT_INIT = 16'hfffe;
    SB_LUT4 i16_4_lut_adj_1642 (.I0(n31_adj_5001), .I1(n1927), .I2(n28_adj_5003), 
            .I3(n1923), .O(n34));
    defparam i16_4_lut_adj_1642.LUT_INIT = 16'hfffe;
    SB_LUT4 i3_4_lut_adj_1643 (.I0(n1940), .I1(n1934), .I2(n1939), .I3(n24797), 
            .O(n21_adj_5029));
    defparam i3_4_lut_adj_1643.LUT_INIT = 16'heccc;
    SB_DFF displacement_i21 (.Q(displacement[21]), .C(clk32MHz), .D(displacement_23__N_58[21]));   // verilog/TinyFPGA_B.v(200[10] 203[6])
    SB_DFF displacement_i20 (.Q(displacement[20]), .C(clk32MHz), .D(displacement_23__N_58[20]));   // verilog/TinyFPGA_B.v(200[10] 203[6])
    SB_DFF displacement_i19 (.Q(displacement[19]), .C(clk32MHz), .D(displacement_23__N_58[19]));   // verilog/TinyFPGA_B.v(200[10] 203[6])
    SB_DFF displacement_i18 (.Q(displacement[18]), .C(clk32MHz), .D(displacement_23__N_58[18]));   // verilog/TinyFPGA_B.v(200[10] 203[6])
    SB_DFF displacement_i17 (.Q(displacement[17]), .C(clk32MHz), .D(displacement_23__N_58[17]));   // verilog/TinyFPGA_B.v(200[10] 203[6])
    SB_DFF displacement_i16 (.Q(displacement[16]), .C(clk32MHz), .D(displacement_23__N_58[16]));   // verilog/TinyFPGA_B.v(200[10] 203[6])
    SB_DFF displacement_i15 (.Q(displacement[15]), .C(clk32MHz), .D(displacement_23__N_58[15]));   // verilog/TinyFPGA_B.v(200[10] 203[6])
    SB_DFF displacement_i14 (.Q(displacement[14]), .C(clk32MHz), .D(displacement_23__N_58[14]));   // verilog/TinyFPGA_B.v(200[10] 203[6])
    SB_DFF displacement_i13 (.Q(displacement[13]), .C(clk32MHz), .D(displacement_23__N_58[13]));   // verilog/TinyFPGA_B.v(200[10] 203[6])
    SB_DFF displacement_i12 (.Q(displacement[12]), .C(clk32MHz), .D(displacement_23__N_58[12]));   // verilog/TinyFPGA_B.v(200[10] 203[6])
    SB_DFF displacement_i11 (.Q(displacement[11]), .C(clk32MHz), .D(displacement_23__N_58[11]));   // verilog/TinyFPGA_B.v(200[10] 203[6])
    SB_DFF displacement_i10 (.Q(displacement[10]), .C(clk32MHz), .D(displacement_23__N_58[10]));   // verilog/TinyFPGA_B.v(200[10] 203[6])
    SB_DFF displacement_i9 (.Q(displacement[9]), .C(clk32MHz), .D(displacement_23__N_58[9]));   // verilog/TinyFPGA_B.v(200[10] 203[6])
    SB_DFF displacement_i8 (.Q(displacement[8]), .C(clk32MHz), .D(displacement_23__N_58[8]));   // verilog/TinyFPGA_B.v(200[10] 203[6])
    SB_DFF displacement_i7 (.Q(displacement[7]), .C(clk32MHz), .D(displacement_23__N_58[7]));   // verilog/TinyFPGA_B.v(200[10] 203[6])
    SB_DFF displacement_i6 (.Q(displacement[6]), .C(clk32MHz), .D(displacement_23__N_58[6]));   // verilog/TinyFPGA_B.v(200[10] 203[6])
    SB_DFF displacement_i5 (.Q(displacement[5]), .C(clk32MHz), .D(displacement_23__N_58[5]));   // verilog/TinyFPGA_B.v(200[10] 203[6])
    SB_DFF displacement_i4 (.Q(displacement[4]), .C(clk32MHz), .D(displacement_23__N_58[4]));   // verilog/TinyFPGA_B.v(200[10] 203[6])
    SB_DFF displacement_i3 (.Q(displacement[3]), .C(clk32MHz), .D(displacement_23__N_58[3]));   // verilog/TinyFPGA_B.v(200[10] 203[6])
    SB_DFF displacement_i2 (.Q(displacement[2]), .C(clk32MHz), .D(displacement_23__N_58[2]));   // verilog/TinyFPGA_B.v(200[10] 203[6])
    SB_DFF displacement_i1 (.Q(displacement[1]), .C(clk32MHz), .D(displacement_23__N_58[1]));   // verilog/TinyFPGA_B.v(200[10] 203[6])
    SB_LUT4 i30805_4_lut (.I0(n21_adj_5029), .I1(n34), .I2(n30_adj_5002), 
            .I3(n22_adj_5028), .O(n1948));
    defparam i30805_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 encoder0_position_23__I_0_i1493_3_lut (.I0(n1948), .I1(n6221), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(encoder0_position_scaled_23__N_34[2]));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1493_3_lut.LUT_INIT = 16'hc5c5;
    SB_LUT4 encoder0_position_23__I_0_i1207_3_lut (.I0(n1769), .I1(n1822), 
            .I2(n1792), .I3(GND_net), .O(n1847));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1207_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1205_3_lut (.I0(n1767), .I1(n1820), 
            .I2(n1792), .I3(GND_net), .O(n1845));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1205_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1204_3_lut (.I0(n1766), .I1(n1819), 
            .I2(n1792), .I3(GND_net), .O(n1844));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1204_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1215_3_lut (.I0(n1777), .I1(n1830), 
            .I2(n1792), .I3(GND_net), .O(n1855));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1215_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1216_3_lut (.I0(n1778), .I1(n1831), 
            .I2(n1792), .I3(GND_net), .O(n1856));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1216_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1206_3_lut (.I0(n1768), .I1(n1821), 
            .I2(n1792), .I3(GND_net), .O(n1846));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1206_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1210_3_lut (.I0(n1772), .I1(n1825), 
            .I2(n1792), .I3(GND_net), .O(n1850));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1210_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1224_3_lut (.I0(n772), .I1(n1839), 
            .I2(n1792), .I3(GND_net), .O(n1864));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1224_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1223_3_lut (.I0(n1785), .I1(n1838), 
            .I2(n1792), .I3(GND_net), .O(n1863));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1223_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mux_3363_i3_3_lut (.I0(encoder0_position[2]), .I1(n23_adj_4904), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n773));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam mux_3363_i3_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_23__I_0_i1219_3_lut (.I0(n1781), .I1(n1834), 
            .I2(n1792), .I3(GND_net), .O(n1859));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1219_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1217_3_lut (.I0(n1779), .I1(n1832), 
            .I2(n1792), .I3(GND_net), .O(n1857));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1217_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1218_3_lut (.I0(n1780), .I1(n1833), 
            .I2(n1792), .I3(GND_net), .O(n1858));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1218_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1214_3_lut (.I0(n1776), .I1(n1829), 
            .I2(n1792), .I3(GND_net), .O(n1854));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1214_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1209_3_lut (.I0(n1771), .I1(n1824), 
            .I2(n1792), .I3(GND_net), .O(n1849));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1209_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1213_3_lut (.I0(n1775), .I1(n1828), 
            .I2(n1792), .I3(GND_net), .O(n1853));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1213_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1212_3_lut (.I0(n1774), .I1(n1827), 
            .I2(n1792), .I3(GND_net), .O(n1852));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1212_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1222_3_lut (.I0(n1784), .I1(n1837), 
            .I2(n1792), .I3(GND_net), .O(n1862));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1222_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1220_3_lut (.I0(n1782), .I1(n1835), 
            .I2(n1792), .I3(GND_net), .O(n1860));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1220_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1221_3_lut (.I0(n1783), .I1(n1836), 
            .I2(n1792), .I3(GND_net), .O(n1861));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1221_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1208_3_lut (.I0(n1770), .I1(n1823), 
            .I2(n1792), .I3(GND_net), .O(n1848));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1208_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1211_3_lut (.I0(n1773), .I1(n1826), 
            .I2(n1792), .I3(GND_net), .O(n1851));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1211_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut (.I0(n1851), .I1(n1848), .I2(GND_net), .I3(GND_net), 
            .O(n18_adj_4899));
    defparam i1_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i19540_3_lut (.I0(n773), .I1(n1863), .I2(n1864), .I3(GND_net), 
            .O(n24683));
    defparam i19540_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i2_4_lut_adj_1644 (.I0(n1861), .I1(n1860), .I2(n24683), .I3(n1862), 
            .O(n34029));
    defparam i2_4_lut_adj_1644.LUT_INIT = 16'h8880;
    SB_LUT4 i13_4_lut_adj_1645 (.I0(n1850), .I1(n1846), .I2(n1856), .I3(n18_adj_4899), 
            .O(n30));
    defparam i13_4_lut_adj_1645.LUT_INIT = 16'hfffe;
    SB_LUT4 i14127_3_lut (.I0(neopxl_color[23]), .I1(\data_in_frame[4] [7]), 
            .I2(n3_adj_4943), .I3(GND_net), .O(n19269));   // verilog/coms.v(127[12] 300[6])
    defparam i14127_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14128_3_lut (.I0(neopxl_color[22]), .I1(\data_in_frame[4] [6]), 
            .I2(n3_adj_4943), .I3(GND_net), .O(n19270));   // verilog/coms.v(127[12] 300[6])
    defparam i14128_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i11_4_lut_adj_1646 (.I0(n1852), .I1(n1853), .I2(n1849), .I3(n1854), 
            .O(n28));
    defparam i11_4_lut_adj_1646.LUT_INIT = 16'hfffe;
    SB_LUT4 i30579_4_lut (.I0(n752), .I1(n755), .I2(n753), .I3(n4_adj_4925), 
            .O(n778));
    defparam i30579_4_lut.LUT_INIT = 16'h0105;
    SB_LUT4 encoder1_position_23__I_0_add_2_19_lut (.I0(GND_net), .I1(encoder1_position[17]), 
            .I2(n8_adj_4948), .I3(n28090), .O(displacement_23__N_58[17])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder1_position_23__I_0_add_2_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i12_4_lut_adj_1647 (.I0(n1858), .I1(n34029), .I2(n1857), .I3(n1859), 
            .O(n29));
    defparam i12_4_lut_adj_1647.LUT_INIT = 16'hfffe;
    SB_LUT4 i10_4_lut_adj_1648 (.I0(n1855), .I1(n1844), .I2(n1845), .I3(n1847), 
            .O(n27));
    defparam i10_4_lut_adj_1648.LUT_INIT = 16'hfffe;
    SB_LUT4 i30778_4_lut (.I0(n27), .I1(n29), .I2(n28), .I3(n30), .O(n1870));
    defparam i30778_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 encoder0_position_23__I_0_i1492_3_lut (.I0(n1870), .I1(n6220), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(encoder0_position_scaled_23__N_34[3]));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1492_3_lut.LUT_INIT = 16'hc5c5;
    SB_CARRY encoder1_position_23__I_0_add_2_19 (.CI(n28090), .I0(encoder1_position[17]), 
            .I1(n8_adj_4948), .CO(n28091));
    SB_LUT4 i14129_3_lut (.I0(neopxl_color[21]), .I1(\data_in_frame[4] [5]), 
            .I2(n3_adj_4943), .I3(GND_net), .O(n19271));   // verilog/coms.v(127[12] 300[6])
    defparam i14129_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i465_3_lut (.I0(n677), .I1(n730), 
            .I2(n700), .I3(GND_net), .O(n755));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i465_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1165_3_lut (.I0(n1702), .I1(n1755), 
            .I2(n1714), .I3(GND_net), .O(n1780));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1165_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1154_3_lut (.I0(n1691), .I1(n1744), 
            .I2(n1714), .I3(GND_net), .O(n1769));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1154_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1161_3_lut (.I0(n1698), .I1(n1751), 
            .I2(n1714), .I3(GND_net), .O(n1776));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1161_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1153_3_lut (.I0(n1690), .I1(n1743), 
            .I2(n1714), .I3(GND_net), .O(n1768));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1153_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder1_position_23__I_0_add_2_18_lut (.I0(GND_net), .I1(encoder1_position[16]), 
            .I2(n9_adj_4949), .I3(n28089), .O(displacement_23__N_58[16])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder1_position_23__I_0_add_2_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_23__I_0_i1159_3_lut (.I0(n1696), .I1(n1749), 
            .I2(n1714), .I3(GND_net), .O(n1774));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1159_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14130_3_lut (.I0(neopxl_color[20]), .I1(\data_in_frame[4] [4]), 
            .I2(n3_adj_4943), .I3(GND_net), .O(n19272));   // verilog/coms.v(127[12] 300[6])
    defparam i14130_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1162_3_lut (.I0(n1699), .I1(n1752), 
            .I2(n1714), .I3(GND_net), .O(n1777));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1162_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1163_3_lut (.I0(n1700), .I1(n1753), 
            .I2(n1714), .I3(GND_net), .O(n1778));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1163_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1170_3_lut (.I0(n771_adj_4968), .I1(n1760), 
            .I2(n1714), .I3(GND_net), .O(n1785));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1170_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14131_3_lut (.I0(neopxl_color[19]), .I1(\data_in_frame[4] [3]), 
            .I2(n3_adj_4943), .I3(GND_net), .O(n19273));   // verilog/coms.v(127[12] 300[6])
    defparam i14131_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1169_3_lut (.I0(n1706), .I1(n1759), 
            .I2(n1714), .I3(GND_net), .O(n1784));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1169_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i518_3_lut (.I0(n755), .I1(n808), 
            .I2(n778), .I3(GND_net), .O(n833));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i518_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mux_3363_i4_3_lut (.I0(encoder0_position[3]), .I1(n22_adj_4905), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n772));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam mux_3363_i4_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_23__I_0_i1156_3_lut (.I0(n1693), .I1(n1746), 
            .I2(n1714), .I3(GND_net), .O(n1771));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1156_3_lut.LUT_INIT = 16'hacac;
    SB_DFFSR encoder0_position_scaled_i22 (.Q(encoder0_position_scaled[22]), 
            .C(clk32MHz), .D(n6202), .R(n2_adj_5004));   // verilog/TinyFPGA_B.v(200[10] 203[6])
    SB_LUT4 encoder0_position_23__I_0_i1151_3_lut (.I0(n1688), .I1(n1741), 
            .I2(n1714), .I3(GND_net), .O(n1766));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1151_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1158_3_lut (.I0(n1695), .I1(n1748), 
            .I2(n1714), .I3(GND_net), .O(n1773));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1158_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1155_3_lut (.I0(n1692), .I1(n1745), 
            .I2(n1714), .I3(GND_net), .O(n1770));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1155_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1164_3_lut (.I0(n1701), .I1(n1754), 
            .I2(n1714), .I3(GND_net), .O(n1779));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1164_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1160_3_lut (.I0(n1697), .I1(n1750), 
            .I2(n1714), .I3(GND_net), .O(n1775));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1160_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1152_3_lut (.I0(n1689), .I1(n1742), 
            .I2(n1714), .I3(GND_net), .O(n1767));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1152_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14132_3_lut (.I0(neopxl_color[18]), .I1(\data_in_frame[4] [2]), 
            .I2(n3_adj_4943), .I3(GND_net), .O(n19274));   // verilog/coms.v(127[12] 300[6])
    defparam i14132_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1157_3_lut (.I0(n1694), .I1(n1747), 
            .I2(n1714), .I3(GND_net), .O(n1772));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1157_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_unary_minus_2_inv_0_i22_1_lut (.I0(encoder0_position[20]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n5_adj_5007));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_unary_minus_2_inv_0_i22_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_23__I_0_unary_minus_2_inv_0_i23_1_lut (.I0(encoder0_position[21]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n4_adj_5006));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_unary_minus_2_inv_0_i23_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_23__I_0_i1168_3_lut (.I0(n1705), .I1(n1758), 
            .I2(n1714), .I3(GND_net), .O(n1783));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1168_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1166_3_lut (.I0(n1703), .I1(n1756), 
            .I2(n1714), .I3(GND_net), .O(n1781));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1166_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1167_3_lut (.I0(n1704), .I1(n1757), 
            .I2(n1714), .I3(GND_net), .O(n1782));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1167_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14133_3_lut (.I0(neopxl_color[17]), .I1(\data_in_frame[4] [1]), 
            .I2(n3_adj_4943), .I3(GND_net), .O(n19275));   // verilog/coms.v(127[12] 300[6])
    defparam i14133_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i19542_3_lut (.I0(n772), .I1(n1784), .I2(n1785), .I3(GND_net), 
            .O(n24685));
    defparam i19542_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i14134_3_lut (.I0(neopxl_color[16]), .I1(\data_in_frame[4] [0]), 
            .I2(n3_adj_4943), .I3(GND_net), .O(n19276));   // verilog/coms.v(127[12] 300[6])
    defparam i14134_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i2_4_lut_adj_1649 (.I0(n1782), .I1(n1781), .I2(n24685), .I3(n1783), 
            .O(n34028));
    defparam i2_4_lut_adj_1649.LUT_INIT = 16'h8880;
    SB_LUT4 i14135_3_lut (.I0(neopxl_color[15]), .I1(\data_in_frame[5] [7]), 
            .I2(n3_adj_4943), .I3(GND_net), .O(n19277));   // verilog/coms.v(127[12] 300[6])
    defparam i14135_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12_4_lut_adj_1650 (.I0(n1772), .I1(n1767), .I2(n1775), .I3(n1779), 
            .O(n28_adj_5072));
    defparam i12_4_lut_adj_1650.LUT_INIT = 16'hfffe;
    SB_LUT4 i10_4_lut_adj_1651 (.I0(n1770), .I1(n1773), .I2(n1766), .I3(n1771), 
            .O(n26_adj_5074));
    defparam i10_4_lut_adj_1651.LUT_INIT = 16'hfffe;
    SB_LUT4 i11_4_lut_adj_1652 (.I0(n1778), .I1(n1777), .I2(n1774), .I3(n1768), 
            .O(n27_adj_5073));
    defparam i11_4_lut_adj_1652.LUT_INIT = 16'hfffe;
    SB_LUT4 i9_4_lut_adj_1653 (.I0(n34028), .I1(n1776), .I2(n1769), .I3(n1780), 
            .O(n25_adj_5075));
    defparam i9_4_lut_adj_1653.LUT_INIT = 16'hfffe;
    SB_LUT4 encoder0_position_23__I_0_unary_minus_2_inv_0_i17_1_lut (.I0(encoder0_position[15]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n10_adj_5012));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_unary_minus_2_inv_0_i17_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i14136_3_lut (.I0(neopxl_color[14]), .I1(\data_in_frame[5] [6]), 
            .I2(n3_adj_4943), .I3(GND_net), .O(n19278));   // verilog/coms.v(127[12] 300[6])
    defparam i14136_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14137_3_lut (.I0(neopxl_color[13]), .I1(\data_in_frame[5] [5]), 
            .I2(n3_adj_4943), .I3(GND_net), .O(n19279));   // verilog/coms.v(127[12] 300[6])
    defparam i14137_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i30752_4_lut (.I0(n25_adj_5075), .I1(n27_adj_5073), .I2(n26_adj_5074), 
            .I3(n28_adj_5072), .O(n1792));
    defparam i30752_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 encoder0_position_23__I_0_i1491_3_lut (.I0(n1792), .I1(n6219), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(encoder0_position_scaled_23__N_34[4]));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1491_3_lut.LUT_INIT = 16'hc5c5;
    SB_LUT4 encoder0_position_23__I_0_i1109_3_lut (.I0(n1621), .I1(n1674), 
            .I2(n1636), .I3(GND_net), .O(n1699));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1109_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1099_3_lut (.I0(n1611), .I1(n1664), 
            .I2(n1636), .I3(GND_net), .O(n1689));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1099_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1101_3_lut (.I0(n1613), .I1(n1666), 
            .I2(n1636), .I3(GND_net), .O(n1691));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1101_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i521_3_lut (.I0(n758), .I1(n811), 
            .I2(n778), .I3(GND_net), .O(n836));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i521_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY add_25_4 (.CI(n27734), .I0(delay_counter[2]), .I1(GND_net), 
            .CO(n27735));
    SB_LUT4 i14138_3_lut (.I0(neopxl_color[12]), .I1(\data_in_frame[5] [4]), 
            .I2(n3_adj_4943), .I3(GND_net), .O(n19280));   // verilog/coms.v(127[12] 300[6])
    defparam i14138_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_unary_minus_2_inv_0_i18_1_lut (.I0(encoder0_position[16]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n9_adj_5011));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_unary_minus_2_inv_0_i18_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_23__I_0_i1104_3_lut (.I0(n1616), .I1(n1669), 
            .I2(n1636), .I3(GND_net), .O(n1694));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1104_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1107_3_lut (.I0(n1619), .I1(n1672), 
            .I2(n1636), .I3(GND_net), .O(n1697));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1107_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1112_3_lut (.I0(n1624), .I1(n1677), 
            .I2(n1636), .I3(GND_net), .O(n1702));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1112_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i520_3_lut (.I0(n757), .I1(n810), 
            .I2(n778), .I3(GND_net), .O(n835));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i520_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14139_3_lut (.I0(neopxl_color[11]), .I1(\data_in_frame[5] [3]), 
            .I2(n3_adj_4943), .I3(GND_net), .O(n19281));   // verilog/coms.v(127[12] 300[6])
    defparam i14139_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i519_3_lut (.I0(n756), .I1(n809), 
            .I2(n778), .I3(GND_net), .O(n834));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i519_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder1_position_23__I_0_add_2_18 (.CI(n28089), .I0(encoder1_position[16]), 
            .I1(n9_adj_4949), .CO(n28090));
    SB_LUT4 encoder1_position_23__I_0_add_2_17_lut (.I0(GND_net), .I1(encoder1_position[15]), 
            .I2(n10_adj_4950), .I3(n28088), .O(displacement_23__N_58[15])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder1_position_23__I_0_add_2_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_25_10_lut (.I0(GND_net), .I1(delay_counter[8]), .I2(GND_net), 
            .I3(n27740), .O(n596)) /* synthesis syn_instantiated=1 */ ;
    defparam add_25_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i14140_3_lut (.I0(neopxl_color[10]), .I1(\data_in_frame[5] [2]), 
            .I2(n3_adj_4943), .I3(GND_net), .O(n19282));   // verilog/coms.v(127[12] 300[6])
    defparam i14140_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1113_3_lut (.I0(n1625), .I1(n1678), 
            .I2(n1636), .I3(GND_net), .O(n1703));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1113_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder1_position_23__I_0_add_2_17 (.CI(n28088), .I0(encoder1_position[15]), 
            .I1(n10_adj_4950), .CO(n28089));
    SB_LUT4 i14141_3_lut (.I0(neopxl_color[9]), .I1(\data_in_frame[5] [1]), 
            .I2(n3_adj_4943), .I3(GND_net), .O(n19283));   // verilog/coms.v(127[12] 300[6])
    defparam i14141_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder1_position_23__I_0_add_2_16_lut (.I0(GND_net), .I1(encoder1_position[14]), 
            .I2(n11_adj_4951), .I3(n28087), .O(displacement_23__N_58[14])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder1_position_23__I_0_add_2_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_23__I_0_i1110_3_lut (.I0(n1622), .I1(n1675), 
            .I2(n1636), .I3(GND_net), .O(n1700));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1110_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1116_3_lut (.I0(n770), .I1(n1681), 
            .I2(n1636), .I3(GND_net), .O(n1706));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1116_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14142_3_lut (.I0(neopxl_color[8]), .I1(\data_in_frame[5] [0]), 
            .I2(n3_adj_4943), .I3(GND_net), .O(n19284));   // verilog/coms.v(127[12] 300[6])
    defparam i14142_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder1_position_23__I_0_add_2_16 (.CI(n28087), .I0(encoder1_position[14]), 
            .I1(n11_adj_4951), .CO(n28088));
    SB_LUT4 add_672_24_lut (.I0(duty[22]), .I1(n37633), .I2(n3), .I3(n27847), 
            .O(pwm_setpoint_22__N_11[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_672_24_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 add_672_23_lut (.I0(duty[21]), .I1(n37633), .I2(n4_adj_4884), 
            .I3(n27846), .O(pwm_setpoint_22__N_11[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_672_23_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 encoder1_position_23__I_0_add_2_15_lut (.I0(GND_net), .I1(encoder1_position[13]), 
            .I2(n12_adj_4952), .I3(n28086), .O(displacement_23__N_58[13])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder1_position_23__I_0_add_2_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_25_10 (.CI(n27740), .I0(delay_counter[8]), .I1(GND_net), 
            .CO(n27741));
    SB_CARRY encoder1_position_23__I_0_add_2_15 (.CI(n28086), .I0(encoder1_position[13]), 
            .I1(n12_adj_4952), .CO(n28087));
    SB_LUT4 encoder1_position_23__I_0_add_2_14_lut (.I0(GND_net), .I1(encoder1_position[12]), 
            .I2(n13_adj_4953), .I3(n28085), .O(displacement_23__N_58[12])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder1_position_23__I_0_add_2_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder1_position_23__I_0_add_2_14 (.CI(n28085), .I0(encoder1_position[12]), 
            .I1(n13_adj_4953), .CO(n28086));
    SB_LUT4 add_25_33_lut (.I0(GND_net), .I1(delay_counter[31]), .I2(GND_net), 
            .I3(n27763), .O(n573)) /* synthesis syn_instantiated=1 */ ;
    defparam add_25_33_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_25_32_lut (.I0(GND_net), .I1(delay_counter[30]), .I2(GND_net), 
            .I3(n27762), .O(n574)) /* synthesis syn_instantiated=1 */ ;
    defparam add_25_32_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder1_position_23__I_0_add_2_13_lut (.I0(GND_net), .I1(encoder1_position[11]), 
            .I2(n14_adj_4954), .I3(n28084), .O(displacement_23__N_58[11])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder1_position_23__I_0_add_2_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder1_position_23__I_0_add_2_13 (.CI(n28084), .I0(encoder1_position[11]), 
            .I1(n14_adj_4954), .CO(n28085));
    SB_LUT4 encoder1_position_23__I_0_add_2_12_lut (.I0(GND_net), .I1(encoder1_position[10]), 
            .I2(n15_adj_4955), .I3(n28083), .O(displacement_23__N_58[10])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder1_position_23__I_0_add_2_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_23__I_0_unary_minus_2_inv_0_i19_1_lut (.I0(encoder0_position[17]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n8_adj_5010));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_unary_minus_2_inv_0_i19_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 RX_I_0_1_lut (.I0(RX_c), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(RX_N_10));   // verilog/TinyFPGA_B.v(143[10:13])
    defparam RX_I_0_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY encoder1_position_23__I_0_add_2_12 (.CI(n28083), .I0(encoder1_position[10]), 
            .I1(n15_adj_4955), .CO(n28084));
    SB_CARRY add_672_23 (.CI(n27846), .I0(n37633), .I1(n4_adj_4884), .CO(n27847));
    SB_LUT4 encoder0_position_23__I_0_i1115_3_lut (.I0(n1627), .I1(n1680), 
            .I2(n1636), .I3(GND_net), .O(n1705));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1115_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14143_3_lut (.I0(neopxl_color[7]), .I1(\data_in_frame[6] [7]), 
            .I2(n3_adj_4943), .I3(GND_net), .O(n19285));   // verilog/coms.v(127[12] 300[6])
    defparam i14143_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1114_3_lut (.I0(n1626), .I1(n1679), 
            .I2(n1636), .I3(GND_net), .O(n1704));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1114_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY add_25_32 (.CI(n27762), .I0(delay_counter[30]), .I1(GND_net), 
            .CO(n27763));
    SB_LUT4 encoder0_position_23__I_0_unary_minus_2_inv_0_i20_1_lut (.I0(encoder0_position[18]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n7_adj_5009));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_unary_minus_2_inv_0_i20_1_lut.LUT_INIT = 16'h5555;
    SB_DFFSR encoder0_position_scaled_i20 (.Q(encoder0_position_scaled[20]), 
            .C(clk32MHz), .D(n6203), .R(n2_adj_5004));   // verilog/TinyFPGA_B.v(200[10] 203[6])
    SB_LUT4 mux_3363_i5_3_lut (.I0(encoder0_position[4]), .I1(n21_adj_4906), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n771_adj_4968));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam mux_3363_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF encoder0_position_scaled_i19 (.Q(encoder0_position_scaled[19]), 
           .C(clk32MHz), .D(encoder0_position_scaled_23__N_34[19]));   // verilog/TinyFPGA_B.v(200[10] 203[6])
    SB_DFF encoder0_position_scaled_i18 (.Q(encoder0_position_scaled[18]), 
           .C(clk32MHz), .D(encoder0_position_scaled_23__N_34[18]));   // verilog/TinyFPGA_B.v(200[10] 203[6])
    SB_DFF encoder0_position_scaled_i17 (.Q(encoder0_position_scaled[17]), 
           .C(clk32MHz), .D(encoder0_position_scaled_23__N_34[17]));   // verilog/TinyFPGA_B.v(200[10] 203[6])
    SB_DFF encoder0_position_scaled_i16 (.Q(encoder0_position_scaled[16]), 
           .C(clk32MHz), .D(encoder0_position_scaled_23__N_34[16]));   // verilog/TinyFPGA_B.v(200[10] 203[6])
    SB_DFF encoder0_position_scaled_i15 (.Q(encoder0_position_scaled[15]), 
           .C(clk32MHz), .D(encoder0_position_scaled_23__N_34[15]));   // verilog/TinyFPGA_B.v(200[10] 203[6])
    SB_DFF encoder0_position_scaled_i14 (.Q(encoder0_position_scaled[14]), 
           .C(clk32MHz), .D(encoder0_position_scaled_23__N_34[14]));   // verilog/TinyFPGA_B.v(200[10] 203[6])
    SB_DFF encoder0_position_scaled_i13 (.Q(encoder0_position_scaled[13]), 
           .C(clk32MHz), .D(encoder0_position_scaled_23__N_34[13]));   // verilog/TinyFPGA_B.v(200[10] 203[6])
    SB_DFF encoder0_position_scaled_i12 (.Q(encoder0_position_scaled[12]), 
           .C(clk32MHz), .D(encoder0_position_scaled_23__N_34[12]));   // verilog/TinyFPGA_B.v(200[10] 203[6])
    SB_DFF encoder0_position_scaled_i11 (.Q(encoder0_position_scaled[11]), 
           .C(clk32MHz), .D(encoder0_position_scaled_23__N_34[11]));   // verilog/TinyFPGA_B.v(200[10] 203[6])
    SB_DFF encoder0_position_scaled_i10 (.Q(encoder0_position_scaled[10]), 
           .C(clk32MHz), .D(encoder0_position_scaled_23__N_34[10]));   // verilog/TinyFPGA_B.v(200[10] 203[6])
    SB_DFF encoder0_position_scaled_i9 (.Q(encoder0_position_scaled[9]), .C(clk32MHz), 
           .D(encoder0_position_scaled_23__N_34[9]));   // verilog/TinyFPGA_B.v(200[10] 203[6])
    SB_DFF encoder0_position_scaled_i8 (.Q(encoder0_position_scaled[8]), .C(clk32MHz), 
           .D(encoder0_position_scaled_23__N_34[8]));   // verilog/TinyFPGA_B.v(200[10] 203[6])
    SB_DFF encoder0_position_scaled_i7 (.Q(encoder0_position_scaled[7]), .C(clk32MHz), 
           .D(encoder0_position_scaled_23__N_34[7]));   // verilog/TinyFPGA_B.v(200[10] 203[6])
    SB_DFF encoder0_position_scaled_i6 (.Q(encoder0_position_scaled[6]), .C(clk32MHz), 
           .D(encoder0_position_scaled_23__N_34[6]));   // verilog/TinyFPGA_B.v(200[10] 203[6])
    SB_DFF encoder0_position_scaled_i5 (.Q(encoder0_position_scaled[5]), .C(clk32MHz), 
           .D(encoder0_position_scaled_23__N_34[5]));   // verilog/TinyFPGA_B.v(200[10] 203[6])
    SB_DFF encoder0_position_scaled_i4 (.Q(encoder0_position_scaled[4]), .C(clk32MHz), 
           .D(encoder0_position_scaled_23__N_34[4]));   // verilog/TinyFPGA_B.v(200[10] 203[6])
    SB_DFF encoder0_position_scaled_i3 (.Q(encoder0_position_scaled[3]), .C(clk32MHz), 
           .D(encoder0_position_scaled_23__N_34[3]));   // verilog/TinyFPGA_B.v(200[10] 203[6])
    SB_DFF encoder0_position_scaled_i2 (.Q(encoder0_position_scaled[2]), .C(clk32MHz), 
           .D(encoder0_position_scaled_23__N_34[2]));   // verilog/TinyFPGA_B.v(200[10] 203[6])
    SB_DFF encoder0_position_scaled_i1 (.Q(encoder0_position_scaled[1]), .C(clk32MHz), 
           .D(encoder0_position_scaled_23__N_34[1]));   // verilog/TinyFPGA_B.v(200[10] 203[6])
    SB_DFF pwm_setpoint_i22 (.Q(pwm_setpoint[22]), .C(clk32MHz), .D(pwm_setpoint_22__N_11[22]));   // verilog/TinyFPGA_B.v(96[10] 109[6])
    SB_DFF pwm_setpoint_i21 (.Q(pwm_setpoint[21]), .C(clk32MHz), .D(pwm_setpoint_22__N_11[21]));   // verilog/TinyFPGA_B.v(96[10] 109[6])
    SB_DFF pwm_setpoint_i20 (.Q(pwm_setpoint[20]), .C(clk32MHz), .D(pwm_setpoint_22__N_11[20]));   // verilog/TinyFPGA_B.v(96[10] 109[6])
    SB_DFF pwm_setpoint_i19 (.Q(pwm_setpoint[19]), .C(clk32MHz), .D(pwm_setpoint_22__N_11[19]));   // verilog/TinyFPGA_B.v(96[10] 109[6])
    SB_DFF pwm_setpoint_i18 (.Q(pwm_setpoint[18]), .C(clk32MHz), .D(pwm_setpoint_22__N_11[18]));   // verilog/TinyFPGA_B.v(96[10] 109[6])
    SB_DFF pwm_setpoint_i17 (.Q(pwm_setpoint[17]), .C(clk32MHz), .D(pwm_setpoint_22__N_11[17]));   // verilog/TinyFPGA_B.v(96[10] 109[6])
    SB_DFF pwm_setpoint_i16 (.Q(pwm_setpoint[16]), .C(clk32MHz), .D(pwm_setpoint_22__N_11[16]));   // verilog/TinyFPGA_B.v(96[10] 109[6])
    SB_DFF pwm_setpoint_i15 (.Q(pwm_setpoint[15]), .C(clk32MHz), .D(pwm_setpoint_22__N_11[15]));   // verilog/TinyFPGA_B.v(96[10] 109[6])
    SB_DFF pwm_setpoint_i14 (.Q(pwm_setpoint[14]), .C(clk32MHz), .D(pwm_setpoint_22__N_11[14]));   // verilog/TinyFPGA_B.v(96[10] 109[6])
    SB_DFF pwm_setpoint_i13 (.Q(pwm_setpoint[13]), .C(clk32MHz), .D(pwm_setpoint_22__N_11[13]));   // verilog/TinyFPGA_B.v(96[10] 109[6])
    SB_DFF pwm_setpoint_i12 (.Q(pwm_setpoint[12]), .C(clk32MHz), .D(pwm_setpoint_22__N_11[12]));   // verilog/TinyFPGA_B.v(96[10] 109[6])
    SB_DFF pwm_setpoint_i11 (.Q(pwm_setpoint[11]), .C(clk32MHz), .D(pwm_setpoint_22__N_11[11]));   // verilog/TinyFPGA_B.v(96[10] 109[6])
    SB_DFF pwm_setpoint_i10 (.Q(pwm_setpoint[10]), .C(clk32MHz), .D(pwm_setpoint_22__N_11[10]));   // verilog/TinyFPGA_B.v(96[10] 109[6])
    SB_DFF pwm_setpoint_i9 (.Q(pwm_setpoint[9]), .C(clk32MHz), .D(pwm_setpoint_22__N_11[9]));   // verilog/TinyFPGA_B.v(96[10] 109[6])
    SB_DFF pwm_setpoint_i8 (.Q(pwm_setpoint[8]), .C(clk32MHz), .D(pwm_setpoint_22__N_11[8]));   // verilog/TinyFPGA_B.v(96[10] 109[6])
    SB_DFF pwm_setpoint_i7 (.Q(pwm_setpoint[7]), .C(clk32MHz), .D(pwm_setpoint_22__N_11[7]));   // verilog/TinyFPGA_B.v(96[10] 109[6])
    SB_DFF pwm_setpoint_i6 (.Q(pwm_setpoint[6]), .C(clk32MHz), .D(pwm_setpoint_22__N_11[6]));   // verilog/TinyFPGA_B.v(96[10] 109[6])
    SB_DFF pwm_setpoint_i5 (.Q(pwm_setpoint[5]), .C(clk32MHz), .D(pwm_setpoint_22__N_11[5]));   // verilog/TinyFPGA_B.v(96[10] 109[6])
    SB_DFF pwm_setpoint_i4 (.Q(pwm_setpoint[4]), .C(clk32MHz), .D(pwm_setpoint_22__N_11[4]));   // verilog/TinyFPGA_B.v(96[10] 109[6])
    SB_DFF pwm_setpoint_i3 (.Q(pwm_setpoint[3]), .C(clk32MHz), .D(pwm_setpoint_22__N_11[3]));   // verilog/TinyFPGA_B.v(96[10] 109[6])
    SB_DFF pwm_setpoint_i2 (.Q(pwm_setpoint[2]), .C(clk32MHz), .D(pwm_setpoint_22__N_11[2]));   // verilog/TinyFPGA_B.v(96[10] 109[6])
    SB_DFF pwm_setpoint_i1 (.Q(pwm_setpoint[1]), .C(clk32MHz), .D(pwm_setpoint_22__N_11[1]));   // verilog/TinyFPGA_B.v(96[10] 109[6])
    SB_LUT4 encoder0_position_23__I_0_i1106_3_lut (.I0(n1618), .I1(n1671), 
            .I2(n1636), .I3(GND_net), .O(n1696));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1106_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14144_3_lut (.I0(neopxl_color[6]), .I1(\data_in_frame[6] [6]), 
            .I2(n3_adj_4943), .I3(GND_net), .O(n19286));   // verilog/coms.v(127[12] 300[6])
    defparam i14144_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 add_25_31_lut (.I0(GND_net), .I1(delay_counter[29]), .I2(GND_net), 
            .I3(n27761), .O(n575)) /* synthesis syn_instantiated=1 */ ;
    defparam add_25_31_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_23__I_0_i1100_3_lut (.I0(n1612), .I1(n1665), 
            .I2(n1636), .I3(GND_net), .O(n1690));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1100_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 add_672_22_lut (.I0(duty[20]), .I1(n37633), .I2(n5), .I3(n27845), 
            .O(pwm_setpoint_22__N_11[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_672_22_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_25_31 (.CI(n27761), .I0(delay_counter[29]), .I1(GND_net), 
            .CO(n27762));
    SB_LUT4 encoder0_position_23__I_0_i1103_3_lut (.I0(n1615), .I1(n1668), 
            .I2(n1636), .I3(GND_net), .O(n1693));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1103_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1108_3_lut (.I0(n1620), .I1(n1673), 
            .I2(n1636), .I3(GND_net), .O(n1698));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1108_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder1_position_23__I_0_add_2_11_lut (.I0(GND_net), .I1(encoder1_position[9]), 
            .I2(n16_adj_4956), .I3(n28082), .O(displacement_23__N_58[9])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder1_position_23__I_0_add_2_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_672_22 (.CI(n27845), .I0(n37633), .I1(n5), .CO(n27846));
    SB_LUT4 i14145_3_lut (.I0(neopxl_color[5]), .I1(\data_in_frame[6] [5]), 
            .I2(n3_adj_4943), .I3(GND_net), .O(n19287));   // verilog/coms.v(127[12] 300[6])
    defparam i14145_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14146_3_lut (.I0(neopxl_color[4]), .I1(\data_in_frame[6] [4]), 
            .I2(n3_adj_4943), .I3(GND_net), .O(n19288));   // verilog/coms.v(127[12] 300[6])
    defparam i14146_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1111_3_lut (.I0(n1623), .I1(n1676), 
            .I2(n1636), .I3(GND_net), .O(n1701));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1111_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1102_3_lut (.I0(n1614), .I1(n1667), 
            .I2(n1636), .I3(GND_net), .O(n1692));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1102_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_unary_minus_2_inv_0_i2_1_lut (.I0(encoder0_position[0]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n25_adj_5027));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_unary_minus_2_inv_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_23__I_0_unary_minus_2_inv_0_i3_1_lut (.I0(encoder0_position[1]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n24_adj_5026));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_unary_minus_2_inv_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_23__I_0_unary_minus_2_inv_0_i4_1_lut (.I0(encoder0_position[2]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n23_adj_5025));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_unary_minus_2_inv_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_23__I_0_unary_minus_2_inv_0_i5_1_lut (.I0(encoder0_position[3]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n22_adj_5024));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_unary_minus_2_inv_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_25_30_lut (.I0(GND_net), .I1(delay_counter[28]), .I2(GND_net), 
            .I3(n27760), .O(n576)) /* synthesis syn_instantiated=1 */ ;
    defparam add_25_30_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_23__I_0_i1105_3_lut (.I0(n1617), .I1(n1670), 
            .I2(n1636), .I3(GND_net), .O(n1695));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1105_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1098_3_lut (.I0(n1610), .I1(n1663), 
            .I2(n1636), .I3(GND_net), .O(n1688));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1098_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i19663_4_lut (.I0(n771_adj_4968), .I1(n1704), .I2(n1705), 
            .I3(n1706), .O(n24807));
    defparam i19663_4_lut.LUT_INIT = 16'hfcec;
    SB_LUT4 i11_4_lut_adj_1654 (.I0(n1688), .I1(n1695), .I2(n1692), .I3(n1701), 
            .O(n26_adj_5078));
    defparam i11_4_lut_adj_1654.LUT_INIT = 16'hfffe;
    SB_LUT4 i14147_3_lut (.I0(neopxl_color[3]), .I1(\data_in_frame[6] [3]), 
            .I2(n3_adj_4943), .I3(GND_net), .O(n19289));   // verilog/coms.v(127[12] 300[6])
    defparam i14147_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i4_4_lut_adj_1655 (.I0(n1700), .I1(n1703), .I2(n1702), .I3(n24807), 
            .O(n19_adj_5080));
    defparam i4_4_lut_adj_1655.LUT_INIT = 16'heaaa;
    SB_LUT4 i1424_4_lut_4_lut (.I0(\ID_READOUT_FSM.state [0]), .I1(\ID_READOUT_FSM.state [1]), 
            .I2(n691), .I3(n17358), .O(n5523));   // verilog/TinyFPGA_B.v(240[5] 264[12])
    defparam i1424_4_lut_4_lut.LUT_INIT = 16'hcc8c;
    SB_LUT4 i2_3_lut_4_lut (.I0(data_ready), .I1(n62), .I2(delay_counter[31]), 
            .I3(\ID_READOUT_FSM.state [0]), .O(n6_adj_5030));   // verilog/TinyFPGA_B.v(237[10] 265[6])
    defparam i2_3_lut_4_lut.LUT_INIT = 16'h080c;
    SB_LUT4 encoder0_position_23__I_0_unary_minus_2_inv_0_i6_1_lut (.I0(encoder0_position[4]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n21_adj_5023));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_unary_minus_2_inv_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_23__I_0_unary_minus_2_inv_0_i7_1_lut (.I0(encoder0_position[5]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n20_adj_5022));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_unary_minus_2_inv_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1_2_lut_4_lut (.I0(control_mode[0]), .I1(control_mode[6]), 
            .I2(n10_adj_5066), .I3(control_mode[2]), .O(n17355));   // verilog/TinyFPGA_B.v(165[5:22])
    defparam i1_2_lut_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 encoder0_position_23__I_0_unary_minus_2_inv_0_i8_1_lut (.I0(encoder0_position[6]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n19_adj_5021));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_unary_minus_2_inv_0_i8_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_23__I_0_unary_minus_2_inv_0_i9_1_lut (.I0(encoder0_position[7]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n18_adj_5020));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_unary_minus_2_inv_0_i9_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mux_3363_i16_3_lut (.I0(encoder0_position[15]), .I1(n10_adj_4917), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n517));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam mux_3363_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_23__I_0_unary_minus_2_inv_0_i10_1_lut (.I0(encoder0_position[8]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n17_adj_5019));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_unary_minus_2_inv_0_i10_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_23__I_0_unary_minus_2_inv_0_i11_1_lut (.I0(encoder0_position[9]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n16_adj_5018));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_unary_minus_2_inv_0_i11_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_23__I_0_unary_minus_2_inv_0_i12_1_lut (.I0(encoder0_position[10]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n15_adj_5017));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_unary_minus_2_inv_0_i12_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1_2_lut_adj_1656 (.I0(n1698), .I1(n1693), .I2(GND_net), .I3(GND_net), 
            .O(n16_adj_5081));
    defparam i1_2_lut_adj_1656.LUT_INIT = 16'heeee;
    SB_CARRY encoder1_position_23__I_0_add_2_11 (.CI(n28082), .I0(encoder1_position[9]), 
            .I1(n16_adj_4956), .CO(n28083));
    SB_LUT4 i14148_3_lut (.I0(neopxl_color[2]), .I1(\data_in_frame[6] [2]), 
            .I2(n3_adj_4943), .I3(GND_net), .O(n19290));   // verilog/coms.v(127[12] 300[6])
    defparam i14148_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14149_3_lut (.I0(neopxl_color[1]), .I1(\data_in_frame[6] [1]), 
            .I2(n3_adj_4943), .I3(GND_net), .O(n19291));   // verilog/coms.v(127[12] 300[6])
    defparam i14149_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i9_4_lut_adj_1657 (.I0(n1697), .I1(n1694), .I2(n1691), .I3(n1689), 
            .O(n24_adj_5079));
    defparam i9_4_lut_adj_1657.LUT_INIT = 16'hfffe;
    SB_LUT4 i13_4_lut_adj_1658 (.I0(n19_adj_5080), .I1(n26_adj_5078), .I2(n1690), 
            .I3(n1696), .O(n28_adj_5077));
    defparam i13_4_lut_adj_1658.LUT_INIT = 16'hfffe;
    SB_CARRY add_25_30 (.CI(n27760), .I0(delay_counter[28]), .I1(GND_net), 
            .CO(n27761));
    SB_LUT4 i30727_4_lut (.I0(n1699), .I1(n28_adj_5077), .I2(n24_adj_5079), 
            .I3(n16_adj_5081), .O(n1714));
    defparam i30727_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 encoder0_position_23__I_0_i1490_3_lut (.I0(n1714), .I1(n6218), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(encoder0_position_scaled_23__N_34[5]));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1490_3_lut.LUT_INIT = 16'hc5c5;
    SB_LUT4 i14150_3_lut (.I0(\data_out_frame[25] [7]), .I1(neopxl_color[7]), 
            .I2(n14867), .I3(GND_net), .O(n19292));   // verilog/coms.v(127[12] 300[6])
    defparam i14150_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14151_3_lut (.I0(\data_out_frame[25] [6]), .I1(neopxl_color[6]), 
            .I2(n14867), .I3(GND_net), .O(n19293));   // verilog/coms.v(127[12] 300[6])
    defparam i14151_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_672_21_lut (.I0(duty[19]), .I1(n37633), .I2(n6_adj_4885), 
            .I3(n27844), .O(pwm_setpoint_22__N_11[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_672_21_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 encoder0_position_23__I_0_i1054_3_lut (.I0(n1541), .I1(n1594), 
            .I2(n1558), .I3(GND_net), .O(n1619));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1054_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1056_3_lut (.I0(n1543), .I1(n1596), 
            .I2(n1558), .I3(GND_net), .O(n1621));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1056_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1055_3_lut (.I0(n1542), .I1(n1595), 
            .I2(n1558), .I3(GND_net), .O(n1620));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1055_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14152_3_lut (.I0(\data_out_frame[25] [5]), .I1(neopxl_color[5]), 
            .I2(n14867), .I3(GND_net), .O(n19294));   // verilog/coms.v(127[12] 300[6])
    defparam i14152_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_23__I_0_unary_minus_2_inv_0_i13_1_lut (.I0(encoder0_position[11]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n14_adj_5016));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_unary_minus_2_inv_0_i13_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder1_position_23__I_0_add_2_10_lut (.I0(GND_net), .I1(encoder1_position[8]), 
            .I2(n17_adj_4957), .I3(n28081), .O(displacement_23__N_58[8])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder1_position_23__I_0_add_2_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i14153_3_lut (.I0(\data_out_frame[25] [4]), .I1(neopxl_color[4]), 
            .I2(n14867), .I3(GND_net), .O(n19295));   // verilog/coms.v(127[12] 300[6])
    defparam i14153_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_23__I_0_unary_minus_2_inv_0_i14_1_lut (.I0(encoder0_position[12]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n13_adj_5015));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_unary_minus_2_inv_0_i14_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_23__I_0_unary_minus_2_inv_0_i15_1_lut (.I0(encoder0_position[13]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n12_adj_5014));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_unary_minus_2_inv_0_i15_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_23__I_0_i522_3_lut (.I0(n516), .I1(n812), 
            .I2(n778), .I3(GND_net), .O(n837));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i522_3_lut.LUT_INIT = 16'hacac;
    SB_IO NEOPXL_pad (.PACKAGE_PIN(NEOPXL), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(NEOPXL_c));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam NEOPXL_pad.PIN_TYPE = 6'b011001;
    defparam NEOPXL_pad.PULLUP = 1'b0;
    defparam NEOPXL_pad.NEG_TRIGGER = 1'b0;
    defparam NEOPXL_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO USBPU_pad (.PACKAGE_PIN(USBPU), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(GND_net));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam USBPU_pad.PIN_TYPE = 6'b011001;
    defparam USBPU_pad.PULLUP = 1'b0;
    defparam USBPU_pad.NEG_TRIGGER = 1'b0;
    defparam USBPU_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO LED_pad (.PACKAGE_PIN(LED), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(LED_c));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam LED_pad.PIN_TYPE = 6'b011001;
    defparam LED_pad.PULLUP = 1'b0;
    defparam LED_pad.NEG_TRIGGER = 1'b0;
    defparam LED_pad.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 i14154_3_lut (.I0(\data_out_frame[25] [3]), .I1(neopxl_color[3]), 
            .I2(n14867), .I3(GND_net), .O(n19296));   // verilog/coms.v(127[12] 300[6])
    defparam i14154_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_23__I_0_i1057_3_lut (.I0(n1544), .I1(n1597), 
            .I2(n1558), .I3(GND_net), .O(n1622));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1057_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1045_3_lut (.I0(n1532), .I1(n1585), 
            .I2(n1558), .I3(GND_net), .O(n1610));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1045_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1053_3_lut (.I0(n1540), .I1(n1593), 
            .I2(n1558), .I3(GND_net), .O(n1618));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1053_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1046_3_lut (.I0(n1533), .I1(n1586), 
            .I2(n1558), .I3(GND_net), .O(n1611));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1046_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14155_3_lut (.I0(\data_out_frame[25] [2]), .I1(neopxl_color[2]), 
            .I2(n14867), .I3(GND_net), .O(n19297));   // verilog/coms.v(127[12] 300[6])
    defparam i14155_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14156_3_lut (.I0(\data_out_frame[25] [1]), .I1(neopxl_color[1]), 
            .I2(n14867), .I3(GND_net), .O(n19298));   // verilog/coms.v(127[12] 300[6])
    defparam i14156_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14157_3_lut (.I0(\data_out_frame[25] [0]), .I1(neopxl_color[0]), 
            .I2(n14867), .I3(GND_net), .O(n19299));   // verilog/coms.v(127[12] 300[6])
    defparam i14157_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_23__I_0_i1062_3_lut (.I0(n526), .I1(n1602), 
            .I2(n1558), .I3(GND_net), .O(n1627));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1062_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1061_3_lut (.I0(n1548), .I1(n1601), 
            .I2(n1558), .I3(GND_net), .O(n1626));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1061_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_unary_minus_2_inv_0_i16_1_lut (.I0(encoder0_position[14]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n11_adj_5013));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_unary_minus_2_inv_0_i16_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i14158_3_lut (.I0(\data_out_frame[24] [7]), .I1(neopxl_color[15]), 
            .I2(n14867), .I3(GND_net), .O(n19300));   // verilog/coms.v(127[12] 300[6])
    defparam i14158_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_3363_i6_3_lut (.I0(encoder0_position[5]), .I1(n20_adj_4907), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n770));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam mux_3363_i6_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14159_3_lut (.I0(\data_out_frame[24] [6]), .I1(neopxl_color[14]), 
            .I2(n14867), .I3(GND_net), .O(n19301));   // verilog/coms.v(127[12] 300[6])
    defparam i14159_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_23__I_0_i1048_3_lut (.I0(n1535), .I1(n1588), 
            .I2(n1558), .I3(GND_net), .O(n1613));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1048_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14160_3_lut (.I0(\data_out_frame[24] [5]), .I1(neopxl_color[13]), 
            .I2(n14867), .I3(GND_net), .O(n19302));   // verilog/coms.v(127[12] 300[6])
    defparam i14160_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14161_3_lut (.I0(\data_out_frame[24] [4]), .I1(neopxl_color[12]), 
            .I2(n14867), .I3(GND_net), .O(n19303));   // verilog/coms.v(127[12] 300[6])
    defparam i14161_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_25_29_lut (.I0(GND_net), .I1(delay_counter[27]), .I2(GND_net), 
            .I3(n27759), .O(n577)) /* synthesis syn_instantiated=1 */ ;
    defparam add_25_29_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i14162_3_lut (.I0(\data_out_frame[24] [3]), .I1(neopxl_color[11]), 
            .I2(n14867), .I3(GND_net), .O(n19304));   // verilog/coms.v(127[12] 300[6])
    defparam i14162_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14163_3_lut (.I0(\data_out_frame[24] [2]), .I1(neopxl_color[10]), 
            .I2(n14867), .I3(GND_net), .O(n19305));   // verilog/coms.v(127[12] 300[6])
    defparam i14163_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14164_3_lut (.I0(\data_out_frame[24] [1]), .I1(neopxl_color[9]), 
            .I2(n14867), .I3(GND_net), .O(n19306));   // verilog/coms.v(127[12] 300[6])
    defparam i14164_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_25_29 (.CI(n27759), .I0(delay_counter[27]), .I1(GND_net), 
            .CO(n27760));
    SB_LUT4 i1_3_lut_3_lut (.I0(\ID_READOUT_FSM.state [0]), .I1(\ID_READOUT_FSM.state [1]), 
            .I2(n17358), .I3(GND_net), .O(n5410));
    defparam i1_3_lut_3_lut.LUT_INIT = 16'h1515;
    SB_LUT4 i14165_3_lut (.I0(\data_out_frame[24] [0]), .I1(neopxl_color[8]), 
            .I2(n14867), .I3(GND_net), .O(n19307));   // verilog/coms.v(127[12] 300[6])
    defparam i14165_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_23__I_0_i1051_3_lut (.I0(n1538), .I1(n1591), 
            .I2(n1558), .I3(GND_net), .O(n1616));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1051_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14166_3_lut (.I0(\data_out_frame[23] [7]), .I1(neopxl_color[23]), 
            .I2(n14867), .I3(GND_net), .O(n19308));   // verilog/coms.v(127[12] 300[6])
    defparam i14166_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_25_3_lut (.I0(GND_net), .I1(delay_counter[1]), .I2(GND_net), 
            .I3(n27733), .O(n603)) /* synthesis syn_instantiated=1 */ ;
    defparam add_25_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_23__I_0_i1050_3_lut (.I0(n1537), .I1(n1590), 
            .I2(n1558), .I3(GND_net), .O(n1615));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1050_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 add_25_28_lut (.I0(GND_net), .I1(delay_counter[26]), .I2(GND_net), 
            .I3(n27758), .O(n578)) /* synthesis syn_instantiated=1 */ ;
    defparam add_25_28_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_672_21 (.CI(n27844), .I0(n37633), .I1(n6_adj_4885), .CO(n27845));
    SB_CARRY encoder1_position_23__I_0_add_2_10 (.CI(n28081), .I0(encoder1_position[8]), 
            .I1(n17_adj_4957), .CO(n28082));
    SB_LUT4 encoder0_position_23__I_0_i1052_3_lut (.I0(n1539), .I1(n1592), 
            .I2(n1558), .I3(GND_net), .O(n1617));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1052_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14167_3_lut (.I0(\data_out_frame[23] [6]), .I1(neopxl_color[22]), 
            .I2(n14867), .I3(GND_net), .O(n19309));   // verilog/coms.v(127[12] 300[6])
    defparam i14167_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder1_position_23__I_0_add_2_9_lut (.I0(GND_net), .I1(encoder1_position[7]), 
            .I2(n18_adj_4958), .I3(n28080), .O(displacement_23__N_58[7])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder1_position_23__I_0_add_2_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_672_20_lut (.I0(duty[18]), .I1(n37633), .I2(n7_adj_4886), 
            .I3(n27843), .O(pwm_setpoint_22__N_11[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_672_20_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 i14168_3_lut (.I0(\data_out_frame[23] [5]), .I1(neopxl_color[21]), 
            .I2(n14867), .I3(GND_net), .O(n19310));   // verilog/coms.v(127[12] 300[6])
    defparam i14168_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_23__I_0_i1047_3_lut (.I0(n1534), .I1(n1587), 
            .I2(n1558), .I3(GND_net), .O(n1612));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1047_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder1_position_23__I_0_add_2_9 (.CI(n28080), .I0(encoder1_position[7]), 
            .I1(n18_adj_4958), .CO(n28081));
    SB_CARRY add_672_20 (.CI(n27843), .I0(n37633), .I1(n7_adj_4886), .CO(n27844));
    SB_LUT4 i14169_3_lut (.I0(\data_out_frame[23] [4]), .I1(neopxl_color[20]), 
            .I2(n14867), .I3(GND_net), .O(n19311));   // verilog/coms.v(127[12] 300[6])
    defparam i14169_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder1_position_23__I_0_add_2_8_lut (.I0(GND_net), .I1(encoder1_position[6]), 
            .I2(n19_adj_4959), .I3(n28079), .O(displacement_23__N_58[6])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder1_position_23__I_0_add_2_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_672_19_lut (.I0(duty[17]), .I1(n37633), .I2(n8), .I3(n27842), 
            .O(pwm_setpoint_22__N_11[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_672_19_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 encoder0_position_23__I_0_i1049_3_lut (.I0(n1536), .I1(n1589), 
            .I2(n1558), .I3(GND_net), .O(n1614));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1049_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder1_position_23__I_0_add_2_8 (.CI(n28079), .I0(encoder1_position[6]), 
            .I1(n19_adj_4959), .CO(n28080));
    SB_LUT4 i13880_3_lut (.I0(\neo_pixel_transmitter.t0 [0]), .I1(timer[0]), 
            .I2(n34265), .I3(GND_net), .O(n19022));   // verilog/neopixel.v(35[12] 117[6])
    defparam i13880_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1060_3_lut (.I0(n1547), .I1(n1600), 
            .I2(n1558), .I3(GND_net), .O(n1625));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1060_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_unary_minus_2_add_3_26_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n2_adj_5004), .I3(n28716), .O(n2)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_unary_minus_2_add_3_26_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_23__I_0_i1058_3_lut (.I0(n1545), .I1(n1598), 
            .I2(n1558), .I3(GND_net), .O(n1623));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1058_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY add_672_19 (.CI(n27842), .I0(n37633), .I1(n8), .CO(n27843));
    SB_LUT4 i13881_3_lut (.I0(IntegralLimit[0]), .I1(\data_in_frame[13] [0]), 
            .I2(n33567), .I3(GND_net), .O(n19023));   // verilog/coms.v(127[12] 300[6])
    defparam i13881_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1059_3_lut (.I0(n1546), .I1(n1599), 
            .I2(n1558), .I3(GND_net), .O(n1624));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1059_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1495_3_lut (.I0(n24787), .I1(n6223), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(encoder0_position_scaled_23__N_34[0]));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1495_3_lut.LUT_INIT = 16'hc5c5;
    SB_LUT4 i19564_3_lut (.I0(n770), .I1(n1626), .I2(n1627), .I3(GND_net), 
            .O(n24707));
    defparam i19564_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i29841_2_lut (.I0(start), .I1(n14_adj_4896), .I2(GND_net), 
            .I3(GND_net), .O(n36208));   // verilog/neopixel.v(35[12] 117[6])
    defparam i29841_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i2_4_lut_adj_1659 (.I0(n1624), .I1(n1623), .I2(n24707), .I3(n1625), 
            .O(n34021));
    defparam i2_4_lut_adj_1659.LUT_INIT = 16'h8880;
    SB_LUT4 i4_2_lut_adj_1660 (.I0(n1611), .I1(n1618), .I2(GND_net), .I3(GND_net), 
            .O(n18_adj_5086));
    defparam i4_2_lut_adj_1660.LUT_INIT = 16'heeee;
    SB_LUT4 encoder1_position_23__I_0_add_2_7_lut (.I0(GND_net), .I1(encoder1_position[5]), 
            .I2(n20_adj_4960), .I3(n28078), .O(displacement_23__N_58[5])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder1_position_23__I_0_add_2_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder1_position_23__I_0_add_2_7 (.CI(n28078), .I0(encoder1_position[5]), 
            .I1(n20_adj_4960), .CO(n28079));
    SB_LUT4 add_672_18_lut (.I0(duty[16]), .I1(n37633), .I2(n9), .I3(n27841), 
            .O(pwm_setpoint_22__N_11[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_672_18_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 i10_4_lut_adj_1661 (.I0(n1614), .I1(n1612), .I2(n1617), .I3(n1615), 
            .O(n24_adj_5084));
    defparam i10_4_lut_adj_1661.LUT_INIT = 16'hfffe;
    SB_LUT4 i8_4_lut_adj_1662 (.I0(n1610), .I1(n1622), .I2(n1620), .I3(n34021), 
            .O(n22_adj_5085));
    defparam i8_4_lut_adj_1662.LUT_INIT = 16'hfffe;
    SB_LUT4 i31_4_lut (.I0(n36208), .I1(n36206), .I2(state[1]), .I3(\neo_pixel_transmitter.done ), 
            .O(n31453));   // verilog/neopixel.v(35[12] 117[6])
    defparam i31_4_lut.LUT_INIT = 16'hcac0;
    SB_LUT4 encoder1_position_23__I_0_add_2_6_lut (.I0(GND_net), .I1(encoder1_position[4]), 
            .I2(n21_adj_4961), .I3(n28077), .O(displacement_23__N_58[4])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder1_position_23__I_0_add_2_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder1_position_23__I_0_add_2_6 (.CI(n28077), .I0(encoder1_position[4]), 
            .I1(n21_adj_4961), .CO(n28078));
    SB_LUT4 i12_4_lut_adj_1663 (.I0(n1616), .I1(n24_adj_5084), .I2(n18_adj_5086), 
            .I3(n1613), .O(n26_adj_5083));
    defparam i12_4_lut_adj_1663.LUT_INIT = 16'hfffe;
    SB_LUT4 i13887_4_lut (.I0(r_Rx_Data), .I1(rx_data[7]), .I2(n23879), 
            .I3(n17539), .O(n19029));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i13887_4_lut.LUT_INIT = 16'hccac;
    SB_LUT4 i30703_4_lut (.I0(n1621), .I1(n26_adj_5083), .I2(n22_adj_5085), 
            .I3(n1619), .O(n1636));
    defparam i30703_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 i14170_3_lut (.I0(\data_out_frame[23] [3]), .I1(neopxl_color[19]), 
            .I2(n14867), .I3(GND_net), .O(n19312));   // verilog/coms.v(127[12] 300[6])
    defparam i14170_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_23__I_0_i1489_3_lut (.I0(n1636), .I1(n6217), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(encoder0_position_scaled_23__N_34[6]));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1489_3_lut.LUT_INIT = 16'hc5c5;
    SB_LUT4 encoder0_position_23__I_0_i1001_3_lut (.I0(n1463), .I1(n1516), 
            .I2(n1480), .I3(GND_net), .O(n1541));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1001_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder1_position_23__I_0_add_2_5_lut (.I0(GND_net), .I1(encoder1_position[3]), 
            .I2(n22_adj_4962), .I3(n28076), .O(displacement_23__N_58[3])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder1_position_23__I_0_add_2_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i14171_3_lut (.I0(\data_out_frame[23] [2]), .I1(neopxl_color[18]), 
            .I2(n14867), .I3(GND_net), .O(n19313));   // verilog/coms.v(127[12] 300[6])
    defparam i14171_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_23__I_0_i995_3_lut (.I0(n1457), .I1(n1510), 
            .I2(n1480), .I3(GND_net), .O(n1535));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i995_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder1_position_23__I_0_add_2_5 (.CI(n28076), .I0(encoder1_position[3]), 
            .I1(n22_adj_4962), .CO(n28077));
    SB_LUT4 encoder0_position_23__I_0_i1003_3_lut (.I0(n1465), .I1(n1518), 
            .I2(n1480), .I3(GND_net), .O(n1543));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1003_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_unary_minus_2_inv_0_i21_1_lut (.I0(encoder0_position[19]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n6_adj_5008));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_unary_minus_2_inv_0_i21_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i14172_3_lut (.I0(\data_out_frame[23] [1]), .I1(neopxl_color[17]), 
            .I2(n14867), .I3(GND_net), .O(n19314));   // verilog/coms.v(127[12] 300[6])
    defparam i14172_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_adj_1664 (.I0(delay_counter[12]), .I1(delay_counter[11]), 
            .I2(GND_net), .I3(GND_net), .O(n4_adj_5082));
    defparam i1_2_lut_adj_1664.LUT_INIT = 16'heeee;
    SB_LUT4 encoder0_position_23__I_0_i996_3_lut (.I0(n1458), .I1(n1511), 
            .I2(n1480), .I3(GND_net), .O(n1536));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i996_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i999_3_lut (.I0(n1461), .I1(n1514), 
            .I2(n1480), .I3(GND_net), .O(n1539));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i999_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1000_3_lut (.I0(n1462), .I1(n1515), 
            .I2(n1480), .I3(GND_net), .O(n1540));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1000_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14173_3_lut (.I0(\data_out_frame[23] [0]), .I1(neopxl_color[16]), 
            .I2(n14867), .I3(GND_net), .O(n19315));   // verilog/coms.v(127[12] 300[6])
    defparam i14173_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_672_18 (.CI(n27841), .I0(n37633), .I1(n9), .CO(n27842));
    SB_LUT4 i14174_3_lut (.I0(\data_out_frame[20] [7]), .I1(displacement[7]), 
            .I2(n14867), .I3(GND_net), .O(n19316));   // verilog/coms.v(127[12] 300[6])
    defparam i14174_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder1_position_23__I_0_add_2_4_lut (.I0(GND_net), .I1(encoder1_position[2]), 
            .I2(n23_adj_4963), .I3(n28075), .O(displacement_23__N_58[2])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder1_position_23__I_0_add_2_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_23__I_0_i998_3_lut (.I0(n1460), .I1(n1513), 
            .I2(n1480), .I3(GND_net), .O(n1538));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i998_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder1_position_23__I_0_add_2_4 (.CI(n28075), .I0(encoder1_position[2]), 
            .I1(n23_adj_4963), .CO(n28076));
    SB_LUT4 i14175_3_lut (.I0(\data_out_frame[20] [6]), .I1(displacement[6]), 
            .I2(n14867), .I3(GND_net), .O(n19317));   // verilog/coms.v(127[12] 300[6])
    defparam i14175_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_23__I_0_i1002_3_lut (.I0(n1464), .I1(n1517), 
            .I2(n1480), .I3(GND_net), .O(n1542));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1002_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder1_position_23__I_0_add_2_3_lut (.I0(GND_net), .I1(encoder1_position[1]), 
            .I2(n24_adj_4964), .I3(n28074), .O(displacement_23__N_58[1])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder1_position_23__I_0_add_2_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_23__I_0_add_1361_26_lut (.I0(GND_net), .I1(n2000), 
            .I2(VCC_net), .I3(n28403), .O(n2053)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1361_26_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_23__I_0_add_1361_25_lut (.I0(GND_net), .I1(n2001), 
            .I2(VCC_net), .I3(n28402), .O(n2054)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1361_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1361_25 (.CI(n28402), .I0(n2001), 
            .I1(VCC_net), .CO(n28403));
    SB_LUT4 encoder0_position_23__I_0_add_1361_24_lut (.I0(GND_net), .I1(n2002), 
            .I2(VCC_net), .I3(n28401), .O(n2055)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1361_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_23__I_0_i993_3_lut (.I0(n1455), .I1(n1508), 
            .I2(n1480), .I3(GND_net), .O(n1533));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i993_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_23__I_0_add_1361_24 (.CI(n28401), .I0(n2002), 
            .I1(VCC_net), .CO(n28402));
    SB_LUT4 add_672_17_lut (.I0(duty[15]), .I1(n37633), .I2(n10_adj_4887), 
            .I3(n27840), .O(pwm_setpoint_22__N_11[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_672_17_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 encoder0_position_23__I_0_add_1361_23_lut (.I0(GND_net), .I1(n2003), 
            .I2(VCC_net), .I3(n28400), .O(n2056)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1361_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_23__I_0_i1008_3_lut (.I0(n768), .I1(n1523), 
            .I2(n1480), .I3(GND_net), .O(n1548));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1008_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_23__I_0_add_1361_23 (.CI(n28400), .I0(n2003), 
            .I1(VCC_net), .CO(n28401));
    SB_CARRY encoder1_position_23__I_0_add_2_3 (.CI(n28074), .I0(encoder1_position[1]), 
            .I1(n24_adj_4964), .CO(n28075));
    SB_LUT4 encoder0_position_23__I_0_i1007_3_lut (.I0(n1469), .I1(n1522), 
            .I2(n1480), .I3(GND_net), .O(n1547));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1007_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_add_1361_22_lut (.I0(GND_net), .I1(n2004), 
            .I2(VCC_net), .I3(n28399), .O(n2057)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1361_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder1_position_23__I_0_add_2_2_lut (.I0(GND_net), .I1(encoder1_position[0]), 
            .I2(n25_adj_4965), .I3(VCC_net), .O(displacement_23__N_58[0])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder1_position_23__I_0_add_2_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i14176_3_lut (.I0(\data_out_frame[20] [5]), .I1(displacement[5]), 
            .I2(n14867), .I3(GND_net), .O(n19318));   // verilog/coms.v(127[12] 300[6])
    defparam i14176_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_23__I_0_add_1361_22 (.CI(n28399), .I0(n2004), 
            .I1(VCC_net), .CO(n28400));
    SB_LUT4 i2_4_lut_adj_1665 (.I0(delay_counter[9]), .I1(n4_adj_5082), 
            .I2(delay_counter[10]), .I3(n17382), .O(n34901));
    defparam i2_4_lut_adj_1665.LUT_INIT = 16'hfcec;
    SB_LUT4 encoder0_position_23__I_0_add_1361_21_lut (.I0(GND_net), .I1(n2005), 
            .I2(VCC_net), .I3(n28398), .O(n2058)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1361_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i2_4_lut_adj_1666 (.I0(n34901), .I1(n17376), .I2(delay_counter[13]), 
            .I3(delay_counter[14]), .O(n34429));
    defparam i2_4_lut_adj_1666.LUT_INIT = 16'hffec;
    SB_CARRY encoder0_position_23__I_0_add_1361_21 (.CI(n28398), .I0(n2005), 
            .I1(VCC_net), .CO(n28399));
    SB_LUT4 encoder0_position_23__I_0_add_1361_20_lut (.I0(GND_net), .I1(n2006), 
            .I2(VCC_net), .I3(n28397), .O(n2059)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1361_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1361_20 (.CI(n28397), .I0(n2006), 
            .I1(VCC_net), .CO(n28398));
    SB_LUT4 i3_3_lut (.I0(delay_counter[20]), .I1(delay_counter[21]), .I2(delay_counter[23]), 
            .I3(GND_net), .O(n8_adj_5087));
    defparam i3_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 encoder0_position_23__I_0_i1006_3_lut (.I0(n1468), .I1(n1521), 
            .I2(n1480), .I3(GND_net), .O(n1546));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1006_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder1_position_23__I_0_add_2_2 (.CI(VCC_net), .I0(encoder1_position[0]), 
            .I1(n25_adj_4965), .CO(n28074));
    SB_LUT4 mux_3363_i7_3_lut (.I0(encoder0_position[6]), .I1(n19_adj_4908), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n526));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam mux_3363_i7_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2_4_lut_adj_1667 (.I0(delay_counter[22]), .I1(n34429), .I2(delay_counter[19]), 
            .I3(delay_counter[18]), .O(n7_adj_5088));
    defparam i2_4_lut_adj_1667.LUT_INIT = 16'ha8a0;
    SB_LUT4 i14177_3_lut (.I0(\data_out_frame[20] [4]), .I1(displacement[4]), 
            .I2(n14867), .I3(GND_net), .O(n19319));   // verilog/coms.v(127[12] 300[6])
    defparam i14177_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_23__I_0_i992_3_lut (.I0(n1454), .I1(n1507), 
            .I2(n1480), .I3(GND_net), .O(n1532));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i992_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14178_3_lut (.I0(\data_out_frame[20] [3]), .I1(displacement[3]), 
            .I2(n14867), .I3(GND_net), .O(n19320));   // verilog/coms.v(127[12] 300[6])
    defparam i14178_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_23__I_0_i997_3_lut (.I0(n1459), .I1(n1512), 
            .I2(n1480), .I3(GND_net), .O(n1537));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i997_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1004_3_lut (.I0(n1466), .I1(n1519), 
            .I2(n1480), .I3(GND_net), .O(n1544));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1004_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_add_1361_19_lut (.I0(GND_net), .I1(n2007), 
            .I2(VCC_net), .I3(n28396), .O(n2060)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1361_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1361_19 (.CI(n28396), .I0(n2007), 
            .I1(VCC_net), .CO(n28397));
    SB_LUT4 encoder0_position_23__I_0_add_1361_18_lut (.I0(GND_net), .I1(n2008), 
            .I2(VCC_net), .I3(n28395), .O(n2061)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1361_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1361_18 (.CI(n28395), .I0(n2008), 
            .I1(VCC_net), .CO(n28396));
    SB_LUT4 encoder0_position_23__I_0_add_1361_17_lut (.I0(GND_net), .I1(n2009), 
            .I2(VCC_net), .I3(n28394), .O(n2062)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1361_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_23__I_0_i994_3_lut (.I0(n1456), .I1(n1509), 
            .I2(n1480), .I3(GND_net), .O(n1534));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i994_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_23__I_0_add_1361_17 (.CI(n28394), .I0(n2009), 
            .I1(VCC_net), .CO(n28395));
    SB_LUT4 i14179_3_lut (.I0(\data_out_frame[20] [2]), .I1(displacement[2]), 
            .I2(n14867), .I3(GND_net), .O(n19321));   // verilog/coms.v(127[12] 300[6])
    defparam i14179_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_23__I_0_add_1361_16_lut (.I0(GND_net), .I1(n2010), 
            .I2(VCC_net), .I3(n28393), .O(n2063)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1361_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1361_16 (.CI(n28393), .I0(n2010), 
            .I1(VCC_net), .CO(n28394));
    SB_LUT4 encoder0_position_23__I_0_i1005_3_lut (.I0(n1467), .I1(n1520), 
            .I2(n1480), .I3(GND_net), .O(n1545));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1005_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_add_1361_15_lut (.I0(GND_net), .I1(n2011), 
            .I2(VCC_net), .I3(n28392), .O(n2064)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1361_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i19673_4_lut (.I0(n526), .I1(n1546), .I2(n1547), .I3(n1548), 
            .O(n24817));
    defparam i19673_4_lut.LUT_INIT = 16'hfcec;
    SB_CARRY encoder0_position_23__I_0_add_1361_15 (.CI(n28392), .I0(n2011), 
            .I1(VCC_net), .CO(n28393));
    SB_LUT4 i4_4_lut_adj_1668 (.I0(n1545), .I1(n1534), .I2(n1544), .I3(n24817), 
            .O(n17_adj_4893));
    defparam i4_4_lut_adj_1668.LUT_INIT = 16'heccc;
    SB_LUT4 encoder0_position_23__I_0_add_1361_14_lut (.I0(GND_net), .I1(n2012), 
            .I2(VCC_net), .I3(n28391), .O(n2065)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1361_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1361_14 (.CI(n28391), .I0(n2012), 
            .I1(VCC_net), .CO(n28392));
    SB_LUT4 i8_4_lut_adj_1669 (.I0(n1533), .I1(n1542), .I2(n1538), .I3(n1540), 
            .O(n21_adj_4891));
    defparam i8_4_lut_adj_1669.LUT_INIT = 16'hfffe;
    SB_LUT4 encoder0_position_23__I_0_add_1361_13_lut (.I0(GND_net), .I1(n2013), 
            .I2(VCC_net), .I3(n28390), .O(n2066)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1361_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1361_13 (.CI(n28390), .I0(n2013), 
            .I1(VCC_net), .CO(n28391));
    SB_LUT4 encoder0_position_23__I_0_add_1361_12_lut (.I0(GND_net), .I1(n2014), 
            .I2(VCC_net), .I3(n28389), .O(n2067)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1361_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i14180_3_lut (.I0(\data_out_frame[20] [1]), .I1(displacement[1]), 
            .I2(n14867), .I3(GND_net), .O(n19322));   // verilog/coms.v(127[12] 300[6])
    defparam i14180_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_23__I_0_add_1361_12 (.CI(n28389), .I0(n2014), 
            .I1(VCC_net), .CO(n28390));
    SB_LUT4 i7_3_lut (.I0(n1539), .I1(n1536), .I2(n1543), .I3(GND_net), 
            .O(n20_adj_4892));
    defparam i7_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 encoder0_position_23__I_0_add_1361_11_lut (.I0(GND_net), .I1(n2015), 
            .I2(VCC_net), .I3(n28388), .O(n2068)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1361_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1361_11 (.CI(n28388), .I0(n2015), 
            .I1(VCC_net), .CO(n28389));
    SB_LUT4 encoder0_position_23__I_0_add_1361_10_lut (.I0(GND_net), .I1(n2016), 
            .I2(VCC_net), .I3(n28387), .O(n2069)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1361_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i18768_4_lut (.I0(n7_adj_5088), .I1(delay_counter[31]), .I2(n17379), 
            .I3(n8_adj_5087), .O(n691));   // verilog/TinyFPGA_B.v(258[14:38])
    defparam i18768_4_lut.LUT_INIT = 16'h3230;
    SB_CARRY encoder0_position_23__I_0_add_1361_10 (.CI(n28387), .I0(n2016), 
            .I1(VCC_net), .CO(n28388));
    SB_LUT4 i5_4_lut_adj_1670 (.I0(delay_counter[27]), .I1(delay_counter[29]), 
            .I2(delay_counter[24]), .I3(delay_counter[26]), .O(n12_adj_5031));
    defparam i5_4_lut_adj_1670.LUT_INIT = 16'hfffe;
    SB_LUT4 encoder0_position_23__I_0_add_1361_9_lut (.I0(GND_net), .I1(n2017), 
            .I2(VCC_net), .I3(n28386), .O(n2070)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1361_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1361_9 (.CI(n28386), .I0(n2017), 
            .I1(VCC_net), .CO(n28387));
    SB_LUT4 encoder0_position_23__I_0_add_1361_8_lut (.I0(GND_net), .I1(n2018), 
            .I2(GND_net), .I3(n28385), .O(n2071)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1361_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i6_4_lut_adj_1671 (.I0(delay_counter[28]), .I1(n12_adj_5031), 
            .I2(delay_counter[25]), .I3(delay_counter[30]), .O(n17379));
    defparam i6_4_lut_adj_1671.LUT_INIT = 16'hfffe;
    SB_LUT4 i2_3_lut (.I0(delay_counter[17]), .I1(delay_counter[16]), .I2(delay_counter[15]), 
            .I3(GND_net), .O(n17376));
    defparam i2_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i5_3_lut (.I0(delay_counter[3]), .I1(delay_counter[5]), .I2(delay_counter[4]), 
            .I3(GND_net), .O(n14_adj_5058));
    defparam i5_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i14181_3_lut (.I0(\data_out_frame[20] [0]), .I1(displacement[0]), 
            .I2(n14867), .I3(GND_net), .O(n19323));   // verilog/coms.v(127[12] 300[6])
    defparam i14181_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11_4_lut_adj_1672 (.I0(n21_adj_4891), .I1(n17_adj_4893), .I2(n1537), 
            .I3(n1532), .O(n24_adj_4890));
    defparam i11_4_lut_adj_1672.LUT_INIT = 16'hfffe;
    SB_LUT4 i30680_4_lut (.I0(n1535), .I1(n24_adj_4890), .I2(n20_adj_4892), 
            .I3(n1541), .O(n1558));
    defparam i30680_4_lut.LUT_INIT = 16'h0001;
    SB_CARRY encoder0_position_23__I_0_add_1361_8 (.CI(n28385), .I0(n2018), 
            .I1(GND_net), .CO(n28386));
    SB_LUT4 i14182_3_lut (.I0(\data_out_frame[19] [7]), .I1(displacement[15]), 
            .I2(n14867), .I3(GND_net), .O(n19324));   // verilog/coms.v(127[12] 300[6])
    defparam i14182_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_23__I_0_add_1361_7_lut (.I0(n2073), .I1(n2019), 
            .I2(GND_net), .I3(n28384), .O(n36224)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1361_7_lut.LUT_INIT = 16'h8228;
    SB_CARRY encoder0_position_23__I_0_add_1361_7 (.CI(n28384), .I0(n2019), 
            .I1(GND_net), .CO(n28385));
    SB_LUT4 i14183_3_lut (.I0(\data_out_frame[19] [6]), .I1(displacement[14]), 
            .I2(n14867), .I3(GND_net), .O(n19325));   // verilog/coms.v(127[12] 300[6])
    defparam i14183_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_23__I_0_i1488_3_lut (.I0(n1558), .I1(n6216), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(encoder0_position_scaled_23__N_34[7]));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1488_3_lut.LUT_INIT = 16'hc5c5;
    SB_LUT4 encoder0_position_23__I_0_i940_3_lut (.I0(n1377), .I1(n1430), 
            .I2(n1402), .I3(GND_net), .O(n1455));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i940_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14184_3_lut (.I0(\data_out_frame[19] [5]), .I1(displacement[13]), 
            .I2(n14867), .I3(GND_net), .O(n19326));   // verilog/coms.v(127[12] 300[6])
    defparam i14184_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_23__I_0_i947_3_lut (.I0(n1384), .I1(n1437), 
            .I2(n1402), .I3(GND_net), .O(n1462));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i947_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14185_3_lut (.I0(\data_out_frame[19] [4]), .I1(displacement[12]), 
            .I2(n14867), .I3(GND_net), .O(n19327));   // verilog/coms.v(127[12] 300[6])
    defparam i14185_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14186_3_lut (.I0(\data_out_frame[19] [3]), .I1(displacement[11]), 
            .I2(n14867), .I3(GND_net), .O(n19328));   // verilog/coms.v(127[12] 300[6])
    defparam i14186_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_23__I_0_add_1361_6_lut (.I0(GND_net), .I1(n2020), 
            .I2(VCC_net), .I3(n28383), .O(n2073)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1361_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_23__I_0_i944_3_lut (.I0(n1381), .I1(n1434), 
            .I2(n1402), .I3(GND_net), .O(n1459));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i944_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i946_3_lut (.I0(n1383), .I1(n1436), 
            .I2(n1402), .I3(GND_net), .O(n1461));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i946_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_23__I_0_add_1361_6 (.CI(n28383), .I0(n2020), 
            .I1(VCC_net), .CO(n28384));
    SB_LUT4 encoder0_position_23__I_0_add_1361_5_lut (.I0(n6_adj_4898), .I1(n2021), 
            .I2(GND_net), .I3(n28382), .O(n36277)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1361_5_lut.LUT_INIT = 16'hebbe;
    SB_CARRY encoder0_position_23__I_0_add_1361_5 (.CI(n28382), .I0(n2021), 
            .I1(GND_net), .CO(n28383));
    SB_LUT4 encoder0_position_23__I_0_add_1361_4_lut (.I0(n2076), .I1(n2022), 
            .I2(VCC_net), .I3(n28381), .O(n6_adj_4898)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1361_4_lut.LUT_INIT = 16'h8228;
    SB_CARRY encoder0_position_23__I_0_add_1361_4 (.CI(n28381), .I0(n2022), 
            .I1(VCC_net), .CO(n28382));
    SB_LUT4 i6_4_lut_adj_1673 (.I0(delay_counter[8]), .I1(delay_counter[7]), 
            .I2(delay_counter[1]), .I3(delay_counter[0]), .O(n15_adj_5057));
    defparam i6_4_lut_adj_1673.LUT_INIT = 16'hfffe;
    SB_LUT4 i8_4_lut_adj_1674 (.I0(n15_adj_5057), .I1(delay_counter[2]), 
            .I2(n14_adj_5058), .I3(delay_counter[6]), .O(n17382));
    defparam i8_4_lut_adj_1674.LUT_INIT = 16'hfffe;
    SB_LUT4 i3396_4_lut (.I0(n17382), .I1(delay_counter[11]), .I2(delay_counter[10]), 
            .I3(delay_counter[9]), .O(n24_adj_4969));
    defparam i3396_4_lut.LUT_INIT = 16'hc8c0;
    SB_LUT4 i2_4_lut_adj_1675 (.I0(n24_adj_4969), .I1(delay_counter[14]), 
            .I2(delay_counter[12]), .I3(delay_counter[13]), .O(n34503));
    defparam i2_4_lut_adj_1675.LUT_INIT = 16'hc800;
    SB_LUT4 encoder0_position_23__I_0_i950_3_lut (.I0(n1387), .I1(n1440), 
            .I2(n1402), .I3(GND_net), .O(n1465));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i950_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_add_1361_3_lut (.I0(GND_net), .I1(n775), 
            .I2(GND_net), .I3(n28380), .O(n2076)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1361_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1361_3 (.CI(n28380), .I0(n775), 
            .I1(GND_net), .CO(n28381));
    SB_CARRY encoder0_position_23__I_0_add_1361_2 (.CI(VCC_net), .I0(GND_net), 
            .I1(VCC_net), .CO(n28380));
    SB_LUT4 add_1918_23_lut (.I0(GND_net), .I1(GND_net), .I2(VCC_net), 
            .I3(n28379), .O(n6202)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1918_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_1918_22_lut (.I0(GND_net), .I1(GND_net), .I2(VCC_net), 
            .I3(n28378), .O(n6203)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1918_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1918_22 (.CI(n28378), .I0(GND_net), .I1(VCC_net), .CO(n28379));
    SB_LUT4 add_1918_21_lut (.I0(encoder0_position[23]), .I1(GND_net), .I2(n619), 
            .I3(n28377), .O(encoder0_position_scaled_23__N_34[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1918_21_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_1918_21 (.CI(n28377), .I0(GND_net), .I1(n619), .CO(n28378));
    SB_LUT4 add_1918_20_lut (.I0(GND_net), .I1(GND_net), .I2(n700), .I3(n28376), 
            .O(n6205)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1918_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1918_20 (.CI(n28376), .I0(GND_net), .I1(n700), .CO(n28377));
    SB_LUT4 add_1918_19_lut (.I0(GND_net), .I1(GND_net), .I2(n778), .I3(n28375), 
            .O(n6206)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1918_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1918_19 (.CI(n28375), .I0(GND_net), .I1(n778), .CO(n28376));
    SB_LUT4 add_1918_18_lut (.I0(GND_net), .I1(GND_net), .I2(n856), .I3(n28374), 
            .O(n6207)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1918_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1918_18 (.CI(n28374), .I0(GND_net), .I1(n856), .CO(n28375));
    SB_LUT4 add_1918_17_lut (.I0(GND_net), .I1(GND_net), .I2(n934), .I3(n28373), 
            .O(n6208)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1918_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i2_3_lut_adj_1676 (.I0(n34503), .I1(delay_counter[18]), .I2(n17376), 
            .I3(GND_net), .O(n34410));
    defparam i2_3_lut_adj_1676.LUT_INIT = 16'hfefe;
    SB_LUT4 i2_4_lut_adj_1677 (.I0(delay_counter[23]), .I1(n34410), .I2(delay_counter[20]), 
            .I3(delay_counter[19]), .O(n7_adj_4889));
    defparam i2_4_lut_adj_1677.LUT_INIT = 16'heaaa;
    SB_LUT4 i4_4_lut_adj_1678 (.I0(n7_adj_4889), .I1(delay_counter[21]), 
            .I2(delay_counter[22]), .I3(n17379), .O(n62));
    defparam i4_4_lut_adj_1678.LUT_INIT = 16'hfffe;
    SB_CARRY add_1918_17 (.CI(n28373), .I0(GND_net), .I1(n934), .CO(n28374));
    SB_LUT4 encoder0_position_23__I_0_i951_3_lut (.I0(n1388), .I1(n1441), 
            .I2(n1402), .I3(GND_net), .O(n1466));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i951_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 add_1918_16_lut (.I0(GND_net), .I1(GND_net), .I2(n1012), .I3(n28372), 
            .O(n6209)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1918_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1918_16 (.CI(n28372), .I0(GND_net), .I1(n1012), .CO(n28373));
    SB_LUT4 i14187_3_lut (.I0(\data_out_frame[19] [2]), .I1(displacement[10]), 
            .I2(n14867), .I3(GND_net), .O(n19329));   // verilog/coms.v(127[12] 300[6])
    defparam i14187_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_23__I_0_i942_3_lut (.I0(n1379), .I1(n1432), 
            .I2(n1402), .I3(GND_net), .O(n1457));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i942_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14188_3_lut (.I0(\data_out_frame[19] [1]), .I1(displacement[9]), 
            .I2(n14867), .I3(GND_net), .O(n19330));   // verilog/coms.v(127[12] 300[6])
    defparam i14188_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_23__I_0_i954_3_lut (.I0(n767), .I1(n1444), 
            .I2(n1402), .I3(GND_net), .O(n1469));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i954_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i953_3_lut (.I0(n1390), .I1(n1443), 
            .I2(n1402), .I3(GND_net), .O(n1468));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i953_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14189_3_lut (.I0(\data_out_frame[19] [0]), .I1(displacement[8]), 
            .I2(n14867), .I3(GND_net), .O(n19331));   // verilog/coms.v(127[12] 300[6])
    defparam i14189_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_23__I_0_i952_3_lut (.I0(n1389), .I1(n1442), 
            .I2(n1402), .I3(GND_net), .O(n1467));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i952_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mux_3363_i8_3_lut (.I0(encoder0_position[7]), .I1(n18_adj_4909), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n768));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam mux_3363_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14190_3_lut (.I0(\data_out_frame[18] [7]), .I1(displacement[23]), 
            .I2(n14867), .I3(GND_net), .O(n19332));   // verilog/coms.v(127[12] 300[6])
    defparam i14190_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_1918_15_lut (.I0(GND_net), .I1(GND_net), .I2(n1090), .I3(n28371), 
            .O(n6210)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1918_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1918_15 (.CI(n28371), .I0(GND_net), .I1(n1090), .CO(n28372));
    SB_LUT4 add_1918_14_lut (.I0(GND_net), .I1(GND_net), .I2(n1168), .I3(n28370), 
            .O(n6211)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1918_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_23__I_0_i939_3_lut (.I0(n1376), .I1(n1429), 
            .I2(n1402), .I3(GND_net), .O(n1454));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i939_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i945_3_lut (.I0(n1382), .I1(n1435), 
            .I2(n1402), .I3(GND_net), .O(n1460));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i945_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13888_4_lut (.I0(r_Rx_Data), .I1(rx_data[6]), .I2(n23879), 
            .I3(n17534), .O(n19030));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i13888_4_lut.LUT_INIT = 16'hccac;
    SB_LUT4 encoder0_position_23__I_0_i941_3_lut (.I0(n1378), .I1(n1431), 
            .I2(n1402), .I3(GND_net), .O(n1456));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i941_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13889_4_lut (.I0(r_Rx_Data), .I1(rx_data[5]), .I2(n4), .I3(n17539), 
            .O(n19031));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i13889_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 encoder0_position_23__I_0_i948_3_lut (.I0(n1385), .I1(n1438), 
            .I2(n1402), .I3(GND_net), .O(n1463));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i948_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i943_3_lut (.I0(n1380), .I1(n1433), 
            .I2(n1402), .I3(GND_net), .O(n1458));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i943_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i949_3_lut (.I0(n1386), .I1(n1439), 
            .I2(n1402), .I3(GND_net), .O(n1464));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i949_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i19675_4_lut (.I0(n768), .I1(n1467), .I2(n1468), .I3(n1469), 
            .O(n24819));
    defparam i19675_4_lut.LUT_INIT = 16'hfcec;
    SB_LUT4 i18767_2_lut (.I0(n62), .I1(delay_counter[31]), .I2(GND_net), 
            .I3(GND_net), .O(read_N_295));   // verilog/TinyFPGA_B.v(243[12:35])
    defparam i18767_2_lut.LUT_INIT = 16'h2222;
    SB_CARRY add_1918_14 (.CI(n28370), .I0(GND_net), .I1(n1168), .CO(n28371));
    SB_LUT4 i13890_4_lut (.I0(r_Rx_Data), .I1(rx_data[4]), .I2(n4), .I3(n17534), 
            .O(n19032));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i13890_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i8_4_lut_adj_1679 (.I0(n1464), .I1(n1458), .I2(n1463), .I3(n1456), 
            .O(n20_adj_5054));
    defparam i8_4_lut_adj_1679.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1680 (.I0(n1457), .I1(n1466), .I2(n1465), .I3(n24819), 
            .O(n13_adj_5056));
    defparam i1_4_lut_adj_1680.LUT_INIT = 16'heaaa;
    SB_LUT4 i13891_4_lut (.I0(r_Rx_Data), .I1(rx_data[3]), .I2(n4_adj_4931), 
            .I3(n17539), .O(n19033));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i13891_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i6_2_lut (.I0(n1461), .I1(n1459), .I2(GND_net), .I3(GND_net), 
            .O(n18_adj_5055));
    defparam i6_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i13892_4_lut (.I0(r_Rx_Data), .I1(rx_data[2]), .I2(n4_adj_4931), 
            .I3(n17534), .O(n19034));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i13892_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i10_4_lut_adj_1681 (.I0(n13_adj_5056), .I1(n20_adj_5054), .I2(n1460), 
            .I3(n1454), .O(n22_adj_5053));
    defparam i10_4_lut_adj_1681.LUT_INIT = 16'hfffe;
    SB_LUT4 i30658_4_lut (.I0(n1462), .I1(n22_adj_5053), .I2(n18_adj_5055), 
            .I3(n1455), .O(n1480));
    defparam i30658_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 add_1918_13_lut (.I0(GND_net), .I1(GND_net), .I2(n1246), .I3(n28369), 
            .O(n6212)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1918_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_23__I_0_i1487_3_lut (.I0(n1480), .I1(n6215), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(encoder0_position_scaled_23__N_34[8]));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1487_3_lut.LUT_INIT = 16'hc5c5;
    SB_CARRY add_1918_13 (.CI(n28369), .I0(GND_net), .I1(n1246), .CO(n28370));
    SB_LUT4 encoder0_position_23__I_0_i892_3_lut (.I0(n1304), .I1(n1357), 
            .I2(n1324), .I3(GND_net), .O(n1382));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i892_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 add_1918_12_lut (.I0(GND_net), .I1(GND_net), .I2(n1324), .I3(n28368), 
            .O(n6213)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1918_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1918_12 (.CI(n28368), .I0(GND_net), .I1(n1324), .CO(n28369));
    SB_CARRY add_672_17 (.CI(n27840), .I0(n37633), .I1(n10_adj_4887), 
            .CO(n27841));
    SB_LUT4 encoder0_position_23__I_0_i886_3_lut (.I0(n1298), .I1(n1351), 
            .I2(n1324), .I3(GND_net), .O(n1376));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i886_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 add_672_16_lut (.I0(duty[14]), .I1(n37633), .I2(n11), .I3(n27839), 
            .O(pwm_setpoint_22__N_11[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_672_16_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 i13893_4_lut (.I0(r_Rx_Data), .I1(rx_data[1]), .I2(n4_adj_4928), 
            .I3(n17539), .O(n19035));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i13893_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 encoder0_position_23__I_0_i891_3_lut (.I0(n1303), .I1(n1356), 
            .I2(n1324), .I3(GND_net), .O(n1381));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i891_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i895_3_lut (.I0(n1307), .I1(n1360), 
            .I2(n1324), .I3(GND_net), .O(n1385));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i895_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14191_3_lut (.I0(\data_out_frame[18] [6]), .I1(displacement[22]), 
            .I2(n14867), .I3(GND_net), .O(n19333));   // verilog/coms.v(127[12] 300[6])
    defparam i14191_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_23__I_0_i898_3_lut (.I0(n1310), .I1(n1363), 
            .I2(n1324), .I3(GND_net), .O(n1388));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i898_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14192_3_lut (.I0(\data_out_frame[18] [5]), .I1(displacement[21]), 
            .I2(n14867), .I3(GND_net), .O(n19334));   // verilog/coms.v(127[12] 300[6])
    defparam i14192_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14193_3_lut (.I0(\data_out_frame[18] [4]), .I1(displacement[20]), 
            .I2(n14867), .I3(GND_net), .O(n19335));   // verilog/coms.v(127[12] 300[6])
    defparam i14193_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_23__I_0_i896_3_lut (.I0(n1308), .I1(n1361), 
            .I2(n1324), .I3(GND_net), .O(n1386));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i896_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14194_3_lut (.I0(\data_out_frame[18] [3]), .I1(displacement[19]), 
            .I2(n14867), .I3(GND_net), .O(n19336));   // verilog/coms.v(127[12] 300[6])
    defparam i14194_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_1918_11_lut (.I0(GND_net), .I1(GND_net), .I2(n1402), .I3(n28367), 
            .O(n6214)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1918_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i14195_3_lut (.I0(\data_out_frame[18] [2]), .I1(displacement[18]), 
            .I2(n14867), .I3(GND_net), .O(n19337));   // verilog/coms.v(127[12] 300[6])
    defparam i14195_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_1918_11 (.CI(n28367), .I0(GND_net), .I1(n1402), .CO(n28368));
    SB_LUT4 encoder0_position_23__I_0_i897_3_lut (.I0(n1309), .I1(n1362), 
            .I2(n1324), .I3(GND_net), .O(n1387));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i897_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14196_3_lut (.I0(\data_out_frame[18] [1]), .I1(displacement[17]), 
            .I2(n14867), .I3(GND_net), .O(n19338));   // verilog/coms.v(127[12] 300[6])
    defparam i14196_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_23__I_0_i900_3_lut (.I0(n523), .I1(n1365), 
            .I2(n1324), .I3(GND_net), .O(n1390));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i900_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY add_25_28 (.CI(n27758), .I0(delay_counter[26]), .I1(GND_net), 
            .CO(n27759));
    SB_LUT4 add_25_27_lut (.I0(GND_net), .I1(delay_counter[25]), .I2(GND_net), 
            .I3(n27757), .O(n579)) /* synthesis syn_instantiated=1 */ ;
    defparam add_25_27_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_23__I_0_i899_3_lut (.I0(n1311), .I1(n1364), 
            .I2(n1324), .I3(GND_net), .O(n1389));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i899_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14197_3_lut (.I0(\data_out_frame[18] [0]), .I1(displacement[16]), 
            .I2(n14867), .I3(GND_net), .O(n19339));   // verilog/coms.v(127[12] 300[6])
    defparam i14197_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_1918_10_lut (.I0(GND_net), .I1(GND_net), .I2(n1480), .I3(n28366), 
            .O(n6215)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1918_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mux_3363_i9_3_lut (.I0(encoder0_position[8]), .I1(n17_adj_4910), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n767));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam mux_3363_i9_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_23__I_0_i888_3_lut (.I0(n1300), .I1(n1353), 
            .I2(n1324), .I3(GND_net), .O(n1378));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i888_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14198_3_lut (.I0(\data_out_frame[17] [7]), .I1(duty[7]), .I2(n14867), 
            .I3(GND_net), .O(n19340));   // verilog/coms.v(127[12] 300[6])
    defparam i14198_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_1918_10 (.CI(n28366), .I0(GND_net), .I1(n1480), .CO(n28367));
    SB_LUT4 add_1918_9_lut (.I0(GND_net), .I1(GND_net), .I2(n1558), .I3(n28365), 
            .O(n6216)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1918_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_25_27 (.CI(n27757), .I0(delay_counter[25]), .I1(GND_net), 
            .CO(n27758));
    SB_CARRY add_1918_9 (.CI(n28365), .I0(GND_net), .I1(n1558), .CO(n28366));
    SB_LUT4 add_25_26_lut (.I0(GND_net), .I1(delay_counter[24]), .I2(GND_net), 
            .I3(n27756), .O(n580)) /* synthesis syn_instantiated=1 */ ;
    defparam add_25_26_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_1918_8_lut (.I0(GND_net), .I1(GND_net), .I2(n1636), .I3(n28364), 
            .O(n6217)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1918_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1918_8 (.CI(n28364), .I0(GND_net), .I1(n1636), .CO(n28365));
    SB_LUT4 add_1918_7_lut (.I0(GND_net), .I1(GND_net), .I2(n1714), .I3(n28363), 
            .O(n6218)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1918_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_25_26 (.CI(n27756), .I0(delay_counter[24]), .I1(GND_net), 
            .CO(n27757));
    SB_LUT4 encoder0_position_23__I_0_i894_3_lut (.I0(n1306), .I1(n1359), 
            .I2(n1324), .I3(GND_net), .O(n1384));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i894_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY add_1918_7 (.CI(n28363), .I0(GND_net), .I1(n1714), .CO(n28364));
    SB_LUT4 add_1918_6_lut (.I0(GND_net), .I1(GND_net), .I2(n1792), .I3(n28362), 
            .O(n6219)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1918_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1918_6 (.CI(n28362), .I0(GND_net), .I1(n1792), .CO(n28363));
    SB_LUT4 add_25_25_lut (.I0(GND_net), .I1(delay_counter[23]), .I2(GND_net), 
            .I3(n27755), .O(n581)) /* synthesis syn_instantiated=1 */ ;
    defparam add_25_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_1918_5_lut (.I0(GND_net), .I1(GND_net), .I2(n1870), .I3(n28361), 
            .O(n6220)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1918_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1918_5 (.CI(n28361), .I0(GND_net), .I1(n1870), .CO(n28362));
    SB_LUT4 add_1918_4_lut (.I0(GND_net), .I1(GND_net), .I2(n1948), .I3(n28360), 
            .O(n6221)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1918_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1918_4 (.CI(n28360), .I0(GND_net), .I1(n1948), .CO(n28361));
    SB_LUT4 add_1918_3_lut (.I0(GND_net), .I1(GND_net), .I2(n2026), .I3(n28359), 
            .O(n6222)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1918_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1918_3 (.CI(n28359), .I0(GND_net), .I1(n2026), .CO(n28360));
    SB_LUT4 add_1918_2_lut (.I0(GND_net), .I1(GND_net), .I2(n24787), .I3(VCC_net), 
            .O(n6223)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1918_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1918_2 (.CI(VCC_net), .I0(GND_net), .I1(n24787), .CO(n28359));
    SB_CARRY add_672_16 (.CI(n27839), .I0(n37633), .I1(n11), .CO(n27840));
    SB_LUT4 encoder0_position_23__I_0_add_1308_24_lut (.I0(GND_net), .I1(n1922), 
            .I2(VCC_net), .I3(n28358), .O(n1975)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1308_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_23__I_0_add_1308_23_lut (.I0(GND_net), .I1(n1923), 
            .I2(VCC_net), .I3(n28357), .O(n1976)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1308_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1308_23 (.CI(n28357), .I0(n1923), 
            .I1(VCC_net), .CO(n28358));
    SB_LUT4 encoder0_position_23__I_0_add_1308_22_lut (.I0(GND_net), .I1(n1924), 
            .I2(VCC_net), .I3(n28356), .O(n1977)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1308_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1308_22 (.CI(n28356), .I0(n1924), 
            .I1(VCC_net), .CO(n28357));
    SB_LUT4 encoder0_position_23__I_0_add_1308_21_lut (.I0(GND_net), .I1(n1925), 
            .I2(VCC_net), .I3(n28355), .O(n1978)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1308_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1308_21 (.CI(n28355), .I0(n1925), 
            .I1(VCC_net), .CO(n28356));
    SB_LUT4 encoder0_position_23__I_0_add_1308_20_lut (.I0(GND_net), .I1(n1926), 
            .I2(VCC_net), .I3(n28354), .O(n1979)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1308_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1308_20 (.CI(n28354), .I0(n1926), 
            .I1(VCC_net), .CO(n28355));
    SB_LUT4 add_672_15_lut (.I0(duty[13]), .I1(n37633), .I2(n12), .I3(n27838), 
            .O(pwm_setpoint_22__N_11[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_672_15_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 encoder0_position_23__I_0_add_1308_19_lut (.I0(GND_net), .I1(n1927), 
            .I2(VCC_net), .I3(n28353), .O(n1980)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1308_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1308_19 (.CI(n28353), .I0(n1927), 
            .I1(VCC_net), .CO(n28354));
    SB_LUT4 encoder0_position_23__I_0_add_1308_18_lut (.I0(GND_net), .I1(n1928), 
            .I2(VCC_net), .I3(n28352), .O(n1981)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1308_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1308_18 (.CI(n28352), .I0(n1928), 
            .I1(VCC_net), .CO(n28353));
    SB_LUT4 encoder0_position_23__I_0_add_1308_17_lut (.I0(GND_net), .I1(n1929), 
            .I2(VCC_net), .I3(n28351), .O(n1982)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1308_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_25_9_lut (.I0(GND_net), .I1(delay_counter[7]), .I2(GND_net), 
            .I3(n27739), .O(n597)) /* synthesis syn_instantiated=1 */ ;
    defparam add_25_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1308_17 (.CI(n28351), .I0(n1929), 
            .I1(VCC_net), .CO(n28352));
    SB_LUT4 encoder0_position_23__I_0_add_1308_16_lut (.I0(GND_net), .I1(n1930), 
            .I2(VCC_net), .I3(n28350), .O(n1983)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1308_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1308_16 (.CI(n28350), .I0(n1930), 
            .I1(VCC_net), .CO(n28351));
    SB_LUT4 encoder0_position_23__I_0_add_1308_15_lut (.I0(GND_net), .I1(n1931), 
            .I2(VCC_net), .I3(n28349), .O(n1984)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1308_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1308_15 (.CI(n28349), .I0(n1931), 
            .I1(VCC_net), .CO(n28350));
    SB_LUT4 encoder0_position_23__I_0_add_1308_14_lut (.I0(GND_net), .I1(n1932), 
            .I2(VCC_net), .I3(n28348), .O(n1985)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1308_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1308_14 (.CI(n28348), .I0(n1932), 
            .I1(VCC_net), .CO(n28349));
    SB_LUT4 encoder0_position_23__I_0_add_1308_13_lut (.I0(GND_net), .I1(n1933), 
            .I2(VCC_net), .I3(n28347), .O(n1986)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1308_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_23__I_0_i889_3_lut (.I0(n1301), .I1(n1354), 
            .I2(n1324), .I3(GND_net), .O(n1379));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i889_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_23__I_0_add_1308_13 (.CI(n28347), .I0(n1933), 
            .I1(VCC_net), .CO(n28348));
    SB_LUT4 encoder0_position_23__I_0_add_1308_12_lut (.I0(GND_net), .I1(n1934), 
            .I2(VCC_net), .I3(n28346), .O(n1987)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1308_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1308_12 (.CI(n28346), .I0(n1934), 
            .I1(VCC_net), .CO(n28347));
    SB_CARRY add_672_15 (.CI(n27838), .I0(n37633), .I1(n12), .CO(n27839));
    SB_LUT4 i14199_3_lut (.I0(\data_out_frame[17] [6]), .I1(duty[6]), .I2(n14867), 
            .I3(GND_net), .O(n19341));   // verilog/coms.v(127[12] 300[6])
    defparam i14199_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_23__I_0_i887_3_lut (.I0(n1299), .I1(n1352), 
            .I2(n1324), .I3(GND_net), .O(n1377));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i887_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i890_3_lut (.I0(n1302), .I1(n1355), 
            .I2(n1324), .I3(GND_net), .O(n1380));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i890_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_add_1308_11_lut (.I0(GND_net), .I1(n1935), 
            .I2(VCC_net), .I3(n28345), .O(n1988)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1308_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1308_11 (.CI(n28345), .I0(n1935), 
            .I1(VCC_net), .CO(n28346));
    SB_LUT4 encoder0_position_23__I_0_i893_3_lut (.I0(n1305), .I1(n1358), 
            .I2(n1324), .I3(GND_net), .O(n1383));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i893_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_add_1308_10_lut (.I0(GND_net), .I1(n1936), 
            .I2(VCC_net), .I3(n28344), .O(n1989)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1308_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i14200_3_lut (.I0(\data_out_frame[17] [5]), .I1(duty[5]), .I2(n14867), 
            .I3(GND_net), .O(n19342));   // verilog/coms.v(127[12] 300[6])
    defparam i14200_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14201_3_lut (.I0(\data_out_frame[17] [4]), .I1(duty[4]), .I2(n14867), 
            .I3(GND_net), .O(n19343));   // verilog/coms.v(127[12] 300[6])
    defparam i14201_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14202_3_lut (.I0(\data_out_frame[17] [3]), .I1(duty[3]), .I2(n14867), 
            .I3(GND_net), .O(n19344));   // verilog/coms.v(127[12] 300[6])
    defparam i14202_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14203_3_lut (.I0(\data_out_frame[17] [2]), .I1(duty[2]), .I2(n14867), 
            .I3(GND_net), .O(n19345));   // verilog/coms.v(127[12] 300[6])
    defparam i14203_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i19574_3_lut (.I0(n767), .I1(n1389), .I2(n1390), .I3(GND_net), 
            .O(n24717));
    defparam i19574_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i14204_3_lut (.I0(\data_out_frame[17] [1]), .I1(duty[1]), .I2(n14867), 
            .I3(GND_net), .O(n19346));   // verilog/coms.v(127[12] 300[6])
    defparam i14204_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2_4_lut_adj_1682 (.I0(n1387), .I1(n1386), .I2(n24717), .I3(n1388), 
            .O(n33923));
    defparam i2_4_lut_adj_1682.LUT_INIT = 16'h8880;
    SB_LUT4 i7_4_lut_adj_1683 (.I0(n1383), .I1(n1380), .I2(n1377), .I3(n33923), 
            .O(n18_adj_4996));
    defparam i7_4_lut_adj_1683.LUT_INIT = 16'hfffe;
    SB_LUT4 i5_2_lut (.I0(n1385), .I1(n1381), .I2(GND_net), .I3(GND_net), 
            .O(n16_adj_4997));
    defparam i5_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i14205_3_lut (.I0(\data_out_frame[17] [0]), .I1(duty[0]), .I2(n14867), 
            .I3(GND_net), .O(n19347));   // verilog/coms.v(127[12] 300[6])
    defparam i14205_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14206_3_lut (.I0(\data_out_frame[16] [7]), .I1(duty[15]), .I2(n14867), 
            .I3(GND_net), .O(n19348));   // verilog/coms.v(127[12] 300[6])
    defparam i14206_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14207_3_lut (.I0(\data_out_frame[16] [6]), .I1(duty[14]), .I2(n14867), 
            .I3(GND_net), .O(n19349));   // verilog/coms.v(127[12] 300[6])
    defparam i14207_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9_4_lut_adj_1684 (.I0(n1379), .I1(n18_adj_4996), .I2(n1384), 
            .I3(n1378), .O(n20_adj_4995));
    defparam i9_4_lut_adj_1684.LUT_INIT = 16'hfffe;
    SB_LUT4 i30447_4_lut (.I0(n1376), .I1(n20_adj_4995), .I2(n16_adj_4997), 
            .I3(n1382), .O(n1402));
    defparam i30447_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 encoder0_position_23__I_0_i1486_3_lut (.I0(n1402), .I1(n6214), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(encoder0_position_scaled_23__N_34[9]));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1486_3_lut.LUT_INIT = 16'hc5c5;
    SB_LUT4 encoder0_position_23__I_0_i834_3_lut (.I0(n1221), .I1(n1274), 
            .I2(n1246), .I3(GND_net), .O(n1299));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i834_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14208_3_lut (.I0(\data_out_frame[16] [5]), .I1(duty[13]), .I2(n14867), 
            .I3(GND_net), .O(n19350));   // verilog/coms.v(127[12] 300[6])
    defparam i14208_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_23__I_0_i836_3_lut (.I0(n1223), .I1(n1276), 
            .I2(n1246), .I3(GND_net), .O(n1301));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i836_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14209_3_lut (.I0(\data_out_frame[16] [4]), .I1(duty[12]), .I2(n14867), 
            .I3(GND_net), .O(n19351));   // verilog/coms.v(127[12] 300[6])
    defparam i14209_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_23__I_0_i839_3_lut (.I0(n1226), .I1(n1279), 
            .I2(n1246), .I3(GND_net), .O(n1304));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i839_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i841_3_lut (.I0(n1228), .I1(n1281), 
            .I2(n1246), .I3(GND_net), .O(n1306));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i841_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14210_3_lut (.I0(\data_out_frame[16] [3]), .I1(duty[11]), .I2(n14867), 
            .I3(GND_net), .O(n19352));   // verilog/coms.v(127[12] 300[6])
    defparam i14210_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14211_3_lut (.I0(\data_out_frame[16] [2]), .I1(duty[10]), .I2(n14867), 
            .I3(GND_net), .O(n19353));   // verilog/coms.v(127[12] 300[6])
    defparam i14211_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_23__I_0_i835_3_lut (.I0(n1222), .I1(n1275), 
            .I2(n1246), .I3(GND_net), .O(n1300));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i835_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i844_3_lut (.I0(n1231), .I1(n1284), 
            .I2(n1246), .I3(GND_net), .O(n1309));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i844_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14212_3_lut (.I0(\data_out_frame[16] [1]), .I1(duty[9]), .I2(n14867), 
            .I3(GND_net), .O(n19354));   // verilog/coms.v(127[12] 300[6])
    defparam i14212_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14213_3_lut (.I0(\data_out_frame[16] [0]), .I1(duty[8]), .I2(n14867), 
            .I3(GND_net), .O(n19355));   // verilog/coms.v(127[12] 300[6])
    defparam i14213_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_23__I_0_i842_3_lut (.I0(n1229), .I1(n1282), 
            .I2(n1246), .I3(GND_net), .O(n1307));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i842_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14214_3_lut (.I0(\data_out_frame[15] [7]), .I1(duty[23]), .I2(n14867), 
            .I3(GND_net), .O(n19356));   // verilog/coms.v(127[12] 300[6])
    defparam i14214_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_23__I_0_i843_3_lut (.I0(n1230), .I1(n1283), 
            .I2(n1246), .I3(GND_net), .O(n1308));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i843_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i840_3_lut (.I0(n1227), .I1(n1280), 
            .I2(n1246), .I3(GND_net), .O(n1305));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i840_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 add_672_14_lut (.I0(duty[12]), .I1(n37633), .I2(n13), .I3(n27837), 
            .O(pwm_setpoint_22__N_11[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_672_14_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 i14215_3_lut (.I0(\data_out_frame[15] [6]), .I1(duty[22]), .I2(n14867), 
            .I3(GND_net), .O(n19357));   // verilog/coms.v(127[12] 300[6])
    defparam i14215_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_25_25 (.CI(n27755), .I0(delay_counter[23]), .I1(GND_net), 
            .CO(n27756));
    SB_CARRY encoder0_position_23__I_0_add_1308_10 (.CI(n28344), .I0(n1936), 
            .I1(VCC_net), .CO(n28345));
    SB_LUT4 encoder0_position_23__I_0_add_1308_9_lut (.I0(GND_net), .I1(n1937), 
            .I2(VCC_net), .I3(n28343), .O(n1990)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1308_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1308_9 (.CI(n28343), .I0(n1937), 
            .I1(VCC_net), .CO(n28344));
    SB_LUT4 encoder0_position_23__I_0_add_1308_8_lut (.I0(GND_net), .I1(n1938), 
            .I2(VCC_net), .I3(n28342), .O(n1991)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1308_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1308_8 (.CI(n28342), .I0(n1938), 
            .I1(VCC_net), .CO(n28343));
    SB_LUT4 encoder0_position_23__I_0_add_1308_7_lut (.I0(GND_net), .I1(n1939), 
            .I2(GND_net), .I3(n28341), .O(n1992)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1308_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1308_7 (.CI(n28341), .I0(n1939), 
            .I1(GND_net), .CO(n28342));
    SB_LUT4 encoder0_position_23__I_0_add_1308_6_lut (.I0(GND_net), .I1(n1940), 
            .I2(GND_net), .I3(n28340), .O(n1993)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1308_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_23__I_0_i833_3_lut (.I0(n1220), .I1(n1273), 
            .I2(n1246), .I3(GND_net), .O(n1298));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i833_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14216_3_lut (.I0(\data_out_frame[15] [5]), .I1(duty[21]), .I2(n14867), 
            .I3(GND_net), .O(n19358));   // verilog/coms.v(127[12] 300[6])
    defparam i14216_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_23__I_0_i837_3_lut (.I0(n1224), .I1(n1277), 
            .I2(n1246), .I3(GND_net), .O(n1302));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i837_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i838_3_lut (.I0(n1225), .I1(n1278), 
            .I2(n1246), .I3(GND_net), .O(n1303));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i838_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i846_3_lut (.I0(n765), .I1(n1286), 
            .I2(n1246), .I3(GND_net), .O(n1311));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i846_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i845_3_lut (.I0(n1232), .I1(n1285), 
            .I2(n1246), .I3(GND_net), .O(n1310));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i845_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mux_3363_i10_3_lut (.I0(encoder0_position[9]), .I1(n16_adj_4911), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n523));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam mux_3363_i10_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14217_3_lut (.I0(\data_out_frame[15] [4]), .I1(duty[20]), .I2(n14867), 
            .I3(GND_net), .O(n19359));   // verilog/coms.v(127[12] 300[6])
    defparam i14217_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14218_3_lut (.I0(\data_out_frame[15] [3]), .I1(duty[19]), .I2(n14867), 
            .I3(GND_net), .O(n19360));   // verilog/coms.v(127[12] 300[6])
    defparam i14218_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14219_3_lut (.I0(\data_out_frame[15] [2]), .I1(duty[18]), .I2(n14867), 
            .I3(GND_net), .O(n19361));   // verilog/coms.v(127[12] 300[6])
    defparam i14219_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_23__I_0_add_1308_6 (.CI(n28340), .I0(n1940), 
            .I1(GND_net), .CO(n28341));
    SB_LUT4 encoder0_position_23__I_0_add_1308_5_lut (.I0(GND_net), .I1(n1941), 
            .I2(VCC_net), .I3(n28339), .O(n1994)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1308_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i19578_3_lut (.I0(n523), .I1(n1310), .I2(n1311), .I3(GND_net), 
            .O(n24721));
    defparam i19578_3_lut.LUT_INIT = 16'hc8c8;
    SB_CARRY encoder0_position_23__I_0_add_1308_5 (.CI(n28339), .I0(n1941), 
            .I1(VCC_net), .CO(n28340));
    SB_LUT4 encoder0_position_23__I_0_add_1308_4_lut (.I0(GND_net), .I1(n1942), 
            .I2(GND_net), .I3(n28338), .O(n1995)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1308_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1308_4 (.CI(n28338), .I0(n1942), 
            .I1(GND_net), .CO(n28339));
    SB_LUT4 encoder0_position_23__I_0_add_1308_3_lut (.I0(GND_net), .I1(n1943), 
            .I2(VCC_net), .I3(n28337), .O(n1996)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1308_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_672_14 (.CI(n27837), .I0(n37633), .I1(n13), .CO(n27838));
    SB_CARRY encoder0_position_23__I_0_add_1308_3 (.CI(n28337), .I0(n1943), 
            .I1(VCC_net), .CO(n28338));
    SB_LUT4 encoder0_position_23__I_0_add_1308_2_lut (.I0(GND_net), .I1(n774), 
            .I2(GND_net), .I3(VCC_net), .O(n1997)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1308_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1308_2 (.CI(VCC_net), .I0(n774), 
            .I1(GND_net), .CO(n28337));
    SB_LUT4 i2_4_lut_adj_1685 (.I0(n1308), .I1(n1307), .I2(n24721), .I3(n1309), 
            .O(n34006));
    defparam i2_4_lut_adj_1685.LUT_INIT = 16'h8880;
    SB_LUT4 encoder0_position_23__I_0_add_1255_23_lut (.I0(GND_net), .I1(n1844), 
            .I2(VCC_net), .I3(n28336), .O(n1897)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1255_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i6_4_lut_adj_1686 (.I0(n1300), .I1(n34006), .I2(n1306), .I3(n1304), 
            .O(n16_adj_5064));
    defparam i6_4_lut_adj_1686.LUT_INIT = 16'hfffe;
    SB_LUT4 i14220_3_lut (.I0(\data_out_frame[15] [1]), .I1(duty[17]), .I2(n14867), 
            .I3(GND_net), .O(n19362));   // verilog/coms.v(127[12] 300[6])
    defparam i14220_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_23__I_0_add_1255_22_lut (.I0(GND_net), .I1(n1845), 
            .I2(VCC_net), .I3(n28335), .O(n1898)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1255_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_25_24_lut (.I0(GND_net), .I1(delay_counter[22]), .I2(GND_net), 
            .I3(n27754), .O(n582)) /* synthesis syn_instantiated=1 */ ;
    defparam add_25_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i7_4_lut_adj_1687 (.I0(n1303), .I1(n1302), .I2(n1298), .I3(n1305), 
            .O(n17_adj_5063));
    defparam i7_4_lut_adj_1687.LUT_INIT = 16'hfffe;
    SB_LUT4 i30856_4_lut (.I0(n17_adj_5063), .I1(n1301), .I2(n16_adj_5064), 
            .I3(n1299), .O(n1324));
    defparam i30856_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 i14221_3_lut (.I0(\data_out_frame[15] [0]), .I1(duty[16]), .I2(n14867), 
            .I3(GND_net), .O(n19363));   // verilog/coms.v(127[12] 300[6])
    defparam i14221_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_23__I_0_i1485_3_lut (.I0(n1324), .I1(n6213), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(encoder0_position_scaled_23__N_34[10]));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1485_3_lut.LUT_INIT = 16'hc5c5;
    SB_CARRY encoder0_position_23__I_0_add_1255_22 (.CI(n28335), .I0(n1845), 
            .I1(VCC_net), .CO(n28336));
    SB_LUT4 i14222_3_lut (.I0(\data_out_frame[14] [7]), .I1(setpoint[7]), 
            .I2(n14867), .I3(GND_net), .O(n19364));   // verilog/coms.v(127[12] 300[6])
    defparam i14222_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_23__I_0_i785_3_lut (.I0(n1147), .I1(n1200), 
            .I2(n1168), .I3(GND_net), .O(n1225));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i785_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i780_3_lut (.I0(n1142), .I1(n1195), 
            .I2(n1168), .I3(GND_net), .O(n1220));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i780_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14223_3_lut (.I0(\data_out_frame[14] [6]), .I1(setpoint[6]), 
            .I2(n14867), .I3(GND_net), .O(n19365));   // verilog/coms.v(127[12] 300[6])
    defparam i14223_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_23__I_0_i786_3_lut (.I0(n1148), .I1(n1201), 
            .I2(n1168), .I3(GND_net), .O(n1226));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i786_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i781_3_lut (.I0(n1143), .I1(n1196), 
            .I2(n1168), .I3(GND_net), .O(n1221));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i781_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14224_3_lut (.I0(\data_out_frame[14] [5]), .I1(setpoint[5]), 
            .I2(n14867), .I3(GND_net), .O(n19366));   // verilog/coms.v(127[12] 300[6])
    defparam i14224_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2_2_lut_adj_1688 (.I0(ID[2]), .I1(ID[4]), .I2(GND_net), .I3(GND_net), 
            .O(n10_adj_5069));   // verilog/TinyFPGA_B.v(256[12:17])
    defparam i2_2_lut_adj_1688.LUT_INIT = 16'heeee;
    SB_LUT4 i6_4_lut_adj_1689 (.I0(ID[7]), .I1(ID[5]), .I2(ID[1]), .I3(ID[0]), 
            .O(n14_adj_5068));   // verilog/TinyFPGA_B.v(256[12:17])
    defparam i6_4_lut_adj_1689.LUT_INIT = 16'hfffe;
    SB_LUT4 encoder0_position_23__I_0_i784_3_lut (.I0(n1146), .I1(n1199), 
            .I2(n1168), .I3(GND_net), .O(n1224));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i784_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14225_3_lut (.I0(\data_out_frame[14] [4]), .I1(setpoint[4]), 
            .I2(n14867), .I3(GND_net), .O(n19367));   // verilog/coms.v(127[12] 300[6])
    defparam i14225_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_23__I_0_i783_3_lut (.I0(n1145), .I1(n1198), 
            .I2(n1168), .I3(GND_net), .O(n1223));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i783_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_add_1255_21_lut (.I0(GND_net), .I1(n1846), 
            .I2(VCC_net), .I3(n28334), .O(n1899)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1255_21_lut.LUT_INIT = 16'hC33C;
    SB_DFFESR delay_counter_i0_i31 (.Q(delay_counter[31]), .C(CLK_c), .E(n5410), 
            .D(n573), .R(n18963));   // verilog/TinyFPGA_B.v(237[10] 265[6])
    SB_LUT4 i7_4_lut_adj_1690 (.I0(ID[3]), .I1(n14_adj_5068), .I2(n10_adj_5069), 
            .I3(ID[6]), .O(n17358));   // verilog/TinyFPGA_B.v(256[12:17])
    defparam i7_4_lut_adj_1690.LUT_INIT = 16'hfffe;
    SB_LUT4 encoder0_position_23__I_0_i787_3_lut (.I0(n1149), .I1(n1202), 
            .I2(n1168), .I3(GND_net), .O(n1227));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i787_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i788_3_lut (.I0(n1150), .I1(n1203), 
            .I2(n1168), .I3(GND_net), .O(n1228));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i788_3_lut.LUT_INIT = 16'hacac;
    SB_DFFESR delay_counter_i0_i16 (.Q(delay_counter[16]), .C(CLK_c), .E(n5410), 
            .D(n588), .R(n18963));   // verilog/TinyFPGA_B.v(237[10] 265[6])
    SB_CARRY encoder0_position_23__I_0_add_1255_21 (.CI(n28334), .I0(n1846), 
            .I1(VCC_net), .CO(n28335));
    SB_DFFESR delay_counter_i0_i15 (.Q(delay_counter[15]), .C(CLK_c), .E(n5410), 
            .D(n589), .R(n18963));   // verilog/TinyFPGA_B.v(237[10] 265[6])
    SB_DFFESR delay_counter_i0_i30 (.Q(delay_counter[30]), .C(CLK_c), .E(n5410), 
            .D(n574), .R(n18963));   // verilog/TinyFPGA_B.v(237[10] 265[6])
    SB_LUT4 encoder0_position_23__I_0_i789_3_lut (.I0(n1151), .I1(n1204), 
            .I2(n1168), .I3(GND_net), .O(n1229));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i789_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i782_3_lut (.I0(n1144), .I1(n1197), 
            .I2(n1168), .I3(GND_net), .O(n1222));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i782_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i792_3_lut (.I0(n521), .I1(n1207), 
            .I2(n1168), .I3(GND_net), .O(n1232));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i792_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i791_3_lut (.I0(n1153), .I1(n1206), 
            .I2(n1168), .I3(GND_net), .O(n1231));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i791_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i790_3_lut (.I0(n1152), .I1(n1205), 
            .I2(n1168), .I3(GND_net), .O(n1230));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i790_3_lut.LUT_INIT = 16'hacac;
    SB_DFFESR delay_counter_i0_i29 (.Q(delay_counter[29]), .C(CLK_c), .E(n5410), 
            .D(n575), .R(n18963));   // verilog/TinyFPGA_B.v(237[10] 265[6])
    SB_DFFESR delay_counter_i0_i14 (.Q(delay_counter[14]), .C(CLK_c), .E(n5410), 
            .D(n590), .R(n18963));   // verilog/TinyFPGA_B.v(237[10] 265[6])
    SB_LUT4 mux_3363_i11_3_lut (.I0(encoder0_position[10]), .I1(n15_adj_4912), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n765));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam mux_3363_i11_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i19682_4_lut (.I0(n765), .I1(n1230), .I2(n1231), .I3(n1232), 
            .O(n24827));
    defparam i19682_4_lut.LUT_INIT = 16'hfcec;
    SB_LUT4 encoder0_position_23__I_0_add_1255_20_lut (.I0(GND_net), .I1(n1847), 
            .I2(VCC_net), .I3(n28333), .O(n1900)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1255_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1255_20 (.CI(n28333), .I0(n1847), 
            .I1(VCC_net), .CO(n28334));
    SB_LUT4 encoder0_position_23__I_0_add_1255_19_lut (.I0(GND_net), .I1(n1848), 
            .I2(VCC_net), .I3(n28332), .O(n1901)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1255_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1255_19 (.CI(n28332), .I0(n1848), 
            .I1(VCC_net), .CO(n28333));
    SB_LUT4 encoder0_position_23__I_0_add_1255_18_lut (.I0(GND_net), .I1(n1849), 
            .I2(VCC_net), .I3(n28331), .O(n1902)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1255_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1255_18 (.CI(n28331), .I0(n1849), 
            .I1(VCC_net), .CO(n28332));
    SB_LUT4 i4_4_lut_adj_1691 (.I0(n1222), .I1(n1229), .I2(n1228), .I3(n24827), 
            .O(n13_adj_4993));
    defparam i4_4_lut_adj_1691.LUT_INIT = 16'heaaa;
    SB_LUT4 encoder0_position_23__I_0_add_1255_17_lut (.I0(GND_net), .I1(n1850), 
            .I2(VCC_net), .I3(n28330), .O(n1903)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1255_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1255_17 (.CI(n28330), .I0(n1850), 
            .I1(VCC_net), .CO(n28331));
    SB_LUT4 encoder0_position_23__I_0_add_1255_16_lut (.I0(GND_net), .I1(n1851), 
            .I2(VCC_net), .I3(n28329), .O(n1904)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1255_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1255_16 (.CI(n28329), .I0(n1851), 
            .I1(VCC_net), .CO(n28330));
    SB_DFFESR delay_counter_i0_i13 (.Q(delay_counter[13]), .C(CLK_c), .E(n5410), 
            .D(n591), .R(n18963));   // verilog/TinyFPGA_B.v(237[10] 265[6])
    SB_DFFESR delay_counter_i0_i12 (.Q(delay_counter[12]), .C(CLK_c), .E(n5410), 
            .D(n592), .R(n18963));   // verilog/TinyFPGA_B.v(237[10] 265[6])
    SB_DFFESR delay_counter_i0_i28 (.Q(delay_counter[28]), .C(CLK_c), .E(n5410), 
            .D(n576), .R(n18963));   // verilog/TinyFPGA_B.v(237[10] 265[6])
    SB_DFFESR delay_counter_i0_i27 (.Q(delay_counter[27]), .C(CLK_c), .E(n5410), 
            .D(n577), .R(n18963));   // verilog/TinyFPGA_B.v(237[10] 265[6])
    SB_LUT4 encoder0_position_23__I_0_add_1255_15_lut (.I0(GND_net), .I1(n1852), 
            .I2(VCC_net), .I3(n28328), .O(n1905)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1255_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i3_2_lut (.I0(n1221), .I1(n1226), .I2(GND_net), .I3(GND_net), 
            .O(n12_adj_4994));
    defparam i3_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i7_4_lut_adj_1692 (.I0(n13_adj_4993), .I1(n1227), .I2(n1223), 
            .I3(n1224), .O(n16_adj_4992));
    defparam i7_4_lut_adj_1692.LUT_INIT = 16'hfffe;
    SB_LUT4 i30525_4_lut (.I0(n1220), .I1(n16_adj_4992), .I2(n12_adj_4994), 
            .I3(n1225), .O(n1246));
    defparam i30525_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 i14226_3_lut (.I0(\data_out_frame[14] [3]), .I1(setpoint[3]), 
            .I2(n14867), .I3(GND_net), .O(n19368));   // verilog/coms.v(127[12] 300[6])
    defparam i14226_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14227_3_lut (.I0(\data_out_frame[14] [2]), .I1(setpoint[2]), 
            .I2(n14867), .I3(GND_net), .O(n19369));   // verilog/coms.v(127[12] 300[6])
    defparam i14227_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14228_3_lut (.I0(\data_out_frame[14] [1]), .I1(setpoint[1]), 
            .I2(n14867), .I3(GND_net), .O(n19370));   // verilog/coms.v(127[12] 300[6])
    defparam i14228_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_23__I_0_add_1255_15 (.CI(n28328), .I0(n1852), 
            .I1(VCC_net), .CO(n28329));
    SB_LUT4 encoder0_position_23__I_0_i1484_3_lut (.I0(n1246), .I1(n6212), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(encoder0_position_scaled_23__N_34[11]));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1484_3_lut.LUT_INIT = 16'hc5c5;
    SB_LUT4 add_672_13_lut (.I0(duty[11]), .I1(n37633), .I2(n14), .I3(n27836), 
            .O(pwm_setpoint_22__N_11[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_672_13_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 encoder0_position_23__I_0_add_1255_14_lut (.I0(GND_net), .I1(n1853), 
            .I2(VCC_net), .I3(n28327), .O(n1906)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1255_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1255_14 (.CI(n28327), .I0(n1853), 
            .I1(VCC_net), .CO(n28328));
    SB_LUT4 encoder0_position_23__I_0_add_1255_13_lut (.I0(GND_net), .I1(n1854), 
            .I2(VCC_net), .I3(n28326), .O(n1907)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1255_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1255_13 (.CI(n28326), .I0(n1854), 
            .I1(VCC_net), .CO(n28327));
    SB_LUT4 encoder0_position_23__I_0_add_1255_12_lut (.I0(GND_net), .I1(n1855), 
            .I2(VCC_net), .I3(n28325), .O(n1908)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1255_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1255_12 (.CI(n28325), .I0(n1855), 
            .I1(VCC_net), .CO(n28326));
    SB_LUT4 encoder0_position_23__I_0_add_1255_11_lut (.I0(GND_net), .I1(n1856), 
            .I2(VCC_net), .I3(n28324), .O(n1909)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1255_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_672_13 (.CI(n27836), .I0(n37633), .I1(n14), .CO(n27837));
    SB_CARRY encoder0_position_23__I_0_add_1255_11 (.CI(n28324), .I0(n1856), 
            .I1(VCC_net), .CO(n28325));
    SB_LUT4 encoder0_position_23__I_0_add_1255_10_lut (.I0(GND_net), .I1(n1857), 
            .I2(VCC_net), .I3(n28323), .O(n1910)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1255_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1255_10 (.CI(n28323), .I0(n1857), 
            .I1(VCC_net), .CO(n28324));
    SB_LUT4 encoder0_position_23__I_0_add_1255_9_lut (.I0(GND_net), .I1(n1858), 
            .I2(VCC_net), .I3(n28322), .O(n1911)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1255_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1255_9 (.CI(n28322), .I0(n1858), 
            .I1(VCC_net), .CO(n28323));
    SB_LUT4 encoder0_position_23__I_0_add_1255_8_lut (.I0(GND_net), .I1(n1859), 
            .I2(VCC_net), .I3(n28321), .O(n1912)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1255_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1255_8 (.CI(n28321), .I0(n1859), 
            .I1(VCC_net), .CO(n28322));
    SB_LUT4 add_672_12_lut (.I0(duty[10]), .I1(n37633), .I2(n15), .I3(n27835), 
            .O(pwm_setpoint_22__N_11[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_672_12_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_672_12 (.CI(n27835), .I0(n37633), .I1(n15), .CO(n27836));
    SB_LUT4 add_672_11_lut (.I0(duty[9]), .I1(n37633), .I2(n16), .I3(n27834), 
            .O(pwm_setpoint_22__N_11[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_672_11_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 encoder0_position_23__I_0_add_1255_7_lut (.I0(GND_net), .I1(n1860), 
            .I2(GND_net), .I3(n28320), .O(n1913)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1255_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1255_7 (.CI(n28320), .I0(n1860), 
            .I1(GND_net), .CO(n28321));
    SB_LUT4 encoder0_position_23__I_0_add_1255_6_lut (.I0(GND_net), .I1(n1861), 
            .I2(GND_net), .I3(n28319), .O(n1914)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1255_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1255_6 (.CI(n28319), .I0(n1861), 
            .I1(GND_net), .CO(n28320));
    SB_LUT4 encoder0_position_23__I_0_add_1255_5_lut (.I0(GND_net), .I1(n1862), 
            .I2(VCC_net), .I3(n28318), .O(n1915)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1255_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1255_5 (.CI(n28318), .I0(n1862), 
            .I1(VCC_net), .CO(n28319));
    SB_LUT4 encoder0_position_23__I_0_add_1255_4_lut (.I0(GND_net), .I1(n1863), 
            .I2(GND_net), .I3(n28317), .O(n1916)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1255_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1255_4 (.CI(n28317), .I0(n1863), 
            .I1(GND_net), .CO(n28318));
    SB_LUT4 encoder0_position_23__I_0_add_1255_3_lut (.I0(GND_net), .I1(n1864), 
            .I2(VCC_net), .I3(n28316), .O(n1917)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1255_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1255_3 (.CI(n28316), .I0(n1864), 
            .I1(VCC_net), .CO(n28317));
    SB_LUT4 encoder0_position_23__I_0_add_1255_2_lut (.I0(GND_net), .I1(n773), 
            .I2(GND_net), .I3(VCC_net), .O(n1918)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1255_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 \ID_READOUT_FSM.state_2__I_0_i5_2_lut  (.I0(\ID_READOUT_FSM.state [0]), 
            .I1(\ID_READOUT_FSM.state [1]), .I2(GND_net), .I3(GND_net), 
            .O(n5_adj_4966));   // verilog/TinyFPGA_B.v(255[7:11])
    defparam \ID_READOUT_FSM.state_2__I_0_i5_2_lut .LUT_INIT = 16'hbbbb;
    SB_CARRY encoder0_position_23__I_0_add_1255_2 (.CI(VCC_net), .I0(n773), 
            .I1(GND_net), .CO(n28316));
    SB_LUT4 encoder0_position_23__I_0_add_1202_22_lut (.I0(GND_net), .I1(n1766), 
            .I2(VCC_net), .I3(n28315), .O(n1819)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1202_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_23__I_0_add_1202_21_lut (.I0(GND_net), .I1(n1767), 
            .I2(VCC_net), .I3(n28314), .O(n1820)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1202_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_25_24 (.CI(n27754), .I0(delay_counter[22]), .I1(GND_net), 
            .CO(n27755));
    SB_CARRY add_672_11 (.CI(n27834), .I0(n37633), .I1(n16), .CO(n27835));
    SB_CARRY encoder0_position_23__I_0_add_1202_21 (.CI(n28314), .I0(n1767), 
            .I1(VCC_net), .CO(n28315));
    SB_LUT4 encoder0_position_23__I_0_add_1202_20_lut (.I0(GND_net), .I1(n1768), 
            .I2(VCC_net), .I3(n28313), .O(n1821)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1202_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i14229_3_lut (.I0(\data_out_frame[14] [0]), .I1(setpoint[0]), 
            .I2(n14867), .I3(GND_net), .O(n19371));   // verilog/coms.v(127[12] 300[6])
    defparam i14229_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14230_3_lut (.I0(\data_out_frame[13] [7]), .I1(setpoint[15]), 
            .I2(n14867), .I3(GND_net), .O(n19372));   // verilog/coms.v(127[12] 300[6])
    defparam i14230_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_23__I_0_i728_3_lut (.I0(n1065), .I1(n1118), 
            .I2(n1090), .I3(GND_net), .O(n1143));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i728_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i727_3_lut (.I0(n1064), .I1(n1117), 
            .I2(n1090), .I3(GND_net), .O(n1142));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i727_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14231_3_lut (.I0(\data_out_frame[13] [6]), .I1(setpoint[14]), 
            .I2(n14867), .I3(GND_net), .O(n19373));   // verilog/coms.v(127[12] 300[6])
    defparam i14231_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_23__I_0_i738_3_lut (.I0(n763), .I1(n1128), 
            .I2(n1090), .I3(GND_net), .O(n1153));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i738_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i737_3_lut (.I0(n1074), .I1(n1127), 
            .I2(n1090), .I3(GND_net), .O(n1152));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i737_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i736_3_lut (.I0(n1073), .I1(n1126), 
            .I2(n1090), .I3(GND_net), .O(n1151));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i736_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mux_3363_i12_3_lut (.I0(encoder0_position[11]), .I1(n14_adj_4913), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n521));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam mux_3363_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14232_3_lut (.I0(\data_out_frame[13] [5]), .I1(setpoint[13]), 
            .I2(n14867), .I3(GND_net), .O(n19374));   // verilog/coms.v(127[12] 300[6])
    defparam i14232_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_23__I_0_i734_3_lut (.I0(n1071), .I1(n1124), 
            .I2(n1090), .I3(GND_net), .O(n1149));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i734_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i730_3_lut (.I0(n1067), .I1(n1120), 
            .I2(n1090), .I3(GND_net), .O(n1145));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i730_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i735_3_lut (.I0(n1072), .I1(n1125), 
            .I2(n1090), .I3(GND_net), .O(n1150));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i735_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i732_3_lut (.I0(n1069), .I1(n1122), 
            .I2(n1090), .I3(GND_net), .O(n1147));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i732_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i729_3_lut (.I0(n1066), .I1(n1119), 
            .I2(n1090), .I3(GND_net), .O(n1144));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i729_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i733_3_lut (.I0(n1070), .I1(n1123), 
            .I2(n1090), .I3(GND_net), .O(n1148));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i733_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i731_3_lut (.I0(n1068), .I1(n1121), 
            .I2(n1090), .I3(GND_net), .O(n1146));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i731_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i19684_4_lut (.I0(n521), .I1(n1151), .I2(n1152), .I3(n1153), 
            .O(n24829));
    defparam i19684_4_lut.LUT_INIT = 16'hfcec;
    SB_LUT4 i6_4_lut_adj_1693 (.I0(n1146), .I1(n1148), .I2(n1144), .I3(n1147), 
            .O(n14_adj_5061));
    defparam i6_4_lut_adj_1693.LUT_INIT = 16'hfffe;
    SB_LUT4 i14233_3_lut (.I0(\data_out_frame[13] [4]), .I1(setpoint[12]), 
            .I2(n14867), .I3(GND_net), .O(n19375));   // verilog/coms.v(127[12] 300[6])
    defparam i14233_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14234_3_lut (.I0(\data_out_frame[13] [3]), .I1(setpoint[11]), 
            .I2(n14867), .I3(GND_net), .O(n19376));   // verilog/coms.v(127[12] 300[6])
    defparam i14234_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_1694 (.I0(n1150), .I1(n1145), .I2(n1149), .I3(n24829), 
            .O(n9_adj_5062));
    defparam i1_4_lut_adj_1694.LUT_INIT = 16'heccc;
    SB_LUT4 i30559_4_lut (.I0(n9_adj_5062), .I1(n14_adj_5061), .I2(n1142), 
            .I3(n1143), .O(n1168));
    defparam i30559_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 encoder0_position_23__I_0_i1483_3_lut (.I0(n1168), .I1(n6211), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(encoder0_position_scaled_23__N_34[12]));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1483_3_lut.LUT_INIT = 16'hc5c5;
    SB_LUT4 encoder0_position_23__I_0_i679_3_lut (.I0(n991), .I1(n1044), 
            .I2(n1012), .I3(GND_net), .O(n1069));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i679_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i676_3_lut (.I0(n988), .I1(n1041), 
            .I2(n1012), .I3(GND_net), .O(n1066));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i676_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i677_3_lut (.I0(n989), .I1(n1042), 
            .I2(n1012), .I3(GND_net), .O(n1067));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i677_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i682_3_lut (.I0(n994), .I1(n1047), 
            .I2(n1012), .I3(GND_net), .O(n1072));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i682_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 LessThan_744_i6_3_lut_3_lut (.I0(pwm_setpoint[2]), .I1(pwm_setpoint[3]), 
            .I2(pwm_counter[3]), .I3(GND_net), .O(n6_adj_4974));   // verilog/pwm.v(21[8:24])
    defparam LessThan_744_i6_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 LessThan_744_i10_3_lut_3_lut (.I0(pwm_setpoint[5]), .I1(pwm_setpoint[6]), 
            .I2(pwm_counter[6]), .I3(GND_net), .O(n10_adj_4978));   // verilog/pwm.v(21[8:24])
    defparam LessThan_744_i10_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 encoder0_position_23__I_0_i680_3_lut (.I0(n992), .I1(n1045), 
            .I2(n1012), .I3(GND_net), .O(n1070));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i680_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i681_3_lut (.I0(n993), .I1(n1046), 
            .I2(n1012), .I3(GND_net), .O(n1071));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i681_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i678_3_lut (.I0(n990), .I1(n1043), 
            .I2(n1012), .I3(GND_net), .O(n1068));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i678_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i674_3_lut (.I0(n986), .I1(n1039), 
            .I2(n1012), .I3(GND_net), .O(n1064));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i674_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i675_3_lut (.I0(n987), .I1(n1040), 
            .I2(n1012), .I3(GND_net), .O(n1065));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i675_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i684_3_lut (.I0(n519), .I1(n1049), 
            .I2(n1012), .I3(GND_net), .O(n1074));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i684_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i683_3_lut (.I0(n995), .I1(n1048), 
            .I2(n1012), .I3(GND_net), .O(n1073));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i683_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mux_3363_i13_3_lut (.I0(encoder0_position[12]), .I1(n13_adj_4914), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n763));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam mux_3363_i13_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i19586_3_lut (.I0(n763), .I1(n1073), .I2(n1074), .I3(GND_net), 
            .O(n24729));
    defparam i19586_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i2_4_lut_adj_1695 (.I0(n1071), .I1(n1070), .I2(n24729), .I3(n1072), 
            .O(n34263));
    defparam i2_4_lut_adj_1695.LUT_INIT = 16'h8880;
    SB_LUT4 i5_4_lut_adj_1696 (.I0(n1065), .I1(n1064), .I2(n34263), .I3(n1068), 
            .O(n12_adj_5000));
    defparam i5_4_lut_adj_1696.LUT_INIT = 16'hfffe;
    SB_LUT4 i30637_4_lut (.I0(n1067), .I1(n12_adj_5000), .I2(n1066), .I3(n1069), 
            .O(n1090));
    defparam i30637_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 i14235_3_lut (.I0(\data_out_frame[13] [2]), .I1(setpoint[10]), 
            .I2(n14867), .I3(GND_net), .O(n19377));   // verilog/coms.v(127[12] 300[6])
    defparam i14235_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_23__I_0_i1482_3_lut (.I0(n1090), .I1(n6210), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(encoder0_position_scaled_23__N_34[13]));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1482_3_lut.LUT_INIT = 16'hc5c5;
    SB_LUT4 encoder0_position_23__I_0_i622_3_lut (.I0(n909), .I1(n962), 
            .I2(n934), .I3(GND_net), .O(n987));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i622_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14236_3_lut (.I0(\data_out_frame[13] [1]), .I1(setpoint[9]), 
            .I2(n14867), .I3(GND_net), .O(n19378));   // verilog/coms.v(127[12] 300[6])
    defparam i14236_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_23__I_0_i623_3_lut (.I0(n910), .I1(n963), 
            .I2(n934), .I3(GND_net), .O(n988));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i623_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i630_3_lut (.I0(n518), .I1(n970), 
            .I2(n934), .I3(GND_net), .O(n995));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i630_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14237_3_lut (.I0(\data_out_frame[13] [0]), .I1(setpoint[8]), 
            .I2(n14867), .I3(GND_net), .O(n19379));   // verilog/coms.v(127[12] 300[6])
    defparam i14237_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_23__I_0_i629_3_lut (.I0(n916), .I1(n969), 
            .I2(n934), .I3(GND_net), .O(n994));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i629_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i628_3_lut (.I0(n915), .I1(n968), 
            .I2(n934), .I3(GND_net), .O(n993));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i628_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mux_3363_i14_3_lut (.I0(encoder0_position[13]), .I1(n12_adj_4915), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n519));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam mux_3363_i14_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14238_3_lut (.I0(\data_out_frame[12] [7]), .I1(setpoint[23]), 
            .I2(n14867), .I3(GND_net), .O(n19380));   // verilog/coms.v(127[12] 300[6])
    defparam i14238_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_23__I_0_i626_3_lut (.I0(n913), .I1(n966), 
            .I2(n934), .I3(GND_net), .O(n991));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i626_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i627_3_lut (.I0(n914), .I1(n967), 
            .I2(n934), .I3(GND_net), .O(n992));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i627_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i625_3_lut (.I0(n912), .I1(n965), 
            .I2(n934), .I3(GND_net), .O(n990));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i625_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i621_3_lut (.I0(n908), .I1(n961), 
            .I2(n934), .I3(GND_net), .O(n986));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i621_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i624_3_lut (.I0(n911), .I1(n964), 
            .I2(n934), .I3(GND_net), .O(n989));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i624_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i19688_4_lut (.I0(n519), .I1(n993), .I2(n994), .I3(n995), 
            .O(n24833));
    defparam i19688_4_lut.LUT_INIT = 16'hfcec;
    SB_LUT4 i2_2_lut_adj_1697 (.I0(n989), .I1(n986), .I2(GND_net), .I3(GND_net), 
            .O(n8_adj_4998));
    defparam i2_2_lut_adj_1697.LUT_INIT = 16'heeee;
    SB_LUT4 i1_4_lut_adj_1698 (.I0(n990), .I1(n992), .I2(n991), .I3(n24833), 
            .O(n7_adj_4999));
    defparam i1_4_lut_adj_1698.LUT_INIT = 16'heaaa;
    SB_LUT4 i30621_4_lut (.I0(n988), .I1(n7_adj_4999), .I2(n987), .I3(n8_adj_4998), 
            .O(n1012));
    defparam i30621_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 i14239_3_lut (.I0(\data_out_frame[12] [6]), .I1(setpoint[22]), 
            .I2(n14867), .I3(GND_net), .O(n19381));   // verilog/coms.v(127[12] 300[6])
    defparam i14239_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_23__I_0_add_1202_20 (.CI(n28313), .I0(n1768), 
            .I1(VCC_net), .CO(n28314));
    SB_LUT4 encoder0_position_23__I_0_add_1202_19_lut (.I0(GND_net), .I1(n1769), 
            .I2(VCC_net), .I3(n28312), .O(n1822)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1202_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1202_19 (.CI(n28312), .I0(n1769), 
            .I1(VCC_net), .CO(n28313));
    SB_LUT4 encoder0_position_23__I_0_add_1202_18_lut (.I0(GND_net), .I1(n1770), 
            .I2(VCC_net), .I3(n28311), .O(n1823)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1202_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1202_18 (.CI(n28311), .I0(n1770), 
            .I1(VCC_net), .CO(n28312));
    SB_LUT4 add_672_10_lut (.I0(duty[8]), .I1(n37633), .I2(n17), .I3(n27833), 
            .O(pwm_setpoint_22__N_11[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_672_10_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 encoder0_position_23__I_0_add_1202_17_lut (.I0(GND_net), .I1(n1771), 
            .I2(VCC_net), .I3(n28310), .O(n1824)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1202_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1202_17 (.CI(n28310), .I0(n1771), 
            .I1(VCC_net), .CO(n28311));
    SB_LUT4 encoder0_position_23__I_0_add_1202_16_lut (.I0(GND_net), .I1(n1772), 
            .I2(VCC_net), .I3(n28309), .O(n1825)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1202_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1202_16 (.CI(n28309), .I0(n1772), 
            .I1(VCC_net), .CO(n28310));
    SB_LUT4 encoder0_position_23__I_0_add_1202_15_lut (.I0(GND_net), .I1(n1773), 
            .I2(VCC_net), .I3(n28308), .O(n1826)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1202_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1202_15 (.CI(n28308), .I0(n1773), 
            .I1(VCC_net), .CO(n28309));
    SB_LUT4 encoder0_position_23__I_0_add_1202_14_lut (.I0(GND_net), .I1(n1774), 
            .I2(VCC_net), .I3(n28307), .O(n1827)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1202_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1202_14 (.CI(n28307), .I0(n1774), 
            .I1(VCC_net), .CO(n28308));
    SB_CARRY add_672_10 (.CI(n27833), .I0(n37633), .I1(n17), .CO(n27834));
    SB_LUT4 encoder0_position_23__I_0_add_1202_13_lut (.I0(GND_net), .I1(n1775), 
            .I2(VCC_net), .I3(n28306), .O(n1828)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1202_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_672_9_lut (.I0(duty[7]), .I1(n37633), .I2(n18), .I3(n27832), 
            .O(pwm_setpoint_22__N_11[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_672_9_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY encoder0_position_23__I_0_add_1202_13 (.CI(n28306), .I0(n1775), 
            .I1(VCC_net), .CO(n28307));
    SB_LUT4 encoder0_position_23__I_0_add_1202_12_lut (.I0(GND_net), .I1(n1776), 
            .I2(VCC_net), .I3(n28305), .O(n1829)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1202_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1202_12 (.CI(n28305), .I0(n1776), 
            .I1(VCC_net), .CO(n28306));
    SB_LUT4 encoder0_position_23__I_0_add_1202_11_lut (.I0(GND_net), .I1(n1777), 
            .I2(VCC_net), .I3(n28304), .O(n1830)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1202_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1202_11 (.CI(n28304), .I0(n1777), 
            .I1(VCC_net), .CO(n28305));
    SB_LUT4 encoder0_position_23__I_0_add_1202_10_lut (.I0(GND_net), .I1(n1778), 
            .I2(VCC_net), .I3(n28303), .O(n1831)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1202_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1202_10 (.CI(n28303), .I0(n1778), 
            .I1(VCC_net), .CO(n28304));
    SB_LUT4 encoder0_position_23__I_0_add_1202_9_lut (.I0(GND_net), .I1(n1779), 
            .I2(VCC_net), .I3(n28302), .O(n1832)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1202_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1202_9 (.CI(n28302), .I0(n1779), 
            .I1(VCC_net), .CO(n28303));
    SB_LUT4 encoder0_position_23__I_0_add_1202_8_lut (.I0(GND_net), .I1(n1780), 
            .I2(VCC_net), .I3(n28301), .O(n1833)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1202_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1202_8 (.CI(n28301), .I0(n1780), 
            .I1(VCC_net), .CO(n28302));
    SB_LUT4 encoder0_position_23__I_0_add_1202_7_lut (.I0(GND_net), .I1(n1781), 
            .I2(GND_net), .I3(n28300), .O(n1834)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1202_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_672_9 (.CI(n27832), .I0(n37633), .I1(n18), .CO(n27833));
    SB_CARRY encoder0_position_23__I_0_add_1202_7 (.CI(n28300), .I0(n1781), 
            .I1(GND_net), .CO(n28301));
    SB_DFF read_61 (.Q(read), .C(CLK_c), .D(n35190));   // verilog/TinyFPGA_B.v(237[10] 265[6])
    SB_DFF ID_i0_i0 (.Q(ID[0]), .C(CLK_c), .D(n19057));   // verilog/TinyFPGA_B.v(237[10] 265[6])
    SB_LUT4 encoder0_position_23__I_0_add_1202_6_lut (.I0(GND_net), .I1(n1782), 
            .I2(GND_net), .I3(n28299), .O(n1835)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1202_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1202_6 (.CI(n28299), .I0(n1782), 
            .I1(GND_net), .CO(n28300));
    SB_LUT4 add_672_8_lut (.I0(duty[6]), .I1(n37633), .I2(n19), .I3(n27831), 
            .O(pwm_setpoint_22__N_11[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_672_8_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 encoder0_position_23__I_0_add_1202_5_lut (.I0(GND_net), .I1(n1783), 
            .I2(VCC_net), .I3(n28298), .O(n1836)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1202_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_25_23_lut (.I0(GND_net), .I1(delay_counter[21]), .I2(GND_net), 
            .I3(n27753), .O(n583)) /* synthesis syn_instantiated=1 */ ;
    defparam add_25_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1202_5 (.CI(n28298), .I0(n1783), 
            .I1(VCC_net), .CO(n28299));
    SB_CARRY add_25_9 (.CI(n27739), .I0(delay_counter[7]), .I1(GND_net), 
            .CO(n27740));
    SB_LUT4 encoder0_position_23__I_0_add_1202_4_lut (.I0(GND_net), .I1(n1784), 
            .I2(GND_net), .I3(n28297), .O(n1837)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1202_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_672_8 (.CI(n27831), .I0(n37633), .I1(n19), .CO(n27832));
    SB_CARRY encoder0_position_23__I_0_add_1202_4 (.CI(n28297), .I0(n1784), 
            .I1(GND_net), .CO(n28298));
    SB_LUT4 encoder0_position_23__I_0_i1481_3_lut (.I0(n1012), .I1(n6209), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(encoder0_position_scaled_23__N_34[14]));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1481_3_lut.LUT_INIT = 16'hc5c5;
    SB_LUT4 encoder0_position_23__I_0_add_1202_3_lut (.I0(GND_net), .I1(n1785), 
            .I2(VCC_net), .I3(n28296), .O(n1838)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1202_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1202_3 (.CI(n28296), .I0(n1785), 
            .I1(VCC_net), .CO(n28297));
    SB_LUT4 encoder0_position_23__I_0_i570_3_lut (.I0(n832), .I1(n885), 
            .I2(n856), .I3(GND_net), .O(n910));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i570_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_add_1202_2_lut (.I0(GND_net), .I1(n772), 
            .I2(GND_net), .I3(VCC_net), .O(n1839)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1202_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1202_2 (.CI(VCC_net), .I0(n772), 
            .I1(GND_net), .CO(n28296));
    SB_LUT4 encoder0_position_23__I_0_i569_3_lut (.I0(n831), .I1(n884), 
            .I2(n856), .I3(GND_net), .O(n909));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i569_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i571_3_lut (.I0(n833), .I1(n886), 
            .I2(n856), .I3(GND_net), .O(n911));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i571_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14240_3_lut (.I0(\data_out_frame[12] [5]), .I1(setpoint[21]), 
            .I2(n14867), .I3(GND_net), .O(n19382));   // verilog/coms.v(127[12] 300[6])
    defparam i14240_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_23__I_0_i576_3_lut (.I0(n517), .I1(n891), 
            .I2(n856), .I3(GND_net), .O(n916));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i576_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_add_1149_21_lut (.I0(GND_net), .I1(n1688), 
            .I2(VCC_net), .I3(n28295), .O(n1741)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1149_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_23__I_0_add_1149_20_lut (.I0(GND_net), .I1(n1689), 
            .I2(VCC_net), .I3(n28294), .O(n1742)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1149_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1149_20 (.CI(n28294), .I0(n1689), 
            .I1(VCC_net), .CO(n28295));
    SB_LUT4 encoder0_position_23__I_0_add_1149_19_lut (.I0(GND_net), .I1(n1690), 
            .I2(VCC_net), .I3(n28293), .O(n1743)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1149_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1149_19 (.CI(n28293), .I0(n1690), 
            .I1(VCC_net), .CO(n28294));
    SB_LUT4 encoder0_position_23__I_0_add_1149_18_lut (.I0(GND_net), .I1(n1691), 
            .I2(VCC_net), .I3(n28292), .O(n1744)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1149_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1149_18 (.CI(n28292), .I0(n1691), 
            .I1(VCC_net), .CO(n28293));
    SB_LUT4 encoder0_position_23__I_0_i575_3_lut (.I0(n837), .I1(n890), 
            .I2(n856), .I3(GND_net), .O(n915));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i575_3_lut.LUT_INIT = 16'hacac;
    SB_DFFESR delay_counter_i0_i26 (.Q(delay_counter[26]), .C(CLK_c), .E(n5410), 
            .D(n578), .R(n18963));   // verilog/TinyFPGA_B.v(237[10] 265[6])
    SB_LUT4 encoder0_position_23__I_0_add_1149_17_lut (.I0(GND_net), .I1(n1692), 
            .I2(VCC_net), .I3(n28291), .O(n1745)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1149_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_4_inv_0_i2_1_lut (.I0(duty[1]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n24));   // verilog/TinyFPGA_B.v(106[23:28])
    defparam unary_minus_4_inv_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY encoder0_position_23__I_0_add_1149_17 (.CI(n28291), .I0(n1692), 
            .I1(VCC_net), .CO(n28292));
    SB_LUT4 encoder0_position_23__I_0_add_1149_16_lut (.I0(GND_net), .I1(n1693), 
            .I2(VCC_net), .I3(n28290), .O(n1746)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1149_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_23__I_0_i409_3_lut_4_lut (.I0(n2), .I1(encoder0_position[23]), 
            .I2(n619), .I3(n6024), .O(n674));
    defparam encoder0_position_23__I_0_i409_3_lut_4_lut.LUT_INIT = 16'h8f80;
    SB_LUT4 mux_75_i1_3_lut_4_lut (.I0(n17355), .I1(control_mode[1]), .I2(motor_state_23__N_82[0]), 
            .I3(encoder0_position_scaled[0]), .O(motor_state[0]));   // verilog/TinyFPGA_B.v(165[5:22])
    defparam mux_75_i1_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 mux_75_i2_3_lut_4_lut (.I0(n17355), .I1(control_mode[1]), .I2(motor_state_23__N_82[1]), 
            .I3(encoder0_position_scaled[1]), .O(motor_state[1]));   // verilog/TinyFPGA_B.v(165[5:22])
    defparam mux_75_i2_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 mux_75_i3_3_lut_4_lut (.I0(n17355), .I1(control_mode[1]), .I2(motor_state_23__N_82[2]), 
            .I3(encoder0_position_scaled[2]), .O(motor_state[2]));   // verilog/TinyFPGA_B.v(165[5:22])
    defparam mux_75_i3_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 mux_75_i4_3_lut_4_lut (.I0(n17355), .I1(control_mode[1]), .I2(motor_state_23__N_82[3]), 
            .I3(encoder0_position_scaled[3]), .O(motor_state[3]));   // verilog/TinyFPGA_B.v(165[5:22])
    defparam mux_75_i4_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 add_25_8_lut (.I0(GND_net), .I1(delay_counter[6]), .I2(GND_net), 
            .I3(n27738), .O(n598)) /* synthesis syn_instantiated=1 */ ;
    defparam add_25_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1149_16 (.CI(n28290), .I0(n1693), 
            .I1(VCC_net), .CO(n28291));
    SB_LUT4 mux_75_i5_3_lut_4_lut (.I0(n17355), .I1(control_mode[1]), .I2(motor_state_23__N_82[4]), 
            .I3(encoder0_position_scaled[4]), .O(motor_state[4]));   // verilog/TinyFPGA_B.v(165[5:22])
    defparam mux_75_i5_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 encoder0_position_23__I_0_add_1149_15_lut (.I0(GND_net), .I1(n1694), 
            .I2(VCC_net), .I3(n28289), .O(n1747)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1149_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mux_75_i6_3_lut_4_lut (.I0(n17355), .I1(control_mode[1]), .I2(motor_state_23__N_82[5]), 
            .I3(encoder0_position_scaled[5]), .O(motor_state[5]));   // verilog/TinyFPGA_B.v(165[5:22])
    defparam mux_75_i6_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 encoder0_position_23__I_0_i574_3_lut (.I0(n836), .I1(n889), 
            .I2(n856), .I3(GND_net), .O(n914));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i574_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_23__I_0_add_1149_15 (.CI(n28289), .I0(n1694), 
            .I1(VCC_net), .CO(n28290));
    SB_LUT4 mux_75_i7_3_lut_4_lut (.I0(n17355), .I1(control_mode[1]), .I2(motor_state_23__N_82[6]), 
            .I3(encoder0_position_scaled[6]), .O(motor_state[6]));   // verilog/TinyFPGA_B.v(165[5:22])
    defparam mux_75_i7_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_CARRY add_25_3 (.CI(n27733), .I0(delay_counter[1]), .I1(GND_net), 
            .CO(n27734));
    SB_LUT4 encoder0_position_23__I_0_add_1149_14_lut (.I0(GND_net), .I1(n1695), 
            .I2(VCC_net), .I3(n28288), .O(n1748)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1149_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mux_75_i8_3_lut_4_lut (.I0(n17355), .I1(control_mode[1]), .I2(motor_state_23__N_82[7]), 
            .I3(encoder0_position_scaled[7]), .O(motor_state[7]));   // verilog/TinyFPGA_B.v(165[5:22])
    defparam mux_75_i8_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_CARRY encoder0_position_23__I_0_add_1149_14 (.CI(n28288), .I0(n1695), 
            .I1(VCC_net), .CO(n28289));
    SB_LUT4 mux_75_i9_3_lut_4_lut (.I0(n17355), .I1(control_mode[1]), .I2(motor_state_23__N_82[8]), 
            .I3(encoder0_position_scaled[8]), .O(motor_state[8]));   // verilog/TinyFPGA_B.v(165[5:22])
    defparam mux_75_i9_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_CARRY add_25_8 (.CI(n27738), .I0(delay_counter[6]), .I1(GND_net), 
            .CO(n27739));
    SB_LUT4 encoder0_position_23__I_0_add_1149_13_lut (.I0(GND_net), .I1(n1696), 
            .I2(VCC_net), .I3(n28287), .O(n1749)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1149_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mux_3363_i15_3_lut (.I0(encoder0_position[14]), .I1(n11_adj_4916), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n518));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam mux_3363_i15_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_23__I_0_add_1149_13 (.CI(n28287), .I0(n1696), 
            .I1(VCC_net), .CO(n28288));
    SB_LUT4 i29594_2_lut_4_lut (.I0(pwm_counter[16]), .I1(pwm_setpoint[16]), 
            .I2(pwm_counter[7]), .I3(pwm_setpoint[7]), .O(n36349));
    defparam i29594_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 encoder0_position_23__I_0_add_1149_12_lut (.I0(GND_net), .I1(n1697), 
            .I2(VCC_net), .I3(n28286), .O(n1750)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1149_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1149_12 (.CI(n28286), .I0(n1697), 
            .I1(VCC_net), .CO(n28287));
    SB_LUT4 encoder0_position_23__I_0_add_1149_11_lut (.I0(GND_net), .I1(n1698), 
            .I2(VCC_net), .I3(n28285), .O(n1751)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1149_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1149_11 (.CI(n28285), .I0(n1698), 
            .I1(VCC_net), .CO(n28286));
    SB_LUT4 encoder0_position_23__I_0_add_1149_10_lut (.I0(GND_net), .I1(n1699), 
            .I2(VCC_net), .I3(n28284), .O(n1752)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1149_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1149_10 (.CI(n28284), .I0(n1699), 
            .I1(VCC_net), .CO(n28285));
    SB_LUT4 encoder0_position_23__I_0_add_1149_9_lut (.I0(GND_net), .I1(n1700), 
            .I2(VCC_net), .I3(n28283), .O(n1753)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1149_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1149_9 (.CI(n28283), .I0(n1700), 
            .I1(VCC_net), .CO(n28284));
    SB_LUT4 encoder0_position_23__I_0_add_1149_8_lut (.I0(GND_net), .I1(n1701), 
            .I2(VCC_net), .I3(n28282), .O(n1754)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1149_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1149_8 (.CI(n28282), .I0(n1701), 
            .I1(VCC_net), .CO(n28283));
    SB_LUT4 encoder0_position_23__I_0_add_1149_7_lut (.I0(GND_net), .I1(n1702), 
            .I2(GND_net), .I3(n28281), .O(n1755)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1149_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1149_7 (.CI(n28281), .I0(n1702), 
            .I1(GND_net), .CO(n28282));
    SB_LUT4 encoder0_position_23__I_0_add_1149_6_lut (.I0(GND_net), .I1(n1703), 
            .I2(GND_net), .I3(n28280), .O(n1756)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1149_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1149_6 (.CI(n28280), .I0(n1703), 
            .I1(GND_net), .CO(n28281));
    SB_LUT4 encoder0_position_23__I_0_add_1149_5_lut (.I0(GND_net), .I1(n1704), 
            .I2(VCC_net), .I3(n28279), .O(n1757)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1149_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1149_5 (.CI(n28279), .I0(n1704), 
            .I1(VCC_net), .CO(n28280));
    SB_LUT4 encoder0_position_23__I_0_add_1149_4_lut (.I0(GND_net), .I1(n1705), 
            .I2(GND_net), .I3(n28278), .O(n1758)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1149_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1149_4 (.CI(n28278), .I0(n1705), 
            .I1(GND_net), .CO(n28279));
    SB_LUT4 encoder0_position_23__I_0_add_1149_3_lut (.I0(GND_net), .I1(n1706), 
            .I2(VCC_net), .I3(n28277), .O(n1759)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1149_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1149_3 (.CI(n28277), .I0(n1706), 
            .I1(VCC_net), .CO(n28278));
    SB_LUT4 encoder0_position_23__I_0_add_1149_2_lut (.I0(GND_net), .I1(n771_adj_4968), 
            .I2(GND_net), .I3(VCC_net), .O(n1760)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1149_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1149_2 (.CI(VCC_net), .I0(n771_adj_4968), 
            .I1(GND_net), .CO(n28277));
    SB_LUT4 encoder0_position_23__I_0_add_1096_20_lut (.I0(GND_net), .I1(n1610), 
            .I2(VCC_net), .I3(n28276), .O(n1663)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1096_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_23__I_0_add_1096_19_lut (.I0(GND_net), .I1(n1611), 
            .I2(VCC_net), .I3(n28275), .O(n1664)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1096_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1096_19 (.CI(n28275), .I0(n1611), 
            .I1(VCC_net), .CO(n28276));
    SB_LUT4 encoder0_position_23__I_0_add_1096_18_lut (.I0(GND_net), .I1(n1612), 
            .I2(VCC_net), .I3(n28274), .O(n1665)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1096_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1096_18 (.CI(n28274), .I0(n1612), 
            .I1(VCC_net), .CO(n28275));
    SB_LUT4 mux_75_i10_3_lut_4_lut (.I0(n17355), .I1(control_mode[1]), .I2(motor_state_23__N_82[9]), 
            .I3(encoder0_position_scaled[9]), .O(motor_state[9]));   // verilog/TinyFPGA_B.v(165[5:22])
    defparam mux_75_i10_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 mux_75_i11_3_lut_4_lut (.I0(n17355), .I1(control_mode[1]), .I2(motor_state_23__N_82[10]), 
            .I3(encoder0_position_scaled[10]), .O(motor_state[10]));   // verilog/TinyFPGA_B.v(165[5:22])
    defparam mux_75_i11_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 encoder0_position_23__I_0_i572_3_lut (.I0(n834), .I1(n887), 
            .I2(n856), .I3(GND_net), .O(n912));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i572_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i568_3_lut (.I0(n830), .I1(n883), 
            .I2(n856), .I3(GND_net), .O(n908));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i568_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i573_3_lut (.I0(n835), .I1(n888), 
            .I2(n856), .I3(GND_net), .O(n913));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i573_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i19690_4_lut (.I0(n518), .I1(n914), .I2(n915), .I3(n916), 
            .O(n24835));
    defparam i19690_4_lut.LUT_INIT = 16'hfcec;
    SB_LUT4 i2_4_lut_adj_1699 (.I0(n913), .I1(n908), .I2(n912), .I3(n24835), 
            .O(n7_adj_5065));
    defparam i2_4_lut_adj_1699.LUT_INIT = 16'heccc;
    SB_LUT4 i30606_4_lut (.I0(n7_adj_5065), .I1(n911), .I2(n909), .I3(n910), 
            .O(n934));
    defparam i30606_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 encoder0_position_23__I_0_i1480_3_lut (.I0(n934), .I1(n6208), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(encoder0_position_scaled_23__N_34[15]));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1480_3_lut.LUT_INIT = 16'hc5c5;
    SB_LUT4 encoder0_position_23__I_0_i516_3_lut (.I0(n753), .I1(n806), 
            .I2(n778), .I3(GND_net), .O(n831));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i516_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i517_3_lut (.I0(n754), .I1(n807), 
            .I2(n778), .I3(GND_net), .O(n832));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i517_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 unary_minus_4_inv_0_i3_1_lut (.I0(duty[2]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n23));   // verilog/TinyFPGA_B.v(106[23:28])
    defparam unary_minus_4_inv_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i19437_3_lut (.I0(n517), .I1(n836), .I2(n837), .I3(GND_net), 
            .O(n24577));
    defparam i19437_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i2_4_lut_adj_1700 (.I0(n834), .I1(n833), .I2(n24577), .I3(n835), 
            .O(n34039));
    defparam i2_4_lut_adj_1700.LUT_INIT = 16'h8880;
    SB_LUT4 unary_minus_4_inv_0_i4_1_lut (.I0(duty[3]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n22));   // verilog/TinyFPGA_B.v(106[23:28])
    defparam unary_minus_4_inv_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i30592_4_lut (.I0(n34039), .I1(n830), .I2(n832), .I3(n831), 
            .O(n856));
    defparam i30592_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 encoder0_position_23__I_0_i1479_3_lut (.I0(n856), .I1(n6207), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(encoder0_position_scaled_23__N_34[16]));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1479_3_lut.LUT_INIT = 16'hc5c5;
    SB_LUT4 encoder0_position_23__I_0_i1478_3_lut (.I0(n778), .I1(n6206), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(encoder0_position_scaled_23__N_34[17]));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1478_3_lut.LUT_INIT = 16'hc5c5;
    SB_LUT4 encoder0_position_23__I_0_i1477_3_lut (.I0(n700), .I1(n6205), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(encoder0_position_scaled_23__N_34[18]));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1477_3_lut.LUT_INIT = 16'hc5c5;
    SB_LUT4 mux_75_i12_3_lut_4_lut (.I0(n17355), .I1(control_mode[1]), .I2(motor_state_23__N_82[11]), 
            .I3(encoder0_position_scaled[11]), .O(motor_state[11]));   // verilog/TinyFPGA_B.v(165[5:22])
    defparam mux_75_i12_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 mux_77_i2_4_lut (.I0(encoder1_position[1]), .I1(displacement[1]), 
            .I2(n15_adj_4934), .I3(n15_adj_4940), .O(motor_state_23__N_82[1]));   // verilog/TinyFPGA_B.v(166[5] 168[10])
    defparam mux_77_i2_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 LessThan_744_i12_3_lut_3_lut (.I0(pwm_setpoint[7]), .I1(pwm_setpoint[16]), 
            .I2(pwm_counter[16]), .I3(GND_net), .O(n12_adj_4980));   // verilog/pwm.v(21[8:24])
    defparam LessThan_744_i12_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i29828_2_lut_3_lut (.I0(n62), .I1(delay_counter[31]), .I2(\ID_READOUT_FSM.state [0]), 
            .I3(GND_net), .O(n36275));
    defparam i29828_2_lut_3_lut.LUT_INIT = 16'hf2f2;
    SB_LUT4 i14241_3_lut (.I0(\data_out_frame[12] [4]), .I1(setpoint[20]), 
            .I2(n14867), .I3(GND_net), .O(n19383));   // verilog/coms.v(127[12] 300[6])
    defparam i14241_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_75_i13_3_lut_4_lut (.I0(n17355), .I1(control_mode[1]), .I2(motor_state_23__N_82[12]), 
            .I3(encoder0_position_scaled[12]), .O(motor_state[12]));   // verilog/TinyFPGA_B.v(165[5:22])
    defparam mux_75_i13_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 mux_75_i14_3_lut_4_lut (.I0(n17355), .I1(control_mode[1]), .I2(motor_state_23__N_82[13]), 
            .I3(encoder0_position_scaled[13]), .O(motor_state[13]));   // verilog/TinyFPGA_B.v(165[5:22])
    defparam mux_75_i14_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 mux_75_i15_3_lut_4_lut (.I0(n17355), .I1(control_mode[1]), .I2(motor_state_23__N_82[14]), 
            .I3(encoder0_position_scaled[14]), .O(motor_state[14]));   // verilog/TinyFPGA_B.v(165[5:22])
    defparam mux_75_i15_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 i14242_3_lut (.I0(\data_out_frame[12] [3]), .I1(setpoint[19]), 
            .I2(n14867), .I3(GND_net), .O(n19384));   // verilog/coms.v(127[12] 300[6])
    defparam i14242_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14243_3_lut (.I0(\data_out_frame[12] [2]), .I1(setpoint[18]), 
            .I2(n14867), .I3(GND_net), .O(n19385));   // verilog/coms.v(127[12] 300[6])
    defparam i14243_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_75_i16_3_lut_4_lut (.I0(n17355), .I1(control_mode[1]), .I2(motor_state_23__N_82[15]), 
            .I3(encoder0_position_scaled[15]), .O(motor_state[15]));   // verilog/TinyFPGA_B.v(165[5:22])
    defparam mux_75_i16_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 i14244_3_lut (.I0(\data_out_frame[12] [1]), .I1(setpoint[17]), 
            .I2(n14867), .I3(GND_net), .O(n19386));   // verilog/coms.v(127[12] 300[6])
    defparam i14244_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14245_3_lut (.I0(\data_out_frame[12] [0]), .I1(setpoint[16]), 
            .I2(n14867), .I3(GND_net), .O(n19387));   // verilog/coms.v(127[12] 300[6])
    defparam i14245_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14246_3_lut (.I0(\data_out_frame[11] [7]), .I1(encoder1_position[7]), 
            .I2(n14867), .I3(GND_net), .O(n19388));   // verilog/coms.v(127[12] 300[6])
    defparam i14246_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14247_3_lut (.I0(\data_out_frame[11] [6]), .I1(encoder1_position[6]), 
            .I2(n14867), .I3(GND_net), .O(n19389));   // verilog/coms.v(127[12] 300[6])
    defparam i14247_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_75_i17_3_lut_4_lut (.I0(n17355), .I1(control_mode[1]), .I2(motor_state_23__N_82[16]), 
            .I3(encoder0_position_scaled[16]), .O(motor_state[16]));   // verilog/TinyFPGA_B.v(165[5:22])
    defparam mux_75_i17_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 mux_75_i18_3_lut_4_lut (.I0(n17355), .I1(control_mode[1]), .I2(motor_state_23__N_82[17]), 
            .I3(encoder0_position_scaled[17]), .O(motor_state[17]));   // verilog/TinyFPGA_B.v(165[5:22])
    defparam mux_75_i18_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 i14248_3_lut (.I0(\data_out_frame[11] [5]), .I1(encoder1_position[5]), 
            .I2(n14867), .I3(GND_net), .O(n19390));   // verilog/coms.v(127[12] 300[6])
    defparam i14248_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14249_3_lut (.I0(\data_out_frame[11] [4]), .I1(encoder1_position[4]), 
            .I2(n14867), .I3(GND_net), .O(n19391));   // verilog/coms.v(127[12] 300[6])
    defparam i14249_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14250_3_lut (.I0(\data_out_frame[11] [3]), .I1(encoder1_position[3]), 
            .I2(n14867), .I3(GND_net), .O(n19392));   // verilog/coms.v(127[12] 300[6])
    defparam i14250_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14251_3_lut (.I0(\data_out_frame[11] [2]), .I1(encoder1_position[2]), 
            .I2(n14867), .I3(GND_net), .O(n19393));   // verilog/coms.v(127[12] 300[6])
    defparam i14251_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14252_3_lut (.I0(\data_out_frame[11] [1]), .I1(encoder1_position[1]), 
            .I2(n14867), .I3(GND_net), .O(n19394));   // verilog/coms.v(127[12] 300[6])
    defparam i14252_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14253_3_lut (.I0(\data_out_frame[11] [0]), .I1(encoder1_position[0]), 
            .I2(n14867), .I3(GND_net), .O(n19395));   // verilog/coms.v(127[12] 300[6])
    defparam i14253_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_75_i19_3_lut_4_lut (.I0(n17355), .I1(control_mode[1]), .I2(motor_state_23__N_82[18]), 
            .I3(encoder0_position_scaled[18]), .O(motor_state[18]));   // verilog/TinyFPGA_B.v(165[5:22])
    defparam mux_75_i19_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 encoder1_position_23__I_0_inv_0_i11_1_lut (.I0(encoder0_position_scaled[10]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n15_adj_4955));   // verilog/TinyFPGA_B.v(202[21:65])
    defparam encoder1_position_23__I_0_inv_0_i11_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i14254_3_lut (.I0(\data_out_frame[10] [7]), .I1(encoder1_position[15]), 
            .I2(n14867), .I3(GND_net), .O(n19396));   // verilog/coms.v(127[12] 300[6])
    defparam i14254_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder1_position_23__I_0_inv_0_i12_1_lut (.I0(encoder0_position_scaled[11]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n14_adj_4954));   // verilog/TinyFPGA_B.v(202[21:65])
    defparam encoder1_position_23__I_0_inv_0_i12_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mux_75_i20_3_lut_4_lut (.I0(n17355), .I1(control_mode[1]), .I2(motor_state_23__N_82[19]), 
            .I3(encoder0_position_scaled[19]), .O(motor_state[19]));   // verilog/TinyFPGA_B.v(165[5:22])
    defparam mux_75_i20_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 encoder1_position_23__I_0_inv_0_i13_1_lut (.I0(encoder0_position_scaled[12]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n13_adj_4953));   // verilog/TinyFPGA_B.v(202[21:65])
    defparam encoder1_position_23__I_0_inv_0_i13_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i14255_3_lut (.I0(\data_out_frame[10] [6]), .I1(encoder1_position[14]), 
            .I2(n14867), .I3(GND_net), .O(n19397));   // verilog/coms.v(127[12] 300[6])
    defparam i14255_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14256_3_lut (.I0(\data_out_frame[10] [5]), .I1(encoder1_position[13]), 
            .I2(n14867), .I3(GND_net), .O(n19398));   // verilog/coms.v(127[12] 300[6])
    defparam i14256_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_77_i3_4_lut (.I0(encoder1_position[2]), .I1(displacement[2]), 
            .I2(n15_adj_4934), .I3(n15_adj_4940), .O(motor_state_23__N_82[2]));   // verilog/TinyFPGA_B.v(166[5] 168[10])
    defparam mux_77_i3_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i14257_3_lut (.I0(\data_out_frame[10] [4]), .I1(encoder1_position[12]), 
            .I2(n14867), .I3(GND_net), .O(n19399));   // verilog/coms.v(127[12] 300[6])
    defparam i14257_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_744_i8_3_lut_3_lut (.I0(pwm_setpoint[4]), .I1(pwm_setpoint[8]), 
            .I2(pwm_counter[8]), .I3(GND_net), .O(n8_adj_4976));   // verilog/pwm.v(21[8:24])
    defparam LessThan_744_i8_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i14258_3_lut (.I0(\data_out_frame[10] [3]), .I1(encoder1_position[11]), 
            .I2(n14867), .I3(GND_net), .O(n19400));   // verilog/coms.v(127[12] 300[6])
    defparam i14258_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_75_i21_3_lut_4_lut (.I0(n17355), .I1(control_mode[1]), .I2(motor_state_23__N_82[20]), 
            .I3(encoder0_position_scaled[20]), .O(motor_state[20]));   // verilog/TinyFPGA_B.v(165[5:22])
    defparam mux_75_i21_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 i14259_3_lut (.I0(\data_out_frame[10] [2]), .I1(encoder1_position[10]), 
            .I2(n14867), .I3(GND_net), .O(n19401));   // verilog/coms.v(127[12] 300[6])
    defparam i14259_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_23__I_0_add_1096_17_lut (.I0(GND_net), .I1(n1613), 
            .I2(VCC_net), .I3(n28273), .O(n1666)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1096_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1096_17 (.CI(n28273), .I0(n1613), 
            .I1(VCC_net), .CO(n28274));
    SB_LUT4 encoder0_position_23__I_0_add_1096_16_lut (.I0(GND_net), .I1(n1614), 
            .I2(VCC_net), .I3(n28272), .O(n1667)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1096_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1096_16 (.CI(n28272), .I0(n1614), 
            .I1(VCC_net), .CO(n28273));
    SB_LUT4 encoder0_position_23__I_0_add_1096_15_lut (.I0(GND_net), .I1(n1615), 
            .I2(VCC_net), .I3(n28271), .O(n1668)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1096_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1096_15 (.CI(n28271), .I0(n1615), 
            .I1(VCC_net), .CO(n28272));
    SB_LUT4 encoder1_position_23__I_0_inv_0_i14_1_lut (.I0(encoder0_position_scaled[13]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n12_adj_4952));   // verilog/TinyFPGA_B.v(202[21:65])
    defparam encoder1_position_23__I_0_inv_0_i14_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_23__I_0_add_1096_14_lut (.I0(GND_net), .I1(n1616), 
            .I2(VCC_net), .I3(n28270), .O(n1669)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1096_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1096_14 (.CI(n28270), .I0(n1616), 
            .I1(VCC_net), .CO(n28271));
    SB_LUT4 encoder0_position_23__I_0_add_1096_13_lut (.I0(GND_net), .I1(n1617), 
            .I2(VCC_net), .I3(n28269), .O(n1670)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1096_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1096_13 (.CI(n28269), .I0(n1617), 
            .I1(VCC_net), .CO(n28270));
    SB_LUT4 encoder0_position_23__I_0_add_1096_12_lut (.I0(GND_net), .I1(n1618), 
            .I2(VCC_net), .I3(n28268), .O(n1671)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1096_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1096_12 (.CI(n28268), .I0(n1618), 
            .I1(VCC_net), .CO(n28269));
    SB_LUT4 encoder0_position_23__I_0_add_1096_11_lut (.I0(GND_net), .I1(n1619), 
            .I2(VCC_net), .I3(n28267), .O(n1672)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1096_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mux_75_i22_3_lut_4_lut (.I0(n17355), .I1(control_mode[1]), .I2(motor_state_23__N_82[21]), 
            .I3(encoder0_position_scaled[22]), .O(motor_state[21]));   // verilog/TinyFPGA_B.v(165[5:22])
    defparam mux_75_i22_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_CARRY encoder0_position_23__I_0_add_1096_11 (.CI(n28267), .I0(n1619), 
            .I1(VCC_net), .CO(n28268));
    SB_CARRY add_25_23 (.CI(n27753), .I0(delay_counter[21]), .I1(GND_net), 
            .CO(n27754));
    SB_LUT4 mux_77_i4_4_lut (.I0(encoder1_position[3]), .I1(displacement[3]), 
            .I2(n15_adj_4934), .I3(n15_adj_4940), .O(motor_state_23__N_82[3]));   // verilog/TinyFPGA_B.v(166[5] 168[10])
    defparam mux_77_i4_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 add_672_7_lut (.I0(duty[5]), .I1(n37633), .I2(n20), .I3(n27830), 
            .O(pwm_setpoint_22__N_11[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_672_7_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 i29608_2_lut_4_lut (.I0(pwm_counter[8]), .I1(pwm_setpoint[8]), 
            .I2(pwm_counter[4]), .I3(pwm_setpoint[4]), .O(n36363));
    defparam i29608_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 mux_75_i23_3_lut_4_lut (.I0(n17355), .I1(control_mode[1]), .I2(motor_state_23__N_82[22]), 
            .I3(encoder0_position_scaled[22]), .O(motor_state[22]));   // verilog/TinyFPGA_B.v(165[5:22])
    defparam mux_75_i23_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 unary_minus_4_inv_0_i22_1_lut (.I0(duty[21]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n4_adj_4884));   // verilog/TinyFPGA_B.v(106[23:28])
    defparam unary_minus_4_inv_0_i22_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i14260_3_lut (.I0(\data_out_frame[10] [1]), .I1(encoder1_position[9]), 
            .I2(n14867), .I3(GND_net), .O(n19402));   // verilog/coms.v(127[12] 300[6])
    defparam i14260_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14261_3_lut (.I0(\data_out_frame[10] [0]), .I1(encoder1_position[8]), 
            .I2(n14867), .I3(GND_net), .O(n19403));   // verilog/coms.v(127[12] 300[6])
    defparam i14261_3_lut.LUT_INIT = 16'hcaca;
    SB_DFFESR delay_counter_i0_i25 (.Q(delay_counter[25]), .C(CLK_c), .E(n5410), 
            .D(n579), .R(n18963));   // verilog/TinyFPGA_B.v(237[10] 265[6])
    SB_LUT4 i14262_3_lut (.I0(\data_out_frame[9] [7]), .I1(encoder1_position[23]), 
            .I2(n14867), .I3(GND_net), .O(n19404));   // verilog/coms.v(127[12] 300[6])
    defparam i14262_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 unary_minus_4_inv_0_i23_1_lut (.I0(duty[22]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n3));   // verilog/TinyFPGA_B.v(106[23:28])
    defparam unary_minus_4_inv_0_i23_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i14263_3_lut (.I0(\data_out_frame[9] [6]), .I1(encoder1_position[22]), 
            .I2(n14867), .I3(GND_net), .O(n19405));   // verilog/coms.v(127[12] 300[6])
    defparam i14263_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14264_3_lut (.I0(\data_out_frame[9] [5]), .I1(encoder1_position[21]), 
            .I2(n14867), .I3(GND_net), .O(n19406));   // verilog/coms.v(127[12] 300[6])
    defparam i14264_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_75_i24_3_lut_4_lut (.I0(n17355), .I1(control_mode[1]), .I2(motor_state_23__N_82[23]), 
            .I3(encoder0_position_scaled[22]), .O(motor_state[23]));   // verilog/TinyFPGA_B.v(165[5:22])
    defparam mux_75_i24_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 mux_77_i5_4_lut (.I0(encoder1_position[4]), .I1(displacement[4]), 
            .I2(n15_adj_4934), .I3(n15_adj_4940), .O(motor_state_23__N_82[4]));   // verilog/TinyFPGA_B.v(166[5] 168[10])
    defparam mux_77_i5_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 encoder0_position_23__I_0_add_1096_10_lut (.I0(GND_net), .I1(n1620), 
            .I2(VCC_net), .I3(n28266), .O(n1673)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1096_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1096_10 (.CI(n28266), .I0(n1620), 
            .I1(VCC_net), .CO(n28267));
    SB_DFF \ID_READOUT_FSM.state__i1  (.Q(\ID_READOUT_FSM.state [1]), .C(CLK_c), 
           .D(n17_adj_4895));   // verilog/TinyFPGA_B.v(237[10] 265[6])
    SB_DFF \ID_READOUT_FSM.state__i0  (.Q(\ID_READOUT_FSM.state [0]), .C(CLK_c), 
           .D(n31783));   // verilog/TinyFPGA_B.v(237[10] 265[6])
    SB_DFF ID_i0_i7 (.Q(ID[7]), .C(CLK_c), .D(n19600));   // verilog/TinyFPGA_B.v(237[10] 265[6])
    SB_DFF ID_i0_i6 (.Q(ID[6]), .C(CLK_c), .D(n19599));   // verilog/TinyFPGA_B.v(237[10] 265[6])
    SB_DFF ID_i0_i5 (.Q(ID[5]), .C(CLK_c), .D(n19598));   // verilog/TinyFPGA_B.v(237[10] 265[6])
    SB_DFF ID_i0_i4 (.Q(ID[4]), .C(CLK_c), .D(n19597));   // verilog/TinyFPGA_B.v(237[10] 265[6])
    SB_DFF ID_i0_i3 (.Q(ID[3]), .C(CLK_c), .D(n19596));   // verilog/TinyFPGA_B.v(237[10] 265[6])
    SB_DFF ID_i0_i2 (.Q(ID[2]), .C(CLK_c), .D(n19595));   // verilog/TinyFPGA_B.v(237[10] 265[6])
    SB_DFF ID_i0_i1 (.Q(ID[1]), .C(CLK_c), .D(n19594));   // verilog/TinyFPGA_B.v(237[10] 265[6])
    SB_CARRY add_672_7 (.CI(n27830), .I0(n37633), .I1(n20), .CO(n27831));
    SB_LUT4 encoder0_position_23__I_0_add_1096_9_lut (.I0(GND_net), .I1(n1621), 
            .I2(VCC_net), .I3(n28265), .O(n1674)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1096_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1096_9 (.CI(n28265), .I0(n1621), 
            .I1(VCC_net), .CO(n28266));
    SB_LUT4 encoder0_position_23__I_0_add_1096_8_lut (.I0(GND_net), .I1(n1622), 
            .I2(VCC_net), .I3(n28264), .O(n1675)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1096_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i14265_3_lut (.I0(\data_out_frame[9] [4]), .I1(encoder1_position[20]), 
            .I2(n14867), .I3(GND_net), .O(n19407));   // verilog/coms.v(127[12] 300[6])
    defparam i14265_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder1_position_23__I_0_inv_0_i15_1_lut (.I0(encoder0_position_scaled[14]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n11_adj_4951));   // verilog/TinyFPGA_B.v(202[21:65])
    defparam encoder1_position_23__I_0_inv_0_i15_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder1_position_23__I_0_inv_0_i16_1_lut (.I0(encoder0_position_scaled[15]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n10_adj_4950));   // verilog/TinyFPGA_B.v(202[21:65])
    defparam encoder1_position_23__I_0_inv_0_i16_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mux_77_i6_4_lut (.I0(encoder1_position[5]), .I1(displacement[5]), 
            .I2(n15_adj_4934), .I3(n15_adj_4940), .O(motor_state_23__N_82[5]));   // verilog/TinyFPGA_B.v(166[5] 168[10])
    defparam mux_77_i6_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i14266_3_lut (.I0(\data_out_frame[9] [3]), .I1(encoder1_position[19]), 
            .I2(n14867), .I3(GND_net), .O(n19408));   // verilog/coms.v(127[12] 300[6])
    defparam i14266_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_3_lut (.I0(\ID_READOUT_FSM.state [0]), .I1(\ID_READOUT_FSM.state [1]), 
            .I2(n17358), .I3(GND_net), .O(n17359));   // verilog/TinyFPGA_B.v(255[7:11])
    defparam i1_2_lut_3_lut.LUT_INIT = 16'hfbfb;
    SB_CARRY encoder0_position_23__I_0_add_1096_8 (.CI(n28264), .I0(n1622), 
            .I1(VCC_net), .CO(n28265));
    SB_LUT4 i14267_3_lut (.I0(\data_out_frame[9] [2]), .I1(encoder1_position[18]), 
            .I2(n14867), .I3(GND_net), .O(n19409));   // verilog/coms.v(127[12] 300[6])
    defparam i14267_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14268_3_lut (.I0(\data_out_frame[9] [1]), .I1(encoder1_position[17]), 
            .I2(n14867), .I3(GND_net), .O(n19410));   // verilog/coms.v(127[12] 300[6])
    defparam i14268_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14269_3_lut (.I0(\data_out_frame[9] [0]), .I1(encoder1_position[16]), 
            .I2(n14867), .I3(GND_net), .O(n19411));   // verilog/coms.v(127[12] 300[6])
    defparam i14269_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14270_3_lut (.I0(\data_out_frame[8] [7]), .I1(encoder0_position_scaled[7]), 
            .I2(n14867), .I3(GND_net), .O(n19412));   // verilog/coms.v(127[12] 300[6])
    defparam i14270_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_23__I_0_add_1096_7_lut (.I0(GND_net), .I1(n1623), 
            .I2(GND_net), .I3(n28263), .O(n1676)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1096_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i14271_3_lut (.I0(\data_out_frame[8] [6]), .I1(encoder0_position_scaled[6]), 
            .I2(n14867), .I3(GND_net), .O(n19413));   // verilog/coms.v(127[12] 300[6])
    defparam i14271_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14272_3_lut (.I0(\data_out_frame[8] [5]), .I1(encoder0_position_scaled[5]), 
            .I2(n14867), .I3(GND_net), .O(n19414));   // verilog/coms.v(127[12] 300[6])
    defparam i14272_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14273_3_lut (.I0(\data_out_frame[8] [4]), .I1(encoder0_position_scaled[4]), 
            .I2(n14867), .I3(GND_net), .O(n19415));   // verilog/coms.v(127[12] 300[6])
    defparam i14273_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14274_3_lut (.I0(\data_out_frame[8] [3]), .I1(encoder0_position_scaled[3]), 
            .I2(n14867), .I3(GND_net), .O(n19416));   // verilog/coms.v(127[12] 300[6])
    defparam i14274_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_23__I_0_add_1096_7 (.CI(n28263), .I0(n1623), 
            .I1(GND_net), .CO(n28264));
    SB_LUT4 i14275_3_lut (.I0(\data_out_frame[8] [2]), .I1(encoder0_position_scaled[2]), 
            .I2(n14867), .I3(GND_net), .O(n19417));   // verilog/coms.v(127[12] 300[6])
    defparam i14275_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_23__I_0_add_1096_6_lut (.I0(GND_net), .I1(n1624), 
            .I2(GND_net), .I3(n28262), .O(n1677)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1096_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1096_6 (.CI(n28262), .I0(n1624), 
            .I1(GND_net), .CO(n28263));
    SB_LUT4 encoder0_position_23__I_0_add_1096_5_lut (.I0(GND_net), .I1(n1625), 
            .I2(VCC_net), .I3(n28261), .O(n1678)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1096_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1096_5 (.CI(n28261), .I0(n1625), 
            .I1(VCC_net), .CO(n28262));
    SB_LUT4 add_25_22_lut (.I0(GND_net), .I1(delay_counter[20]), .I2(GND_net), 
            .I3(n27752), .O(n584)) /* synthesis syn_instantiated=1 */ ;
    defparam add_25_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_25_7_lut (.I0(GND_net), .I1(delay_counter[5]), .I2(GND_net), 
            .I3(n27737), .O(n599)) /* synthesis syn_instantiated=1 */ ;
    defparam add_25_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_23__I_0_add_1096_4_lut (.I0(GND_net), .I1(n1626), 
            .I2(GND_net), .I3(n28260), .O(n1679)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1096_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1096_4 (.CI(n28260), .I0(n1626), 
            .I1(GND_net), .CO(n28261));
    SB_LUT4 encoder0_position_23__I_0_add_1096_3_lut (.I0(GND_net), .I1(n1627), 
            .I2(VCC_net), .I3(n28259), .O(n1680)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1096_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1096_3 (.CI(n28259), .I0(n1627), 
            .I1(VCC_net), .CO(n28260));
    SB_LUT4 encoder0_position_23__I_0_add_1096_2_lut (.I0(GND_net), .I1(n770), 
            .I2(GND_net), .I3(VCC_net), .O(n1681)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1096_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1096_2 (.CI(VCC_net), .I0(n770), 
            .I1(GND_net), .CO(n28259));
    SB_LUT4 add_672_6_lut (.I0(duty[4]), .I1(n37633), .I2(n21), .I3(n27829), 
            .O(pwm_setpoint_22__N_11[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_672_6_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 unary_minus_4_inv_0_i5_1_lut (.I0(duty[4]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n21));   // verilog/TinyFPGA_B.v(106[23:28])
    defparam unary_minus_4_inv_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_672_6 (.CI(n27829), .I0(n37633), .I1(n21), .CO(n27830));
    SB_LUT4 encoder0_position_23__I_0_add_1043_19_lut (.I0(GND_net), .I1(n1532), 
            .I2(VCC_net), .I3(n28258), .O(n1585)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1043_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_23__I_0_add_1043_18_lut (.I0(GND_net), .I1(n1533), 
            .I2(VCC_net), .I3(n28257), .O(n1586)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1043_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1043_18 (.CI(n28257), .I0(n1533), 
            .I1(VCC_net), .CO(n28258));
    SB_LUT4 encoder0_position_23__I_0_add_1043_17_lut (.I0(GND_net), .I1(n1534), 
            .I2(VCC_net), .I3(n28256), .O(n1587)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1043_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1043_17 (.CI(n28256), .I0(n1534), 
            .I1(VCC_net), .CO(n28257));
    SB_LUT4 encoder0_position_23__I_0_add_1043_16_lut (.I0(GND_net), .I1(n1535), 
            .I2(VCC_net), .I3(n28255), .O(n1588)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1043_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1043_16 (.CI(n28255), .I0(n1535), 
            .I1(VCC_net), .CO(n28256));
    SB_LUT4 encoder0_position_23__I_0_add_1043_15_lut (.I0(GND_net), .I1(n1536), 
            .I2(VCC_net), .I3(n28254), .O(n1589)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1043_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1043_15 (.CI(n28254), .I0(n1536), 
            .I1(VCC_net), .CO(n28255));
    SB_LUT4 encoder0_position_23__I_0_add_1043_14_lut (.I0(GND_net), .I1(n1537), 
            .I2(VCC_net), .I3(n28253), .O(n1590)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1043_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_25_22 (.CI(n27752), .I0(delay_counter[20]), .I1(GND_net), 
            .CO(n27753));
    SB_LUT4 add_25_2_lut (.I0(GND_net), .I1(delay_counter[0]), .I2(GND_net), 
            .I3(VCC_net), .O(n604)) /* synthesis syn_instantiated=1 */ ;
    defparam add_25_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1043_14 (.CI(n28253), .I0(n1537), 
            .I1(VCC_net), .CO(n28254));
    SB_LUT4 encoder0_position_23__I_0_add_1043_13_lut (.I0(GND_net), .I1(n1538), 
            .I2(VCC_net), .I3(n28252), .O(n1591)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1043_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1043_13 (.CI(n28252), .I0(n1538), 
            .I1(VCC_net), .CO(n28253));
    SB_LUT4 encoder0_position_23__I_0_add_1043_12_lut (.I0(GND_net), .I1(n1539), 
            .I2(VCC_net), .I3(n28251), .O(n1592)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1043_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_25_7 (.CI(n27737), .I0(delay_counter[5]), .I1(GND_net), 
            .CO(n27738));
    SB_CARRY encoder0_position_23__I_0_add_1043_12 (.CI(n28251), .I0(n1539), 
            .I1(VCC_net), .CO(n28252));
    SB_LUT4 encoder0_position_23__I_0_add_1043_11_lut (.I0(GND_net), .I1(n1540), 
            .I2(VCC_net), .I3(n28250), .O(n1593)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1043_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1043_11 (.CI(n28250), .I0(n1540), 
            .I1(VCC_net), .CO(n28251));
    SB_LUT4 encoder0_position_23__I_0_add_1043_10_lut (.I0(GND_net), .I1(n1541), 
            .I2(VCC_net), .I3(n28249), .O(n1594)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1043_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1043_10 (.CI(n28249), .I0(n1541), 
            .I1(VCC_net), .CO(n28250));
    SB_LUT4 add_25_21_lut (.I0(GND_net), .I1(delay_counter[19]), .I2(GND_net), 
            .I3(n27751), .O(n585)) /* synthesis syn_instantiated=1 */ ;
    defparam add_25_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_672_5_lut (.I0(duty[3]), .I1(n37633), .I2(n22), .I3(n27828), 
            .O(pwm_setpoint_22__N_11[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_672_5_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_25_21 (.CI(n27751), .I0(delay_counter[19]), .I1(GND_net), 
            .CO(n27752));
    SB_CARRY add_25_2 (.CI(VCC_net), .I0(delay_counter[0]), .I1(GND_net), 
            .CO(n27733));
    SB_LUT4 encoder0_position_23__I_0_add_1043_9_lut (.I0(GND_net), .I1(n1542), 
            .I2(VCC_net), .I3(n28248), .O(n1595)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1043_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1043_9 (.CI(n28248), .I0(n1542), 
            .I1(VCC_net), .CO(n28249));
    SB_LUT4 encoder0_position_23__I_0_add_1043_8_lut (.I0(GND_net), .I1(n1543), 
            .I2(VCC_net), .I3(n28247), .O(n1596)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1043_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_672_5 (.CI(n27828), .I0(n37633), .I1(n22), .CO(n27829));
    SB_LUT4 add_672_4_lut (.I0(duty[2]), .I1(n37633), .I2(n23), .I3(n27827), 
            .O(pwm_setpoint_22__N_11[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_672_4_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY encoder0_position_23__I_0_add_1043_8 (.CI(n28247), .I0(n1543), 
            .I1(VCC_net), .CO(n28248));
    SB_LUT4 encoder0_position_23__I_0_add_1043_7_lut (.I0(GND_net), .I1(n1544), 
            .I2(GND_net), .I3(n28246), .O(n1597)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1043_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_672_4 (.CI(n27827), .I0(n37633), .I1(n23), .CO(n27828));
    SB_CARRY encoder0_position_23__I_0_add_1043_7 (.CI(n28246), .I0(n1544), 
            .I1(GND_net), .CO(n28247));
    SB_LUT4 encoder0_position_23__I_0_add_1043_6_lut (.I0(GND_net), .I1(n1545), 
            .I2(GND_net), .I3(n28245), .O(n1598)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1043_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1043_6 (.CI(n28245), .I0(n1545), 
            .I1(GND_net), .CO(n28246));
    SB_LUT4 encoder0_position_23__I_0_add_1043_5_lut (.I0(GND_net), .I1(n1546), 
            .I2(VCC_net), .I3(n28244), .O(n1599)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1043_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_23__I_0_unary_minus_2_inv_0_i24_1_lut (.I0(encoder0_position[22]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n3_adj_5005));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_unary_minus_2_inv_0_i24_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY encoder0_position_23__I_0_add_1043_5 (.CI(n28244), .I0(n1546), 
            .I1(VCC_net), .CO(n28245));
    SB_LUT4 encoder0_position_23__I_0_add_1043_4_lut (.I0(GND_net), .I1(n1547), 
            .I2(GND_net), .I3(n28243), .O(n1600)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1043_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1043_4 (.CI(n28243), .I0(n1547), 
            .I1(GND_net), .CO(n28244));
    SB_LUT4 encoder0_position_23__I_0_add_1043_3_lut (.I0(GND_net), .I1(n1548), 
            .I2(VCC_net), .I3(n28242), .O(n1601)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1043_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1043_3 (.CI(n28242), .I0(n1548), 
            .I1(VCC_net), .CO(n28243));
    SB_LUT4 LessThan_744_i35_2_lut (.I0(pwm_counter[17]), .I1(pwm_setpoint[17]), 
            .I2(GND_net), .I3(GND_net), .O(n35));   // verilog/pwm.v(21[8:24])
    defparam LessThan_744_i35_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 encoder0_position_23__I_0_add_1043_2_lut (.I0(GND_net), .I1(n526), 
            .I2(GND_net), .I3(VCC_net), .O(n1602)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1043_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_2_lut_adj_1701 (.I0(n17360), .I1(pwm_counter[31]), .I2(GND_net), 
            .I3(GND_net), .O(n17362));
    defparam i1_2_lut_adj_1701.LUT_INIT = 16'heeee;
    SB_CARRY encoder0_position_23__I_0_add_1043_2 (.CI(VCC_net), .I0(n526), 
            .I1(GND_net), .CO(n28242));
    SB_LUT4 encoder0_position_23__I_0_add_990_18_lut (.I0(GND_net), .I1(n1454), 
            .I2(VCC_net), .I3(n28241), .O(n1507)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_990_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_23__I_0_add_990_17_lut (.I0(GND_net), .I1(n1455), 
            .I2(VCC_net), .I3(n28240), .O(n1508)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_990_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_990_17 (.CI(n28240), .I0(n1455), 
            .I1(VCC_net), .CO(n28241));
    SB_LUT4 encoder0_position_23__I_0_add_990_16_lut (.I0(GND_net), .I1(n1456), 
            .I2(VCC_net), .I3(n28239), .O(n1509)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_990_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i29600_4_lut (.I0(n27_adj_4988), .I1(n15_adj_4982), .I2(n13_adj_4981), 
            .I3(n11_adj_4979), .O(n36355));
    defparam i29600_4_lut.LUT_INIT = 16'haaab;
    SB_CARRY encoder0_position_23__I_0_add_990_16 (.CI(n28239), .I0(n1456), 
            .I1(VCC_net), .CO(n28240));
    SB_LUT4 encoder0_position_23__I_0_add_990_15_lut (.I0(GND_net), .I1(n1457), 
            .I2(VCC_net), .I3(n28238), .O(n1510)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_990_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i29889_4_lut (.I0(n9_adj_4977), .I1(n7_adj_4975), .I2(pwm_counter[2]), 
            .I3(pwm_setpoint[2]), .O(n36644));
    defparam i29889_4_lut.LUT_INIT = 16'heffe;
    SB_CARRY encoder0_position_23__I_0_add_990_15 (.CI(n28238), .I0(n1457), 
            .I1(VCC_net), .CO(n28239));
    SB_LUT4 encoder0_position_23__I_0_add_990_14_lut (.I0(GND_net), .I1(n1458), 
            .I2(VCC_net), .I3(n28237), .O(n1511)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_990_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_990_14 (.CI(n28237), .I0(n1458), 
            .I1(VCC_net), .CO(n28238));
    SB_LUT4 i30061_4_lut (.I0(n15_adj_4982), .I1(n13_adj_4981), .I2(n11_adj_4979), 
            .I3(n36644), .O(n36816));
    defparam i30061_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 encoder0_position_23__I_0_add_990_13_lut (.I0(GND_net), .I1(n1459), 
            .I2(VCC_net), .I3(n28236), .O(n1512)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_990_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i30059_4_lut (.I0(n21_adj_4985), .I1(n19_adj_4984), .I2(n17_adj_4983), 
            .I3(n36816), .O(n36814));
    defparam i30059_4_lut.LUT_INIT = 16'hfeff;
    SB_CARRY encoder0_position_23__I_0_add_990_13 (.CI(n28236), .I0(n1459), 
            .I1(VCC_net), .CO(n28237));
    SB_LUT4 i29602_4_lut (.I0(n27_adj_4988), .I1(n25_adj_4987), .I2(n23_adj_4986), 
            .I3(n36814), .O(n36357));
    defparam i29602_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 encoder0_position_23__I_0_add_990_12_lut (.I0(GND_net), .I1(n1460), 
            .I2(VCC_net), .I3(n28235), .O(n1513)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_990_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_990_12 (.CI(n28235), .I0(n1460), 
            .I1(VCC_net), .CO(n28236));
    SB_LUT4 LessThan_744_i4_4_lut (.I0(pwm_setpoint[0]), .I1(pwm_setpoint[1]), 
            .I2(pwm_counter[1]), .I3(pwm_counter[0]), .O(n4_adj_4973));   // verilog/pwm.v(21[8:24])
    defparam LessThan_744_i4_4_lut.LUT_INIT = 16'h0c8e;
    SB_LUT4 encoder0_position_23__I_0_add_990_11_lut (.I0(GND_net), .I1(n1461), 
            .I2(VCC_net), .I3(n28234), .O(n1514)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_990_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i30209_3_lut (.I0(n4_adj_4973), .I1(pwm_setpoint[13]), .I2(n27_adj_4988), 
            .I3(GND_net), .O(n36964));   // verilog/pwm.v(21[8:24])
    defparam i30209_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_23__I_0_add_990_11 (.CI(n28234), .I0(n1461), 
            .I1(VCC_net), .CO(n28235));
    SB_LUT4 encoder0_position_23__I_0_add_990_10_lut (.I0(GND_net), .I1(n1462), 
            .I2(VCC_net), .I3(n28233), .O(n1515)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_990_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_990_10 (.CI(n28233), .I0(n1462), 
            .I1(VCC_net), .CO(n28234));
    SB_LUT4 encoder0_position_23__I_0_add_990_9_lut (.I0(GND_net), .I1(n1463), 
            .I2(VCC_net), .I3(n28232), .O(n1516)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_990_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_990_9 (.CI(n28232), .I0(n1463), 
            .I1(VCC_net), .CO(n28233));
    SB_LUT4 encoder0_position_23__I_0_add_990_8_lut (.I0(GND_net), .I1(n1464), 
            .I2(VCC_net), .I3(n28231), .O(n1517)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_990_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_990_8 (.CI(n28231), .I0(n1464), 
            .I1(VCC_net), .CO(n28232));
    SB_LUT4 LessThan_744_i30_3_lut (.I0(n12_adj_4980), .I1(pwm_setpoint[17]), 
            .I2(n35), .I3(GND_net), .O(n30_adj_4990));   // verilog/pwm.v(21[8:24])
    defparam LessThan_744_i30_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i30210_3_lut (.I0(n36964), .I1(pwm_setpoint[14]), .I2(n29_adj_4989), 
            .I3(GND_net), .O(n36965));   // verilog/pwm.v(21[8:24])
    defparam i30210_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_23__I_0_add_990_7_lut (.I0(GND_net), .I1(n1465), 
            .I2(GND_net), .I3(n28230), .O(n1518)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_990_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_990_7 (.CI(n28230), .I0(n1465), 
            .I1(GND_net), .CO(n28231));
    SB_LUT4 i29596_4_lut (.I0(n33), .I1(n31), .I2(n29_adj_4989), .I3(n36355), 
            .O(n36351));
    defparam i29596_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i30322_4_lut (.I0(n30_adj_4990), .I1(n10_adj_4978), .I2(n35), 
            .I3(n36349), .O(n37077));   // verilog/pwm.v(21[8:24])
    defparam i30322_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 encoder0_position_23__I_0_add_990_6_lut (.I0(GND_net), .I1(n1466), 
            .I2(GND_net), .I3(n28229), .O(n1519)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_990_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i30190_3_lut (.I0(n36965), .I1(pwm_setpoint[15]), .I2(n31), 
            .I3(GND_net), .O(n36945));   // verilog/pwm.v(21[8:24])
    defparam i30190_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_23__I_0_add_990_6 (.CI(n28229), .I0(n1466), 
            .I1(GND_net), .CO(n28230));
    SB_LUT4 encoder0_position_23__I_0_add_990_5_lut (.I0(GND_net), .I1(n1467), 
            .I2(VCC_net), .I3(n28228), .O(n1520)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_990_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i30211_3_lut (.I0(n6_adj_4974), .I1(pwm_setpoint[10]), .I2(n21_adj_4985), 
            .I3(GND_net), .O(n36966));   // verilog/pwm.v(21[8:24])
    defparam i30211_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_23__I_0_add_990_5 (.CI(n28228), .I0(n1467), 
            .I1(VCC_net), .CO(n28229));
    SB_LUT4 i30212_3_lut (.I0(n36966), .I1(pwm_setpoint[11]), .I2(n23_adj_4986), 
            .I3(GND_net), .O(n36967));   // verilog/pwm.v(21[8:24])
    defparam i30212_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_23__I_0_add_990_4_lut (.I0(GND_net), .I1(n1468), 
            .I2(GND_net), .I3(n28227), .O(n1521)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_990_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_990_4 (.CI(n28227), .I0(n1468), 
            .I1(GND_net), .CO(n28228));
    SB_LUT4 encoder0_position_23__I_0_add_990_3_lut (.I0(GND_net), .I1(n1469), 
            .I2(VCC_net), .I3(n28226), .O(n1522)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_990_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i29879_4_lut (.I0(n23_adj_4986), .I1(n21_adj_4985), .I2(n19_adj_4984), 
            .I3(n36363), .O(n36634));
    defparam i29879_4_lut.LUT_INIT = 16'heeef;
    SB_CARRY encoder0_position_23__I_0_add_990_3 (.CI(n28226), .I0(n1469), 
            .I1(VCC_net), .CO(n28227));
    SB_LUT4 encoder0_position_23__I_0_add_990_2_lut (.I0(GND_net), .I1(n768), 
            .I2(GND_net), .I3(VCC_net), .O(n1523)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_990_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i30123_3_lut (.I0(n8_adj_4976), .I1(pwm_setpoint[9]), .I2(n19_adj_4984), 
            .I3(GND_net), .O(n36878));   // verilog/pwm.v(21[8:24])
    defparam i30123_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_23__I_0_add_990_2 (.CI(VCC_net), .I0(n768), 
            .I1(GND_net), .CO(n28226));
    SB_LUT4 i30188_3_lut (.I0(n36967), .I1(pwm_setpoint[12]), .I2(n25_adj_4987), 
            .I3(GND_net), .O(n36943));   // verilog/pwm.v(21[8:24])
    defparam i30188_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i30145_4_lut (.I0(n33), .I1(n31), .I2(n29_adj_4989), .I3(n36357), 
            .O(n36900));
    defparam i30145_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 encoder0_position_23__I_0_add_937_17_lut (.I0(GND_net), .I1(n1376), 
            .I2(VCC_net), .I3(n28225), .O(n1429)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_937_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i30371_4_lut (.I0(n36945), .I1(n37077), .I2(n35), .I3(n36351), 
            .O(n37126));   // verilog/pwm.v(21[8:24])
    defparam i30371_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i30205_4_lut (.I0(n36943), .I1(n36878), .I2(n25_adj_4987), 
            .I3(n36634), .O(n36960));   // verilog/pwm.v(21[8:24])
    defparam i30205_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 encoder0_position_23__I_0_add_937_16_lut (.I0(GND_net), .I1(n1377), 
            .I2(VCC_net), .I3(n28224), .O(n1430)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_937_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_937_16 (.CI(n28224), .I0(n1377), 
            .I1(VCC_net), .CO(n28225));
    SB_LUT4 i30375_4_lut (.I0(n36960), .I1(n37126), .I2(n35), .I3(n36900), 
            .O(n37130));   // verilog/pwm.v(21[8:24])
    defparam i30375_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 encoder0_position_23__I_0_add_937_15_lut (.I0(GND_net), .I1(n1378), 
            .I2(VCC_net), .I3(n28223), .O(n1431)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_937_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i30376_3_lut (.I0(n37130), .I1(pwm_setpoint[18]), .I2(pwm_counter[18]), 
            .I3(GND_net), .O(n37131));   // verilog/pwm.v(21[8:24])
    defparam i30376_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i30374_3_lut (.I0(n37131), .I1(pwm_setpoint[19]), .I2(pwm_counter[19]), 
            .I3(GND_net), .O(n37129));   // verilog/pwm.v(21[8:24])
    defparam i30374_3_lut.LUT_INIT = 16'h8e8e;
    SB_CARRY encoder0_position_23__I_0_add_937_15 (.CI(n28223), .I0(n1378), 
            .I1(VCC_net), .CO(n28224));
    SB_LUT4 encoder0_position_23__I_0_add_937_14_lut (.I0(GND_net), .I1(n1379), 
            .I2(VCC_net), .I3(n28222), .O(n1432)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_937_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i30302_3_lut (.I0(n37129), .I1(pwm_setpoint[20]), .I2(pwm_counter[20]), 
            .I3(GND_net), .O(n37057));   // verilog/pwm.v(21[8:24])
    defparam i30302_3_lut.LUT_INIT = 16'h8e8e;
    SB_CARRY encoder0_position_23__I_0_add_937_14 (.CI(n28222), .I0(n1379), 
            .I1(VCC_net), .CO(n28223));
    SB_LUT4 encoder0_position_23__I_0_add_937_13_lut (.I0(GND_net), .I1(n1380), 
            .I2(VCC_net), .I3(n28221), .O(n1433)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_937_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_937_13 (.CI(n28221), .I0(n1380), 
            .I1(VCC_net), .CO(n28222));
    SB_LUT4 encoder0_position_23__I_0_add_937_12_lut (.I0(GND_net), .I1(n1381), 
            .I2(VCC_net), .I3(n28220), .O(n1434)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_937_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_937_12 (.CI(n28220), .I0(n1381), 
            .I1(VCC_net), .CO(n28221));
    SB_LUT4 encoder0_position_23__I_0_add_937_11_lut (.I0(GND_net), .I1(n1382), 
            .I2(VCC_net), .I3(n28219), .O(n1435)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_937_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_937_11 (.CI(n28219), .I0(n1382), 
            .I1(VCC_net), .CO(n28220));
    SB_LUT4 encoder0_position_23__I_0_add_937_10_lut (.I0(GND_net), .I1(n1383), 
            .I2(VCC_net), .I3(n28218), .O(n1436)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_937_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_937_10 (.CI(n28218), .I0(n1383), 
            .I1(VCC_net), .CO(n28219));
    SB_LUT4 i30303_3_lut (.I0(n37057), .I1(pwm_setpoint[21]), .I2(pwm_counter[21]), 
            .I3(GND_net), .O(n37058));   // verilog/pwm.v(21[8:24])
    defparam i30303_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 encoder0_position_23__I_0_add_937_9_lut (.I0(GND_net), .I1(n1384), 
            .I2(VCC_net), .I3(n28217), .O(n1437)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_937_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_25_20_lut (.I0(GND_net), .I1(delay_counter[18]), .I2(GND_net), 
            .I3(n27750), .O(n586)) /* synthesis syn_instantiated=1 */ ;
    defparam add_25_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_937_9 (.CI(n28217), .I0(n1384), 
            .I1(VCC_net), .CO(n28218));
    SB_LUT4 encoder0_position_23__I_0_add_937_8_lut (.I0(GND_net), .I1(n1385), 
            .I2(VCC_net), .I3(n28216), .O(n1438)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_937_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_937_8 (.CI(n28216), .I0(n1385), 
            .I1(VCC_net), .CO(n28217));
    SB_LUT4 encoder0_position_23__I_0_add_937_7_lut (.I0(GND_net), .I1(n1386), 
            .I2(GND_net), .I3(n28215), .O(n1439)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_937_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_937_7 (.CI(n28215), .I0(n1386), 
            .I1(GND_net), .CO(n28216));
    SB_LUT4 encoder0_position_23__I_0_add_937_6_lut (.I0(GND_net), .I1(n1387), 
            .I2(GND_net), .I3(n28214), .O(n1440)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_937_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_937_6 (.CI(n28214), .I0(n1387), 
            .I1(GND_net), .CO(n28215));
    SB_LUT4 encoder0_position_23__I_0_add_937_5_lut (.I0(GND_net), .I1(n1388), 
            .I2(VCC_net), .I3(n28213), .O(n1441)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_937_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_937_5 (.CI(n28213), .I0(n1388), 
            .I1(VCC_net), .CO(n28214));
    SB_LUT4 encoder0_position_23__I_0_add_937_4_lut (.I0(GND_net), .I1(n1389), 
            .I2(GND_net), .I3(n28212), .O(n1442)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_937_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_937_4 (.CI(n28212), .I0(n1389), 
            .I1(GND_net), .CO(n28213));
    SB_LUT4 encoder0_position_23__I_0_add_937_3_lut (.I0(GND_net), .I1(n1390), 
            .I2(VCC_net), .I3(n28211), .O(n1443)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_937_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_937_3 (.CI(n28211), .I0(n1390), 
            .I1(VCC_net), .CO(n28212));
    SB_LUT4 encoder0_position_23__I_0_add_937_2_lut (.I0(GND_net), .I1(n767), 
            .I2(GND_net), .I3(VCC_net), .O(n1444)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_937_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_937_2 (.CI(VCC_net), .I0(n767), 
            .I1(GND_net), .CO(n28211));
    SB_LUT4 encoder0_position_23__I_0_add_884_16_lut (.I0(GND_net), .I1(n1298), 
            .I2(VCC_net), .I3(n28210), .O(n1351)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_884_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_23__I_0_add_884_15_lut (.I0(GND_net), .I1(n1299), 
            .I2(VCC_net), .I3(n28209), .O(n1352)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_884_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_884_15 (.CI(n28209), .I0(n1299), 
            .I1(VCC_net), .CO(n28210));
    SB_CARRY add_25_20 (.CI(n27750), .I0(delay_counter[18]), .I1(GND_net), 
            .CO(n27751));
    SB_LUT4 encoder0_position_23__I_0_add_884_14_lut (.I0(GND_net), .I1(n1300), 
            .I2(VCC_net), .I3(n28208), .O(n1353)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_884_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_884_14 (.CI(n28208), .I0(n1300), 
            .I1(VCC_net), .CO(n28209));
    SB_LUT4 encoder0_position_23__I_0_add_884_13_lut (.I0(GND_net), .I1(n1301), 
            .I2(VCC_net), .I3(n28207), .O(n1354)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_884_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_25_19_lut (.I0(GND_net), .I1(delay_counter[17]), .I2(GND_net), 
            .I3(n27749), .O(n587)) /* synthesis syn_instantiated=1 */ ;
    defparam add_25_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_884_13 (.CI(n28207), .I0(n1301), 
            .I1(VCC_net), .CO(n28208));
    SB_LUT4 add_25_6_lut (.I0(GND_net), .I1(delay_counter[4]), .I2(GND_net), 
            .I3(n27736), .O(n600)) /* synthesis syn_instantiated=1 */ ;
    defparam add_25_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_25_19 (.CI(n27749), .I0(delay_counter[17]), .I1(GND_net), 
            .CO(n27750));
    SB_LUT4 add_25_18_lut (.I0(GND_net), .I1(delay_counter[16]), .I2(GND_net), 
            .I3(n27748), .O(n588)) /* synthesis syn_instantiated=1 */ ;
    defparam add_25_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_25_18 (.CI(n27748), .I0(delay_counter[16]), .I1(GND_net), 
            .CO(n27749));
    SB_LUT4 i3_4_lut_4_lut (.I0(r_SM_Main_adj_5135[1]), .I1(r_SM_Main_adj_5135[0]), 
            .I2(r_SM_Main_adj_5135[2]), .I3(r_SM_Main_2__N_3487[1]), .O(n38214));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i3_4_lut_4_lut.LUT_INIT = 16'h0800;
    SB_LUT4 encoder0_position_23__I_0_add_884_12_lut (.I0(GND_net), .I1(n1302), 
            .I2(VCC_net), .I3(n28206), .O(n1355)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_884_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_884_12 (.CI(n28206), .I0(n1302), 
            .I1(VCC_net), .CO(n28207));
    SB_LUT4 encoder0_position_23__I_0_add_884_11_lut (.I0(GND_net), .I1(n1303), 
            .I2(VCC_net), .I3(n28205), .O(n1356)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_884_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_884_11 (.CI(n28205), .I0(n1303), 
            .I1(VCC_net), .CO(n28206));
    SB_DFFESR delay_counter_i0_i24 (.Q(delay_counter[24]), .C(CLK_c), .E(n5410), 
            .D(n580), .R(n18963));   // verilog/TinyFPGA_B.v(237[10] 265[6])
    SB_LUT4 encoder0_position_23__I_0_add_884_10_lut (.I0(GND_net), .I1(n1304), 
            .I2(VCC_net), .I3(n28204), .O(n1357)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_884_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_884_10 (.CI(n28204), .I0(n1304), 
            .I1(VCC_net), .CO(n28205));
    SB_LUT4 add_672_3_lut (.I0(duty[1]), .I1(n37633), .I2(n24), .I3(n27826), 
            .O(pwm_setpoint_22__N_11[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_672_3_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 encoder0_position_23__I_0_add_884_9_lut (.I0(GND_net), .I1(n1305), 
            .I2(VCC_net), .I3(n28203), .O(n1358)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_884_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_884_9 (.CI(n28203), .I0(n1305), 
            .I1(VCC_net), .CO(n28204));
    SB_LUT4 encoder0_position_23__I_0_unary_minus_2_inv_0_i25_1_lut (.I0(encoder0_position[23]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n2_adj_5004));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_unary_minus_2_inv_0_i25_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_23__I_0_add_884_8_lut (.I0(GND_net), .I1(n1306), 
            .I2(VCC_net), .I3(n28202), .O(n1359)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_884_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_884_8 (.CI(n28202), .I0(n1306), 
            .I1(VCC_net), .CO(n28203));
    SB_DFFESR delay_counter_i0_i23 (.Q(delay_counter[23]), .C(CLK_c), .E(n5410), 
            .D(n581), .R(n18963));   // verilog/TinyFPGA_B.v(237[10] 265[6])
    SB_LUT4 encoder0_position_23__I_0_add_884_7_lut (.I0(GND_net), .I1(n1307), 
            .I2(GND_net), .I3(n28201), .O(n1360)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_884_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_884_7 (.CI(n28201), .I0(n1307), 
            .I1(GND_net), .CO(n28202));
    SB_DFFESR delay_counter_i0_i22 (.Q(delay_counter[22]), .C(CLK_c), .E(n5410), 
            .D(n582), .R(n18963));   // verilog/TinyFPGA_B.v(237[10] 265[6])
    SB_LUT4 encoder0_position_23__I_0_add_884_6_lut (.I0(GND_net), .I1(n1308), 
            .I2(GND_net), .I3(n28200), .O(n1361)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_884_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_884_6 (.CI(n28200), .I0(n1308), 
            .I1(GND_net), .CO(n28201));
    SB_LUT4 encoder0_position_23__I_0_add_884_5_lut (.I0(GND_net), .I1(n1309), 
            .I2(VCC_net), .I3(n28199), .O(n1362)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_884_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_884_5 (.CI(n28199), .I0(n1309), 
            .I1(VCC_net), .CO(n28200));
    SB_LUT4 encoder0_position_23__I_0_add_884_4_lut (.I0(GND_net), .I1(n1310), 
            .I2(GND_net), .I3(n28198), .O(n1363)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_884_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_884_4 (.CI(n28198), .I0(n1310), 
            .I1(GND_net), .CO(n28199));
    SB_LUT4 encoder0_position_23__I_0_add_884_3_lut (.I0(GND_net), .I1(n1311), 
            .I2(VCC_net), .I3(n28197), .O(n1364)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_884_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_884_3 (.CI(n28197), .I0(n1311), 
            .I1(VCC_net), .CO(n28198));
    SB_LUT4 encoder0_position_23__I_0_add_884_2_lut (.I0(GND_net), .I1(n523), 
            .I2(GND_net), .I3(VCC_net), .O(n1365)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_884_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_884_2 (.CI(VCC_net), .I0(n523), 
            .I1(GND_net), .CO(n28197));
    SB_CARRY add_672_3 (.CI(n27826), .I0(n37633), .I1(n24), .CO(n27827));
    SB_DFFESR delay_counter_i0_i21 (.Q(delay_counter[21]), .C(CLK_c), .E(n5410), 
            .D(n583), .R(n18963));   // verilog/TinyFPGA_B.v(237[10] 265[6])
    SB_LUT4 add_25_17_lut (.I0(GND_net), .I1(delay_counter[15]), .I2(GND_net), 
            .I3(n27747), .O(n589)) /* synthesis syn_instantiated=1 */ ;
    defparam add_25_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i14276_3_lut (.I0(\data_out_frame[8] [1]), .I1(encoder0_position_scaled[1]), 
            .I2(n14867), .I3(GND_net), .O(n19418));   // verilog/coms.v(127[12] 300[6])
    defparam i14276_3_lut.LUT_INIT = 16'hcaca;
    SB_DFFESR delay_counter_i0_i20 (.Q(delay_counter[20]), .C(CLK_c), .E(n5410), 
            .D(n584), .R(n18963));   // verilog/TinyFPGA_B.v(237[10] 265[6])
    SB_CARRY add_25_17 (.CI(n27747), .I0(delay_counter[15]), .I1(GND_net), 
            .CO(n27748));
    SB_LUT4 i14277_3_lut (.I0(\data_out_frame[8] [0]), .I1(encoder0_position_scaled[0]), 
            .I2(n14867), .I3(GND_net), .O(n19419));   // verilog/coms.v(127[12] 300[6])
    defparam i14277_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14278_3_lut (.I0(\data_out_frame[7] [7]), .I1(encoder0_position_scaled[15]), 
            .I2(n14867), .I3(GND_net), .O(n19420));   // verilog/coms.v(127[12] 300[6])
    defparam i14278_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14279_3_lut (.I0(\data_out_frame[7] [6]), .I1(encoder0_position_scaled[14]), 
            .I2(n14867), .I3(GND_net), .O(n19421));   // verilog/coms.v(127[12] 300[6])
    defparam i14279_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_23__I_0_add_831_15_lut (.I0(GND_net), .I1(n1220), 
            .I2(VCC_net), .I3(n28188), .O(n1273)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_831_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_23__I_0_add_831_14_lut (.I0(GND_net), .I1(n1221), 
            .I2(VCC_net), .I3(n28187), .O(n1274)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_831_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_831_14 (.CI(n28187), .I0(n1221), 
            .I1(VCC_net), .CO(n28188));
    SB_LUT4 encoder0_position_23__I_0_add_831_13_lut (.I0(GND_net), .I1(n1222), 
            .I2(VCC_net), .I3(n28186), .O(n1275)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_831_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i14280_3_lut (.I0(\data_out_frame[7] [5]), .I1(encoder0_position_scaled[13]), 
            .I2(n14867), .I3(GND_net), .O(n19422));   // verilog/coms.v(127[12] 300[6])
    defparam i14280_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_23__I_0_add_831_13 (.CI(n28186), .I0(n1222), 
            .I1(VCC_net), .CO(n28187));
    SB_LUT4 i14281_3_lut (.I0(\data_out_frame[7] [4]), .I1(encoder0_position_scaled[12]), 
            .I2(n14867), .I3(GND_net), .O(n19423));   // verilog/coms.v(127[12] 300[6])
    defparam i14281_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14282_3_lut (.I0(\data_out_frame[7] [3]), .I1(encoder0_position_scaled[11]), 
            .I2(n14867), .I3(GND_net), .O(n19424));   // verilog/coms.v(127[12] 300[6])
    defparam i14282_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14283_3_lut (.I0(\data_out_frame[7] [2]), .I1(encoder0_position_scaled[10]), 
            .I2(n14867), .I3(GND_net), .O(n19425));   // verilog/coms.v(127[12] 300[6])
    defparam i14283_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_77_i7_4_lut (.I0(encoder1_position[6]), .I1(displacement[6]), 
            .I2(n15_adj_4934), .I3(n15_adj_4940), .O(motor_state_23__N_82[6]));   // verilog/TinyFPGA_B.v(166[5] 168[10])
    defparam mux_77_i7_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i14284_3_lut (.I0(\data_out_frame[7] [1]), .I1(encoder0_position_scaled[9]), 
            .I2(n14867), .I3(GND_net), .O(n19426));   // verilog/coms.v(127[12] 300[6])
    defparam i14284_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14285_3_lut (.I0(\data_out_frame[7] [0]), .I1(encoder0_position_scaled[8]), 
            .I2(n14867), .I3(GND_net), .O(n19427));   // verilog/coms.v(127[12] 300[6])
    defparam i14285_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14286_3_lut (.I0(\data_out_frame[6] [7]), .I1(encoder0_position_scaled[22]), 
            .I2(n14867), .I3(GND_net), .O(n19428));   // verilog/coms.v(127[12] 300[6])
    defparam i14286_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14287_3_lut (.I0(\data_out_frame[6] [6]), .I1(encoder0_position_scaled[22]), 
            .I2(n14867), .I3(GND_net), .O(n19429));   // verilog/coms.v(127[12] 300[6])
    defparam i14287_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder1_position_23__I_0_inv_0_i17_1_lut (.I0(encoder0_position_scaled[16]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n9_adj_4949));   // verilog/TinyFPGA_B.v(202[21:65])
    defparam encoder1_position_23__I_0_inv_0_i17_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i14288_3_lut (.I0(\data_out_frame[6] [5]), .I1(encoder0_position_scaled[22]), 
            .I2(n14867), .I3(GND_net), .O(n19430));   // verilog/coms.v(127[12] 300[6])
    defparam i14288_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14289_3_lut (.I0(\data_out_frame[6] [4]), .I1(encoder0_position_scaled[20]), 
            .I2(n14867), .I3(GND_net), .O(n19431));   // verilog/coms.v(127[12] 300[6])
    defparam i14289_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_23__I_0_add_831_12_lut (.I0(GND_net), .I1(n1223), 
            .I2(VCC_net), .I3(n28185), .O(n1276)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_831_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder1_position_23__I_0_inv_0_i18_1_lut (.I0(encoder0_position_scaled[17]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n8_adj_4948));   // verilog/TinyFPGA_B.v(202[21:65])
    defparam encoder1_position_23__I_0_inv_0_i18_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i14290_3_lut (.I0(\data_out_frame[6] [3]), .I1(encoder0_position_scaled[19]), 
            .I2(n14867), .I3(GND_net), .O(n19432));   // verilog/coms.v(127[12] 300[6])
    defparam i14290_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14291_3_lut (.I0(\data_out_frame[6] [2]), .I1(encoder0_position_scaled[18]), 
            .I2(n14867), .I3(GND_net), .O(n19433));   // verilog/coms.v(127[12] 300[6])
    defparam i14291_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14292_3_lut (.I0(\data_out_frame[6] [1]), .I1(encoder0_position_scaled[17]), 
            .I2(n14867), .I3(GND_net), .O(n19434));   // verilog/coms.v(127[12] 300[6])
    defparam i14292_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14293_3_lut (.I0(\data_out_frame[6] [0]), .I1(encoder0_position_scaled[16]), 
            .I2(n14867), .I3(GND_net), .O(n19435));   // verilog/coms.v(127[12] 300[6])
    defparam i14293_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_23__I_0_add_831_12 (.CI(n28185), .I0(n1223), 
            .I1(VCC_net), .CO(n28186));
    SB_LUT4 i14294_3_lut (.I0(\data_out_frame[5] [7]), .I1(control_mode[7]), 
            .I2(n14867), .I3(GND_net), .O(n19436));   // verilog/coms.v(127[12] 300[6])
    defparam i14294_3_lut.LUT_INIT = 16'hcaca;
    SB_DFFESR delay_counter_i0_i19 (.Q(delay_counter[19]), .C(CLK_c), .E(n5410), 
            .D(n585), .R(n18963));   // verilog/TinyFPGA_B.v(237[10] 265[6])
    SB_LUT4 encoder0_position_23__I_0_add_831_11_lut (.I0(GND_net), .I1(n1224), 
            .I2(VCC_net), .I3(n28184), .O(n1277)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_831_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_831_11 (.CI(n28184), .I0(n1224), 
            .I1(VCC_net), .CO(n28185));
    SB_LUT4 encoder0_position_23__I_0_add_831_10_lut (.I0(GND_net), .I1(n1225), 
            .I2(VCC_net), .I3(n28183), .O(n1278)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_831_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i14295_3_lut (.I0(\data_out_frame[5] [6]), .I1(control_mode[6]), 
            .I2(n14867), .I3(GND_net), .O(n19437));   // verilog/coms.v(127[12] 300[6])
    defparam i14295_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14296_3_lut (.I0(\data_out_frame[5] [5]), .I1(control_mode[5]), 
            .I2(n14867), .I3(GND_net), .O(n19438));   // verilog/coms.v(127[12] 300[6])
    defparam i14296_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_25_16_lut (.I0(GND_net), .I1(delay_counter[14]), .I2(GND_net), 
            .I3(n27746), .O(n590)) /* synthesis syn_instantiated=1 */ ;
    defparam add_25_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_831_10 (.CI(n28183), .I0(n1225), 
            .I1(VCC_net), .CO(n28184));
    SB_LUT4 i14297_3_lut (.I0(\data_out_frame[5] [4]), .I1(control_mode[4]), 
            .I2(n14867), .I3(GND_net), .O(n19439));   // verilog/coms.v(127[12] 300[6])
    defparam i14297_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_23__I_0_add_831_9_lut (.I0(GND_net), .I1(n1226), 
            .I2(VCC_net), .I3(n28182), .O(n1279)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_831_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_831_9 (.CI(n28182), .I0(n1226), 
            .I1(VCC_net), .CO(n28183));
    SB_LUT4 i14298_3_lut (.I0(\data_out_frame[5] [3]), .I1(control_mode[3]), 
            .I2(n14867), .I3(GND_net), .O(n19440));   // verilog/coms.v(127[12] 300[6])
    defparam i14298_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_23__I_0_add_831_8_lut (.I0(GND_net), .I1(n1227), 
            .I2(VCC_net), .I3(n28181), .O(n1280)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_831_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_831_8 (.CI(n28181), .I0(n1227), 
            .I1(VCC_net), .CO(n28182));
    SB_LUT4 encoder0_position_23__I_0_add_831_7_lut (.I0(GND_net), .I1(n1228), 
            .I2(GND_net), .I3(n28180), .O(n1281)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_831_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_831_7 (.CI(n28180), .I0(n1228), 
            .I1(GND_net), .CO(n28181));
    SB_LUT4 encoder0_position_23__I_0_add_831_6_lut (.I0(GND_net), .I1(n1229), 
            .I2(GND_net), .I3(n28179), .O(n1282)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_831_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_831_6 (.CI(n28179), .I0(n1229), 
            .I1(GND_net), .CO(n28180));
    SB_LUT4 encoder0_position_23__I_0_add_831_5_lut (.I0(GND_net), .I1(n1230), 
            .I2(VCC_net), .I3(n28178), .O(n1283)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_831_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i14299_3_lut (.I0(\data_out_frame[5] [2]), .I1(control_mode[2]), 
            .I2(n14867), .I3(GND_net), .O(n19441));   // verilog/coms.v(127[12] 300[6])
    defparam i14299_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13850_4_lut (.I0(n5410), .I1(n691), .I2(n36275), .I3(n17359), 
            .O(n18963));   // verilog/TinyFPGA_B.v(237[10] 265[6])
    defparam i13850_4_lut.LUT_INIT = 16'ha088;
    SB_LUT4 i14300_3_lut (.I0(\data_out_frame[5] [1]), .I1(control_mode[1]), 
            .I2(n14867), .I3(GND_net), .O(n19442));   // verilog/coms.v(127[12] 300[6])
    defparam i14300_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14301_3_lut (.I0(\data_out_frame[5] [0]), .I1(control_mode[0]), 
            .I2(n14867), .I3(GND_net), .O(n19443));   // verilog/coms.v(127[12] 300[6])
    defparam i14301_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14302_3_lut (.I0(\data_out_frame[4] [7]), .I1(ID[7]), .I2(n14867), 
            .I3(GND_net), .O(n19444));   // verilog/coms.v(127[12] 300[6])
    defparam i14302_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14303_3_lut (.I0(\data_out_frame[4] [6]), .I1(ID[6]), .I2(n14867), 
            .I3(GND_net), .O(n19445));   // verilog/coms.v(127[12] 300[6])
    defparam i14303_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_23__I_0_add_831_5 (.CI(n28178), .I0(n1230), 
            .I1(VCC_net), .CO(n28179));
    SB_LUT4 encoder0_position_23__I_0_add_831_4_lut (.I0(GND_net), .I1(n1231), 
            .I2(GND_net), .I3(n28177), .O(n1284)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_831_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_831_4 (.CI(n28177), .I0(n1231), 
            .I1(GND_net), .CO(n28178));
    SB_LUT4 encoder0_position_23__I_0_add_831_3_lut (.I0(GND_net), .I1(n1232), 
            .I2(VCC_net), .I3(n28176), .O(n1285)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_831_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i14304_3_lut (.I0(\data_out_frame[4] [5]), .I1(ID[5]), .I2(n14867), 
            .I3(GND_net), .O(n19446));   // verilog/coms.v(127[12] 300[6])
    defparam i14304_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_23__I_0_add_831_3 (.CI(n28176), .I0(n1232), 
            .I1(VCC_net), .CO(n28177));
    SB_LUT4 i14305_3_lut (.I0(\data_out_frame[4] [4]), .I1(ID[4]), .I2(n14867), 
            .I3(GND_net), .O(n19447));   // verilog/coms.v(127[12] 300[6])
    defparam i14305_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14306_3_lut (.I0(\data_out_frame[4] [3]), .I1(ID[3]), .I2(n14867), 
            .I3(GND_net), .O(n19448));   // verilog/coms.v(127[12] 300[6])
    defparam i14306_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14307_3_lut (.I0(\data_out_frame[4] [2]), .I1(ID[2]), .I2(n14867), 
            .I3(GND_net), .O(n19449));   // verilog/coms.v(127[12] 300[6])
    defparam i14307_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF encoder0_position_scaled_i0 (.Q(encoder0_position_scaled[0]), .C(clk32MHz), 
           .D(encoder0_position_scaled_23__N_34[0]));   // verilog/TinyFPGA_B.v(200[10] 203[6])
    SB_LUT4 i14308_3_lut (.I0(\data_out_frame[4] [1]), .I1(ID[1]), .I2(n14867), 
            .I3(GND_net), .O(n19450));   // verilog/coms.v(127[12] 300[6])
    defparam i14308_3_lut.LUT_INIT = 16'hcaca;
    pll32MHz pll32MHz_inst (.GND_net(GND_net), .CLK_c(CLK_c), .VCC_net(VCC_net), 
            .clk32MHz(clk32MHz)) /* synthesis syn_module_defined=1 */ ;   // verilog/TinyFPGA_B.v(34[10] 37[2])
    SB_LUT4 encoder0_position_23__I_0_add_831_2_lut (.I0(GND_net), .I1(n765), 
            .I2(GND_net), .I3(VCC_net), .O(n1286)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_831_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_831_2 (.CI(VCC_net), .I0(n765), 
            .I1(GND_net), .CO(n28176));
    SB_LUT4 encoder0_position_23__I_0_add_778_14_lut (.I0(GND_net), .I1(n1142), 
            .I2(VCC_net), .I3(n28175), .O(n1195)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_778_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i14309_3_lut (.I0(\data_out_frame[4] [0]), .I1(ID[0]), .I2(n14867), 
            .I3(GND_net), .O(n19451));   // verilog/coms.v(127[12] 300[6])
    defparam i14309_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14310_3_lut (.I0(Ki[15]), .I1(\data_in_frame[4] [7]), .I2(n33567), 
            .I3(GND_net), .O(n19452));   // verilog/coms.v(127[12] 300[6])
    defparam i14310_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_add_778_13_lut (.I0(GND_net), .I1(n1143), 
            .I2(VCC_net), .I3(n28174), .O(n1196)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_778_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_778_13 (.CI(n28174), .I0(n1143), 
            .I1(VCC_net), .CO(n28175));
    SB_LUT4 i16_4_lut_adj_1702 (.I0(state_adj_5158[0]), .I1(n36289), .I2(n5212), 
            .I3(n23736), .O(n8_adj_4900));   // verilog/i2c_controller.v(91[8] 173[6])
    defparam i16_4_lut_adj_1702.LUT_INIT = 16'h3afa;
    SB_LUT4 i14319_3_lut (.I0(Ki[14]), .I1(\data_in_frame[4] [6]), .I2(n33567), 
            .I3(GND_net), .O(n19461));   // verilog/coms.v(127[12] 300[6])
    defparam i14319_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_add_778_12_lut (.I0(GND_net), .I1(n1144), 
            .I2(VCC_net), .I3(n28173), .O(n1197)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_778_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_778_12 (.CI(n28173), .I0(n1144), 
            .I1(VCC_net), .CO(n28174));
    SB_CARRY add_25_16 (.CI(n27746), .I0(delay_counter[14]), .I1(GND_net), 
            .CO(n27747));
    SB_LUT4 i14320_3_lut (.I0(Ki[13]), .I1(\data_in_frame[4] [5]), .I2(n33567), 
            .I3(GND_net), .O(n19462));   // verilog/coms.v(127[12] 300[6])
    defparam i14320_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_add_778_11_lut (.I0(GND_net), .I1(n1145), 
            .I2(VCC_net), .I3(n28172), .O(n1198)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_778_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_778_11 (.CI(n28172), .I0(n1145), 
            .I1(VCC_net), .CO(n28173));
    SB_LUT4 i14321_3_lut (.I0(Ki[12]), .I1(\data_in_frame[4] [4]), .I2(n33567), 
            .I3(GND_net), .O(n19463));   // verilog/coms.v(127[12] 300[6])
    defparam i14321_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_add_778_10_lut (.I0(GND_net), .I1(n1146), 
            .I2(VCC_net), .I3(n28171), .O(n1199)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_778_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_778_10 (.CI(n28171), .I0(n1146), 
            .I1(VCC_net), .CO(n28172));
    SB_LUT4 encoder0_position_23__I_0_add_778_9_lut (.I0(GND_net), .I1(n1147), 
            .I2(VCC_net), .I3(n28170), .O(n1200)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_778_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_778_9 (.CI(n28170), .I0(n1147), 
            .I1(VCC_net), .CO(n28171));
    SB_LUT4 encoder0_position_23__I_0_add_778_8_lut (.I0(GND_net), .I1(n1148), 
            .I2(VCC_net), .I3(n28169), .O(n1201)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_778_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_778_8 (.CI(n28169), .I0(n1148), 
            .I1(VCC_net), .CO(n28170));
    SB_LUT4 encoder0_position_23__I_0_add_778_7_lut (.I0(GND_net), .I1(n1149), 
            .I2(GND_net), .I3(n28168), .O(n1202)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_778_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_778_7 (.CI(n28168), .I0(n1149), 
            .I1(GND_net), .CO(n28169));
    SB_LUT4 i14322_3_lut (.I0(Ki[11]), .I1(\data_in_frame[4] [3]), .I2(n33567), 
            .I3(GND_net), .O(n19464));   // verilog/coms.v(127[12] 300[6])
    defparam i14322_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_add_778_6_lut (.I0(GND_net), .I1(n1150), 
            .I2(GND_net), .I3(n28167), .O(n1203)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_778_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_778_6 (.CI(n28167), .I0(n1150), 
            .I1(GND_net), .CO(n28168));
    SB_LUT4 add_672_2_lut (.I0(duty[0]), .I1(n37633), .I2(n25), .I3(VCC_net), 
            .O(pwm_setpoint_22__N_11[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_672_2_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 encoder0_position_23__I_0_add_778_5_lut (.I0(GND_net), .I1(n1151), 
            .I2(VCC_net), .I3(n28166), .O(n1204)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_778_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_778_5 (.CI(n28166), .I0(n1151), 
            .I1(VCC_net), .CO(n28167));
    SB_LUT4 encoder0_position_23__I_0_add_778_4_lut (.I0(GND_net), .I1(n1152), 
            .I2(GND_net), .I3(n28165), .O(n1205)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_778_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_672_2 (.CI(VCC_net), .I0(n37633), .I1(n25), .CO(n27826));
    SB_CARRY encoder0_position_23__I_0_add_778_4 (.CI(n28165), .I0(n1152), 
            .I1(GND_net), .CO(n28166));
    SB_LUT4 encoder0_position_23__I_0_add_778_3_lut (.I0(GND_net), .I1(n1153), 
            .I2(VCC_net), .I3(n28164), .O(n1206)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_778_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_778_3 (.CI(n28164), .I0(n1153), 
            .I1(VCC_net), .CO(n28165));
    SB_LUT4 encoder0_position_23__I_0_add_778_2_lut (.I0(GND_net), .I1(n521), 
            .I2(GND_net), .I3(VCC_net), .O(n1207)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_778_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_778_2 (.CI(VCC_net), .I0(n521), 
            .I1(GND_net), .CO(n28164));
    SB_LUT4 encoder0_position_23__I_0_add_725_13_lut (.I0(GND_net), .I1(n1064), 
            .I2(VCC_net), .I3(n28163), .O(n1117)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_725_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_23__I_0_add_725_12_lut (.I0(GND_net), .I1(n1065), 
            .I2(VCC_net), .I3(n28162), .O(n1118)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_725_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_725_12 (.CI(n28162), .I0(n1065), 
            .I1(VCC_net), .CO(n28163));
    SB_LUT4 i14323_3_lut (.I0(Ki[10]), .I1(\data_in_frame[4] [2]), .I2(n33567), 
            .I3(GND_net), .O(n19465));   // verilog/coms.v(127[12] 300[6])
    defparam i14323_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_add_725_11_lut (.I0(GND_net), .I1(n1066), 
            .I2(VCC_net), .I3(n28161), .O(n1119)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_725_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_725_11 (.CI(n28161), .I0(n1066), 
            .I1(VCC_net), .CO(n28162));
    SB_LUT4 encoder0_position_23__I_0_add_725_10_lut (.I0(GND_net), .I1(n1067), 
            .I2(VCC_net), .I3(n28160), .O(n1120)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_725_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_725_10 (.CI(n28160), .I0(n1067), 
            .I1(VCC_net), .CO(n28161));
    SB_LUT4 encoder0_position_23__I_0_add_725_9_lut (.I0(GND_net), .I1(n1068), 
            .I2(VCC_net), .I3(n28159), .O(n1121)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_725_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_725_9 (.CI(n28159), .I0(n1068), 
            .I1(VCC_net), .CO(n28160));
    SB_LUT4 encoder0_position_23__I_0_add_725_8_lut (.I0(GND_net), .I1(n1069), 
            .I2(VCC_net), .I3(n28158), .O(n1122)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_725_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_725_8 (.CI(n28158), .I0(n1069), 
            .I1(VCC_net), .CO(n28159));
    SB_LUT4 encoder0_position_23__I_0_add_725_7_lut (.I0(GND_net), .I1(n1070), 
            .I2(GND_net), .I3(n28157), .O(n1123)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_725_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_725_7 (.CI(n28157), .I0(n1070), 
            .I1(GND_net), .CO(n28158));
    SB_LUT4 encoder0_position_23__I_0_add_725_6_lut (.I0(GND_net), .I1(n1071), 
            .I2(GND_net), .I3(n28156), .O(n1124)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_725_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_725_6 (.CI(n28156), .I0(n1071), 
            .I1(GND_net), .CO(n28157));
    SB_LUT4 encoder0_position_23__I_0_add_725_5_lut (.I0(GND_net), .I1(n1072), 
            .I2(VCC_net), .I3(n28155), .O(n1125)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_725_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_725_5 (.CI(n28155), .I0(n1072), 
            .I1(VCC_net), .CO(n28156));
    SB_LUT4 encoder0_position_23__I_0_add_725_4_lut (.I0(GND_net), .I1(n1073), 
            .I2(GND_net), .I3(n28154), .O(n1126)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_725_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_725_4 (.CI(n28154), .I0(n1073), 
            .I1(GND_net), .CO(n28155));
    SB_LUT4 encoder0_position_23__I_0_add_725_3_lut (.I0(GND_net), .I1(n1074), 
            .I2(VCC_net), .I3(n28153), .O(n1127)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_725_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_725_3 (.CI(n28153), .I0(n1074), 
            .I1(VCC_net), .CO(n28154));
    SB_LUT4 encoder0_position_23__I_0_add_725_2_lut (.I0(GND_net), .I1(n763), 
            .I2(GND_net), .I3(VCC_net), .O(n1128)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_725_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_725_2 (.CI(VCC_net), .I0(n763), 
            .I1(GND_net), .CO(n28153));
    SB_LUT4 encoder0_position_23__I_0_add_672_12_lut (.I0(GND_net), .I1(n986), 
            .I2(VCC_net), .I3(n28152), .O(n1039)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_672_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_23__I_0_add_672_11_lut (.I0(GND_net), .I1(n987), 
            .I2(VCC_net), .I3(n28151), .O(n1040)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_672_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_672_11 (.CI(n28151), .I0(n987), 
            .I1(VCC_net), .CO(n28152));
    SB_LUT4 encoder0_position_23__I_0_add_672_10_lut (.I0(GND_net), .I1(n988), 
            .I2(VCC_net), .I3(n28150), .O(n1041)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_672_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_672_10 (.CI(n28150), .I0(n988), 
            .I1(VCC_net), .CO(n28151));
    SB_LUT4 encoder0_position_23__I_0_add_672_9_lut (.I0(GND_net), .I1(n989), 
            .I2(VCC_net), .I3(n28149), .O(n1042)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_672_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_672_9 (.CI(n28149), .I0(n989), 
            .I1(VCC_net), .CO(n28150));
    SB_LUT4 encoder0_position_23__I_0_add_672_8_lut (.I0(GND_net), .I1(n990), 
            .I2(VCC_net), .I3(n28148), .O(n1043)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_672_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_672_8 (.CI(n28148), .I0(n990), 
            .I1(VCC_net), .CO(n28149));
    SB_LUT4 i14324_3_lut (.I0(Ki[9]), .I1(\data_in_frame[4] [1]), .I2(n33567), 
            .I3(GND_net), .O(n19466));   // verilog/coms.v(127[12] 300[6])
    defparam i14324_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mux_77_i8_4_lut (.I0(encoder1_position[7]), .I1(displacement[7]), 
            .I2(n15_adj_4934), .I3(n15_adj_4940), .O(motor_state_23__N_82[7]));   // verilog/TinyFPGA_B.v(166[5] 168[10])
    defparam mux_77_i8_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 encoder0_position_23__I_0_add_672_7_lut (.I0(GND_net), .I1(n991), 
            .I2(GND_net), .I3(n28147), .O(n1044)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_672_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_672_7 (.CI(n28147), .I0(n991), 
            .I1(GND_net), .CO(n28148));
    SB_LUT4 encoder0_position_23__I_0_add_672_6_lut (.I0(GND_net), .I1(n992), 
            .I2(GND_net), .I3(n28146), .O(n1045)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_672_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_25_15_lut (.I0(GND_net), .I1(delay_counter[13]), .I2(GND_net), 
            .I3(n27745), .O(n591)) /* synthesis syn_instantiated=1 */ ;
    defparam add_25_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_672_6 (.CI(n28146), .I0(n992), 
            .I1(GND_net), .CO(n28147));
    SB_LUT4 encoder0_position_23__I_0_add_672_5_lut (.I0(GND_net), .I1(n993), 
            .I2(VCC_net), .I3(n28145), .O(n1046)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_672_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_672_5 (.CI(n28145), .I0(n993), 
            .I1(VCC_net), .CO(n28146));
    SB_LUT4 encoder0_position_23__I_0_add_672_4_lut (.I0(GND_net), .I1(n994), 
            .I2(GND_net), .I3(n28144), .O(n1047)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_672_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i14325_3_lut (.I0(Ki[8]), .I1(\data_in_frame[4] [0]), .I2(n33567), 
            .I3(GND_net), .O(n19467));   // verilog/coms.v(127[12] 300[6])
    defparam i14325_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mux_77_i9_4_lut (.I0(encoder1_position[8]), .I1(displacement[8]), 
            .I2(n15_adj_4934), .I3(n15_adj_4940), .O(motor_state_23__N_82[8]));   // verilog/TinyFPGA_B.v(166[5] 168[10])
    defparam mux_77_i9_4_lut.LUT_INIT = 16'h0aca;
    SB_CARRY encoder0_position_23__I_0_add_672_4 (.CI(n28144), .I0(n994), 
            .I1(GND_net), .CO(n28145));
    SB_LUT4 encoder0_position_23__I_0_add_672_3_lut (.I0(GND_net), .I1(n995), 
            .I2(VCC_net), .I3(n28143), .O(n1048)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_672_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_672_3 (.CI(n28143), .I0(n995), 
            .I1(VCC_net), .CO(n28144));
    SB_LUT4 i14326_3_lut (.I0(Ki[7]), .I1(\data_in_frame[5] [7]), .I2(n33567), 
            .I3(GND_net), .O(n19468));   // verilog/coms.v(127[12] 300[6])
    defparam i14326_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_add_672_2_lut (.I0(GND_net), .I1(n519), 
            .I2(GND_net), .I3(VCC_net), .O(n1049)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_672_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_672_2 (.CI(VCC_net), .I0(n519), 
            .I1(GND_net), .CO(n28143));
    SB_LUT4 encoder0_position_23__I_0_add_619_11_lut (.I0(GND_net), .I1(n908), 
            .I2(VCC_net), .I3(n28142), .O(n961)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_619_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_25_15 (.CI(n27745), .I0(delay_counter[13]), .I1(GND_net), 
            .CO(n27746));
    SB_LUT4 i14327_3_lut (.I0(Ki[6]), .I1(\data_in_frame[5] [6]), .I2(n33567), 
            .I3(GND_net), .O(n19469));   // verilog/coms.v(127[12] 300[6])
    defparam i14327_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14328_3_lut (.I0(Ki[5]), .I1(\data_in_frame[5] [5]), .I2(n33567), 
            .I3(GND_net), .O(n19470));   // verilog/coms.v(127[12] 300[6])
    defparam i14328_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14329_3_lut (.I0(Ki[4]), .I1(\data_in_frame[5] [4]), .I2(n33567), 
            .I3(GND_net), .O(n19471));   // verilog/coms.v(127[12] 300[6])
    defparam i14329_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 add_25_14_lut (.I0(GND_net), .I1(delay_counter[12]), .I2(GND_net), 
            .I3(n27744), .O(n592)) /* synthesis syn_instantiated=1 */ ;
    defparam add_25_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_23__I_0_add_619_10_lut (.I0(GND_net), .I1(n909), 
            .I2(VCC_net), .I3(n28141), .O(n962)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_619_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_619_10 (.CI(n28141), .I0(n909), 
            .I1(VCC_net), .CO(n28142));
    SB_LUT4 i14330_3_lut (.I0(Ki[3]), .I1(\data_in_frame[5] [3]), .I2(n33567), 
            .I3(GND_net), .O(n19472));   // verilog/coms.v(127[12] 300[6])
    defparam i14330_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_add_619_9_lut (.I0(GND_net), .I1(n910), 
            .I2(VCC_net), .I3(n28140), .O(n963)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_619_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_619_9 (.CI(n28140), .I0(n910), 
            .I1(VCC_net), .CO(n28141));
    SB_LUT4 i14331_3_lut (.I0(Ki[2]), .I1(\data_in_frame[5] [2]), .I2(n33567), 
            .I3(GND_net), .O(n19473));   // verilog/coms.v(127[12] 300[6])
    defparam i14331_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i29834_3_lut_4_lut (.I0(\neo_pixel_transmitter.done ), .I1(state[0]), 
            .I2(n24759), .I3(start), .O(n36206));
    defparam i29834_3_lut_4_lut.LUT_INIT = 16'hff10;
    SB_LUT4 encoder1_position_23__I_0_inv_0_i19_1_lut (.I0(encoder0_position_scaled[18]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n7_adj_4947));   // verilog/TinyFPGA_B.v(202[21:65])
    defparam encoder1_position_23__I_0_inv_0_i19_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i14332_3_lut (.I0(Ki[1]), .I1(\data_in_frame[5] [1]), .I2(n33567), 
            .I3(GND_net), .O(n19474));   // verilog/coms.v(127[12] 300[6])
    defparam i14332_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i2_3_lut_4_lut_adj_1703 (.I0(\neo_pixel_transmitter.done ), .I1(state[0]), 
            .I2(n24759), .I3(state[1]), .O(n33926));
    defparam i2_3_lut_4_lut_adj_1703.LUT_INIT = 16'h0100;
    SB_LUT4 encoder1_position_23__I_0_inv_0_i20_1_lut (.I0(encoder0_position_scaled[19]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n6_adj_4946));   // verilog/TinyFPGA_B.v(202[21:65])
    defparam encoder1_position_23__I_0_inv_0_i20_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i14333_3_lut (.I0(Kp[15]), .I1(\data_in_frame[2] [7]), .I2(n33567), 
            .I3(GND_net), .O(n19475));   // verilog/coms.v(127[12] 300[6])
    defparam i14333_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_add_619_8_lut (.I0(GND_net), .I1(n911), 
            .I2(VCC_net), .I3(n28139), .O(n964)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_619_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_619_8 (.CI(n28139), .I0(n911), 
            .I1(VCC_net), .CO(n28140));
    SB_LUT4 i14334_3_lut (.I0(Kp[14]), .I1(\data_in_frame[2] [6]), .I2(n33567), 
            .I3(GND_net), .O(n19476));   // verilog/coms.v(127[12] 300[6])
    defparam i14334_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY add_25_6 (.CI(n27736), .I0(delay_counter[4]), .I1(GND_net), 
            .CO(n27737));
    SB_LUT4 encoder0_position_23__I_0_add_619_7_lut (.I0(GND_net), .I1(n912), 
            .I2(GND_net), .I3(n28138), .O(n965)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_619_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_619_7 (.CI(n28138), .I0(n912), 
            .I1(GND_net), .CO(n28139));
    SB_LUT4 encoder0_position_23__I_0_add_619_6_lut (.I0(GND_net), .I1(n913), 
            .I2(GND_net), .I3(n28137), .O(n966)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_619_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_619_6 (.CI(n28137), .I0(n913), 
            .I1(GND_net), .CO(n28138));
    SB_LUT4 encoder0_position_23__I_0_add_619_5_lut (.I0(GND_net), .I1(n914), 
            .I2(VCC_net), .I3(n28136), .O(n967)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_619_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_619_5 (.CI(n28136), .I0(n914), 
            .I1(VCC_net), .CO(n28137));
    SB_LUT4 encoder0_position_23__I_0_add_619_4_lut (.I0(GND_net), .I1(n915), 
            .I2(GND_net), .I3(n28135), .O(n968)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_619_4_lut.LUT_INIT = 16'hC33C;
    GND i1 (.Y(GND_net));
    SB_LUT4 mux_77_i10_4_lut (.I0(encoder1_position[9]), .I1(displacement[9]), 
            .I2(n15_adj_4934), .I3(n15_adj_4940), .O(motor_state_23__N_82[9]));   // verilog/TinyFPGA_B.v(166[5] 168[10])
    defparam mux_77_i10_4_lut.LUT_INIT = 16'h0aca;
    SB_CARRY add_25_14 (.CI(n27744), .I0(delay_counter[12]), .I1(GND_net), 
            .CO(n27745));
    SB_CARRY encoder0_position_23__I_0_add_619_4 (.CI(n28135), .I0(n915), 
            .I1(GND_net), .CO(n28136));
    SB_LUT4 encoder0_position_23__I_0_add_619_3_lut (.I0(GND_net), .I1(n916), 
            .I2(VCC_net), .I3(n28134), .O(n969)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_619_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_619_3 (.CI(n28134), .I0(n916), 
            .I1(VCC_net), .CO(n28135));
    SB_LUT4 encoder0_position_23__I_0_add_619_2_lut (.I0(GND_net), .I1(n518), 
            .I2(GND_net), .I3(VCC_net), .O(n970)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_619_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_619_2 (.CI(VCC_net), .I0(n518), 
            .I1(GND_net), .CO(n28134));
    SB_LUT4 encoder0_position_23__I_0_add_566_10_lut (.I0(GND_net), .I1(n830), 
            .I2(VCC_net), .I3(n28133), .O(n883)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_566_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_23__I_0_add_566_9_lut (.I0(GND_net), .I1(n831), 
            .I2(VCC_net), .I3(n28132), .O(n884)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_566_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_566_9 (.CI(n28132), .I0(n831), 
            .I1(VCC_net), .CO(n28133));
    SB_LUT4 encoder0_position_23__I_0_add_566_8_lut (.I0(GND_net), .I1(n832), 
            .I2(VCC_net), .I3(n28131), .O(n885)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_566_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_566_8 (.CI(n28131), .I0(n832), 
            .I1(VCC_net), .CO(n28132));
    SB_LUT4 i14335_3_lut (.I0(Kp[13]), .I1(\data_in_frame[2] [5]), .I2(n33567), 
            .I3(GND_net), .O(n19477));   // verilog/coms.v(127[12] 300[6])
    defparam i14335_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14336_3_lut (.I0(Kp[12]), .I1(\data_in_frame[2] [4]), .I2(n33567), 
            .I3(GND_net), .O(n19478));   // verilog/coms.v(127[12] 300[6])
    defparam i14336_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder1_position_23__I_0_inv_0_i21_1_lut (.I0(encoder0_position_scaled[20]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n5_adj_4945));   // verilog/TinyFPGA_B.v(202[21:65])
    defparam encoder1_position_23__I_0_inv_0_i21_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i14337_3_lut (.I0(Kp[11]), .I1(\data_in_frame[2] [3]), .I2(n33567), 
            .I3(GND_net), .O(n19479));   // verilog/coms.v(127[12] 300[6])
    defparam i14337_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14338_3_lut (.I0(Kp[10]), .I1(\data_in_frame[2] [2]), .I2(n33567), 
            .I3(GND_net), .O(n19480));   // verilog/coms.v(127[12] 300[6])
    defparam i14338_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14339_3_lut (.I0(Kp[9]), .I1(\data_in_frame[2] [1]), .I2(n33567), 
            .I3(GND_net), .O(n19481));   // verilog/coms.v(127[12] 300[6])
    defparam i14339_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14340_3_lut (.I0(Kp[8]), .I1(\data_in_frame[2] [0]), .I2(n33567), 
            .I3(GND_net), .O(n19482));   // verilog/coms.v(127[12] 300[6])
    defparam i14340_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14341_3_lut (.I0(Kp[7]), .I1(\data_in_frame[3] [7]), .I2(n33567), 
            .I3(GND_net), .O(n19483));   // verilog/coms.v(127[12] 300[6])
    defparam i14341_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14342_3_lut (.I0(Kp[6]), .I1(\data_in_frame[3] [6]), .I2(n33567), 
            .I3(GND_net), .O(n19484));   // verilog/coms.v(127[12] 300[6])
    defparam i14342_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14343_3_lut (.I0(Kp[5]), .I1(\data_in_frame[3] [5]), .I2(n33567), 
            .I3(GND_net), .O(n19485));   // verilog/coms.v(127[12] 300[6])
    defparam i14343_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14344_3_lut (.I0(Kp[4]), .I1(\data_in_frame[3] [4]), .I2(n33567), 
            .I3(GND_net), .O(n19486));   // verilog/coms.v(127[12] 300[6])
    defparam i14344_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14345_3_lut (.I0(Kp[3]), .I1(\data_in_frame[3] [3]), .I2(n33567), 
            .I3(GND_net), .O(n19487));   // verilog/coms.v(127[12] 300[6])
    defparam i14345_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14346_3_lut (.I0(Kp[2]), .I1(\data_in_frame[3] [2]), .I2(n33567), 
            .I3(GND_net), .O(n19488));   // verilog/coms.v(127[12] 300[6])
    defparam i14346_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14347_3_lut (.I0(Kp[1]), .I1(\data_in_frame[3] [1]), .I2(n33567), 
            .I3(GND_net), .O(n19489));   // verilog/coms.v(127[12] 300[6])
    defparam i14347_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14348_3_lut (.I0(\data_in[3] [7]), .I1(rx_data[7]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n19490));   // verilog/coms.v(127[12] 300[6])
    defparam i14348_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14349_3_lut (.I0(\data_in[3] [6]), .I1(rx_data[6]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n19491));   // verilog/coms.v(127[12] 300[6])
    defparam i14349_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14350_3_lut (.I0(\data_in[3] [5]), .I1(rx_data[5]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n19492));   // verilog/coms.v(127[12] 300[6])
    defparam i14350_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14351_3_lut (.I0(\data_in[3] [4]), .I1(rx_data[4]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n19493));   // verilog/coms.v(127[12] 300[6])
    defparam i14351_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14352_3_lut (.I0(\data_in[3] [3]), .I1(rx_data[3]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n19494));   // verilog/coms.v(127[12] 300[6])
    defparam i14352_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14353_3_lut (.I0(\data_in[3] [2]), .I1(rx_data[2]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n19495));   // verilog/coms.v(127[12] 300[6])
    defparam i14353_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14354_3_lut (.I0(\data_in[3] [1]), .I1(rx_data[1]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n19496));   // verilog/coms.v(127[12] 300[6])
    defparam i14354_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14355_3_lut (.I0(\data_in[3] [0]), .I1(rx_data[0]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n19497));   // verilog/coms.v(127[12] 300[6])
    defparam i14355_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14356_3_lut (.I0(\data_in[2] [7]), .I1(\data_in[3] [7]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n19498));   // verilog/coms.v(127[12] 300[6])
    defparam i14356_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14357_3_lut (.I0(\data_in[2] [6]), .I1(\data_in[3] [6]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n19499));   // verilog/coms.v(127[12] 300[6])
    defparam i14357_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14358_3_lut (.I0(\data_in[2] [5]), .I1(\data_in[3] [5]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n19500));   // verilog/coms.v(127[12] 300[6])
    defparam i14358_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14359_3_lut (.I0(\data_in[2] [4]), .I1(\data_in[3] [4]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n19501));   // verilog/coms.v(127[12] 300[6])
    defparam i14359_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14360_3_lut (.I0(\data_in[2] [3]), .I1(\data_in[3] [3]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n19502));   // verilog/coms.v(127[12] 300[6])
    defparam i14360_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14361_3_lut (.I0(\data_in[2] [2]), .I1(\data_in[3] [2]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n19503));   // verilog/coms.v(127[12] 300[6])
    defparam i14361_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14362_3_lut (.I0(\data_in[2] [1]), .I1(\data_in[3] [1]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n19504));   // verilog/coms.v(127[12] 300[6])
    defparam i14362_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14363_3_lut (.I0(\data_in[2] [0]), .I1(\data_in[3] [0]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n19505));   // verilog/coms.v(127[12] 300[6])
    defparam i14363_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14364_3_lut (.I0(\data_in[1] [7]), .I1(\data_in[2] [7]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n19506));   // verilog/coms.v(127[12] 300[6])
    defparam i14364_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14365_3_lut (.I0(\data_in[1] [6]), .I1(\data_in[2] [6]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n19507));   // verilog/coms.v(127[12] 300[6])
    defparam i14365_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14366_3_lut (.I0(\data_in[1] [5]), .I1(\data_in[2] [5]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n19508));   // verilog/coms.v(127[12] 300[6])
    defparam i14366_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14367_3_lut (.I0(\data_in[1] [4]), .I1(\data_in[2] [4]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n19509));   // verilog/coms.v(127[12] 300[6])
    defparam i14367_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14368_3_lut (.I0(\data_in[1] [3]), .I1(\data_in[2] [3]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n19510));   // verilog/coms.v(127[12] 300[6])
    defparam i14368_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_77_i11_4_lut (.I0(encoder1_position[10]), .I1(displacement[10]), 
            .I2(n15_adj_4934), .I3(n15_adj_4940), .O(motor_state_23__N_82[10]));   // verilog/TinyFPGA_B.v(166[5] 168[10])
    defparam mux_77_i11_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i14369_3_lut (.I0(\data_in[1] [2]), .I1(\data_in[2] [2]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n19511));   // verilog/coms.v(127[12] 300[6])
    defparam i14369_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14370_3_lut (.I0(\data_in[1] [1]), .I1(\data_in[2] [1]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n19512));   // verilog/coms.v(127[12] 300[6])
    defparam i14370_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_77_i12_4_lut (.I0(encoder1_position[11]), .I1(displacement[11]), 
            .I2(n15_adj_4934), .I3(n15_adj_4940), .O(motor_state_23__N_82[11]));   // verilog/TinyFPGA_B.v(166[5] 168[10])
    defparam mux_77_i12_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i14371_3_lut (.I0(\data_in[1] [0]), .I1(\data_in[2] [0]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n19513));   // verilog/coms.v(127[12] 300[6])
    defparam i14371_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14372_3_lut (.I0(\data_in[0] [7]), .I1(\data_in[1] [7]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n19514));   // verilog/coms.v(127[12] 300[6])
    defparam i14372_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14373_3_lut (.I0(\data_in[0] [6]), .I1(\data_in[1] [6]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n19515));   // verilog/coms.v(127[12] 300[6])
    defparam i14373_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14374_3_lut (.I0(\data_in[0] [5]), .I1(\data_in[1] [5]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n19516));   // verilog/coms.v(127[12] 300[6])
    defparam i14374_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14375_3_lut (.I0(\data_in[0] [4]), .I1(\data_in[1] [4]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n19517));   // verilog/coms.v(127[12] 300[6])
    defparam i14375_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder1_position_23__I_0_inv_0_i23_1_lut (.I0(encoder0_position_scaled[22]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n3_adj_4944));   // verilog/TinyFPGA_B.v(202[21:65])
    defparam encoder1_position_23__I_0_inv_0_i23_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mux_77_i13_4_lut (.I0(encoder1_position[12]), .I1(displacement[12]), 
            .I2(n15_adj_4934), .I3(n15_adj_4940), .O(motor_state_23__N_82[12]));   // verilog/TinyFPGA_B.v(166[5] 168[10])
    defparam mux_77_i13_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i14376_3_lut (.I0(\data_in[0] [3]), .I1(\data_in[1] [3]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n19518));   // verilog/coms.v(127[12] 300[6])
    defparam i14376_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14377_3_lut (.I0(\data_in[0] [2]), .I1(\data_in[1] [2]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n19519));   // verilog/coms.v(127[12] 300[6])
    defparam i14377_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14378_3_lut (.I0(\data_in[0] [1]), .I1(\data_in[1] [1]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n19520));   // verilog/coms.v(127[12] 300[6])
    defparam i14378_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14379_3_lut (.I0(\neo_pixel_transmitter.t0 [31]), .I1(timer[31]), 
            .I2(n34265), .I3(GND_net), .O(n19521));   // verilog/neopixel.v(35[12] 117[6])
    defparam i14379_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14383_3_lut (.I0(\neo_pixel_transmitter.t0 [30]), .I1(timer[30]), 
            .I2(n34265), .I3(GND_net), .O(n19525));   // verilog/neopixel.v(35[12] 117[6])
    defparam i14383_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mux_77_i14_4_lut (.I0(encoder1_position[13]), .I1(displacement[13]), 
            .I2(n15_adj_4934), .I3(n15_adj_4940), .O(motor_state_23__N_82[13]));   // verilog/TinyFPGA_B.v(166[5] 168[10])
    defparam mux_77_i14_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i14384_3_lut (.I0(\neo_pixel_transmitter.t0 [29]), .I1(timer[29]), 
            .I2(n34265), .I3(GND_net), .O(n19526));   // verilog/neopixel.v(35[12] 117[6])
    defparam i14384_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14385_3_lut (.I0(\neo_pixel_transmitter.t0 [28]), .I1(timer[28]), 
            .I2(n34265), .I3(GND_net), .O(n19527));   // verilog/neopixel.v(35[12] 117[6])
    defparam i14385_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14386_3_lut (.I0(\neo_pixel_transmitter.t0 [27]), .I1(timer[27]), 
            .I2(n34265), .I3(GND_net), .O(n19528));   // verilog/neopixel.v(35[12] 117[6])
    defparam i14386_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mux_77_i15_4_lut (.I0(encoder1_position[14]), .I1(displacement[14]), 
            .I2(n15_adj_4934), .I3(n15_adj_4940), .O(motor_state_23__N_82[14]));   // verilog/TinyFPGA_B.v(166[5] 168[10])
    defparam mux_77_i15_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i14387_3_lut (.I0(\neo_pixel_transmitter.t0 [26]), .I1(timer[26]), 
            .I2(n34265), .I3(GND_net), .O(n19529));   // verilog/neopixel.v(35[12] 117[6])
    defparam i14387_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14391_3_lut (.I0(\neo_pixel_transmitter.t0 [25]), .I1(timer[25]), 
            .I2(n34265), .I3(GND_net), .O(n19533));   // verilog/neopixel.v(35[12] 117[6])
    defparam i14391_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14392_3_lut (.I0(\neo_pixel_transmitter.t0 [24]), .I1(timer[24]), 
            .I2(n34265), .I3(GND_net), .O(n19534));   // verilog/neopixel.v(35[12] 117[6])
    defparam i14392_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14393_3_lut (.I0(\neo_pixel_transmitter.t0 [23]), .I1(timer[23]), 
            .I2(n34265), .I3(GND_net), .O(n19535));   // verilog/neopixel.v(35[12] 117[6])
    defparam i14393_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14394_3_lut (.I0(\neo_pixel_transmitter.t0 [22]), .I1(timer[22]), 
            .I2(n34265), .I3(GND_net), .O(n19536));   // verilog/neopixel.v(35[12] 117[6])
    defparam i14394_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mux_77_i16_4_lut (.I0(encoder1_position[15]), .I1(displacement[15]), 
            .I2(n15_adj_4934), .I3(n15_adj_4940), .O(motor_state_23__N_82[15]));   // verilog/TinyFPGA_B.v(166[5] 168[10])
    defparam mux_77_i16_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i14395_3_lut (.I0(\neo_pixel_transmitter.t0 [21]), .I1(timer[21]), 
            .I2(n34265), .I3(GND_net), .O(n19537));   // verilog/neopixel.v(35[12] 117[6])
    defparam i14395_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mux_77_i17_4_lut (.I0(encoder1_position[16]), .I1(displacement[16]), 
            .I2(n15_adj_4934), .I3(n15_adj_4940), .O(motor_state_23__N_82[16]));   // verilog/TinyFPGA_B.v(166[5] 168[10])
    defparam mux_77_i17_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i14396_3_lut (.I0(\neo_pixel_transmitter.t0 [20]), .I1(timer[20]), 
            .I2(n34265), .I3(GND_net), .O(n19538));   // verilog/neopixel.v(35[12] 117[6])
    defparam i14396_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14397_3_lut (.I0(\neo_pixel_transmitter.t0 [19]), .I1(timer[19]), 
            .I2(n34265), .I3(GND_net), .O(n19539));   // verilog/neopixel.v(35[12] 117[6])
    defparam i14397_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14398_3_lut (.I0(\neo_pixel_transmitter.t0 [18]), .I1(timer[18]), 
            .I2(n34265), .I3(GND_net), .O(n19540));   // verilog/neopixel.v(35[12] 117[6])
    defparam i14398_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14399_3_lut (.I0(\neo_pixel_transmitter.t0 [17]), .I1(timer[17]), 
            .I2(n34265), .I3(GND_net), .O(n19541));   // verilog/neopixel.v(35[12] 117[6])
    defparam i14399_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14400_3_lut (.I0(\neo_pixel_transmitter.t0 [16]), .I1(timer[16]), 
            .I2(n34265), .I3(GND_net), .O(n19542));   // verilog/neopixel.v(35[12] 117[6])
    defparam i14400_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14401_3_lut (.I0(\neo_pixel_transmitter.t0 [15]), .I1(timer[15]), 
            .I2(n34265), .I3(GND_net), .O(n19543));   // verilog/neopixel.v(35[12] 117[6])
    defparam i14401_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14402_3_lut (.I0(\neo_pixel_transmitter.t0 [14]), .I1(timer[14]), 
            .I2(n34265), .I3(GND_net), .O(n19544));   // verilog/neopixel.v(35[12] 117[6])
    defparam i14402_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14403_3_lut (.I0(\neo_pixel_transmitter.t0 [13]), .I1(timer[13]), 
            .I2(n34265), .I3(GND_net), .O(n19545));   // verilog/neopixel.v(35[12] 117[6])
    defparam i14403_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14404_3_lut (.I0(\neo_pixel_transmitter.t0 [12]), .I1(timer[12]), 
            .I2(n34265), .I3(GND_net), .O(n19546));   // verilog/neopixel.v(35[12] 117[6])
    defparam i14404_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mux_77_i18_4_lut (.I0(encoder1_position[17]), .I1(displacement[17]), 
            .I2(n15_adj_4934), .I3(n15_adj_4940), .O(motor_state_23__N_82[17]));   // verilog/TinyFPGA_B.v(166[5] 168[10])
    defparam mux_77_i18_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i14405_3_lut (.I0(\neo_pixel_transmitter.t0 [11]), .I1(timer[11]), 
            .I2(n34265), .I3(GND_net), .O(n19547));   // verilog/neopixel.v(35[12] 117[6])
    defparam i14405_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14406_3_lut (.I0(\neo_pixel_transmitter.t0 [10]), .I1(timer[10]), 
            .I2(n34265), .I3(GND_net), .O(n19548));   // verilog/neopixel.v(35[12] 117[6])
    defparam i14406_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mux_77_i19_4_lut (.I0(encoder1_position[18]), .I1(displacement[18]), 
            .I2(n15_adj_4934), .I3(n15_adj_4940), .O(motor_state_23__N_82[18]));   // verilog/TinyFPGA_B.v(166[5] 168[10])
    defparam mux_77_i19_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i14407_3_lut (.I0(\neo_pixel_transmitter.t0 [9]), .I1(timer[9]), 
            .I2(n34265), .I3(GND_net), .O(n19549));   // verilog/neopixel.v(35[12] 117[6])
    defparam i14407_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14408_3_lut (.I0(\neo_pixel_transmitter.t0 [8]), .I1(timer[8]), 
            .I2(n34265), .I3(GND_net), .O(n19550));   // verilog/neopixel.v(35[12] 117[6])
    defparam i14408_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14409_3_lut (.I0(\neo_pixel_transmitter.t0 [7]), .I1(timer[7]), 
            .I2(n34265), .I3(GND_net), .O(n19551));   // verilog/neopixel.v(35[12] 117[6])
    defparam i14409_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14410_3_lut (.I0(\neo_pixel_transmitter.t0 [6]), .I1(timer[6]), 
            .I2(n34265), .I3(GND_net), .O(n19552));   // verilog/neopixel.v(35[12] 117[6])
    defparam i14410_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14411_3_lut (.I0(\neo_pixel_transmitter.t0 [5]), .I1(timer[5]), 
            .I2(n34265), .I3(GND_net), .O(n19553));   // verilog/neopixel.v(35[12] 117[6])
    defparam i14411_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14412_3_lut (.I0(\neo_pixel_transmitter.t0 [4]), .I1(timer[4]), 
            .I2(n34265), .I3(GND_net), .O(n19554));   // verilog/neopixel.v(35[12] 117[6])
    defparam i14412_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14413_3_lut (.I0(\neo_pixel_transmitter.t0 [3]), .I1(timer[3]), 
            .I2(n34265), .I3(GND_net), .O(n19555));   // verilog/neopixel.v(35[12] 117[6])
    defparam i14413_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14414_3_lut (.I0(\neo_pixel_transmitter.t0 [2]), .I1(timer[2]), 
            .I2(n34265), .I3(GND_net), .O(n19556));   // verilog/neopixel.v(35[12] 117[6])
    defparam i14414_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mux_77_i20_4_lut (.I0(encoder1_position[19]), .I1(displacement[19]), 
            .I2(n15_adj_4934), .I3(n15_adj_4940), .O(motor_state_23__N_82[19]));   // verilog/TinyFPGA_B.v(166[5] 168[10])
    defparam mux_77_i20_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_77_i21_4_lut (.I0(encoder1_position[20]), .I1(displacement[20]), 
            .I2(n15_adj_4934), .I3(n15_adj_4940), .O(motor_state_23__N_82[20]));   // verilog/TinyFPGA_B.v(166[5] 168[10])
    defparam mux_77_i21_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i14415_3_lut (.I0(\neo_pixel_transmitter.t0 [1]), .I1(timer[1]), 
            .I2(n34265), .I3(GND_net), .O(n19557));   // verilog/neopixel.v(35[12] 117[6])
    defparam i14415_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mux_77_i22_4_lut (.I0(encoder1_position[21]), .I1(displacement[21]), 
            .I2(n15_adj_4934), .I3(n15_adj_4940), .O(motor_state_23__N_82[21]));   // verilog/TinyFPGA_B.v(166[5] 168[10])
    defparam mux_77_i22_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i14416_4_lut (.I0(state_7__N_3914[3]), .I1(data[4]), .I2(n4_adj_4941), 
            .I3(n17513), .O(n19558));   // verilog/i2c_controller.v(91[8] 173[6])
    defparam i14416_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i14417_3_lut (.I0(IntegralLimit[23]), .I1(\data_in_frame[11] [7]), 
            .I2(n33567), .I3(GND_net), .O(n19559));   // verilog/coms.v(127[12] 300[6])
    defparam i14417_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mux_77_i23_4_lut (.I0(encoder1_position[22]), .I1(displacement[22]), 
            .I2(n15_adj_4934), .I3(n15_adj_4940), .O(motor_state_23__N_82[22]));   // verilog/TinyFPGA_B.v(166[5] 168[10])
    defparam mux_77_i23_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i14418_3_lut (.I0(IntegralLimit[22]), .I1(\data_in_frame[11] [6]), 
            .I2(n33567), .I3(GND_net), .O(n19560));   // verilog/coms.v(127[12] 300[6])
    defparam i14418_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14419_3_lut (.I0(IntegralLimit[21]), .I1(\data_in_frame[11] [5]), 
            .I2(n33567), .I3(GND_net), .O(n19561));   // verilog/coms.v(127[12] 300[6])
    defparam i14419_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i4_4_lut_adj_1704 (.I0(control_mode[3]), .I1(control_mode[5]), 
            .I2(control_mode[4]), .I3(control_mode[7]), .O(n10_adj_5066));   // verilog/TinyFPGA_B.v(165[5:22])
    defparam i4_4_lut_adj_1704.LUT_INIT = 16'hfffe;
    SB_LUT4 i5_3_lut_adj_1705 (.I0(control_mode[6]), .I1(n10_adj_5066), 
            .I2(control_mode[2]), .I3(GND_net), .O(n17506));   // verilog/TinyFPGA_B.v(165[5:22])
    defparam i5_3_lut_adj_1705.LUT_INIT = 16'hfefe;
    SB_LUT4 i1_2_lut_adj_1706 (.I0(n17355), .I1(control_mode[1]), .I2(GND_net), 
            .I3(GND_net), .O(n15_adj_4940));   // verilog/TinyFPGA_B.v(167[5:22])
    defparam i1_2_lut_adj_1706.LUT_INIT = 16'hbbbb;
    SB_LUT4 i14420_3_lut (.I0(IntegralLimit[20]), .I1(\data_in_frame[11] [4]), 
            .I2(n33567), .I3(GND_net), .O(n19562));   // verilog/coms.v(127[12] 300[6])
    defparam i14420_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i2_3_lut_adj_1707 (.I0(control_mode[0]), .I1(control_mode[1]), 
            .I2(n17506), .I3(GND_net), .O(n15_adj_4934));   // verilog/TinyFPGA_B.v(166[5:22])
    defparam i2_3_lut_adj_1707.LUT_INIT = 16'hfdfd;
    SB_LUT4 mux_77_i24_4_lut (.I0(encoder1_position[23]), .I1(displacement[23]), 
            .I2(n15_adj_4934), .I3(n15_adj_4940), .O(motor_state_23__N_82[23]));   // verilog/TinyFPGA_B.v(166[5] 168[10])
    defparam mux_77_i24_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i14421_3_lut (.I0(IntegralLimit[19]), .I1(\data_in_frame[11] [3]), 
            .I2(n33567), .I3(GND_net), .O(n19563));   // verilog/coms.v(127[12] 300[6])
    defparam i14421_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14422_3_lut (.I0(IntegralLimit[18]), .I1(\data_in_frame[11] [2]), 
            .I2(n33567), .I3(GND_net), .O(n19564));   // verilog/coms.v(127[12] 300[6])
    defparam i14422_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14423_3_lut (.I0(IntegralLimit[17]), .I1(\data_in_frame[11] [1]), 
            .I2(n33567), .I3(GND_net), .O(n19565));   // verilog/coms.v(127[12] 300[6])
    defparam i14423_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14424_3_lut (.I0(IntegralLimit[16]), .I1(\data_in_frame[11] [0]), 
            .I2(n33567), .I3(GND_net), .O(n19566));   // verilog/coms.v(127[12] 300[6])
    defparam i14424_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14425_3_lut (.I0(IntegralLimit[15]), .I1(\data_in_frame[12] [7]), 
            .I2(n33567), .I3(GND_net), .O(n19567));   // verilog/coms.v(127[12] 300[6])
    defparam i14425_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14426_3_lut (.I0(IntegralLimit[14]), .I1(\data_in_frame[12] [6]), 
            .I2(n33567), .I3(GND_net), .O(n19568));   // verilog/coms.v(127[12] 300[6])
    defparam i14426_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i463_3_lut (.I0(n675), .I1(n728), 
            .I2(n700), .I3(GND_net), .O(n753));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i463_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14427_3_lut (.I0(IntegralLimit[13]), .I1(\data_in_frame[12] [5]), 
            .I2(n33567), .I3(GND_net), .O(n19569));   // verilog/coms.v(127[12] 300[6])
    defparam i14427_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mux_3363_i19_3_lut (.I0(encoder0_position[18]), .I1(n7_adj_4920), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n598_adj_4967));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam mux_3363_i19_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14428_3_lut (.I0(IntegralLimit[12]), .I1(\data_in_frame[12] [4]), 
            .I2(n33567), .I3(GND_net), .O(n19570));   // verilog/coms.v(127[12] 300[6])
    defparam i14428_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_adj_1708 (.I0(n598_adj_4967), .I1(n6_adj_4921), .I2(GND_net), 
            .I3(GND_net), .O(n7));
    defparam i1_2_lut_adj_1708.LUT_INIT = 16'heeee;
    SB_LUT4 i14429_3_lut (.I0(IntegralLimit[11]), .I1(\data_in_frame[12] [3]), 
            .I2(n33567), .I3(GND_net), .O(n19571));   // verilog/coms.v(127[12] 300[6])
    defparam i14429_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_1709 (.I0(n4_adj_4923), .I1(n2), .I2(n5_adj_4922), 
            .I3(n7), .O(n4_adj_4970));
    defparam i1_4_lut_adj_1709.LUT_INIT = 16'hc888;
    SB_LUT4 i14430_3_lut (.I0(IntegralLimit[10]), .I1(\data_in_frame[12] [2]), 
            .I2(n33567), .I3(GND_net), .O(n19572));   // verilog/coms.v(127[12] 300[6])
    defparam i14430_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14431_3_lut (.I0(IntegralLimit[9]), .I1(\data_in_frame[12] [1]), 
            .I2(n33567), .I3(GND_net), .O(n19573));   // verilog/coms.v(127[12] 300[6])
    defparam i14431_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14432_3_lut (.I0(IntegralLimit[8]), .I1(\data_in_frame[12] [0]), 
            .I2(n33567), .I3(GND_net), .O(n19574));   // verilog/coms.v(127[12] 300[6])
    defparam i14432_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14433_3_lut (.I0(IntegralLimit[7]), .I1(\data_in_frame[13] [7]), 
            .I2(n33567), .I3(GND_net), .O(n19575));   // verilog/coms.v(127[12] 300[6])
    defparam i14433_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i30196_3_lut (.I0(n37058), .I1(pwm_setpoint[22]), .I2(pwm_counter[22]), 
            .I3(GND_net), .O(n36951));   // verilog/pwm.v(21[8:24])
    defparam i30196_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i14434_3_lut (.I0(IntegralLimit[6]), .I1(\data_in_frame[13] [6]), 
            .I2(n33567), .I3(GND_net), .O(n19576));   // verilog/coms.v(127[12] 300[6])
    defparam i14434_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14435_3_lut (.I0(IntegralLimit[5]), .I1(\data_in_frame[13] [5]), 
            .I2(n33567), .I3(GND_net), .O(n19577));   // verilog/coms.v(127[12] 300[6])
    defparam i14435_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i3688_2_lut (.I0(n2), .I1(encoder0_position[23]), .I2(GND_net), 
            .I3(GND_net), .O(n509));
    defparam i3688_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i14436_3_lut (.I0(IntegralLimit[4]), .I1(\data_in_frame[13] [4]), 
            .I2(n33567), .I3(GND_net), .O(n19578));   // verilog/coms.v(127[12] 300[6])
    defparam i14436_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i26629_4_lut (.I0(encoder0_position[22]), .I1(n36211), .I2(encoder0_position[23]), 
            .I3(n3_adj_4924), .O(n675));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam i26629_4_lut.LUT_INIT = 16'hca0a;
    SB_LUT4 i14437_3_lut (.I0(IntegralLimit[3]), .I1(\data_in_frame[13] [3]), 
            .I2(n33567), .I3(GND_net), .O(n19579));   // verilog/coms.v(127[12] 300[6])
    defparam i14437_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14438_3_lut (.I0(IntegralLimit[2]), .I1(\data_in_frame[13] [2]), 
            .I2(n33567), .I3(GND_net), .O(n19580));   // verilog/coms.v(127[12] 300[6])
    defparam i14438_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14439_3_lut (.I0(IntegralLimit[1]), .I1(\data_in_frame[13] [1]), 
            .I2(n33567), .I3(GND_net), .O(n19581));   // verilog/coms.v(127[12] 300[6])
    defparam i14439_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14440_4_lut (.I0(state_7__N_3914[3]), .I1(data[3]), .I2(n4_adj_4942), 
            .I3(n17518), .O(n19582));   // verilog/i2c_controller.v(91[8] 173[6])
    defparam i14440_4_lut.LUT_INIT = 16'hccca;
    motorControl control (.GND_net(GND_net), .\Kp[2] (Kp[2]), .\Kp[3] (Kp[3]), 
            .\Ki[0] (Ki[0]), .\Kp[0] (Kp[0]), .\Kp[4] (Kp[4]), .\Kp[5] (Kp[5]), 
            .\Kp[6] (Kp[6]), .\Kp[7] (Kp[7]), .\Kp[8] (Kp[8]), .\Kp[9] (Kp[9]), 
            .\Kp[10] (Kp[10]), .\Kp[11] (Kp[11]), .\Kp[12] (Kp[12]), .\Kp[13] (Kp[13]), 
            .\Kp[14] (Kp[14]), .\Kp[15] (Kp[15]), .\Kp[1] (Kp[1]), .PWMLimit({PWMLimit}), 
            .IntegralLimit({IntegralLimit}), .\Ki[1] (Ki[1]), .\Ki[2] (Ki[2]), 
            .\Ki[3] (Ki[3]), .\Ki[4] (Ki[4]), .\Ki[5] (Ki[5]), .\Ki[6] (Ki[6]), 
            .\Ki[7] (Ki[7]), .\Ki[8] (Ki[8]), .\Ki[9] (Ki[9]), .\Ki[10] (Ki[10]), 
            .\Ki[11] (Ki[11]), .duty({duty}), .clk32MHz(clk32MHz), .\Ki[12] (Ki[12]), 
            .\Ki[13] (Ki[13]), .\Ki[14] (Ki[14]), .\Ki[15] (Ki[15]), .VCC_net(VCC_net), 
            .setpoint({setpoint}), .motor_state({motor_state}), .n37633(n37633)) /* synthesis syn_module_defined=1 */ ;   // verilog/TinyFPGA_B.v(170[16] 182[4])
    SB_LUT4 i14441_4_lut (.I0(r_Rx_Data), .I1(rx_data[0]), .I2(n4_adj_4928), 
            .I3(n17534), .O(n19583));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i14441_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i14442_4_lut (.I0(state_7__N_3914[3]), .I1(data[2]), .I2(n4_adj_4942), 
            .I3(n17513), .O(n19584));   // verilog/i2c_controller.v(91[8] 173[6])
    defparam i14442_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i14446_3_lut (.I0(quadA_debounced), .I1(reg_B[1]), .I2(n35256), 
            .I3(GND_net), .O(n19588));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(186[9] 190[16])
    defparam i14446_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14450_4_lut (.I0(state_7__N_3914[3]), .I1(data[1]), .I2(n10_adj_5076), 
            .I3(n17518), .O(n19592));   // verilog/i2c_controller.v(91[8] 173[6])
    defparam i14450_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i14451_3_lut (.I0(quadA_debounced_adj_4926), .I1(reg_B_adj_5146[1]), 
            .I2(n35209), .I3(GND_net), .O(n19593));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(186[9] 190[16])
    defparam i14451_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14452_3_lut (.I0(ID[1]), .I1(data[1]), .I2(n35211), .I3(GND_net), 
            .O(n19594));   // verilog/TinyFPGA_B.v(237[10] 265[6])
    defparam i14452_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14453_3_lut (.I0(ID[2]), .I1(data[2]), .I2(n35211), .I3(GND_net), 
            .O(n19595));   // verilog/TinyFPGA_B.v(237[10] 265[6])
    defparam i14453_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14454_3_lut (.I0(ID[3]), .I1(data[3]), .I2(n35211), .I3(GND_net), 
            .O(n19596));   // verilog/TinyFPGA_B.v(237[10] 265[6])
    defparam i14454_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14455_3_lut (.I0(ID[4]), .I1(data[4]), .I2(n35211), .I3(GND_net), 
            .O(n19597));   // verilog/TinyFPGA_B.v(237[10] 265[6])
    defparam i14455_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14456_3_lut (.I0(ID[5]), .I1(data[5]), .I2(n35211), .I3(GND_net), 
            .O(n19598));   // verilog/TinyFPGA_B.v(237[10] 265[6])
    defparam i14456_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14457_3_lut (.I0(ID[6]), .I1(data[6]), .I2(n35211), .I3(GND_net), 
            .O(n19599));   // verilog/TinyFPGA_B.v(237[10] 265[6])
    defparam i14457_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14458_3_lut (.I0(ID[7]), .I1(data[7]), .I2(n35211), .I3(GND_net), 
            .O(n19600));   // verilog/TinyFPGA_B.v(237[10] 265[6])
    defparam i14458_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12_4_lut_adj_1710 (.I0(n5592), .I1(DE_c), .I2(n17504), .I3(n17474), 
            .O(n32173));   // verilog/coms.v(127[12] 300[6])
    defparam i12_4_lut_adj_1710.LUT_INIT = 16'hc0ca;
    SB_LUT4 i29801_4_lut (.I0(n5_adj_4966), .I1(n6_adj_5030), .I2(n5523), 
            .I3(n1247), .O(n36263));   // verilog/TinyFPGA_B.v(237[10] 265[6])
    defparam i29801_4_lut.LUT_INIT = 16'h080c;
    SB_LUT4 i49_4_lut (.I0(n36263), .I1(data_ready), .I2(\ID_READOUT_FSM.state [0]), 
            .I3(n5523), .O(n31783));   // verilog/TinyFPGA_B.v(237[10] 265[6])
    defparam i49_4_lut.LUT_INIT = 16'hfa3a;
    SB_LUT4 i14382_3_lut (.I0(n18954), .I1(r_Bit_Index[0]), .I2(n18732), 
            .I3(GND_net), .O(n19524));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i14382_3_lut.LUT_INIT = 16'h1414;
    SB_LUT4 i14318_3_lut (.I0(n18956), .I1(r_Bit_Index_adj_5137[0]), .I2(n18738), 
            .I3(GND_net), .O(n19460));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i14318_3_lut.LUT_INIT = 16'h1414;
    SB_LUT4 i1_4_lut_adj_1711 (.I0(n24036), .I1(n33535), .I2(state_adj_5128[0]), 
            .I3(read), .O(n32323));   // verilog/eeprom.v(26[8] 58[4])
    defparam i1_4_lut_adj_1711.LUT_INIT = 16'h8280;
    SB_LUT4 i266_2_lut (.I0(n691), .I1(n17358), .I2(GND_net), .I3(GND_net), 
            .O(n1247));   // verilog/TinyFPGA_B.v(256[9] 262[12])
    defparam i266_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i1_4_lut_adj_1712 (.I0(n5_adj_4966), .I1(\ID_READOUT_FSM.state [0]), 
            .I2(n1247), .I3(read_N_295), .O(n25_adj_4894));   // verilog/TinyFPGA_B.v(237[10] 265[6])
    defparam i1_4_lut_adj_1712.LUT_INIT = 16'h7350;
    SB_LUT4 i28595_2_lut (.I0(data_ready), .I1(\ID_READOUT_FSM.state [0]), 
            .I2(GND_net), .I3(GND_net), .O(n35348));
    defparam i28595_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i30504_4_lut (.I0(\ID_READOUT_FSM.state [1]), .I1(n5523), .I2(n35348), 
            .I3(n25_adj_4894), .O(n17_adj_4895));   // verilog/TinyFPGA_B.v(237[10] 265[6])
    defparam i30504_4_lut.LUT_INIT = 16'h88ba;
    SB_LUT4 i26723_4_lut (.I0(n7_adj_4972), .I1(state_adj_5128[0]), .I2(n6_adj_4932), 
            .I3(state_adj_5158[0]), .O(n33471));
    defparam i26723_4_lut.LUT_INIT = 16'hccc8;
    SB_LUT4 i1_3_lut_adj_1713 (.I0(state_adj_5128[1]), .I1(read), .I2(n33535), 
            .I3(GND_net), .O(n12_adj_4901));   // verilog/eeprom.v(26[8] 58[4])
    defparam i1_3_lut_adj_1713.LUT_INIT = 16'ha2a2;
    SB_LUT4 i1_4_lut_adj_1714 (.I0(n24036), .I1(n12_adj_4901), .I2(state_adj_5128[0]), 
            .I3(n33535), .O(n32331));   // verilog/eeprom.v(26[8] 58[4])
    defparam i1_4_lut_adj_1714.LUT_INIT = 16'h88a8;
    SB_LUT4 i13898_4_lut (.I0(n33425), .I1(state[1]), .I2(state_3__N_402[1]), 
            .I3(n18685), .O(n19040));   // verilog/neopixel.v(35[12] 117[6])
    defparam i13898_4_lut.LUT_INIT = 16'hfaee;
    SB_LUT4 unary_minus_4_inv_0_i6_1_lut (.I0(duty[5]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n20));   // verilog/TinyFPGA_B.v(106[23:28])
    defparam unary_minus_4_inv_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i13899_3_lut (.I0(\data_in[0] [0]), .I1(\data_in[1] [0]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n19041));   // verilog/coms.v(127[12] 300[6])
    defparam i13899_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13900_3_lut (.I0(Kp[0]), .I1(\data_in_frame[3] [0]), .I2(n33567), 
            .I3(GND_net), .O(n19042));   // verilog/coms.v(127[12] 300[6])
    defparam i13900_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13901_3_lut (.I0(Ki[0]), .I1(\data_in_frame[5] [0]), .I2(n33567), 
            .I3(GND_net), .O(n19043));   // verilog/coms.v(127[12] 300[6])
    defparam i13901_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13902_3_lut (.I0(neopxl_color[0]), .I1(\data_in_frame[6] [0]), 
            .I2(n3_adj_4943), .I3(GND_net), .O(n19044));   // verilog/coms.v(127[12] 300[6])
    defparam i13902_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i26627_3_lut (.I0(encoder0_position[21]), .I1(n33367), .I2(encoder0_position[23]), 
            .I3(GND_net), .O(n676));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam i26627_3_lut.LUT_INIT = 16'hcaca;
    coms neopxl_color_23__I_0 (.n63(n63_adj_4971), .n771(n771), .n10417(n10417), 
         .GND_net(GND_net), .\data_out_frame[19] ({\data_out_frame[19] }), 
         .\data_out_frame[23] ({\data_out_frame[23] }), .\data_out_frame[24] ({\data_out_frame[24] }), 
         .\data_out_frame[17] ({\data_out_frame[17] }), .n3303(n3303), .n123(n123), 
         .\FRAME_MATCHER.state_31__N_2662[1] (\FRAME_MATCHER.state_31__N_2662 [1]), 
         .clk32MHz(clk32MHz), .\data_out_frame[15] ({\data_out_frame[15] }), 
         .\data_out_frame[20] ({\data_out_frame[20] }), .\data_out_frame[13] ({\data_out_frame[13] }), 
         .\data_in_frame[4] ({\data_in_frame[4] }), .\data_in_frame[1] ({\data_in_frame[1] }), 
         .\data_out_frame[18] ({\data_out_frame[18] }), .\data_out_frame[25] ({\data_out_frame[25] }), 
         .\data_out_frame[16] ({\data_out_frame[16] }), .\data_in_frame[3] ({\data_in_frame[3] }), 
         .\data_out_frame[10] ({\data_out_frame[10] }), .\data_out_frame[8] ({\data_out_frame[8] }), 
         .\data_out_frame[6] ({\data_out_frame[6] }), .\data_out_frame[12] ({\data_out_frame[12] }), 
         .n33567(n33567), .\data_out_frame[11] ({\data_out_frame[11] }), 
         .\data_out_frame[5] ({\data_out_frame[5] }), .\data_out_frame[14] ({\data_out_frame[14] }), 
         .\data_out_frame[7] ({\data_out_frame[7] }), .\data_in_frame[13] ({\data_in_frame[13] }), 
         .\data_in_frame[9] ({\data_in_frame[9] }), .\data_out_frame[9] ({\data_out_frame[9] }), 
         .\data_out_frame[4] ({\data_out_frame[4] }), .\data_in_frame[6] ({\data_in_frame[6] }), 
         .\data_in_frame[5] ({\data_in_frame[5] }), .\data_in_frame[8] ({\data_in_frame[8] }), 
         .rx_data({rx_data}), .\data_in_frame[12] ({\data_in_frame[12] }), 
         .\FRAME_MATCHER.state ({Open_0, Open_1, Open_2, Open_3, Open_4, 
         Open_5, Open_6, Open_7, Open_8, Open_9, Open_10, Open_11, 
         Open_12, Open_13, Open_14, Open_15, Open_16, Open_17, Open_18, 
         Open_19, Open_20, Open_21, Open_22, Open_23, Open_24, Open_25, 
         Open_26, Open_27, \FRAME_MATCHER.state [3], Open_28, Open_29, 
         Open_30}), .\data_in_frame[2] ({\data_in_frame[2] }), .\FRAME_MATCHER.state[0] (\FRAME_MATCHER.state [0]), 
         .n63_adj_8(n63), .n2970(n2970), .n14711(n14711), .n39(n39), 
         .\data_in[1] ({\data_in[1] }), .\data_in[0] ({\data_in[0] }), .\data_in[3] ({\data_in[3] }), 
         .\data_in[2] ({\data_in[2] }), .n4452(n4452), .\data_in_frame[10] ({\data_in_frame[10] }), 
         .\data_in_frame[11] ({\data_in_frame[11] }), .rx_data_ready(rx_data_ready), 
         .setpoint({setpoint}), .\state[2] (state_adj_5158[2]), .\state[3] (state_adj_5158[3]), 
         .n10(n10), .\data_in_frame[21] ({\data_in_frame[21] }), .n3(n3_adj_4943), 
         .n7(n7_adj_5045), .ID({ID}), .n17474(n17474), .n17552(n17552), 
         .n17476(n17476), .n5592(n5592), .tx_active(tx_active), .n19101(n19101), 
         .n19100(n19100), .n19099(n19099), .n19098(n19098), .n19097(n19097), 
         .n19096(n19096), .n19095(n19095), .n19094(n19094), .n19093(n19093), 
         .control_mode({control_mode}), .n19092(n19092), .n19091(n19091), 
         .n19090(n19090), .n19089(n19089), .n19088(n19088), .n19087(n19087), 
         .n19086(n19086), .PWMLimit({PWMLimit}), .n19085(n19085), .n19084(n19084), 
         .n19083(n19083), .n19082(n19082), .n19081(n19081), .n19080(n19080), 
         .n19079(n19079), .n19078(n19078), .n19077(n19077), .n19076(n19076), 
         .n19075(n19075), .n19074(n19074), .n19073(n19073), .n19072(n19072), 
         .n19071(n19071), .n19070(n19070), .n19069(n19069), .n19068(n19068), 
         .n19067(n19067), .n19066(n19066), .n19065(n19065), .n19064(n19064), 
         .n38205(n38205), .n38206(n38206), .n32009(n32009), .n19047(n19047), 
         .n19046(n19046), .n19044(n19044), .neopxl_color({neopxl_color}), 
         .LED_c(LED_c), .n19043(n19043), .\Ki[0] (Ki[0]), .n19042(n19042), 
         .\Kp[0] (Kp[0]), .n19041(n19041), .n32173(n32173), .DE_c(DE_c), 
         .n19581(n19581), .IntegralLimit({IntegralLimit}), .n19580(n19580), 
         .n19579(n19579), .n19578(n19578), .n19577(n19577), .n19576(n19576), 
         .n19575(n19575), .n19574(n19574), .n19573(n19573), .n19572(n19572), 
         .n19571(n19571), .n19570(n19570), .n19569(n19569), .n19568(n19568), 
         .n19567(n19567), .n19566(n19566), .n19565(n19565), .n19564(n19564), 
         .n19563(n19563), .n19562(n19562), .n19561(n19561), .n19560(n19560), 
         .n19559(n19559), .n19520(n19520), .n19519(n19519), .n19518(n19518), 
         .n19517(n19517), .n19516(n19516), .n19515(n19515), .n19514(n19514), 
         .n19513(n19513), .n19512(n19512), .n19511(n19511), .n19510(n19510), 
         .n19509(n19509), .n19508(n19508), .n19507(n19507), .n19506(n19506), 
         .n19505(n19505), .n19504(n19504), .n19503(n19503), .n19502(n19502), 
         .n19501(n19501), .n19500(n19500), .n19499(n19499), .n19498(n19498), 
         .n19497(n19497), .n19496(n19496), .n19495(n19495), .n19494(n19494), 
         .n19493(n19493), .n19492(n19492), .n19491(n19491), .n19490(n19490), 
         .n19489(n19489), .\Kp[1] (Kp[1]), .n19488(n19488), .\Kp[2] (Kp[2]), 
         .n19487(n19487), .\Kp[3] (Kp[3]), .n19486(n19486), .\Kp[4] (Kp[4]), 
         .n19485(n19485), .\Kp[5] (Kp[5]), .n19484(n19484), .\Kp[6] (Kp[6]), 
         .n19483(n19483), .\Kp[7] (Kp[7]), .n19482(n19482), .\Kp[8] (Kp[8]), 
         .n19481(n19481), .\Kp[9] (Kp[9]), .n19480(n19480), .\Kp[10] (Kp[10]), 
         .n19479(n19479), .\Kp[11] (Kp[11]), .n19478(n19478), .\Kp[12] (Kp[12]), 
         .n19477(n19477), .\Kp[13] (Kp[13]), .n19476(n19476), .\Kp[14] (Kp[14]), 
         .n19475(n19475), .\Kp[15] (Kp[15]), .n19474(n19474), .\Ki[1] (Ki[1]), 
         .n19473(n19473), .\Ki[2] (Ki[2]), .n19472(n19472), .\Ki[3] (Ki[3]), 
         .n19471(n19471), .\Ki[4] (Ki[4]), .n19470(n19470), .\Ki[5] (Ki[5]), 
         .n19469(n19469), .\Ki[6] (Ki[6]), .n19468(n19468), .\Ki[7] (Ki[7]), 
         .n19467(n19467), .\Ki[8] (Ki[8]), .n19466(n19466), .\Ki[9] (Ki[9]), 
         .n19465(n19465), .\Ki[10] (Ki[10]), .n19464(n19464), .\Ki[11] (Ki[11]), 
         .n19463(n19463), .\Ki[12] (Ki[12]), .n19462(n19462), .\Ki[13] (Ki[13]), 
         .n19461(n19461), .\Ki[14] (Ki[14]), .n19452(n19452), .\Ki[15] (Ki[15]), 
         .n19451(n19451), .n19450(n19450), .n19449(n19449), .n19448(n19448), 
         .n19447(n19447), .n19446(n19446), .n19445(n19445), .n19444(n19444), 
         .n19443(n19443), .n19442(n19442), .n19441(n19441), .n19440(n19440), 
         .n19439(n19439), .n19438(n19438), .n19437(n19437), .n19436(n19436), 
         .n19435(n19435), .n19434(n19434), .n19433(n19433), .n19432(n19432), 
         .n19431(n19431), .n19430(n19430), .n19429(n19429), .n19428(n19428), 
         .n19427(n19427), .n19426(n19426), .n19425(n19425), .n19424(n19424), 
         .n19423(n19423), .n19422(n19422), .n19421(n19421), .n19420(n19420), 
         .n19419(n19419), .n19418(n19418), .n19417(n19417), .n19416(n19416), 
         .n19415(n19415), .n19414(n19414), .n19413(n19413), .n19412(n19412), 
         .n19411(n19411), .n19410(n19410), .n19409(n19409), .n19408(n19408), 
         .n19407(n19407), .n19406(n19406), .n19405(n19405), .n19404(n19404), 
         .n19403(n19403), .n19402(n19402), .n19401(n19401), .n19400(n19400), 
         .n19399(n19399), .n19398(n19398), .n19397(n19397), .n19396(n19396), 
         .n19395(n19395), .n19394(n19394), .n19393(n19393), .n19392(n19392), 
         .n19391(n19391), .n19390(n19390), .n19389(n19389), .n19388(n19388), 
         .n19387(n19387), .n19386(n19386), .n19385(n19385), .n19384(n19384), 
         .n19383(n19383), .\state[0] (state_adj_5158[0]), .n5690(n5690), 
         .n19382(n19382), .n19381(n19381), .n32(n32_adj_5070), .n19380(n19380), 
         .n19379(n19379), .n19378(n19378), .n19377(n19377), .n19376(n19376), 
         .n19375(n19375), .n19374(n19374), .n19373(n19373), .n19372(n19372), 
         .n19371(n19371), .n19370(n19370), .n19369(n19369), .n19368(n19368), 
         .n19367(n19367), .n19366(n19366), .n19365(n19365), .n19364(n19364), 
         .n19363(n19363), .n19362(n19362), .n19361(n19361), .n19360(n19360), 
         .n19359(n19359), .n19358(n19358), .n19357(n19357), .n19356(n19356), 
         .n19355(n19355), .n19354(n19354), .n19353(n19353), .n19352(n19352), 
         .n19351(n19351), .n19350(n19350), .n19349(n19349), .n19348(n19348), 
         .n19347(n19347), .n19346(n19346), .n19345(n19345), .n19344(n19344), 
         .n19343(n19343), .n19342(n19342), .n19341(n19341), .n19340(n19340), 
         .n19339(n19339), .n19338(n19338), .n19337(n19337), .n19336(n19336), 
         .n19335(n19335), .n19334(n19334), .n19333(n19333), .n19332(n19332), 
         .n19331(n19331), .n19330(n19330), .n19329(n19329), .n19328(n19328), 
         .n19327(n19327), .n19326(n19326), .n19325(n19325), .n19324(n19324), 
         .n19323(n19323), .n19322(n19322), .n19321(n19321), .n19320(n19320), 
         .n19319(n19319), .n19318(n19318), .n19317(n19317), .n19316(n19316), 
         .n19315(n19315), .n19314(n19314), .n19313(n19313), .n19312(n19312), 
         .n19023(n19023), .n19311(n19311), .n19310(n19310), .n19309(n19309), 
         .n19308(n19308), .n19307(n19307), .n19306(n19306), .n19305(n19305), 
         .n19304(n19304), .n19303(n19303), .n19302(n19302), .n19301(n19301), 
         .n19300(n19300), .n19299(n19299), .n19298(n19298), .n19297(n19297), 
         .n19296(n19296), .n19295(n19295), .n19294(n19294), .n19293(n19293), 
         .n19292(n19292), .n19291(n19291), .n19290(n19290), .n19289(n19289), 
         .n19288(n19288), .n19287(n19287), .n19286(n19286), .n19285(n19285), 
         .n19284(n19284), .n19283(n19283), .n19282(n19282), .n19281(n19281), 
         .n19280(n19280), .n19279(n19279), .n19278(n19278), .n19277(n19277), 
         .n19276(n19276), .n19275(n19275), .n19274(n19274), .n14867(n14867), 
         .n19273(n19273), .n19272(n19272), .n19271(n19271), .n19270(n19270), 
         .n19269(n19269), .n19229(n19229), .n19228(n19228), .n19227(n19227), 
         .n19226(n19226), .n19225(n19225), .n19224(n19224), .n19223(n19223), 
         .n19222(n19222), .n19165(n19165), .n19164(n19164), .n19163(n19163), 
         .n19162(n19162), .n19161(n19161), .n19160(n19160), .n19159(n19159), 
         .n19158(n19158), .n32667(n32667), .n32679(n32679), .n32660(n32660), 
         .n17504(n17504), .n20830(n20830), .n5(n5_adj_4991), .n38579(n38579), 
         .n18738(n18738), .n18956(n18956), .tx_o(tx_o), .r_SM_Main({r_SM_Main_adj_5135}), 
         .VCC_net(VCC_net), .\r_SM_Main_2__N_3487[1] (r_SM_Main_2__N_3487[1]), 
         .n4(n4_adj_4888), .\r_Bit_Index[0] (r_Bit_Index_adj_5137[0]), .n19052(n19052), 
         .n19460(n19460), .n38214(n38214), .tx_enable(tx_enable), .n10524(n10524), 
         .n18732(n18732), .n18954(n18954), .r_Rx_Data(r_Rx_Data), .RX_N_10(RX_N_10), 
         .\r_Bit_Index[0]_adj_9 (r_Bit_Index[0]), .n23879(n23879), .n4_adj_10(n4), 
         .n4_adj_11(n4_adj_4931), .n17539(n17539), .n19524(n19524), .n19583(n19583), 
         .n19035(n19035), .n19034(n19034), .n19033(n19033), .n19032(n19032), 
         .n19031(n19031), .n19030(n19030), .n19029(n19029), .n17534(n17534), 
         .n4_adj_12(n4_adj_4928)) /* synthesis syn_module_defined=1 */ ;   // verilog/TinyFPGA_B.v(137[8] 160[4])
    SB_LUT4 unary_minus_4_inv_0_i7_1_lut (.I0(duty[6]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n19));   // verilog/TinyFPGA_B.v(106[23:28])
    defparam unary_minus_4_inv_0_i7_1_lut.LUT_INIT = 16'h5555;
    pwm PWM (.n36951(n36951), .VCC_net(VCC_net), .INHA_c(INHA_c), .clk32MHz(clk32MHz), 
        .n17362(n17362), .GND_net(GND_net), .pwm_counter({pwm_counter}), 
        .n17360(n17360)) /* synthesis syn_module_defined=1 */ ;   // verilog/TinyFPGA_B.v(89[6] 94[3])
    SB_LUT4 i13904_3_lut (.I0(control_mode[0]), .I1(\data_in_frame[1] [0]), 
            .I2(n33567), .I3(GND_net), .O(n19046));   // verilog/coms.v(127[12] 300[6])
    defparam i13904_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13905_3_lut (.I0(PWMLimit[0]), .I1(\data_in_frame[10] [0]), 
            .I2(n33567), .I3(GND_net), .O(n19047));   // verilog/coms.v(127[12] 300[6])
    defparam i13905_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i28553_4_lut (.I0(n17476), .I1(n39), .I2(n771), .I3(n3303), 
            .O(n35305));
    defparam i28553_4_lut.LUT_INIT = 16'hfac8;
    SB_LUT4 i1_4_lut_adj_1715 (.I0(n32688), .I1(\FRAME_MATCHER.state [0]), 
            .I2(n35305), .I3(n14711), .O(n48));   // verilog/coms.v(127[12] 300[6])
    defparam i1_4_lut_adj_1715.LUT_INIT = 16'h8caf;
    SB_LUT4 i1_4_lut_adj_1716 (.I0(n7_adj_5045), .I1(n48), .I2(\FRAME_MATCHER.state [3]), 
            .I3(n17474), .O(n32009));   // verilog/coms.v(127[12] 300[6])
    defparam i1_4_lut_adj_1716.LUT_INIT = 16'hccdc;
    SB_LUT4 i13907_3_lut (.I0(quadB_debounced), .I1(reg_B[0]), .I2(n35256), 
            .I3(GND_net), .O(n19049));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(186[9] 190[16])
    defparam i13907_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_1717 (.I0(enable_slow_N_4001), .I1(data_ready), 
            .I2(state_adj_5128[1]), .I3(state_adj_5128[0]), .O(n32425));   // verilog/eeprom.v(26[8] 58[4])
    defparam i1_4_lut_adj_1717.LUT_INIT = 16'hccd0;
    SB_LUT4 i13909_4_lut (.I0(rw), .I1(state_adj_5128[0]), .I2(state_adj_5128[1]), 
            .I3(n3647), .O(n19051));   // verilog/eeprom.v(26[8] 58[4])
    defparam i13909_4_lut.LUT_INIT = 16'hacaa;
    EEPROM eeprom (.CLK_c(CLK_c), .n3646({n3647}), .\state[1] (state_adj_5128[1]), 
           .enable_slow_N_4001(enable_slow_N_4001), .GND_net(GND_net), .read(read), 
           .\state[0] (state_adj_5128[0]), .\state[2] (state_adj_5158[2]), 
           .n7(n7_adj_4972), .n19051(n19051), .rw(rw), .n32425(n32425), 
           .data_ready(data_ready), .n24036(n24036), .n33471(n33471), 
           .n33535(n33535), .n32331(n32331), .n32323(n32323), .\state[3] (state_adj_5158[3]), 
           .n6(n6_adj_4932), .n5212(n5212), .\state_7__N_3914[3] (state_7__N_3914[3]), 
           .\saved_addr[0] (saved_addr[0]), .\state[0]_adj_3 (state_adj_5158[0]), 
           .\state_7__N_3898[0] (state_7__N_3898[0]), .n10(n10_adj_5076), 
           .scl_enable(scl_enable), .VCC_net(VCC_net), .sda_enable(sda_enable), 
           .n23736(n23736), .n10_adj_4(n10), .n5690(n5690), .n19061(n19061), 
           .data({data}), .n19060(n19060), .n19056(n19056), .n19055(n19055), 
           .n19054(n19054), .n19592(n19592), .n19584(n19584), .n19582(n19582), 
           .n19558(n19558), .n8(n8_adj_4900), .scl(scl), .sda_out(sda_out), 
           .n36289(n36289), .n4(n4_adj_4942), .n23836(n23836), .n17518(n17518), 
           .n4_adj_5(n4_adj_4941), .n17513(n17513)) /* synthesis syn_noprune=1, syn_module_defined=1 */ ;   // verilog/TinyFPGA_B.v(267[10] 278[6])
    SB_LUT4 i13910_4_lut (.I0(tx_active), .I1(r_SM_Main_adj_5135[1]), .I2(n10524), 
            .I3(n4_adj_4888), .O(n19052));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i13910_4_lut.LUT_INIT = 16'h32aa;
    SB_LUT4 i13911_3_lut (.I0(quadB_debounced_adj_4927), .I1(reg_B_adj_5146[0]), 
            .I2(n35209), .I3(GND_net), .O(n19053));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(186[9] 190[16])
    defparam i13911_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13912_4_lut (.I0(state_7__N_3914[3]), .I1(data[7]), .I2(n23836), 
            .I3(n17518), .O(n19054));   // verilog/i2c_controller.v(91[8] 173[6])
    defparam i13912_4_lut.LUT_INIT = 16'hccac;
    SB_LUT4 i26656_3_lut (.I0(encoder0_position[19]), .I1(n33399), .I2(encoder0_position[23]), 
            .I3(GND_net), .O(n678));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam i26656_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13913_4_lut (.I0(state_7__N_3914[3]), .I1(data[6]), .I2(n23836), 
            .I3(n17513), .O(n19055));   // verilog/i2c_controller.v(91[8] 173[6])
    defparam i13913_4_lut.LUT_INIT = 16'hccac;
    SB_LUT4 i13914_4_lut (.I0(saved_addr[0]), .I1(rw), .I2(state_7__N_3898[0]), 
            .I3(enable_slow_N_4001), .O(n19056));   // verilog/i2c_controller.v(91[8] 173[6])
    defparam i13914_4_lut.LUT_INIT = 16'haaca;
    SB_LUT4 i2_3_lut_adj_1718 (.I0(data_ready), .I1(\ID_READOUT_FSM.state [1]), 
            .I2(\ID_READOUT_FSM.state [0]), .I3(GND_net), .O(n35211));
    defparam i2_3_lut_adj_1718.LUT_INIT = 16'hdfdf;
    SB_LUT4 i13915_3_lut (.I0(ID[0]), .I1(data[0]), .I2(n35211), .I3(GND_net), 
            .O(n19057));   // verilog/TinyFPGA_B.v(237[10] 265[6])
    defparam i13915_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i3_4_lut_adj_1719 (.I0(\ID_READOUT_FSM.state [1]), .I1(n62), 
            .I2(delay_counter[31]), .I3(\ID_READOUT_FSM.state [0]), .O(n35190));
    defparam i3_4_lut_adj_1719.LUT_INIT = 16'h0004;
    SB_LUT4 i13918_4_lut (.I0(state_7__N_3914[3]), .I1(data[5]), .I2(n4_adj_4941), 
            .I3(n17518), .O(n19060));   // verilog/i2c_controller.v(91[8] 173[6])
    defparam i13918_4_lut.LUT_INIT = 16'hccca;
    \quad(DEBOUNCE_TICKS=100)  quad_counter1 (.encoder1_position({encoder1_position}), 
            .clk32MHz(clk32MHz), .data_o({quadA_debounced_adj_4926, quadB_debounced_adj_4927}), 
            .GND_net(GND_net), .ENCODER1_A_c_1(ENCODER1_A_c_1), .reg_B({reg_B_adj_5146}), 
            .VCC_net(VCC_net), .n35209(n35209), .n19053(n19053), .ENCODER1_B_c_0(ENCODER1_B_c_0), 
            .n19593(n19593)) /* synthesis syn_module_defined=1 */ ;   // verilog/TinyFPGA_B.v(193[15] 198[4])
    SB_LUT4 i13919_4_lut (.I0(state_7__N_3914[3]), .I1(data[0]), .I2(n10_adj_5076), 
            .I3(n17513), .O(n19061));   // verilog/i2c_controller.v(91[8] 173[6])
    defparam i13919_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i1_4_lut_adj_1720 (.I0(n63_adj_4971), .I1(n5_adj_4991), .I2(n2970), 
            .I3(n20830), .O(n6));   // verilog/coms.v(127[12] 300[6])
    defparam i1_4_lut_adj_1720.LUT_INIT = 16'heccc;
    SB_LUT4 i1_4_lut_adj_1721 (.I0(n17476), .I1(n63_adj_4971), .I2(n10417), 
            .I3(n32_adj_5070), .O(n5_adj_5071));   // verilog/coms.v(127[12] 300[6])
    defparam i1_4_lut_adj_1721.LUT_INIT = 16'hdc50;
    SB_LUT4 i3_4_lut_adj_1722 (.I0(n4452), .I1(n6), .I2(n17552), .I3(n38579), 
            .O(n8_adj_4933));   // verilog/coms.v(127[12] 300[6])
    defparam i3_4_lut_adj_1722.LUT_INIT = 16'hcfce;
    SB_LUT4 i4_4_lut_adj_1723 (.I0(n20830), .I1(n8_adj_4933), .I2(n63), 
            .I3(n5_adj_5071), .O(n38206));   // verilog/coms.v(127[12] 300[6])
    defparam i4_4_lut_adj_1723.LUT_INIT = 16'hefcf;
    
endmodule
//
// Verilog Description of module \quad(DEBOUNCE_TICKS=100)_U1 
//

module \quad(DEBOUNCE_TICKS=100)_U1  (encoder0_position, GND_net, data_o, 
            clk32MHz, reg_B, VCC_net, n35256, n19049, ENCODER0_B_c_0, 
            n19588, ENCODER0_A_c_1) /* synthesis syn_module_defined=1 */ ;
    output [23:0]encoder0_position;
    input GND_net;
    output [1:0]data_o;
    input clk32MHz;
    output [1:0]reg_B;
    input VCC_net;
    output n35256;
    input n19049;
    input ENCODER0_B_c_0;
    input n19588;
    input ENCODER0_A_c_1;
    
    wire clk32MHz /* synthesis SET_AS_NETWORK=clk32MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(33[6:14])
    wire [23:0]n3203;
    
    wire n3199, n27933, n27934, B_delayed, count_direction, n27932, 
        count_enable, A_delayed, n27931, n27930, n27929, n27928, 
        n27927, n27926, n27925, n27924, n27923, n27922, n27921, 
        n27944, n27943, n27942, n27941, n27940, n27939, n27938, 
        n27937, n27936, n27935;
    
    SB_LUT4 add_741_14_lut (.I0(GND_net), .I1(encoder0_position[12]), .I2(n3199), 
            .I3(n27933), .O(n3203[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_741_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_741_14 (.CI(n27933), .I0(encoder0_position[12]), .I1(n3199), 
            .CO(n27934));
    SB_LUT4 quadA_debounced_I_0_2_lut (.I0(data_o[1]), .I1(B_delayed), .I2(GND_net), 
            .I3(GND_net), .O(count_direction));   // quad.v(26[26:53])
    defparam quadA_debounced_I_0_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_741_13_lut (.I0(GND_net), .I1(encoder0_position[11]), .I2(n3199), 
            .I3(n27932), .O(n3203[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_741_13_lut.LUT_INIT = 16'hC33C;
    SB_DFFE count_i0_i0 (.Q(encoder0_position[0]), .C(clk32MHz), .E(count_enable), 
            .D(n3203[0]));   // quad.v(35[10] 41[6])
    SB_DFF B_delayed_16 (.Q(B_delayed), .C(clk32MHz), .D(data_o[0]));   // quad.v(23[10:54])
    SB_DFF A_delayed_15 (.Q(A_delayed), .C(clk32MHz), .D(data_o[1]));   // quad.v(22[10:54])
    SB_CARRY add_741_13 (.CI(n27932), .I0(encoder0_position[11]), .I1(n3199), 
            .CO(n27933));
    SB_LUT4 add_741_12_lut (.I0(GND_net), .I1(encoder0_position[10]), .I2(n3199), 
            .I3(n27931), .O(n3203[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_741_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_741_12 (.CI(n27931), .I0(encoder0_position[10]), .I1(n3199), 
            .CO(n27932));
    SB_LUT4 add_741_11_lut (.I0(GND_net), .I1(encoder0_position[9]), .I2(n3199), 
            .I3(n27930), .O(n3203[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_741_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_741_11 (.CI(n27930), .I0(encoder0_position[9]), .I1(n3199), 
            .CO(n27931));
    SB_LUT4 add_741_10_lut (.I0(GND_net), .I1(encoder0_position[8]), .I2(n3199), 
            .I3(n27929), .O(n3203[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_741_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_741_10 (.CI(n27929), .I0(encoder0_position[8]), .I1(n3199), 
            .CO(n27930));
    SB_LUT4 add_741_9_lut (.I0(GND_net), .I1(encoder0_position[7]), .I2(n3199), 
            .I3(n27928), .O(n3203[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_741_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_741_9 (.CI(n27928), .I0(encoder0_position[7]), .I1(n3199), 
            .CO(n27929));
    SB_LUT4 add_741_8_lut (.I0(GND_net), .I1(encoder0_position[6]), .I2(n3199), 
            .I3(n27927), .O(n3203[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_741_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_741_8 (.CI(n27927), .I0(encoder0_position[6]), .I1(n3199), 
            .CO(n27928));
    SB_LUT4 add_741_7_lut (.I0(GND_net), .I1(encoder0_position[5]), .I2(n3199), 
            .I3(n27926), .O(n3203[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_741_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_741_7 (.CI(n27926), .I0(encoder0_position[5]), .I1(n3199), 
            .CO(n27927));
    SB_LUT4 add_741_6_lut (.I0(GND_net), .I1(encoder0_position[4]), .I2(n3199), 
            .I3(n27925), .O(n3203[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_741_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_741_6 (.CI(n27925), .I0(encoder0_position[4]), .I1(n3199), 
            .CO(n27926));
    SB_LUT4 add_741_5_lut (.I0(GND_net), .I1(encoder0_position[3]), .I2(n3199), 
            .I3(n27924), .O(n3203[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_741_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_741_5 (.CI(n27924), .I0(encoder0_position[3]), .I1(n3199), 
            .CO(n27925));
    SB_LUT4 add_741_4_lut (.I0(GND_net), .I1(encoder0_position[2]), .I2(n3199), 
            .I3(n27923), .O(n3203[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_741_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_741_4 (.CI(n27923), .I0(encoder0_position[2]), .I1(n3199), 
            .CO(n27924));
    SB_LUT4 add_741_3_lut (.I0(GND_net), .I1(encoder0_position[1]), .I2(n3199), 
            .I3(n27922), .O(n3203[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_741_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_741_3 (.CI(n27922), .I0(encoder0_position[1]), .I1(n3199), 
            .CO(n27923));
    SB_LUT4 add_741_2_lut (.I0(GND_net), .I1(encoder0_position[0]), .I2(count_direction), 
            .I3(n27921), .O(n3203[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_741_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_741_2 (.CI(n27921), .I0(encoder0_position[0]), .I1(count_direction), 
            .CO(n27922));
    SB_CARRY add_741_1 (.CI(GND_net), .I0(n3199), .I1(n3199), .CO(n27921));
    SB_DFFE count_i0_i23 (.Q(encoder0_position[23]), .C(clk32MHz), .E(count_enable), 
            .D(n3203[23]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i22 (.Q(encoder0_position[22]), .C(clk32MHz), .E(count_enable), 
            .D(n3203[22]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i21 (.Q(encoder0_position[21]), .C(clk32MHz), .E(count_enable), 
            .D(n3203[21]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i20 (.Q(encoder0_position[20]), .C(clk32MHz), .E(count_enable), 
            .D(n3203[20]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i19 (.Q(encoder0_position[19]), .C(clk32MHz), .E(count_enable), 
            .D(n3203[19]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i18 (.Q(encoder0_position[18]), .C(clk32MHz), .E(count_enable), 
            .D(n3203[18]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i17 (.Q(encoder0_position[17]), .C(clk32MHz), .E(count_enable), 
            .D(n3203[17]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i16 (.Q(encoder0_position[16]), .C(clk32MHz), .E(count_enable), 
            .D(n3203[16]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i15 (.Q(encoder0_position[15]), .C(clk32MHz), .E(count_enable), 
            .D(n3203[15]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i14 (.Q(encoder0_position[14]), .C(clk32MHz), .E(count_enable), 
            .D(n3203[14]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i13 (.Q(encoder0_position[13]), .C(clk32MHz), .E(count_enable), 
            .D(n3203[13]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i12 (.Q(encoder0_position[12]), .C(clk32MHz), .E(count_enable), 
            .D(n3203[12]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i11 (.Q(encoder0_position[11]), .C(clk32MHz), .E(count_enable), 
            .D(n3203[11]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i10 (.Q(encoder0_position[10]), .C(clk32MHz), .E(count_enable), 
            .D(n3203[10]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i9 (.Q(encoder0_position[9]), .C(clk32MHz), .E(count_enable), 
            .D(n3203[9]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i8 (.Q(encoder0_position[8]), .C(clk32MHz), .E(count_enable), 
            .D(n3203[8]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i7 (.Q(encoder0_position[7]), .C(clk32MHz), .E(count_enable), 
            .D(n3203[7]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i6 (.Q(encoder0_position[6]), .C(clk32MHz), .E(count_enable), 
            .D(n3203[6]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i5 (.Q(encoder0_position[5]), .C(clk32MHz), .E(count_enable), 
            .D(n3203[5]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i4 (.Q(encoder0_position[4]), .C(clk32MHz), .E(count_enable), 
            .D(n3203[4]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i3 (.Q(encoder0_position[3]), .C(clk32MHz), .E(count_enable), 
            .D(n3203[3]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i2 (.Q(encoder0_position[2]), .C(clk32MHz), .E(count_enable), 
            .D(n3203[2]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i1 (.Q(encoder0_position[1]), .C(clk32MHz), .E(count_enable), 
            .D(n3203[1]));   // quad.v(35[10] 41[6])
    SB_LUT4 i1182_1_lut_2_lut (.I0(data_o[1]), .I1(B_delayed), .I2(GND_net), 
            .I3(GND_net), .O(n3199));   // quad.v(37[5] 40[8])
    defparam i1182_1_lut_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i3_4_lut (.I0(data_o[1]), .I1(A_delayed), .I2(B_delayed), 
            .I3(data_o[0]), .O(count_enable));   // quad.v(25[23:80])
    defparam i3_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 add_741_25_lut (.I0(GND_net), .I1(encoder0_position[23]), .I2(n3199), 
            .I3(n27944), .O(n3203[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_741_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_741_24_lut (.I0(GND_net), .I1(encoder0_position[22]), .I2(n3199), 
            .I3(n27943), .O(n3203[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_741_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_741_24 (.CI(n27943), .I0(encoder0_position[22]), .I1(n3199), 
            .CO(n27944));
    SB_LUT4 add_741_23_lut (.I0(GND_net), .I1(encoder0_position[21]), .I2(n3199), 
            .I3(n27942), .O(n3203[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_741_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_741_23 (.CI(n27942), .I0(encoder0_position[21]), .I1(n3199), 
            .CO(n27943));
    SB_LUT4 add_741_22_lut (.I0(GND_net), .I1(encoder0_position[20]), .I2(n3199), 
            .I3(n27941), .O(n3203[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_741_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_741_22 (.CI(n27941), .I0(encoder0_position[20]), .I1(n3199), 
            .CO(n27942));
    SB_LUT4 add_741_21_lut (.I0(GND_net), .I1(encoder0_position[19]), .I2(n3199), 
            .I3(n27940), .O(n3203[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_741_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_741_21 (.CI(n27940), .I0(encoder0_position[19]), .I1(n3199), 
            .CO(n27941));
    SB_LUT4 add_741_20_lut (.I0(GND_net), .I1(encoder0_position[18]), .I2(n3199), 
            .I3(n27939), .O(n3203[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_741_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_741_20 (.CI(n27939), .I0(encoder0_position[18]), .I1(n3199), 
            .CO(n27940));
    SB_LUT4 add_741_19_lut (.I0(GND_net), .I1(encoder0_position[17]), .I2(n3199), 
            .I3(n27938), .O(n3203[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_741_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_741_19 (.CI(n27938), .I0(encoder0_position[17]), .I1(n3199), 
            .CO(n27939));
    SB_LUT4 add_741_18_lut (.I0(GND_net), .I1(encoder0_position[16]), .I2(n3199), 
            .I3(n27937), .O(n3203[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_741_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_741_18 (.CI(n27937), .I0(encoder0_position[16]), .I1(n3199), 
            .CO(n27938));
    SB_LUT4 add_741_17_lut (.I0(GND_net), .I1(encoder0_position[15]), .I2(n3199), 
            .I3(n27936), .O(n3203[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_741_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_741_17 (.CI(n27936), .I0(encoder0_position[15]), .I1(n3199), 
            .CO(n27937));
    SB_LUT4 add_741_16_lut (.I0(GND_net), .I1(encoder0_position[14]), .I2(n3199), 
            .I3(n27935), .O(n3203[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_741_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_741_16 (.CI(n27935), .I0(encoder0_position[14]), .I1(n3199), 
            .CO(n27936));
    SB_LUT4 add_741_15_lut (.I0(GND_net), .I1(encoder0_position[13]), .I2(n3199), 
            .I3(n27934), .O(n3203[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_741_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_741_15 (.CI(n27934), .I0(encoder0_position[13]), .I1(n3199), 
            .CO(n27935));
    \grp_debouncer(2,100)_U0  debounce (.reg_B({reg_B}), .clk32MHz(clk32MHz), 
            .GND_net(GND_net), .VCC_net(VCC_net), .n35256(n35256), .n19049(n19049), 
            .data_o({data_o}), .ENCODER0_B_c_0(ENCODER0_B_c_0), .n19588(n19588), 
            .ENCODER0_A_c_1(ENCODER0_A_c_1));   // quad.v(15[37] 19[4])
    
endmodule
//
// Verilog Description of module \grp_debouncer(2,100)_U0 
//

module \grp_debouncer(2,100)_U0  (reg_B, clk32MHz, GND_net, VCC_net, 
            n35256, n19049, data_o, ENCODER0_B_c_0, n19588, ENCODER0_A_c_1);
    output [1:0]reg_B;
    input clk32MHz;
    input GND_net;
    input VCC_net;
    output n35256;
    input n19049;
    output [1:0]data_o;
    input ENCODER0_B_c_0;
    input n19588;
    input ENCODER0_A_c_1;
    
    wire clk32MHz /* synthesis SET_AS_NETWORK=clk32MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(33[6:14])
    wire [1:0]reg_A;   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(142[12:17])
    wire [6:0]n33;
    wire [6:0]cnt_reg;   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(149[12:19])
    
    wire n28618, n28617, n28616, n28615, n28614, n28613, n12, 
        n2, cnt_next_6__N_3730;
    
    SB_DFF reg_B_i0 (.Q(reg_B[0]), .C(clk32MHz), .D(reg_A[0]));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(178[9] 184[16])
    SB_LUT4 cnt_reg_1585_add_4_8_lut (.I0(GND_net), .I1(GND_net), .I2(cnt_reg[6]), 
            .I3(n28618), .O(n33[6])) /* synthesis syn_instantiated=1 */ ;
    defparam cnt_reg_1585_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 cnt_reg_1585_add_4_7_lut (.I0(GND_net), .I1(GND_net), .I2(cnt_reg[5]), 
            .I3(n28617), .O(n33[5])) /* synthesis syn_instantiated=1 */ ;
    defparam cnt_reg_1585_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY cnt_reg_1585_add_4_7 (.CI(n28617), .I0(GND_net), .I1(cnt_reg[5]), 
            .CO(n28618));
    SB_LUT4 cnt_reg_1585_add_4_6_lut (.I0(GND_net), .I1(GND_net), .I2(cnt_reg[4]), 
            .I3(n28616), .O(n33[4])) /* synthesis syn_instantiated=1 */ ;
    defparam cnt_reg_1585_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY cnt_reg_1585_add_4_6 (.CI(n28616), .I0(GND_net), .I1(cnt_reg[4]), 
            .CO(n28617));
    SB_LUT4 cnt_reg_1585_add_4_5_lut (.I0(GND_net), .I1(GND_net), .I2(cnt_reg[3]), 
            .I3(n28615), .O(n33[3])) /* synthesis syn_instantiated=1 */ ;
    defparam cnt_reg_1585_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY cnt_reg_1585_add_4_5 (.CI(n28615), .I0(GND_net), .I1(cnt_reg[3]), 
            .CO(n28616));
    SB_LUT4 cnt_reg_1585_add_4_4_lut (.I0(GND_net), .I1(GND_net), .I2(cnt_reg[2]), 
            .I3(n28614), .O(n33[2])) /* synthesis syn_instantiated=1 */ ;
    defparam cnt_reg_1585_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY cnt_reg_1585_add_4_4 (.CI(n28614), .I0(GND_net), .I1(cnt_reg[2]), 
            .CO(n28615));
    SB_LUT4 cnt_reg_1585_add_4_3_lut (.I0(GND_net), .I1(GND_net), .I2(cnt_reg[1]), 
            .I3(n28613), .O(n33[1])) /* synthesis syn_instantiated=1 */ ;
    defparam cnt_reg_1585_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY cnt_reg_1585_add_4_3 (.CI(n28613), .I0(GND_net), .I1(cnt_reg[1]), 
            .CO(n28614));
    SB_LUT4 cnt_reg_1585_add_4_2_lut (.I0(GND_net), .I1(GND_net), .I2(cnt_reg[0]), 
            .I3(VCC_net), .O(n33[0])) /* synthesis syn_instantiated=1 */ ;
    defparam cnt_reg_1585_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY cnt_reg_1585_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(cnt_reg[0]), 
            .CO(n28613));
    SB_LUT4 i5_4_lut (.I0(cnt_reg[1]), .I1(cnt_reg[4]), .I2(cnt_reg[3]), 
            .I3(cnt_reg[6]), .O(n12));
    defparam i5_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i6_4_lut (.I0(cnt_reg[5]), .I1(n12), .I2(cnt_reg[0]), .I3(cnt_reg[2]), 
            .O(n35256));
    defparam i6_4_lut.LUT_INIT = 16'hfdff;
    SB_LUT4 reg_B_1__I_0_i2_2_lut (.I0(reg_B[1]), .I1(reg_A[1]), .I2(GND_net), 
            .I3(GND_net), .O(n2));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(193[46:60])
    defparam reg_B_1__I_0_i2_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i2_4_lut (.I0(reg_B[0]), .I1(n35256), .I2(reg_A[0]), .I3(n2), 
            .O(cnt_next_6__N_3730));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[40:72])
    defparam i2_4_lut.LUT_INIT = 16'hff7b;
    SB_DFFSR cnt_reg_1585__i0 (.Q(cnt_reg[0]), .C(clk32MHz), .D(n33[0]), 
            .R(cnt_next_6__N_3730));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[78:85])
    SB_DFF reg_out_i0_i0 (.Q(data_o[0]), .C(clk32MHz), .D(n19049));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(186[9] 190[16])
    SB_DFF reg_B_i1 (.Q(reg_B[1]), .C(clk32MHz), .D(reg_A[1]));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(178[9] 184[16])
    SB_DFF reg_A_i0 (.Q(reg_A[0]), .C(clk32MHz), .D(ENCODER0_B_c_0));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(178[9] 184[16])
    SB_DFF reg_out_i0_i1 (.Q(data_o[1]), .C(clk32MHz), .D(n19588));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(186[9] 190[16])
    SB_DFF reg_A_i1 (.Q(reg_A[1]), .C(clk32MHz), .D(ENCODER0_A_c_1));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(178[9] 184[16])
    SB_DFFSR cnt_reg_1585__i1 (.Q(cnt_reg[1]), .C(clk32MHz), .D(n33[1]), 
            .R(cnt_next_6__N_3730));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[78:85])
    SB_DFFSR cnt_reg_1585__i2 (.Q(cnt_reg[2]), .C(clk32MHz), .D(n33[2]), 
            .R(cnt_next_6__N_3730));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[78:85])
    SB_DFFSR cnt_reg_1585__i3 (.Q(cnt_reg[3]), .C(clk32MHz), .D(n33[3]), 
            .R(cnt_next_6__N_3730));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[78:85])
    SB_DFFSR cnt_reg_1585__i4 (.Q(cnt_reg[4]), .C(clk32MHz), .D(n33[4]), 
            .R(cnt_next_6__N_3730));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[78:85])
    SB_DFFSR cnt_reg_1585__i5 (.Q(cnt_reg[5]), .C(clk32MHz), .D(n33[5]), 
            .R(cnt_next_6__N_3730));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[78:85])
    SB_DFFSR cnt_reg_1585__i6 (.Q(cnt_reg[6]), .C(clk32MHz), .D(n33[6]), 
            .R(cnt_next_6__N_3730));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[78:85])
    
endmodule
//
// Verilog Description of module neopixel
//

module neopixel (\neo_pixel_transmitter.done , clk32MHz, \neo_pixel_transmitter.t0 , 
            GND_net, VCC_net, timer, start, n14, n24759, \state[0] , 
            \state[1] , \state_3__N_402[1] , LED_c, neopxl_color, n18685, 
            n33425, n19040, n19557, n19556, n19555, n19554, n19553, 
            n19552, n19551, n19550, n19549, n19548, n19547, n19546, 
            n19545, n19544, n19543, n19542, n19541, n19540, n19539, 
            n19538, n19537, n19536, n19535, n19534, n19533, n19529, 
            n19528, n19527, n19526, n19525, n19521, NEOPXL_c, n33926, 
            n31453, n19022, n34265) /* synthesis syn_module_defined=1 */ ;
    output \neo_pixel_transmitter.done ;
    input clk32MHz;
    output [31:0]\neo_pixel_transmitter.t0 ;
    input GND_net;
    input VCC_net;
    output [31:0]timer;
    output start;
    output n14;
    output n24759;
    output \state[0] ;
    output \state[1] ;
    output \state_3__N_402[1] ;
    input LED_c;
    input [23:0]neopxl_color;
    output n18685;
    output n33425;
    input n19040;
    input n19557;
    input n19556;
    input n19555;
    input n19554;
    input n19553;
    input n19552;
    input n19551;
    input n19550;
    input n19549;
    input n19548;
    input n19547;
    input n19546;
    input n19545;
    input n19544;
    input n19543;
    input n19542;
    input n19541;
    input n19540;
    input n19539;
    input n19538;
    input n19537;
    input n19536;
    input n19535;
    input n19534;
    input n19533;
    input n19529;
    input n19528;
    input n19527;
    input n19526;
    input n19525;
    input n19521;
    output NEOPXL_c;
    input n33926;
    input n31453;
    input n19022;
    output n34265;
    
    wire clk32MHz /* synthesis SET_AS_NETWORK=clk32MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(33[6:14])
    
    wire n28793, n1903, n1928, n28794, \neo_pixel_transmitter.done_N_610 , 
        n35264;
    wire [31:0]n1;
    
    wire n2103, n2097, n18;
    wire [31:0]bit_ctr;   // verilog/neopixel.v(18[12:19])
    
    wire n2109, n24625, n2093, n2108, n2100, n30, n2098, n2094, 
        n2099, n28, n2105, n2096, n2095, n2102, n29, n2101, 
        n2107, n2104, n2106, n27, n2126, n1304, n1305, n10, 
        n1303, n1309, n12, n1306, n1308, n1302, n16, n1307, 
        n1301, n1334, n2027, n37625;
    wire [31:0]n255;
    
    wire n18566, n18886, n2003, n1904, n28792, n2004, n1905, n28791, 
        n27769, n27770, n2005, n1906, n28790, n2006, n1907, n28789, 
        n27786, n27768, n27787, n2489, n2390, n2423, n28692, n2490, 
        n2391, n28691, n2491, n2392, n28690, n2492, n2393, n28689, 
        n2493, n2394, n28688, n2494, n2395, n28687, n2495, n2396, 
        n28686, n2496, n2397, n28685, n2497, n2398, n28684, n2007, 
        n1908, n28788, n2498, n2399, n28683, n2008, n1909, n37622, 
        n28787, n2621, n37626, n2591, n2608, n2601, n2605, n36, 
        n2606, n2609, n25, n2593, n2596, n2600, n2590, n34, 
        n2594, n2589, n40, n2602, n2588, n2604, n2607, n38, 
        n2598, n2603, n39, n2592, n2597, n2595, n2599, n37, 
        n2522, n37624, n2499, n2400, n28682, n29627, n30003, n2500, 
        n2401, n28681, n2501, n2402, n28680, n2502, n2403, n28679, 
        n2503, n2404, n28678, n2504, n2405, n28677, n2505, n2406, 
        n28676, n2506, n2407, n28675, n1829, n37644, n2507, n2408, 
        n28674, n2508, n2409, n37623, n28673, n2009, n2509, n1806, 
        n1803, n1798, n1805, n24, n1808, n1804, n1802, n1807, 
        n22, n28672, n1800, n1799, n1797, n1801, n23, n1796, 
        n1809, n21_adj_4738, n1994, n28786, n28671, n28670, n28669, 
        n28668, n1730, n37643, n28667, n1699, n1709, n17_adj_4739, 
        n28666, n1698, n1707, n1703, n1705, n21_adj_4740, n1704, 
        n1701, n1708, n20_adj_4741, n1702, n1697, n24_adj_4742, 
        n1700, n1706, n1631, n37642, n28665, n28664, n28663, n28662, 
        n28661, n1607, n1603, n1598, n1605, n20_adj_4743, n1600, 
        n1609, n13, n28660, n28659, n1604, n1606, n18_adj_4744, 
        n1599, n1602, n22_adj_4745, n1601, n1608, n1532, n37641, 
        n1995, n28785, n28658, n28657, n28656, n28655, n28654, 
        n1506, n1503, n1500, n1501, n18_adj_4746, n1504, n1502, 
        n1499, n20_adj_4747, n1505, n1509, n15_adj_4748, n1508, 
        n1507, n28653, n1433, n37640, n28652, n2687, n28651, n2688, 
        n28650, n27785, n2689, n28649, n2690, n28648, n2691, n28647, 
        n1409, n24609, n2692, n28646, n2693, n28645, n2694, n28644, 
        n2695, n28643, n1405, n1407, n1400, n16_adj_4749, n2696, 
        n28642, n1402, n1403, n1401, n1406, n17_adj_4750, n1408, 
        n1404, n2697, n28641, n1037, n37639, n2698, n28640;
    wire [31:0]n971;
    
    wire n2, n1009, n1007, n1006, n1005, n16024, n1008, n906, 
        n905, n907, n35312, n18794, n36260, n36262, n35358, n38_adj_4751, 
        n4, n2699, n28639, n2700, n28638, n2701, n28637, n1136, 
        n37637, n1109, n24607, n1105, n1103, n1108, n12_adj_4755, 
        n2702, n28636, n1107, n1106, n1104, n3116, n37636, n2703, 
        n28635, n27784, n2704, n28634, n2705, n28633, n2706, n28632, 
        n2707, n28631, n1996, n28784, n2708, n28630, n2709, n1997, 
        n28783, n27783, n3102, n3090, n3103, n3085, n42, n3089, 
        n3094, n3101, n3098, n46, n3099, n3091, n3106, n3100, 
        n44, n3097, n3088, n3104, n3092, n45, n3105, n3083, 
        n3093, n3096, n43, n3108, n3109, n40_adj_4756, n3107, 
        n3087, n3086, n48, n52, n3095, n3084, n39_adj_4757, n3017, 
        n37635, n2324, n37634, n27782, n1998, n28782, n27767, 
        n1999, n28781, n2000, n28780, n27781, n27766, n2001, n28779, 
        n27780, n27765, n2002, n28778, n28777, n28776, n28775, 
        n28774, n27764, n28773, n3007, n2988, n2986, n2993, n42_adj_4759, 
        n3003, n3009, n29_adj_4760, n28772, n28771, n3008, n3002, 
        n3004, n2996, n40_adj_4761, n2994, n2995, n2999, n2985, 
        n45_adj_4762, n2989, n2990, n2984, n3006, n44_adj_4763, 
        n2997, n2998, n2987, n3005, n43_adj_4764, n2991, n2992, 
        n47, n3001, n3000, n49, n28105, n28104, n28103, n2192, 
        n28770, n2918, n37632, n2193, n28769, n2194, n28768, n28102, 
        n2195, n28767, n27779, n2196, n28766, n2197, n28765, n2198, 
        n28764, n28101, n28100, n28099, n28098, n2199, n28763, 
        n2200, n28762, n27778, n37627, n28097, n2786, n2720, n28566, 
        n2787, n28565, n2788, n28564, n2789, n28563, n2790, n28562, 
        n2791, n28561, n2792, n28560, n2793, n28559, n2201, n28761, 
        n2794, n28558, n2795, n28557, n2796, n28556, n27777, n2797, 
        n28555, n2202, n28760, n27776, n2203, n28759, n2798, n28554, 
        n2799, n28553, n2800, n28552, n2204, n28758, n2205, n28757, 
        n2206, n28756, n2801, n28551, n2802, n28550, n2803, n28549, 
        n2804, n28548, n2207, n28755, n2805, n28547, n2806, n28546, 
        n2208, n37628, n28754, n2209, n2807, n28545, n2808, n37629, 
        n28544, n2291, n2225, n28753, n2292, n28752, n2293, n28751, 
        n2809, n2294, n28750, n2885, n2819, n28543, n2886, n28542;
    wire [31:0]n133;
    
    wire n2887, n28541, n2888, n28540, n2295, n28749, n2889, n28539, 
        n2296, n28748, n2890, n28538, n2891, n28537, n2892, n28536, 
        n2893, n28535, n2894, n28534, n2895, n28533, n2297, n28747, 
        n2896, n28532, n2897, n28531, n2898, n28530, n2899, n28529, 
        n2900, n28528, n2901, n28527, n2902, n28526, n2903, n28525, 
        n2298, n28746, n1902, n1897, n26, n2299, n28745, n1899, 
        n1900, n24_adj_4766, n2904, n28524, n1901, n1896, n1895, 
        n25_adj_4767, n1898, n23_adj_4768, n2300, n28744, n2905, 
        n28523, n2906, n28522, n2907, n28521, n2908, n37631, n28520, 
        n2909, n28519, n28518, n2301, n28743, n28517, n28516, 
        n28515, n28514, n2302, n28742, n28513, n28512, n28511, 
        n2303, n28741, n2304, n28740, n28510, n28509, n28508, 
        n18_adj_4769, n28_adj_4770, n26_adj_4771, n27_adj_4772, n2305, 
        n28739, n28507, n2306, n28738, n2307, n28737, n25_adj_4773, 
        n2308, n37630, n28736, n24_adj_4774, n34_adj_4775, n22_adj_4776, 
        n38_adj_4777, n36_adj_4778, n37_adj_4779, n35, n2309, n28506, 
        n28735, n28505, n28734, n28504, n27775, n28503, n28733, 
        n28502, n28732, n28501, n28500, n28731, n27774, n28730, 
        n28499, n28729, n28498, n28497, n28728, n28496, n28495, 
        n24613, n28494, n28493, n28492, n28491, n28490, n28489, 
        n33365, n36222, n27_adj_4781, n33, n32, n31, n35_adj_4782, 
        n37_adj_4783;
    wire [31:0]one_wire_N_553;
    
    wire n17526, n28727, n28488, n28726, n28725, n28487, n28486, 
        n27773, n35064, n28485, n28484, n22_adj_4784, n27975, n28483, 
        n28482, n28481, n28480, n28479, n28478, n46_adj_4785, n44_adj_4786, 
        n45_adj_4787, n43_adj_4788, n42_adj_4789, n40_adj_4790, n48_adj_4791, 
        n52_adj_4792, n51, n29522, n24675, n33371, n14_adj_4793, 
        n28477, n28476, n28475, n28724, n23_adj_4794, n27974, n28474, 
        n28473, n28472, n28471, n10_adj_4795, n17393, n17509, n1251, 
        n24735, n5449, n36280, n28470, n33377, n28723, n28469, 
        n28468, n28467, n28466, n28465, n28722, n28464, n28463, 
        n28462, n28461, n28460, n28_adj_4796, n27973, n28459, n28721, 
        n28458, n28720, n28457, n28456, n28719, n28455, n28454, 
        n26_adj_4797, n27972, n28453, n28452, n28451, n28450, n28449, 
        n8799, n29995, n78, n28448, n28447, n28446, n27772, n28445, 
        n28444, n28443, n28442, n28441, n28440, n28718, n21_adj_4798, 
        n27971, n28717, n28439, n28438, n27970, n33451, n29671, 
        n24_adj_4799, n36_adj_4800, n25_adj_4801, n27_adj_4802, n37_adj_4803, 
        n63, n28437, n61, n28436, n59, n28435, n57, n28434, 
        n708, n55, n28433, n53, n28432, n51_adj_4804, n28431, 
        n49_adj_4805, n28430, n27771, n47_adj_4806, n28429, n45_adj_4807, 
        n28428, n43_adj_4808, n28427, n29_adj_4809, n30_adj_4810, 
        n37880, n37883, n10_adj_4811, n16_adj_4812, n33545, n41, 
        n28426, n32651, n116, n39_adj_4813, n28425, n37_adj_4814, 
        n28424, n35_adj_4815, n28423, n33_adj_4816, n28422, n31_adj_4817, 
        n28421, n29_adj_4818, n28420, n27_adj_4819, n28419, n25_adj_4820, 
        n28418, n23_adj_4821, n28417, n21_adj_4822, n28416, n27969, 
        n19_adj_4823, n28415, n17_adj_4824, n28414, n15_adj_4825, 
        n28413, n13_adj_4826, n28412, n37826, n35482, n11_adj_4827, 
        n28411, n3209, n27968, n1202, n28410, n1203, n28409, n1204, 
        n28408, n1205, n28407, n1206, n28406, n1207, n28405, n1208, 
        n28404, n27967, n1209, n37820, n35485, n37808, n35491, 
        n27966, n27965, n27964, n739, n33419, n60, n27963, n37742, 
        n37745, n37730, n36892, n27962, n27961, n27960, n27959, 
        n608, n33444, n27958, n27957, n33533, n24659, n33551, 
        n103, n32559, n18588, \neo_pixel_transmitter.done_N_616 , n1235, 
        n37638, n14_adj_4829, n9_adj_4830, n27956, n27955;
    wire [3:0]state_3__N_402;
    
    wire n27954, n838, n22_adj_4840, n30_adj_4841, n34_adj_4842, n32_adj_4843, 
        n33_adj_4844, n31_adj_4845, n27794, n27793, n33_adj_4846, 
        n27882, n41_adj_4847, n27881, n27953, n38_adj_4850, n27952, 
        n43_adj_4851, n40_adj_4852, n46_adj_4853, n27792, n39_adj_4854, 
        n27880, n27951, n47_adj_4855, n807, n27950, n27879, n27949, 
        n27948, n27947, n16028, n27878, n27946, n27945, n4_adj_4856, 
        n28196, n28195, n28194, n28193, n28192, n28191, n28190, 
        n28189, n27791, n40_adj_4857, n38_adj_4858, n28867, n27790, 
        n28866, n28865, n28864, n28863, n28862, n28861, n39_adj_4859, 
        n28860, n28859, n28858, n37_adj_4860, n28857, n28856, n28855, 
        n28854, n28853, n28852, n28851, n28850, n28849, n28848, 
        n28847, n28846, n28845, n28844, n28843, n28842, n28841, 
        n28840, n28839, n34_adj_4861, n42_adj_4862, n28838, n46_adj_4863, 
        n28837, n33_adj_4864, n28836, n28835, n28834, n28833, n28832, 
        n28831, n28830, n27789, n28829, n28828, n28827, n28826, 
        n28825, n28824, n28823, n28822, n28821, n28820, n28819, 
        n28818, n27788, n28817, n28816, n28815, n28814, n28813, 
        n28812, n28811, n28810, n28809, n28808, n28807, n28806, 
        n28805, n28804, n28803, n28802, n28_adj_4865, n32_adj_4866, 
        n30_adj_4867, n31_adj_4868, n29_adj_4869, n28801, n28800, 
        n28799, n28798, n28797, n28796, n28795, n28_adj_4870, n38_adj_4871, 
        n24637, n36_adj_4872, n42_adj_4873, n40_adj_4874, n41_adj_4875, 
        n39_adj_4876, n34121, n37664, n37667, n34867, n28_adj_4877, 
        n26_adj_4878, n27_adj_4879, n25_adj_4880, n14_adj_4881, n13_adj_4882, 
        n35175, n15_adj_4883, n1265;
    wire [4:0]color_bit_N_596;
    
    wire n36249;
    
    SB_CARRY mod_5_add_1339_9 (.CI(n28793), .I0(n1903), .I1(n1928), .CO(n28794));
    SB_DFFE \neo_pixel_transmitter.done_104  (.Q(\neo_pixel_transmitter.done ), 
            .C(clk32MHz), .E(n35264), .D(\neo_pixel_transmitter.done_N_610 ));   // verilog/neopixel.v(35[12] 117[6])
    SB_LUT4 sub_14_inv_0_i13_1_lut (.I0(\neo_pixel_transmitter.t0 [12]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[12]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i13_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1_2_lut (.I0(n2103), .I1(n2097), .I2(GND_net), .I3(GND_net), 
            .O(n18));
    defparam i1_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i19482_2_lut (.I0(bit_ctr[14]), .I1(n2109), .I2(GND_net), 
            .I3(GND_net), .O(n24625));
    defparam i19482_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i13_4_lut (.I0(n2093), .I1(n2108), .I2(n2100), .I3(n18), 
            .O(n30));
    defparam i13_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i11_4_lut (.I0(n2098), .I1(n24625), .I2(n2094), .I3(n2099), 
            .O(n28));
    defparam i11_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i12_4_lut (.I0(n2105), .I1(n2096), .I2(n2095), .I3(n2102), 
            .O(n29));
    defparam i12_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i10_4_lut (.I0(n2101), .I1(n2107), .I2(n2104), .I3(n2106), 
            .O(n27));
    defparam i10_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i16_4_lut (.I0(n27), .I1(n29), .I2(n28), .I3(n30), .O(n2126));
    defparam i16_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_adj_1501 (.I0(n1304), .I1(n1305), .I2(GND_net), .I3(GND_net), 
            .O(n10));
    defparam i1_2_lut_adj_1501.LUT_INIT = 16'heeee;
    SB_LUT4 i3_3_lut (.I0(bit_ctr[22]), .I1(n1303), .I2(n1309), .I3(GND_net), 
            .O(n12));
    defparam i3_3_lut.LUT_INIT = 16'hecec;
    SB_LUT4 i7_4_lut (.I0(n1306), .I1(n1308), .I2(n1302), .I3(n10), 
            .O(n16));
    defparam i7_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i8_4_lut (.I0(n1307), .I1(n16), .I2(n12), .I3(n1301), .O(n1334));
    defparam i8_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i30872_1_lut (.I0(n2027), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n37625));
    defparam i30872_1_lut.LUT_INIT = 16'h5555;
    SB_DFFESR bit_ctr_i0_i1 (.Q(bit_ctr[1]), .C(clk32MHz), .E(n18566), 
            .D(n255[1]), .R(n18886));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFESR bit_ctr_i0_i2 (.Q(bit_ctr[2]), .C(clk32MHz), .E(n18566), 
            .D(n255[2]), .R(n18886));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFESR bit_ctr_i0_i3 (.Q(bit_ctr[3]), .C(clk32MHz), .E(n18566), 
            .D(n255[3]), .R(n18886));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFESR bit_ctr_i0_i4 (.Q(bit_ctr[4]), .C(clk32MHz), .E(n18566), 
            .D(n255[4]), .R(n18886));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFESR bit_ctr_i0_i5 (.Q(bit_ctr[5]), .C(clk32MHz), .E(n18566), 
            .D(n255[5]), .R(n18886));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFESR bit_ctr_i0_i6 (.Q(bit_ctr[6]), .C(clk32MHz), .E(n18566), 
            .D(n255[6]), .R(n18886));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFESR bit_ctr_i0_i7 (.Q(bit_ctr[7]), .C(clk32MHz), .E(n18566), 
            .D(n255[7]), .R(n18886));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFESR bit_ctr_i0_i8 (.Q(bit_ctr[8]), .C(clk32MHz), .E(n18566), 
            .D(n255[8]), .R(n18886));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFESR bit_ctr_i0_i9 (.Q(bit_ctr[9]), .C(clk32MHz), .E(n18566), 
            .D(n255[9]), .R(n18886));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFESR bit_ctr_i0_i10 (.Q(bit_ctr[10]), .C(clk32MHz), .E(n18566), 
            .D(n255[10]), .R(n18886));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFESR bit_ctr_i0_i11 (.Q(bit_ctr[11]), .C(clk32MHz), .E(n18566), 
            .D(n255[11]), .R(n18886));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFESR bit_ctr_i0_i12 (.Q(bit_ctr[12]), .C(clk32MHz), .E(n18566), 
            .D(n255[12]), .R(n18886));   // verilog/neopixel.v(35[12] 117[6])
    SB_LUT4 sub_14_inv_0_i14_1_lut (.I0(\neo_pixel_transmitter.t0 [13]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[13]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i14_1_lut.LUT_INIT = 16'h5555;
    SB_DFFESR bit_ctr_i0_i13 (.Q(bit_ctr[13]), .C(clk32MHz), .E(n18566), 
            .D(n255[13]), .R(n18886));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFESR bit_ctr_i0_i14 (.Q(bit_ctr[14]), .C(clk32MHz), .E(n18566), 
            .D(n255[14]), .R(n18886));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFESR bit_ctr_i0_i15 (.Q(bit_ctr[15]), .C(clk32MHz), .E(n18566), 
            .D(n255[15]), .R(n18886));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFESR bit_ctr_i0_i16 (.Q(bit_ctr[16]), .C(clk32MHz), .E(n18566), 
            .D(n255[16]), .R(n18886));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFESR bit_ctr_i0_i17 (.Q(bit_ctr[17]), .C(clk32MHz), .E(n18566), 
            .D(n255[17]), .R(n18886));   // verilog/neopixel.v(35[12] 117[6])
    SB_LUT4 sub_14_inv_0_i15_1_lut (.I0(\neo_pixel_transmitter.t0 [14]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[14]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i15_1_lut.LUT_INIT = 16'h5555;
    SB_DFFESR bit_ctr_i0_i18 (.Q(bit_ctr[18]), .C(clk32MHz), .E(n18566), 
            .D(n255[18]), .R(n18886));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFESR bit_ctr_i0_i19 (.Q(bit_ctr[19]), .C(clk32MHz), .E(n18566), 
            .D(n255[19]), .R(n18886));   // verilog/neopixel.v(35[12] 117[6])
    SB_LUT4 mod_5_add_1339_8_lut (.I0(n1904), .I1(n1904), .I2(n1928), 
            .I3(n28792), .O(n2003)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_8_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1339_8 (.CI(n28792), .I0(n1904), .I1(n1928), .CO(n28793));
    SB_LUT4 mod_5_add_1339_7_lut (.I0(n1905), .I1(n1905), .I2(n1928), 
            .I3(n28791), .O(n2004)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_7_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY add_21_8 (.CI(n27769), .I0(bit_ctr[6]), .I1(GND_net), .CO(n27770));
    SB_CARRY mod_5_add_1339_7 (.CI(n28791), .I0(n1905), .I1(n1928), .CO(n28792));
    SB_LUT4 mod_5_add_1339_6_lut (.I0(n1906), .I1(n1906), .I2(n1928), 
            .I3(n28790), .O(n2005)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_6_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1339_6 (.CI(n28790), .I0(n1906), .I1(n1928), .CO(n28791));
    SB_LUT4 mod_5_add_1339_5_lut (.I0(n1907), .I1(n1907), .I2(n1928), 
            .I3(n28789), .O(n2006)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_5_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 add_21_25_lut (.I0(GND_net), .I1(bit_ctr[23]), .I2(GND_net), 
            .I3(n27786), .O(n255[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_14_inv_0_i16_1_lut (.I0(\neo_pixel_transmitter.t0 [15]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[15]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i16_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_21_7_lut (.I0(GND_net), .I1(bit_ctr[5]), .I2(GND_net), 
            .I3(n27768), .O(n255[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_21_25 (.CI(n27786), .I0(bit_ctr[23]), .I1(GND_net), .CO(n27787));
    SB_LUT4 mod_5_add_1674_22_lut (.I0(n2390), .I1(n2390), .I2(n2423), 
            .I3(n28692), .O(n2489)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_22_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1674_21_lut (.I0(n2391), .I1(n2391), .I2(n2423), 
            .I3(n28691), .O(n2490)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_21_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 sub_14_inv_0_i17_1_lut (.I0(\neo_pixel_transmitter.t0 [16]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[16]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i17_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY mod_5_add_1674_21 (.CI(n28691), .I0(n2391), .I1(n2423), .CO(n28692));
    SB_LUT4 mod_5_add_1674_20_lut (.I0(n2392), .I1(n2392), .I2(n2423), 
            .I3(n28690), .O(n2491)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_20_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1674_20 (.CI(n28690), .I0(n2392), .I1(n2423), .CO(n28691));
    SB_LUT4 mod_5_add_1674_19_lut (.I0(n2393), .I1(n2393), .I2(n2423), 
            .I3(n28689), .O(n2492)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_19_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1674_19 (.CI(n28689), .I0(n2393), .I1(n2423), .CO(n28690));
    SB_LUT4 mod_5_add_1674_18_lut (.I0(n2394), .I1(n2394), .I2(n2423), 
            .I3(n28688), .O(n2493)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_18_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1674_18 (.CI(n28688), .I0(n2394), .I1(n2423), .CO(n28689));
    SB_LUT4 mod_5_add_1674_17_lut (.I0(n2395), .I1(n2395), .I2(n2423), 
            .I3(n28687), .O(n2494)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_17_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1674_17 (.CI(n28687), .I0(n2395), .I1(n2423), .CO(n28688));
    SB_LUT4 mod_5_add_1674_16_lut (.I0(n2396), .I1(n2396), .I2(n2423), 
            .I3(n28686), .O(n2495)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_16_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1674_16 (.CI(n28686), .I0(n2396), .I1(n2423), .CO(n28687));
    SB_LUT4 mod_5_add_1674_15_lut (.I0(n2397), .I1(n2397), .I2(n2423), 
            .I3(n28685), .O(n2496)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_15_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1674_15 (.CI(n28685), .I0(n2397), .I1(n2423), .CO(n28686));
    SB_CARRY mod_5_add_1339_5 (.CI(n28789), .I0(n1907), .I1(n1928), .CO(n28790));
    SB_LUT4 mod_5_add_1674_14_lut (.I0(n2398), .I1(n2398), .I2(n2423), 
            .I3(n28684), .O(n2497)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_14_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1339_4_lut (.I0(n1908), .I1(n1908), .I2(n1928), 
            .I3(n28788), .O(n2007)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_4_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1674_14 (.CI(n28684), .I0(n2398), .I1(n2423), .CO(n28685));
    SB_LUT4 mod_5_add_1674_13_lut (.I0(n2399), .I1(n2399), .I2(n2423), 
            .I3(n28683), .O(n2498)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_13_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1339_4 (.CI(n28788), .I0(n1908), .I1(n1928), .CO(n28789));
    SB_LUT4 mod_5_add_1339_3_lut (.I0(n1909), .I1(n1909), .I2(n37622), 
            .I3(n28787), .O(n2008)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_3_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1674_13 (.CI(n28683), .I0(n2399), .I1(n2423), .CO(n28684));
    SB_LUT4 sub_14_inv_0_i18_1_lut (.I0(\neo_pixel_transmitter.t0 [17]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[17]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i18_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i30873_1_lut (.I0(n2621), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n37626));
    defparam i30873_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i14_4_lut (.I0(n2591), .I1(n2608), .I2(n2601), .I3(n2605), 
            .O(n36));
    defparam i14_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i3_3_lut_adj_1502 (.I0(n2606), .I1(bit_ctr[9]), .I2(n2609), 
            .I3(GND_net), .O(n25));
    defparam i3_3_lut_adj_1502.LUT_INIT = 16'heaea;
    SB_LUT4 i12_4_lut_adj_1503 (.I0(n2593), .I1(n2596), .I2(n2600), .I3(n2590), 
            .O(n34));
    defparam i12_4_lut_adj_1503.LUT_INIT = 16'hfffe;
    SB_LUT4 i18_4_lut (.I0(n25), .I1(n36), .I2(n2594), .I3(n2589), .O(n40));
    defparam i18_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i16_4_lut_adj_1504 (.I0(n2602), .I1(n2588), .I2(n2604), .I3(n2607), 
            .O(n38));
    defparam i16_4_lut_adj_1504.LUT_INIT = 16'hfffe;
    SB_LUT4 i17_3_lut (.I0(n2598), .I1(n34), .I2(n2603), .I3(GND_net), 
            .O(n39));
    defparam i17_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i15_4_lut (.I0(n2592), .I1(n2597), .I2(n2595), .I3(n2599), 
            .O(n37));
    defparam i15_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i21_4_lut (.I0(n37), .I1(n39), .I2(n38), .I3(n40), .O(n2621));
    defparam i21_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i30871_1_lut (.I0(n2522), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n37624));
    defparam i30871_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY mod_5_add_1339_3 (.CI(n28787), .I0(n1909), .I1(n37622), .CO(n28788));
    SB_LUT4 mod_5_add_1674_12_lut (.I0(n2400), .I1(n2400), .I2(n2423), 
            .I3(n28682), .O(n2499)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_12_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1674_12 (.CI(n28682), .I0(n2400), .I1(n2423), .CO(n28683));
    SB_LUT4 i1_2_lut_adj_1505 (.I0(bit_ctr[3]), .I1(n29627), .I2(GND_net), 
            .I3(GND_net), .O(n30003));
    defparam i1_2_lut_adj_1505.LUT_INIT = 16'h6666;
    SB_DFFESR bit_ctr_i0_i20 (.Q(bit_ctr[20]), .C(clk32MHz), .E(n18566), 
            .D(n255[20]), .R(n18886));   // verilog/neopixel.v(35[12] 117[6])
    SB_LUT4 mod_5_add_1674_11_lut (.I0(n2401), .I1(n2401), .I2(n2423), 
            .I3(n28681), .O(n2500)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_11_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1674_11 (.CI(n28681), .I0(n2401), .I1(n2423), .CO(n28682));
    SB_LUT4 sub_14_inv_0_i19_1_lut (.I0(\neo_pixel_transmitter.t0 [18]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[18]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i19_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mod_5_add_1674_10_lut (.I0(n2402), .I1(n2402), .I2(n2423), 
            .I3(n28680), .O(n2501)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_10_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1674_10 (.CI(n28680), .I0(n2402), .I1(n2423), .CO(n28681));
    SB_LUT4 mod_5_add_1674_9_lut (.I0(n2403), .I1(n2403), .I2(n2423), 
            .I3(n28679), .O(n2502)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_9_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1674_9 (.CI(n28679), .I0(n2403), .I1(n2423), .CO(n28680));
    SB_LUT4 mod_5_add_1674_8_lut (.I0(n2404), .I1(n2404), .I2(n2423), 
            .I3(n28678), .O(n2503)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_8_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1674_8 (.CI(n28678), .I0(n2404), .I1(n2423), .CO(n28679));
    SB_LUT4 mod_5_add_1674_7_lut (.I0(n2405), .I1(n2405), .I2(n2423), 
            .I3(n28677), .O(n2504)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_7_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1674_7 (.CI(n28677), .I0(n2405), .I1(n2423), .CO(n28678));
    SB_LUT4 mod_5_add_1674_6_lut (.I0(n2406), .I1(n2406), .I2(n2423), 
            .I3(n28676), .O(n2505)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_6_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1674_6 (.CI(n28676), .I0(n2406), .I1(n2423), .CO(n28677));
    SB_LUT4 mod_5_add_1674_5_lut (.I0(n2407), .I1(n2407), .I2(n2423), 
            .I3(n28675), .O(n2506)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_5_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1674_5 (.CI(n28675), .I0(n2407), .I1(n2423), .CO(n28676));
    SB_LUT4 i30891_1_lut (.I0(n1829), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n37644));
    defparam i30891_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mod_5_add_1674_4_lut (.I0(n2408), .I1(n2408), .I2(n2423), 
            .I3(n28674), .O(n2507)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_4_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1674_4 (.CI(n28674), .I0(n2408), .I1(n2423), .CO(n28675));
    SB_LUT4 mod_5_add_1674_3_lut (.I0(n2409), .I1(n2409), .I2(n37623), 
            .I3(n28673), .O(n2508)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_3_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1674_3 (.CI(n28673), .I0(n2409), .I1(n37623), .CO(n28674));
    SB_LUT4 mod_5_add_1339_2_lut (.I0(bit_ctr[16]), .I1(bit_ctr[16]), .I2(n37622), 
            .I3(VCC_net), .O(n2009)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_2_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 mod_5_add_1674_2_lut (.I0(bit_ctr[11]), .I1(bit_ctr[11]), .I2(n37623), 
            .I3(VCC_net), .O(n2509)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_2_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1674_2 (.CI(VCC_net), .I0(bit_ctr[11]), .I1(n37623), 
            .CO(n28673));
    SB_LUT4 i10_4_lut_adj_1506 (.I0(n1806), .I1(n1803), .I2(n1798), .I3(n1805), 
            .O(n24));
    defparam i10_4_lut_adj_1506.LUT_INIT = 16'hfffe;
    SB_LUT4 i8_4_lut_adj_1507 (.I0(n1808), .I1(n1804), .I2(n1802), .I3(n1807), 
            .O(n22));
    defparam i8_4_lut_adj_1507.LUT_INIT = 16'hfffe;
    SB_LUT4 mod_5_add_1741_23_lut (.I0(n2489), .I1(n2489), .I2(n2522), 
            .I3(n28672), .O(n2588)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_23_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i9_4_lut (.I0(n1800), .I1(n1799), .I2(n1797), .I3(n1801), 
            .O(n23));
    defparam i9_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i7_3_lut (.I0(n1796), .I1(bit_ctr[17]), .I2(n1809), .I3(GND_net), 
            .O(n21_adj_4738));
    defparam i7_3_lut.LUT_INIT = 16'heaea;
    SB_CARRY mod_5_add_1339_2 (.CI(VCC_net), .I0(bit_ctr[16]), .I1(n37622), 
            .CO(n28787));
    SB_LUT4 i13_4_lut_adj_1508 (.I0(n21_adj_4738), .I1(n23), .I2(n22), 
            .I3(n24), .O(n1829));
    defparam i13_4_lut_adj_1508.LUT_INIT = 16'hfffe;
    SB_LUT4 mod_5_add_1406_18_lut (.I0(n1994), .I1(n1994), .I2(n2027), 
            .I3(n28786), .O(n2093)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_18_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1741_22_lut (.I0(n2490), .I1(n2490), .I2(n2522), 
            .I3(n28671), .O(n2589)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_22_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1741_22 (.CI(n28671), .I0(n2490), .I1(n2522), .CO(n28672));
    SB_LUT4 mod_5_add_1741_21_lut (.I0(n2491), .I1(n2491), .I2(n2522), 
            .I3(n28670), .O(n2590)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_21_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1741_21 (.CI(n28670), .I0(n2491), .I1(n2522), .CO(n28671));
    SB_LUT4 mod_5_add_1741_20_lut (.I0(n2492), .I1(n2492), .I2(n2522), 
            .I3(n28669), .O(n2591)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_20_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1741_20 (.CI(n28669), .I0(n2492), .I1(n2522), .CO(n28670));
    SB_LUT4 mod_5_add_1741_19_lut (.I0(n2493), .I1(n2493), .I2(n2522), 
            .I3(n28668), .O(n2592)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_19_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i30890_1_lut (.I0(n1730), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n37643));
    defparam i30890_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY mod_5_add_1741_19 (.CI(n28668), .I0(n2493), .I1(n2522), .CO(n28669));
    SB_LUT4 mod_5_add_1741_18_lut (.I0(n2494), .I1(n2494), .I2(n2522), 
            .I3(n28667), .O(n2593)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_18_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i4_3_lut (.I0(bit_ctr[18]), .I1(n1699), .I2(n1709), .I3(GND_net), 
            .O(n17_adj_4739));
    defparam i4_3_lut.LUT_INIT = 16'hecec;
    SB_CARRY mod_5_add_1741_18 (.CI(n28667), .I0(n2494), .I1(n2522), .CO(n28668));
    SB_LUT4 mod_5_add_1741_17_lut (.I0(n2495), .I1(n2495), .I2(n2522), 
            .I3(n28666), .O(n2594)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_17_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i8_4_lut_adj_1509 (.I0(n1698), .I1(n1707), .I2(n1703), .I3(n1705), 
            .O(n21_adj_4740));
    defparam i8_4_lut_adj_1509.LUT_INIT = 16'hfffe;
    SB_LUT4 i7_3_lut_adj_1510 (.I0(n1704), .I1(n1701), .I2(n1708), .I3(GND_net), 
            .O(n20_adj_4741));
    defparam i7_3_lut_adj_1510.LUT_INIT = 16'hfefe;
    SB_LUT4 i11_4_lut_adj_1511 (.I0(n21_adj_4740), .I1(n17_adj_4739), .I2(n1702), 
            .I3(n1697), .O(n24_adj_4742));
    defparam i11_4_lut_adj_1511.LUT_INIT = 16'hfffe;
    SB_LUT4 i12_4_lut_adj_1512 (.I0(n1700), .I1(n24_adj_4742), .I2(n20_adj_4741), 
            .I3(n1706), .O(n1730));
    defparam i12_4_lut_adj_1512.LUT_INIT = 16'hfffe;
    SB_DFFESR bit_ctr_i0_i21 (.Q(bit_ctr[21]), .C(clk32MHz), .E(n18566), 
            .D(n255[21]), .R(n18886));   // verilog/neopixel.v(35[12] 117[6])
    SB_LUT4 i30889_1_lut (.I0(n1631), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n37642));
    defparam i30889_1_lut.LUT_INIT = 16'h5555;
    SB_DFFESR bit_ctr_i0_i22 (.Q(bit_ctr[22]), .C(clk32MHz), .E(n18566), 
            .D(n255[22]), .R(n18886));   // verilog/neopixel.v(35[12] 117[6])
    SB_CARRY mod_5_add_1741_17 (.CI(n28666), .I0(n2495), .I1(n2522), .CO(n28667));
    SB_LUT4 mod_5_add_1741_16_lut (.I0(n2496), .I1(n2496), .I2(n2522), 
            .I3(n28665), .O(n2595)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_16_lut.LUT_INIT = 16'hCA3A;
    SB_DFFESR bit_ctr_i0_i23 (.Q(bit_ctr[23]), .C(clk32MHz), .E(n18566), 
            .D(n255[23]), .R(n18886));   // verilog/neopixel.v(35[12] 117[6])
    SB_CARRY mod_5_add_1741_16 (.CI(n28665), .I0(n2496), .I1(n2522), .CO(n28666));
    SB_LUT4 mod_5_add_1741_15_lut (.I0(n2497), .I1(n2497), .I2(n2522), 
            .I3(n28664), .O(n2596)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_15_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1741_15 (.CI(n28664), .I0(n2497), .I1(n2522), .CO(n28665));
    SB_LUT4 mod_5_add_1741_14_lut (.I0(n2498), .I1(n2498), .I2(n2522), 
            .I3(n28663), .O(n2597)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_14_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1741_14 (.CI(n28663), .I0(n2498), .I1(n2522), .CO(n28664));
    SB_DFFESR bit_ctr_i0_i24 (.Q(bit_ctr[24]), .C(clk32MHz), .E(n18566), 
            .D(n255[24]), .R(n18886));   // verilog/neopixel.v(35[12] 117[6])
    SB_LUT4 mod_5_add_1741_13_lut (.I0(n2499), .I1(n2499), .I2(n2522), 
            .I3(n28662), .O(n2598)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_13_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1741_13 (.CI(n28662), .I0(n2499), .I1(n2522), .CO(n28663));
    SB_DFFESR bit_ctr_i0_i25 (.Q(bit_ctr[25]), .C(clk32MHz), .E(n18566), 
            .D(n255[25]), .R(n18886));   // verilog/neopixel.v(35[12] 117[6])
    SB_LUT4 mod_5_add_1741_12_lut (.I0(n2500), .I1(n2500), .I2(n2522), 
            .I3(n28661), .O(n2599)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_12_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i8_4_lut_adj_1513 (.I0(n1607), .I1(n1603), .I2(n1598), .I3(n1605), 
            .O(n20_adj_4743));
    defparam i8_4_lut_adj_1513.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_3_lut (.I0(bit_ctr[19]), .I1(n1600), .I2(n1609), .I3(GND_net), 
            .O(n13));
    defparam i1_3_lut.LUT_INIT = 16'hecec;
    SB_CARRY mod_5_add_1741_12 (.CI(n28661), .I0(n2500), .I1(n2522), .CO(n28662));
    SB_LUT4 mod_5_add_1741_11_lut (.I0(n2501), .I1(n2501), .I2(n2522), 
            .I3(n28660), .O(n2600)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_11_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1741_11 (.CI(n28660), .I0(n2501), .I1(n2522), .CO(n28661));
    SB_LUT4 mod_5_add_1741_10_lut (.I0(n2502), .I1(n2502), .I2(n2522), 
            .I3(n28659), .O(n2601)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_10_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 sub_14_inv_0_i20_1_lut (.I0(\neo_pixel_transmitter.t0 [19]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[19]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i20_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i6_2_lut (.I0(n1604), .I1(n1606), .I2(GND_net), .I3(GND_net), 
            .O(n18_adj_4744));
    defparam i6_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i10_4_lut_adj_1514 (.I0(n13), .I1(n20_adj_4743), .I2(n1599), 
            .I3(n1602), .O(n22_adj_4745));
    defparam i10_4_lut_adj_1514.LUT_INIT = 16'hfffe;
    SB_CARRY mod_5_add_1741_10 (.CI(n28659), .I0(n2502), .I1(n2522), .CO(n28660));
    SB_LUT4 i11_4_lut_adj_1515 (.I0(n1601), .I1(n22_adj_4745), .I2(n18_adj_4744), 
            .I3(n1608), .O(n1631));
    defparam i11_4_lut_adj_1515.LUT_INIT = 16'hfffe;
    SB_LUT4 i30888_1_lut (.I0(n1532), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n37641));
    defparam i30888_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mod_5_add_1406_17_lut (.I0(n1995), .I1(n1995), .I2(n2027), 
            .I3(n28785), .O(n2094)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_17_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1741_9_lut (.I0(n2503), .I1(n2503), .I2(n2522), 
            .I3(n28658), .O(n2602)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_9_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1741_9 (.CI(n28658), .I0(n2503), .I1(n2522), .CO(n28659));
    SB_LUT4 mod_5_add_1741_8_lut (.I0(n2504), .I1(n2504), .I2(n2522), 
            .I3(n28657), .O(n2603)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_8_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1741_8 (.CI(n28657), .I0(n2504), .I1(n2522), .CO(n28658));
    SB_LUT4 mod_5_add_1741_7_lut (.I0(n2505), .I1(n2505), .I2(n2522), 
            .I3(n28656), .O(n2604)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_7_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1741_7 (.CI(n28656), .I0(n2505), .I1(n2522), .CO(n28657));
    SB_LUT4 mod_5_add_1741_6_lut (.I0(n2506), .I1(n2506), .I2(n2522), 
            .I3(n28655), .O(n2605)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_6_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1741_6 (.CI(n28655), .I0(n2506), .I1(n2522), .CO(n28656));
    SB_LUT4 mod_5_add_1741_5_lut (.I0(n2507), .I1(n2507), .I2(n2522), 
            .I3(n28654), .O(n2606)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_5_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i7_4_lut_adj_1516 (.I0(n1506), .I1(n1503), .I2(n1500), .I3(n1501), 
            .O(n18_adj_4746));
    defparam i7_4_lut_adj_1516.LUT_INIT = 16'hfffe;
    SB_LUT4 i9_4_lut_adj_1517 (.I0(n1504), .I1(n18_adj_4746), .I2(n1502), 
            .I3(n1499), .O(n20_adj_4747));
    defparam i9_4_lut_adj_1517.LUT_INIT = 16'hfffe;
    SB_LUT4 i4_3_lut_adj_1518 (.I0(bit_ctr[20]), .I1(n1505), .I2(n1509), 
            .I3(GND_net), .O(n15_adj_4748));
    defparam i4_3_lut_adj_1518.LUT_INIT = 16'hecec;
    SB_LUT4 i10_4_lut_adj_1519 (.I0(n15_adj_4748), .I1(n20_adj_4747), .I2(n1508), 
            .I3(n1507), .O(n1532));
    defparam i10_4_lut_adj_1519.LUT_INIT = 16'hfffe;
    SB_CARRY mod_5_add_1406_17 (.CI(n28785), .I0(n1995), .I1(n2027), .CO(n28786));
    SB_CARRY mod_5_add_1741_5 (.CI(n28654), .I0(n2507), .I1(n2522), .CO(n28655));
    SB_LUT4 mod_5_add_1741_4_lut (.I0(n2508), .I1(n2508), .I2(n2522), 
            .I3(n28653), .O(n2607)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_4_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1741_4 (.CI(n28653), .I0(n2508), .I1(n2522), .CO(n28654));
    SB_LUT4 i30887_1_lut (.I0(n1433), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n37640));
    defparam i30887_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mod_5_add_1741_3_lut (.I0(n2509), .I1(n2509), .I2(n37624), 
            .I3(n28652), .O(n2608)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_3_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1741_3 (.CI(n28652), .I0(n2509), .I1(n37624), .CO(n28653));
    SB_LUT4 mod_5_add_1741_2_lut (.I0(bit_ctr[10]), .I1(bit_ctr[10]), .I2(n37624), 
            .I3(VCC_net), .O(n2609)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_2_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1741_2 (.CI(VCC_net), .I0(bit_ctr[10]), .I1(n37624), 
            .CO(n28652));
    SB_LUT4 mod_5_add_1808_24_lut (.I0(n2588), .I1(n2588), .I2(n2621), 
            .I3(n28651), .O(n2687)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_24_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1808_23_lut (.I0(n2589), .I1(n2589), .I2(n2621), 
            .I3(n28650), .O(n2688)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_23_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 add_21_24_lut (.I0(GND_net), .I1(bit_ctr[22]), .I2(GND_net), 
            .I3(n27785), .O(n255[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1808_23 (.CI(n28650), .I0(n2589), .I1(n2621), .CO(n28651));
    SB_LUT4 mod_5_add_1808_22_lut (.I0(n2590), .I1(n2590), .I2(n2621), 
            .I3(n28649), .O(n2689)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_22_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY add_21_24 (.CI(n27785), .I0(bit_ctr[22]), .I1(GND_net), .CO(n27786));
    SB_CARRY mod_5_add_1808_22 (.CI(n28649), .I0(n2590), .I1(n2621), .CO(n28650));
    SB_LUT4 mod_5_add_1808_21_lut (.I0(n2591), .I1(n2591), .I2(n2621), 
            .I3(n28648), .O(n2690)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_21_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1808_21 (.CI(n28648), .I0(n2591), .I1(n2621), .CO(n28649));
    SB_LUT4 mod_5_add_1808_20_lut (.I0(n2592), .I1(n2592), .I2(n2621), 
            .I3(n28647), .O(n2691)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_20_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i19466_2_lut (.I0(bit_ctr[21]), .I1(n1409), .I2(GND_net), 
            .I3(GND_net), .O(n24609));
    defparam i19466_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY mod_5_add_1808_20 (.CI(n28647), .I0(n2592), .I1(n2621), .CO(n28648));
    SB_LUT4 mod_5_add_1808_19_lut (.I0(n2593), .I1(n2593), .I2(n2621), 
            .I3(n28646), .O(n2692)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_19_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1808_19 (.CI(n28646), .I0(n2593), .I1(n2621), .CO(n28647));
    SB_LUT4 mod_5_add_1808_18_lut (.I0(n2594), .I1(n2594), .I2(n2621), 
            .I3(n28645), .O(n2693)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_18_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1808_18 (.CI(n28645), .I0(n2594), .I1(n2621), .CO(n28646));
    SB_LUT4 mod_5_add_1808_17_lut (.I0(n2595), .I1(n2595), .I2(n2621), 
            .I3(n28644), .O(n2694)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_17_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1808_17 (.CI(n28644), .I0(n2595), .I1(n2621), .CO(n28645));
    SB_DFFESR bit_ctr_i0_i26 (.Q(bit_ctr[26]), .C(clk32MHz), .E(n18566), 
            .D(n255[26]), .R(n18886));   // verilog/neopixel.v(35[12] 117[6])
    SB_LUT4 mod_5_add_1808_16_lut (.I0(n2596), .I1(n2596), .I2(n2621), 
            .I3(n28643), .O(n2695)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_16_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i6_4_lut (.I0(n1405), .I1(n24609), .I2(n1407), .I3(n1400), 
            .O(n16_adj_4749));
    defparam i6_4_lut.LUT_INIT = 16'hfffe;
    SB_CARRY mod_5_add_1808_16 (.CI(n28643), .I0(n2596), .I1(n2621), .CO(n28644));
    SB_LUT4 mod_5_add_1808_15_lut (.I0(n2597), .I1(n2597), .I2(n2621), 
            .I3(n28642), .O(n2696)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_15_lut.LUT_INIT = 16'hCA3A;
    SB_DFFESR bit_ctr_i0_i27 (.Q(bit_ctr[27]), .C(clk32MHz), .E(n18566), 
            .D(n255[27]), .R(n18886));   // verilog/neopixel.v(35[12] 117[6])
    SB_LUT4 i7_4_lut_adj_1520 (.I0(n1402), .I1(n1403), .I2(n1401), .I3(n1406), 
            .O(n17_adj_4750));
    defparam i7_4_lut_adj_1520.LUT_INIT = 16'hfffe;
    SB_LUT4 i9_4_lut_adj_1521 (.I0(n17_adj_4750), .I1(n1408), .I2(n16_adj_4749), 
            .I3(n1404), .O(n1433));
    defparam i9_4_lut_adj_1521.LUT_INIT = 16'hfffe;
    SB_CARRY mod_5_add_1808_15 (.CI(n28642), .I0(n2597), .I1(n2621), .CO(n28643));
    SB_LUT4 mod_5_add_1808_14_lut (.I0(n2598), .I1(n2598), .I2(n2621), 
            .I3(n28641), .O(n2697)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_14_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1808_14 (.CI(n28641), .I0(n2598), .I1(n2621), .CO(n28642));
    SB_LUT4 i30886_1_lut (.I0(n1037), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n37639));   // verilog/neopixel.v(18[12:19])
    defparam i30886_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mod_5_add_1808_13_lut (.I0(n2599), .I1(n2599), .I2(n2621), 
            .I3(n28640), .O(n2698)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_13_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i18573_3_lut (.I0(bit_ctr[26]), .I1(n971[26]), .I2(n2), .I3(GND_net), 
            .O(n1009));
    defparam i18573_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i30422_2_lut (.I0(n2), .I1(n971[28]), .I2(GND_net), .I3(GND_net), 
            .O(n1007));   // verilog/neopixel.v(22[26:36])
    defparam i30422_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i30411_2_lut (.I0(n2), .I1(n971[29]), .I2(GND_net), .I3(GND_net), 
            .O(n1006));
    defparam i30411_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i30427_2_lut (.I0(n2), .I1(n971[30]), .I2(GND_net), .I3(GND_net), 
            .O(n1005));   // verilog/neopixel.v(22[26:36])
    defparam i30427_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i18579_3_lut (.I0(n16024), .I1(n971[27]), .I2(n2), .I3(GND_net), 
            .O(n1008));
    defparam i18579_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i28559_3_lut (.I0(n906), .I1(n905), .I2(n907), .I3(GND_net), 
            .O(n35312));
    defparam i28559_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i4_4_lut (.I0(n18794), .I1(n35312), .I2(bit_ctr[26]), .I3(n16024), 
            .O(n2));
    defparam i4_4_lut.LUT_INIT = 16'h0111;
    SB_LUT4 i29800_3_lut (.I0(n971[26]), .I1(n971[29]), .I2(bit_ctr[25]), 
            .I3(GND_net), .O(n36260));
    defparam i29800_3_lut.LUT_INIT = 16'hecec;
    SB_LUT4 i29802_2_lut (.I0(bit_ctr[25]), .I1(bit_ctr[26]), .I2(GND_net), 
            .I3(GND_net), .O(n36262));
    defparam i29802_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i28603_3_lut (.I0(n971[30]), .I1(n971[28]), .I2(n971[31]), 
            .I3(GND_net), .O(n35358));
    defparam i28603_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i41_4_lut (.I0(n36262), .I1(n36260), .I2(n2), .I3(n907), 
            .O(n38_adj_4751));
    defparam i41_4_lut.LUT_INIT = 16'hfcac;
    SB_LUT4 i4_4_lut_adj_1522 (.I0(n38_adj_4751), .I1(n2), .I2(n1008), 
            .I3(n35358), .O(n1037));   // verilog/neopixel.v(18[12:19])
    defparam i4_4_lut_adj_1522.LUT_INIT = 16'hfbfa;
    SB_LUT4 i30451_2_lut (.I0(n2), .I1(n971[31]), .I2(GND_net), .I3(GND_net), 
            .O(n4));   // verilog/neopixel.v(22[26:36])
    defparam i30451_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 sub_14_inv_0_i21_1_lut (.I0(\neo_pixel_transmitter.t0 [20]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[20]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i21_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i22_1_lut (.I0(\neo_pixel_transmitter.t0 [21]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[21]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i22_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY mod_5_add_1808_13 (.CI(n28640), .I0(n2599), .I1(n2621), .CO(n28641));
    SB_LUT4 sub_14_inv_0_i23_1_lut (.I0(\neo_pixel_transmitter.t0 [22]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[22]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i23_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mod_5_add_1808_12_lut (.I0(n2600), .I1(n2600), .I2(n2621), 
            .I3(n28639), .O(n2699)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_12_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1808_12 (.CI(n28639), .I0(n2600), .I1(n2621), .CO(n28640));
    SB_LUT4 mod_5_add_1808_11_lut (.I0(n2601), .I1(n2601), .I2(n2621), 
            .I3(n28638), .O(n2700)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_11_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1808_11 (.CI(n28638), .I0(n2601), .I1(n2621), .CO(n28639));
    SB_LUT4 sub_14_inv_0_i24_1_lut (.I0(\neo_pixel_transmitter.t0 [23]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[23]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i24_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mod_5_add_1808_10_lut (.I0(n2602), .I1(n2602), .I2(n2621), 
            .I3(n28637), .O(n2701)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_10_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i30884_1_lut (.I0(n1136), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n37637));
    defparam i30884_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY mod_5_add_1808_10 (.CI(n28637), .I0(n2602), .I1(n2621), .CO(n28638));
    SB_LUT4 i19464_2_lut (.I0(bit_ctr[24]), .I1(n1109), .I2(GND_net), 
            .I3(GND_net), .O(n24607));
    defparam i19464_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i5_4_lut (.I0(n1105), .I1(n1103), .I2(n24607), .I3(n1108), 
            .O(n12_adj_4755));
    defparam i5_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 mod_5_add_1808_9_lut (.I0(n2603), .I1(n2603), .I2(n2621), 
            .I3(n28636), .O(n2702)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_9_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i6_4_lut_adj_1523 (.I0(n1107), .I1(n12_adj_4755), .I2(n1106), 
            .I3(n1104), .O(n1136));
    defparam i6_4_lut_adj_1523.LUT_INIT = 16'hfffe;
    SB_LUT4 sub_14_inv_0_i25_1_lut (.I0(\neo_pixel_transmitter.t0 [24]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[24]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i25_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY mod_5_add_1808_9 (.CI(n28636), .I0(n2603), .I1(n2621), .CO(n28637));
    SB_LUT4 i30883_1_lut (.I0(n3116), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n37636));
    defparam i30883_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mod_5_add_1808_8_lut (.I0(n2604), .I1(n2604), .I2(n2621), 
            .I3(n28635), .O(n2703)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_8_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1808_8 (.CI(n28635), .I0(n2604), .I1(n2621), .CO(n28636));
    SB_LUT4 add_21_23_lut (.I0(GND_net), .I1(bit_ctr[21]), .I2(GND_net), 
            .I3(n27784), .O(n255[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_14_inv_0_i26_1_lut (.I0(\neo_pixel_transmitter.t0 [25]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[25]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i26_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mod_5_add_1808_7_lut (.I0(n2605), .I1(n2605), .I2(n2621), 
            .I3(n28634), .O(n2704)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_7_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1808_7 (.CI(n28634), .I0(n2605), .I1(n2621), .CO(n28635));
    SB_LUT4 mod_5_add_1808_6_lut (.I0(n2606), .I1(n2606), .I2(n2621), 
            .I3(n28633), .O(n2705)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_6_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1808_6 (.CI(n28633), .I0(n2606), .I1(n2621), .CO(n28634));
    SB_LUT4 mod_5_add_1808_5_lut (.I0(n2607), .I1(n2607), .I2(n2621), 
            .I3(n28632), .O(n2706)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_5_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1808_5 (.CI(n28632), .I0(n2607), .I1(n2621), .CO(n28633));
    SB_LUT4 mod_5_add_1808_4_lut (.I0(n2608), .I1(n2608), .I2(n2621), 
            .I3(n28631), .O(n2707)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_4_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1808_4 (.CI(n28631), .I0(n2608), .I1(n2621), .CO(n28632));
    SB_LUT4 mod_5_add_1406_16_lut (.I0(n1996), .I1(n1996), .I2(n2027), 
            .I3(n28784), .O(n2095)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_16_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1808_3_lut (.I0(n2609), .I1(n2609), .I2(n37626), 
            .I3(n28630), .O(n2708)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_3_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1808_3 (.CI(n28630), .I0(n2609), .I1(n37626), .CO(n28631));
    SB_DFFESR bit_ctr_i0_i28 (.Q(bit_ctr[28]), .C(clk32MHz), .E(n18566), 
            .D(n255[28]), .R(n18886));   // verilog/neopixel.v(35[12] 117[6])
    SB_LUT4 mod_5_add_1808_2_lut (.I0(bit_ctr[9]), .I1(bit_ctr[9]), .I2(n37626), 
            .I3(VCC_net), .O(n2709)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_2_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1406_16 (.CI(n28784), .I0(n1996), .I1(n2027), .CO(n28785));
    SB_CARRY add_21_23 (.CI(n27784), .I0(bit_ctr[21]), .I1(GND_net), .CO(n27785));
    SB_CARRY mod_5_add_1808_2 (.CI(VCC_net), .I0(bit_ctr[9]), .I1(n37626), 
            .CO(n28630));
    SB_LUT4 mod_5_add_1406_15_lut (.I0(n1997), .I1(n1997), .I2(n2027), 
            .I3(n28783), .O(n2096)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_15_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 add_21_22_lut (.I0(GND_net), .I1(bit_ctr[20]), .I2(GND_net), 
            .I3(n27783), .O(n255[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i15_4_lut_adj_1524 (.I0(n3102), .I1(n3090), .I2(n3103), .I3(n3085), 
            .O(n42));
    defparam i15_4_lut_adj_1524.LUT_INIT = 16'hfffe;
    SB_LUT4 i19_4_lut (.I0(n3089), .I1(n3094), .I2(n3101), .I3(n3098), 
            .O(n46));
    defparam i19_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i17_4_lut (.I0(n3099), .I1(n3091), .I2(n3106), .I3(n3100), 
            .O(n44));
    defparam i17_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i18_4_lut_adj_1525 (.I0(n3097), .I1(n3088), .I2(n3104), .I3(n3092), 
            .O(n45));
    defparam i18_4_lut_adj_1525.LUT_INIT = 16'hfffe;
    SB_LUT4 i16_4_lut_adj_1526 (.I0(n3105), .I1(n3083), .I2(n3093), .I3(n3096), 
            .O(n43));
    defparam i16_4_lut_adj_1526.LUT_INIT = 16'hfffe;
    SB_LUT4 i13_3_lut (.I0(bit_ctr[4]), .I1(n3108), .I2(n3109), .I3(GND_net), 
            .O(n40_adj_4756));
    defparam i13_3_lut.LUT_INIT = 16'hecec;
    SB_CARRY mod_5_add_1406_15 (.CI(n28783), .I0(n1997), .I1(n2027), .CO(n28784));
    SB_LUT4 i21_4_lut_adj_1527 (.I0(n3107), .I1(n42), .I2(n3087), .I3(n3086), 
            .O(n48));
    defparam i21_4_lut_adj_1527.LUT_INIT = 16'hfffe;
    SB_LUT4 i25_4_lut (.I0(n43), .I1(n45), .I2(n44), .I3(n46), .O(n52));
    defparam i25_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i12_2_lut (.I0(n3095), .I1(n3084), .I2(GND_net), .I3(GND_net), 
            .O(n39_adj_4757));
    defparam i12_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i26_4_lut (.I0(n39_adj_4757), .I1(n52), .I2(n48), .I3(n40_adj_4756), 
            .O(n3116));
    defparam i26_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 sub_14_inv_0_i27_1_lut (.I0(\neo_pixel_transmitter.t0 [26]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[26]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i27_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i30882_1_lut (.I0(n3017), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n37635));
    defparam i30882_1_lut.LUT_INIT = 16'h5555;
    SB_DFFESR bit_ctr_i0_i29 (.Q(bit_ctr[29]), .C(clk32MHz), .E(n18566), 
            .D(n255[29]), .R(n18886));   // verilog/neopixel.v(35[12] 117[6])
    SB_LUT4 i30881_1_lut (.I0(n2324), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n37634));
    defparam i30881_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i28_1_lut (.I0(\neo_pixel_transmitter.t0 [27]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[27]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i28_1_lut.LUT_INIT = 16'h5555;
    SB_DFFESR bit_ctr_i0_i30 (.Q(bit_ctr[30]), .C(clk32MHz), .E(n18566), 
            .D(n255[30]), .R(n18886));   // verilog/neopixel.v(35[12] 117[6])
    SB_CARRY add_21_22 (.CI(n27783), .I0(bit_ctr[20]), .I1(GND_net), .CO(n27784));
    SB_LUT4 add_21_21_lut (.I0(GND_net), .I1(bit_ctr[19]), .I2(GND_net), 
            .I3(n27782), .O(n255[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_1406_14_lut (.I0(n1998), .I1(n1998), .I2(n2027), 
            .I3(n28782), .O(n2097)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_14_lut.LUT_INIT = 16'hCA3A;
    SB_DFFESR bit_ctr_i0_i31 (.Q(bit_ctr[31]), .C(clk32MHz), .E(n18566), 
            .D(n255[31]), .R(n18886));   // verilog/neopixel.v(35[12] 117[6])
    SB_CARRY add_21_7 (.CI(n27768), .I0(bit_ctr[5]), .I1(GND_net), .CO(n27769));
    SB_LUT4 add_21_6_lut (.I0(GND_net), .I1(bit_ctr[4]), .I2(GND_net), 
            .I3(n27767), .O(n255[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1406_14 (.CI(n28782), .I0(n1998), .I1(n2027), .CO(n28783));
    SB_CARRY add_21_6 (.CI(n27767), .I0(bit_ctr[4]), .I1(GND_net), .CO(n27768));
    SB_LUT4 mod_5_add_1406_13_lut (.I0(n1999), .I1(n1999), .I2(n2027), 
            .I3(n28781), .O(n2098)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_13_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1406_13 (.CI(n28781), .I0(n1999), .I1(n2027), .CO(n28782));
    SB_LUT4 mod_5_add_1406_12_lut (.I0(n2000), .I1(n2000), .I2(n2027), 
            .I3(n28780), .O(n2099)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_12_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY add_21_21 (.CI(n27782), .I0(bit_ctr[19]), .I1(GND_net), .CO(n27783));
    SB_LUT4 add_21_20_lut (.I0(GND_net), .I1(bit_ctr[18]), .I2(GND_net), 
            .I3(n27781), .O(n255[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1406_12 (.CI(n28780), .I0(n2000), .I1(n2027), .CO(n28781));
    SB_LUT4 add_21_5_lut (.I0(GND_net), .I1(bit_ctr[3]), .I2(GND_net), 
            .I3(n27766), .O(n255[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_21_5 (.CI(n27766), .I0(bit_ctr[3]), .I1(GND_net), .CO(n27767));
    SB_LUT4 mod_5_add_1406_11_lut (.I0(n2001), .I1(n2001), .I2(n2027), 
            .I3(n28779), .O(n2100)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_11_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY add_21_20 (.CI(n27781), .I0(bit_ctr[18]), .I1(GND_net), .CO(n27782));
    SB_LUT4 add_21_19_lut (.I0(GND_net), .I1(bit_ctr[17]), .I2(GND_net), 
            .I3(n27780), .O(n255[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_14_inv_0_i29_1_lut (.I0(\neo_pixel_transmitter.t0 [28]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[28]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i29_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_21_4_lut (.I0(GND_net), .I1(bit_ctr[2]), .I2(GND_net), 
            .I3(n27765), .O(n255[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1406_11 (.CI(n28779), .I0(n2001), .I1(n2027), .CO(n28780));
    SB_LUT4 mod_5_add_1406_10_lut (.I0(n2002), .I1(n2002), .I2(n2027), 
            .I3(n28778), .O(n2101)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_10_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1406_10 (.CI(n28778), .I0(n2002), .I1(n2027), .CO(n28779));
    SB_LUT4 mod_5_add_1406_9_lut (.I0(n2003), .I1(n2003), .I2(n2027), 
            .I3(n28777), .O(n2102)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_9_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1406_9 (.CI(n28777), .I0(n2003), .I1(n2027), .CO(n28778));
    SB_CARRY add_21_4 (.CI(n27765), .I0(bit_ctr[2]), .I1(GND_net), .CO(n27766));
    SB_LUT4 mod_5_add_1406_8_lut (.I0(n2004), .I1(n2004), .I2(n2027), 
            .I3(n28776), .O(n2103)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_8_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1406_8 (.CI(n28776), .I0(n2004), .I1(n2027), .CO(n28777));
    SB_LUT4 sub_14_inv_0_i30_1_lut (.I0(\neo_pixel_transmitter.t0 [29]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[29]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i30_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_21_19 (.CI(n27780), .I0(bit_ctr[17]), .I1(GND_net), .CO(n27781));
    SB_LUT4 mod_5_add_1406_7_lut (.I0(n2005), .I1(n2005), .I2(n2027), 
            .I3(n28775), .O(n2104)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_7_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1406_7 (.CI(n28775), .I0(n2005), .I1(n2027), .CO(n28776));
    SB_LUT4 mod_5_add_1406_6_lut (.I0(n2006), .I1(n2006), .I2(n2027), 
            .I3(n28774), .O(n2105)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_6_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1406_6 (.CI(n28774), .I0(n2006), .I1(n2027), .CO(n28775));
    SB_LUT4 add_21_3_lut (.I0(GND_net), .I1(bit_ctr[1]), .I2(GND_net), 
            .I3(n27764), .O(n255[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_1406_5_lut (.I0(n2007), .I1(n2007), .I2(n2027), 
            .I3(n28773), .O(n2106)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_5_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1406_5 (.CI(n28773), .I0(n2007), .I1(n2027), .CO(n28774));
    SB_LUT4 i16_4_lut_adj_1528 (.I0(n3007), .I1(n2988), .I2(n2986), .I3(n2993), 
            .O(n42_adj_4759));
    defparam i16_4_lut_adj_1528.LUT_INIT = 16'hfffe;
    SB_LUT4 i3_3_lut_adj_1529 (.I0(bit_ctr[5]), .I1(n3003), .I2(n3009), 
            .I3(GND_net), .O(n29_adj_4760));
    defparam i3_3_lut_adj_1529.LUT_INIT = 16'hecec;
    SB_LUT4 mod_5_add_1406_4_lut (.I0(n2008), .I1(n2008), .I2(n2027), 
            .I3(n28772), .O(n2107)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_4_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1406_4 (.CI(n28772), .I0(n2008), .I1(n2027), .CO(n28773));
    SB_LUT4 mod_5_add_1406_3_lut (.I0(n2009), .I1(n2009), .I2(n37625), 
            .I3(n28771), .O(n2108)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_3_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 i14_4_lut_adj_1530 (.I0(n3008), .I1(n3002), .I2(n3004), .I3(n2996), 
            .O(n40_adj_4761));
    defparam i14_4_lut_adj_1530.LUT_INIT = 16'hfffe;
    SB_LUT4 i19_4_lut_adj_1531 (.I0(n2994), .I1(n2995), .I2(n2999), .I3(n2985), 
            .O(n45_adj_4762));
    defparam i19_4_lut_adj_1531.LUT_INIT = 16'hfffe;
    SB_CARRY mod_5_add_1406_3 (.CI(n28771), .I0(n2009), .I1(n37625), .CO(n28772));
    SB_LUT4 mod_5_add_1406_2_lut (.I0(bit_ctr[15]), .I1(bit_ctr[15]), .I2(n37625), 
            .I3(VCC_net), .O(n2109)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_2_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 i18_4_lut_adj_1532 (.I0(n2989), .I1(n2990), .I2(n2984), .I3(n3006), 
            .O(n44_adj_4763));
    defparam i18_4_lut_adj_1532.LUT_INIT = 16'hfffe;
    SB_LUT4 i17_4_lut_adj_1533 (.I0(n2997), .I1(n2998), .I2(n2987), .I3(n3005), 
            .O(n43_adj_4764));
    defparam i17_4_lut_adj_1533.LUT_INIT = 16'hfffe;
    SB_LUT4 i21_4_lut_adj_1534 (.I0(n29_adj_4760), .I1(n42_adj_4759), .I2(n2991), 
            .I3(n2992), .O(n47));
    defparam i21_4_lut_adj_1534.LUT_INIT = 16'hfffe;
    SB_LUT4 i23_4_lut (.I0(n45_adj_4762), .I1(n3001), .I2(n40_adj_4761), 
            .I3(n3000), .O(n49));
    defparam i23_4_lut.LUT_INIT = 16'hfffe;
    SB_CARRY mod_5_add_1406_2 (.CI(VCC_net), .I0(bit_ctr[15]), .I1(n37625), 
            .CO(n28771));
    SB_CARRY add_21_3 (.CI(n27764), .I0(bit_ctr[1]), .I1(GND_net), .CO(n27765));
    SB_LUT4 i25_4_lut_adj_1535 (.I0(n49), .I1(n47), .I2(n43_adj_4764), 
            .I3(n44_adj_4763), .O(n3017));
    defparam i25_4_lut_adj_1535.LUT_INIT = 16'hfffe;
    SB_LUT4 mod_5_add_937_11_lut (.I0(n1301), .I1(n1301), .I2(n1334), 
            .I3(n28105), .O(n1400)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_937_11_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_937_10_lut (.I0(n1302), .I1(n1302), .I2(n1334), 
            .I3(n28104), .O(n1401)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_937_10_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_937_10 (.CI(n28104), .I0(n1302), .I1(n1334), .CO(n28105));
    SB_LUT4 sub_14_inv_0_i31_1_lut (.I0(\neo_pixel_transmitter.t0 [30]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[30]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i31_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i32_1_lut (.I0(\neo_pixel_transmitter.t0 [31]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[31]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i32_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mod_5_add_937_9_lut (.I0(n1303), .I1(n1303), .I2(n1334), .I3(n28103), 
            .O(n1402)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_937_9_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1473_19_lut (.I0(n2093), .I1(n2093), .I2(n2126), 
            .I3(n28770), .O(n2192)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_19_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i30879_1_lut (.I0(n2918), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n37632));
    defparam i30879_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY mod_5_add_937_9 (.CI(n28103), .I0(n1303), .I1(n1334), .CO(n28104));
    SB_LUT4 mod_5_add_1473_18_lut (.I0(n2094), .I1(n2094), .I2(n2126), 
            .I3(n28769), .O(n2193)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_18_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1473_18 (.CI(n28769), .I0(n2094), .I1(n2126), .CO(n28770));
    SB_LUT4 mod_5_add_1473_17_lut (.I0(n2095), .I1(n2095), .I2(n2126), 
            .I3(n28768), .O(n2194)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_17_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_937_8_lut (.I0(n1304), .I1(n1304), .I2(n1334), .I3(n28102), 
            .O(n1403)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_937_8_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1473_17 (.CI(n28768), .I0(n2095), .I1(n2126), .CO(n28769));
    SB_LUT4 mod_5_add_1473_16_lut (.I0(n2096), .I1(n2096), .I2(n2126), 
            .I3(n28767), .O(n2195)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_16_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 add_21_18_lut (.I0(GND_net), .I1(bit_ctr[16]), .I2(GND_net), 
            .I3(n27779), .O(n255[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1473_16 (.CI(n28767), .I0(n2096), .I1(n2126), .CO(n28768));
    SB_LUT4 mod_5_add_1473_15_lut (.I0(n2097), .I1(n2097), .I2(n2126), 
            .I3(n28766), .O(n2196)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_15_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_937_8 (.CI(n28102), .I0(n1304), .I1(n1334), .CO(n28103));
    SB_CARRY mod_5_add_1473_15 (.CI(n28766), .I0(n2097), .I1(n2126), .CO(n28767));
    SB_LUT4 mod_5_add_1473_14_lut (.I0(n2098), .I1(n2098), .I2(n2126), 
            .I3(n28765), .O(n2197)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_14_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1473_14 (.CI(n28765), .I0(n2098), .I1(n2126), .CO(n28766));
    SB_LUT4 mod_5_add_1473_13_lut (.I0(n2099), .I1(n2099), .I2(n2126), 
            .I3(n28764), .O(n2198)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_13_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_937_7_lut (.I0(n1305), .I1(n1305), .I2(n1334), .I3(n28101), 
            .O(n1404)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_937_7_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_937_7 (.CI(n28101), .I0(n1305), .I1(n1334), .CO(n28102));
    SB_LUT4 mod_5_add_937_6_lut (.I0(n1306), .I1(n1306), .I2(n1334), .I3(n28100), 
            .O(n1405)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_937_6_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_937_6 (.CI(n28100), .I0(n1306), .I1(n1334), .CO(n28101));
    SB_LUT4 mod_5_add_937_5_lut (.I0(n1307), .I1(n1307), .I2(n1334), .I3(n28099), 
            .O(n1406)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_937_5_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_937_5 (.CI(n28099), .I0(n1307), .I1(n1334), .CO(n28100));
    SB_LUT4 mod_5_add_937_4_lut (.I0(n1308), .I1(n1308), .I2(n1334), .I3(n28098), 
            .O(n1407)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_937_4_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY add_21_18 (.CI(n27779), .I0(bit_ctr[16]), .I1(GND_net), .CO(n27780));
    SB_CARRY mod_5_add_1473_13 (.CI(n28764), .I0(n2099), .I1(n2126), .CO(n28765));
    SB_LUT4 mod_5_add_1473_12_lut (.I0(n2100), .I1(n2100), .I2(n2126), 
            .I3(n28763), .O(n2199)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_12_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_937_4 (.CI(n28098), .I0(n1308), .I1(n1334), .CO(n28099));
    SB_CARRY mod_5_add_1473_12 (.CI(n28763), .I0(n2100), .I1(n2126), .CO(n28764));
    SB_LUT4 mod_5_add_1473_11_lut (.I0(n2101), .I1(n2101), .I2(n2126), 
            .I3(n28762), .O(n2200)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_11_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 add_21_17_lut (.I0(GND_net), .I1(bit_ctr[15]), .I2(GND_net), 
            .I3(n27778), .O(n255[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_937_3_lut (.I0(n1309), .I1(n1309), .I2(n37627), 
            .I3(n28097), .O(n1408)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_937_3_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 mod_5_add_1875_25_lut (.I0(n2687), .I1(n2687), .I2(n2720), 
            .I3(n28566), .O(n2786)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_25_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1875_24_lut (.I0(n2688), .I1(n2688), .I2(n2720), 
            .I3(n28565), .O(n2787)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_24_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1875_24 (.CI(n28565), .I0(n2688), .I1(n2720), .CO(n28566));
    SB_LUT4 mod_5_add_1875_23_lut (.I0(n2689), .I1(n2689), .I2(n2720), 
            .I3(n28564), .O(n2788)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_23_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1875_23 (.CI(n28564), .I0(n2689), .I1(n2720), .CO(n28565));
    SB_LUT4 mod_5_add_1875_22_lut (.I0(n2690), .I1(n2690), .I2(n2720), 
            .I3(n28563), .O(n2789)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_22_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1875_22 (.CI(n28563), .I0(n2690), .I1(n2720), .CO(n28564));
    SB_LUT4 mod_5_add_1875_21_lut (.I0(n2691), .I1(n2691), .I2(n2720), 
            .I3(n28562), .O(n2790)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_21_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1875_21 (.CI(n28562), .I0(n2691), .I1(n2720), .CO(n28563));
    SB_LUT4 mod_5_add_1875_20_lut (.I0(n2692), .I1(n2692), .I2(n2720), 
            .I3(n28561), .O(n2791)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_20_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1875_20 (.CI(n28561), .I0(n2692), .I1(n2720), .CO(n28562));
    SB_LUT4 mod_5_add_1875_19_lut (.I0(n2693), .I1(n2693), .I2(n2720), 
            .I3(n28560), .O(n2792)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_19_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY add_21_17 (.CI(n27778), .I0(bit_ctr[15]), .I1(GND_net), .CO(n27779));
    SB_CARRY mod_5_add_1473_11 (.CI(n28762), .I0(n2101), .I1(n2126), .CO(n28763));
    SB_CARRY mod_5_add_1875_19 (.CI(n28560), .I0(n2693), .I1(n2720), .CO(n28561));
    SB_LUT4 mod_5_add_1875_18_lut (.I0(n2694), .I1(n2694), .I2(n2720), 
            .I3(n28559), .O(n2793)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_18_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1473_10_lut (.I0(n2102), .I1(n2102), .I2(n2126), 
            .I3(n28761), .O(n2201)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_10_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1875_18 (.CI(n28559), .I0(n2694), .I1(n2720), .CO(n28560));
    SB_LUT4 mod_5_add_1875_17_lut (.I0(n2695), .I1(n2695), .I2(n2720), 
            .I3(n28558), .O(n2794)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_17_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1875_17 (.CI(n28558), .I0(n2695), .I1(n2720), .CO(n28559));
    SB_CARRY mod_5_add_937_3 (.CI(n28097), .I0(n1309), .I1(n37627), .CO(n28098));
    SB_CARRY mod_5_add_1473_10 (.CI(n28761), .I0(n2102), .I1(n2126), .CO(n28762));
    SB_LUT4 mod_5_add_1875_16_lut (.I0(n2696), .I1(n2696), .I2(n2720), 
            .I3(n28557), .O(n2795)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_16_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1875_16 (.CI(n28557), .I0(n2696), .I1(n2720), .CO(n28558));
    SB_LUT4 mod_5_add_937_2_lut (.I0(bit_ctr[22]), .I1(bit_ctr[22]), .I2(n37627), 
            .I3(VCC_net), .O(n1409)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_937_2_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 mod_5_add_1875_15_lut (.I0(n2697), .I1(n2697), .I2(n2720), 
            .I3(n28556), .O(n2796)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_15_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_937_2 (.CI(VCC_net), .I0(bit_ctr[22]), .I1(n37627), 
            .CO(n28097));
    SB_LUT4 add_21_16_lut (.I0(GND_net), .I1(bit_ctr[14]), .I2(GND_net), 
            .I3(n27777), .O(n255[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1875_15 (.CI(n28556), .I0(n2697), .I1(n2720), .CO(n28557));
    SB_CARRY add_21_16 (.CI(n27777), .I0(bit_ctr[14]), .I1(GND_net), .CO(n27778));
    SB_LUT4 mod_5_add_1875_14_lut (.I0(n2698), .I1(n2698), .I2(n2720), 
            .I3(n28555), .O(n2797)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_14_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1473_9_lut (.I0(n2103), .I1(n2103), .I2(n2126), 
            .I3(n28760), .O(n2202)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_9_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1875_14 (.CI(n28555), .I0(n2698), .I1(n2720), .CO(n28556));
    SB_CARRY mod_5_add_1473_9 (.CI(n28760), .I0(n2103), .I1(n2126), .CO(n28761));
    SB_LUT4 add_21_15_lut (.I0(GND_net), .I1(bit_ctr[13]), .I2(GND_net), 
            .I3(n27776), .O(n255[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_21_15 (.CI(n27776), .I0(bit_ctr[13]), .I1(GND_net), .CO(n27777));
    SB_LUT4 mod_5_add_1473_8_lut (.I0(n2104), .I1(n2104), .I2(n2126), 
            .I3(n28759), .O(n2203)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_8_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1875_13_lut (.I0(n2699), .I1(n2699), .I2(n2720), 
            .I3(n28554), .O(n2798)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_13_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1875_13 (.CI(n28554), .I0(n2699), .I1(n2720), .CO(n28555));
    SB_LUT4 mod_5_add_1875_12_lut (.I0(n2700), .I1(n2700), .I2(n2720), 
            .I3(n28553), .O(n2799)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_12_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1875_12 (.CI(n28553), .I0(n2700), .I1(n2720), .CO(n28554));
    SB_CARRY mod_5_add_1473_8 (.CI(n28759), .I0(n2104), .I1(n2126), .CO(n28760));
    SB_LUT4 mod_5_add_1875_11_lut (.I0(n2701), .I1(n2701), .I2(n2720), 
            .I3(n28552), .O(n2800)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_11_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1473_7_lut (.I0(n2105), .I1(n2105), .I2(n2126), 
            .I3(n28758), .O(n2204)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_7_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1473_7 (.CI(n28758), .I0(n2105), .I1(n2126), .CO(n28759));
    SB_LUT4 mod_5_add_1473_6_lut (.I0(n2106), .I1(n2106), .I2(n2126), 
            .I3(n28757), .O(n2205)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_6_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1473_6 (.CI(n28757), .I0(n2106), .I1(n2126), .CO(n28758));
    SB_LUT4 mod_5_add_1473_5_lut (.I0(n2107), .I1(n2107), .I2(n2126), 
            .I3(n28756), .O(n2206)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_5_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1875_11 (.CI(n28552), .I0(n2701), .I1(n2720), .CO(n28553));
    SB_CARRY mod_5_add_1473_5 (.CI(n28756), .I0(n2107), .I1(n2126), .CO(n28757));
    SB_LUT4 mod_5_add_1875_10_lut (.I0(n2702), .I1(n2702), .I2(n2720), 
            .I3(n28551), .O(n2801)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_10_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1875_10 (.CI(n28551), .I0(n2702), .I1(n2720), .CO(n28552));
    SB_LUT4 mod_5_add_1875_9_lut (.I0(n2703), .I1(n2703), .I2(n2720), 
            .I3(n28550), .O(n2802)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_9_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1875_9 (.CI(n28550), .I0(n2703), .I1(n2720), .CO(n28551));
    SB_LUT4 mod_5_add_1875_8_lut (.I0(n2704), .I1(n2704), .I2(n2720), 
            .I3(n28549), .O(n2803)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_8_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1875_8 (.CI(n28549), .I0(n2704), .I1(n2720), .CO(n28550));
    SB_LUT4 mod_5_add_1875_7_lut (.I0(n2705), .I1(n2705), .I2(n2720), 
            .I3(n28548), .O(n2804)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_7_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1875_7 (.CI(n28548), .I0(n2705), .I1(n2720), .CO(n28549));
    SB_LUT4 mod_5_add_1473_4_lut (.I0(n2108), .I1(n2108), .I2(n2126), 
            .I3(n28755), .O(n2207)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_4_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1875_6_lut (.I0(n2706), .I1(n2706), .I2(n2720), 
            .I3(n28547), .O(n2805)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_6_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1875_6 (.CI(n28547), .I0(n2706), .I1(n2720), .CO(n28548));
    SB_LUT4 mod_5_add_1875_5_lut (.I0(n2707), .I1(n2707), .I2(n2720), 
            .I3(n28546), .O(n2806)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_5_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1473_4 (.CI(n28755), .I0(n2108), .I1(n2126), .CO(n28756));
    SB_LUT4 mod_5_add_1473_3_lut (.I0(n2109), .I1(n2109), .I2(n37628), 
            .I3(n28754), .O(n2208)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_3_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1875_5 (.CI(n28546), .I0(n2707), .I1(n2720), .CO(n28547));
    SB_CARRY mod_5_add_1473_3 (.CI(n28754), .I0(n2109), .I1(n37628), .CO(n28755));
    SB_LUT4 mod_5_add_1473_2_lut (.I0(bit_ctr[14]), .I1(bit_ctr[14]), .I2(n37628), 
            .I3(VCC_net), .O(n2209)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_2_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 mod_5_add_1875_4_lut (.I0(n2708), .I1(n2708), .I2(n2720), 
            .I3(n28545), .O(n2807)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_4_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1473_2 (.CI(VCC_net), .I0(bit_ctr[14]), .I1(n37628), 
            .CO(n28754));
    SB_CARRY mod_5_add_1875_4 (.CI(n28545), .I0(n2708), .I1(n2720), .CO(n28546));
    SB_LUT4 mod_5_add_1875_3_lut (.I0(n2709), .I1(n2709), .I2(n37629), 
            .I3(n28544), .O(n2808)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_3_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 mod_5_add_1540_20_lut (.I0(n2192), .I1(n2192), .I2(n2225), 
            .I3(n28753), .O(n2291)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_20_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1875_3 (.CI(n28544), .I0(n2709), .I1(n37629), .CO(n28545));
    SB_LUT4 mod_5_add_1540_19_lut (.I0(n2193), .I1(n2193), .I2(n2225), 
            .I3(n28752), .O(n2292)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_19_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1540_19 (.CI(n28752), .I0(n2193), .I1(n2225), .CO(n28753));
    SB_LUT4 mod_5_add_1540_18_lut (.I0(n2194), .I1(n2194), .I2(n2225), 
            .I3(n28751), .O(n2293)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_18_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1875_2_lut (.I0(bit_ctr[8]), .I1(bit_ctr[8]), .I2(n37629), 
            .I3(VCC_net), .O(n2809)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_2_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1540_18 (.CI(n28751), .I0(n2194), .I1(n2225), .CO(n28752));
    SB_LUT4 mod_5_add_1540_17_lut (.I0(n2195), .I1(n2195), .I2(n2225), 
            .I3(n28750), .O(n2294)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_17_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1875_2 (.CI(VCC_net), .I0(bit_ctr[8]), .I1(n37629), 
            .CO(n28544));
    SB_LUT4 mod_5_add_1942_26_lut (.I0(n2786), .I1(n2786), .I2(n2819), 
            .I3(n28543), .O(n2885)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_26_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1942_25_lut (.I0(n2787), .I1(n2787), .I2(n2819), 
            .I3(n28542), .O(n2886)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_25_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1942_25 (.CI(n28542), .I0(n2787), .I1(n2819), .CO(n28543));
    SB_DFF timer_1579__i0 (.Q(timer[0]), .C(clk32MHz), .D(n133[0]));   // verilog/neopixel.v(12[12:21])
    SB_LUT4 mod_5_add_1942_24_lut (.I0(n2788), .I1(n2788), .I2(n2819), 
            .I3(n28541), .O(n2887)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_24_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1942_24 (.CI(n28541), .I0(n2788), .I1(n2819), .CO(n28542));
    SB_LUT4 mod_5_add_1942_23_lut (.I0(n2789), .I1(n2789), .I2(n2819), 
            .I3(n28540), .O(n2888)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_23_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1942_23 (.CI(n28540), .I0(n2789), .I1(n2819), .CO(n28541));
    SB_CARRY mod_5_add_1540_17 (.CI(n28750), .I0(n2195), .I1(n2225), .CO(n28751));
    SB_LUT4 mod_5_add_1540_16_lut (.I0(n2196), .I1(n2196), .I2(n2225), 
            .I3(n28749), .O(n2295)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_16_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1942_22_lut (.I0(n2790), .I1(n2790), .I2(n2819), 
            .I3(n28539), .O(n2889)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_22_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1540_16 (.CI(n28749), .I0(n2196), .I1(n2225), .CO(n28750));
    SB_LUT4 mod_5_add_1540_15_lut (.I0(n2197), .I1(n2197), .I2(n2225), 
            .I3(n28748), .O(n2296)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_15_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1942_22 (.CI(n28539), .I0(n2790), .I1(n2819), .CO(n28540));
    SB_LUT4 mod_5_add_1942_21_lut (.I0(n2791), .I1(n2791), .I2(n2819), 
            .I3(n28538), .O(n2890)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_21_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1942_21 (.CI(n28538), .I0(n2791), .I1(n2819), .CO(n28539));
    SB_LUT4 mod_5_add_1942_20_lut (.I0(n2792), .I1(n2792), .I2(n2819), 
            .I3(n28537), .O(n2891)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_20_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1942_20 (.CI(n28537), .I0(n2792), .I1(n2819), .CO(n28538));
    SB_CARRY mod_5_add_1540_15 (.CI(n28748), .I0(n2197), .I1(n2225), .CO(n28749));
    SB_LUT4 mod_5_add_1942_19_lut (.I0(n2793), .I1(n2793), .I2(n2819), 
            .I3(n28536), .O(n2892)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_19_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1942_19 (.CI(n28536), .I0(n2793), .I1(n2819), .CO(n28537));
    SB_LUT4 mod_5_add_1942_18_lut (.I0(n2794), .I1(n2794), .I2(n2819), 
            .I3(n28535), .O(n2893)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_18_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1942_18 (.CI(n28535), .I0(n2794), .I1(n2819), .CO(n28536));
    SB_LUT4 mod_5_add_1942_17_lut (.I0(n2795), .I1(n2795), .I2(n2819), 
            .I3(n28534), .O(n2894)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_17_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1942_17 (.CI(n28534), .I0(n2795), .I1(n2819), .CO(n28535));
    SB_LUT4 mod_5_add_1942_16_lut (.I0(n2796), .I1(n2796), .I2(n2819), 
            .I3(n28533), .O(n2895)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_16_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1540_14_lut (.I0(n2198), .I1(n2198), .I2(n2225), 
            .I3(n28747), .O(n2297)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_14_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1942_16 (.CI(n28533), .I0(n2796), .I1(n2819), .CO(n28534));
    SB_LUT4 mod_5_add_1942_15_lut (.I0(n2797), .I1(n2797), .I2(n2819), 
            .I3(n28532), .O(n2896)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_15_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1942_15 (.CI(n28532), .I0(n2797), .I1(n2819), .CO(n28533));
    SB_LUT4 mod_5_add_1942_14_lut (.I0(n2798), .I1(n2798), .I2(n2819), 
            .I3(n28531), .O(n2897)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_14_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1942_14 (.CI(n28531), .I0(n2798), .I1(n2819), .CO(n28532));
    SB_LUT4 mod_5_add_1942_13_lut (.I0(n2799), .I1(n2799), .I2(n2819), 
            .I3(n28530), .O(n2898)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_13_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1942_13 (.CI(n28530), .I0(n2799), .I1(n2819), .CO(n28531));
    SB_LUT4 mod_5_add_1942_12_lut (.I0(n2800), .I1(n2800), .I2(n2819), 
            .I3(n28529), .O(n2899)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_12_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1942_12 (.CI(n28529), .I0(n2800), .I1(n2819), .CO(n28530));
    SB_LUT4 mod_5_add_1942_11_lut (.I0(n2801), .I1(n2801), .I2(n2819), 
            .I3(n28528), .O(n2900)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_11_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1942_11 (.CI(n28528), .I0(n2801), .I1(n2819), .CO(n28529));
    SB_CARRY mod_5_add_1540_14 (.CI(n28747), .I0(n2198), .I1(n2225), .CO(n28748));
    SB_LUT4 mod_5_add_1942_10_lut (.I0(n2802), .I1(n2802), .I2(n2819), 
            .I3(n28527), .O(n2901)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_10_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1942_10 (.CI(n28527), .I0(n2802), .I1(n2819), .CO(n28528));
    SB_LUT4 mod_5_add_1942_9_lut (.I0(n2803), .I1(n2803), .I2(n2819), 
            .I3(n28526), .O(n2902)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_9_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1942_9 (.CI(n28526), .I0(n2803), .I1(n2819), .CO(n28527));
    SB_LUT4 mod_5_add_1942_8_lut (.I0(n2804), .I1(n2804), .I2(n2819), 
            .I3(n28525), .O(n2903)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_8_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1942_8 (.CI(n28525), .I0(n2804), .I1(n2819), .CO(n28526));
    SB_LUT4 mod_5_add_1540_13_lut (.I0(n2199), .I1(n2199), .I2(n2225), 
            .I3(n28746), .O(n2298)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_13_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i11_4_lut_adj_1536 (.I0(n1903), .I1(n1905), .I2(n1902), .I3(n1897), 
            .O(n26));
    defparam i11_4_lut_adj_1536.LUT_INIT = 16'hfffe;
    SB_CARRY mod_5_add_1540_13 (.CI(n28746), .I0(n2199), .I1(n2225), .CO(n28747));
    SB_LUT4 mod_5_add_1540_12_lut (.I0(n2200), .I1(n2200), .I2(n2225), 
            .I3(n28745), .O(n2299)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_12_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i9_4_lut_adj_1537 (.I0(n1899), .I1(n1906), .I2(n1904), .I3(n1900), 
            .O(n24_adj_4766));
    defparam i9_4_lut_adj_1537.LUT_INIT = 16'hfffe;
    SB_CARRY mod_5_add_1540_12 (.CI(n28745), .I0(n2200), .I1(n2225), .CO(n28746));
    SB_LUT4 mod_5_add_1942_7_lut (.I0(n2805), .I1(n2805), .I2(n2819), 
            .I3(n28524), .O(n2904)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_7_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i10_4_lut_adj_1538 (.I0(n1901), .I1(n1896), .I2(n1895), .I3(n1908), 
            .O(n25_adj_4767));
    defparam i10_4_lut_adj_1538.LUT_INIT = 16'hfffe;
    SB_LUT4 i8_4_lut_adj_1539 (.I0(n1898), .I1(bit_ctr[16]), .I2(n1907), 
            .I3(n1909), .O(n23_adj_4768));
    defparam i8_4_lut_adj_1539.LUT_INIT = 16'hfefa;
    SB_LUT4 i14_4_lut_adj_1540 (.I0(n23_adj_4768), .I1(n25_adj_4767), .I2(n24_adj_4766), 
            .I3(n26), .O(n1928));
    defparam i14_4_lut_adj_1540.LUT_INIT = 16'hfffe;
    SB_CARRY mod_5_add_1942_7 (.CI(n28524), .I0(n2805), .I1(n2819), .CO(n28525));
    SB_LUT4 mod_5_add_1540_11_lut (.I0(n2201), .I1(n2201), .I2(n2225), 
            .I3(n28744), .O(n2300)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_11_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1540_11 (.CI(n28744), .I0(n2201), .I1(n2225), .CO(n28745));
    SB_LUT4 mod_5_add_1942_6_lut (.I0(n2806), .I1(n2806), .I2(n2819), 
            .I3(n28523), .O(n2905)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_6_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1942_6 (.CI(n28523), .I0(n2806), .I1(n2819), .CO(n28524));
    SB_LUT4 mod_5_add_1942_5_lut (.I0(n2807), .I1(n2807), .I2(n2819), 
            .I3(n28522), .O(n2906)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_5_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1942_5 (.CI(n28522), .I0(n2807), .I1(n2819), .CO(n28523));
    SB_LUT4 mod_5_add_1942_4_lut (.I0(n2808), .I1(n2808), .I2(n2819), 
            .I3(n28521), .O(n2907)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_4_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1942_4 (.CI(n28521), .I0(n2808), .I1(n2819), .CO(n28522));
    SB_LUT4 mod_5_add_1942_3_lut (.I0(n2809), .I1(n2809), .I2(n37631), 
            .I3(n28520), .O(n2908)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_3_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1942_3 (.CI(n28520), .I0(n2809), .I1(n37631), .CO(n28521));
    SB_LUT4 mod_5_add_1942_2_lut (.I0(bit_ctr[7]), .I1(bit_ctr[7]), .I2(n37631), 
            .I3(VCC_net), .O(n2909)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_2_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1942_2 (.CI(VCC_net), .I0(bit_ctr[7]), .I1(n37631), 
            .CO(n28520));
    SB_LUT4 mod_5_add_2009_27_lut (.I0(n2885), .I1(n2885), .I2(n2918), 
            .I3(n28519), .O(n2984)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_27_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_2009_26_lut (.I0(n2886), .I1(n2886), .I2(n2918), 
            .I3(n28518), .O(n2985)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_26_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2009_26 (.CI(n28518), .I0(n2886), .I1(n2918), .CO(n28519));
    SB_LUT4 mod_5_add_1540_10_lut (.I0(n2202), .I1(n2202), .I2(n2225), 
            .I3(n28743), .O(n2301)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_10_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1540_10 (.CI(n28743), .I0(n2202), .I1(n2225), .CO(n28744));
    SB_LUT4 mod_5_add_2009_25_lut (.I0(n2887), .I1(n2887), .I2(n2918), 
            .I3(n28517), .O(n2986)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_25_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2009_25 (.CI(n28517), .I0(n2887), .I1(n2918), .CO(n28518));
    SB_LUT4 mod_5_add_2009_24_lut (.I0(n2888), .I1(n2888), .I2(n2918), 
            .I3(n28516), .O(n2987)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_24_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2009_24 (.CI(n28516), .I0(n2888), .I1(n2918), .CO(n28517));
    SB_LUT4 mod_5_add_2009_23_lut (.I0(n2889), .I1(n2889), .I2(n2918), 
            .I3(n28515), .O(n2988)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_23_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2009_23 (.CI(n28515), .I0(n2889), .I1(n2918), .CO(n28516));
    SB_LUT4 mod_5_add_2009_22_lut (.I0(n2890), .I1(n2890), .I2(n2918), 
            .I3(n28514), .O(n2989)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_22_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1540_9_lut (.I0(n2203), .I1(n2203), .I2(n2225), 
            .I3(n28742), .O(n2302)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_9_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 add_21_2_lut (.I0(GND_net), .I1(bit_ctr[0]), .I2(GND_net), 
            .I3(VCC_net), .O(n255[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_2009_22 (.CI(n28514), .I0(n2890), .I1(n2918), .CO(n28515));
    SB_LUT4 mod_5_add_2009_21_lut (.I0(n2891), .I1(n2891), .I2(n2918), 
            .I3(n28513), .O(n2990)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_21_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2009_21 (.CI(n28513), .I0(n2891), .I1(n2918), .CO(n28514));
    SB_LUT4 mod_5_add_2009_20_lut (.I0(n2892), .I1(n2892), .I2(n2918), 
            .I3(n28512), .O(n2991)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_20_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2009_20 (.CI(n28512), .I0(n2892), .I1(n2918), .CO(n28513));
    SB_CARRY mod_5_add_1540_9 (.CI(n28742), .I0(n2203), .I1(n2225), .CO(n28743));
    SB_LUT4 mod_5_add_2009_19_lut (.I0(n2893), .I1(n2893), .I2(n2918), 
            .I3(n28511), .O(n2992)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_19_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1540_8_lut (.I0(n2204), .I1(n2204), .I2(n2225), 
            .I3(n28741), .O(n2303)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_8_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1540_8 (.CI(n28741), .I0(n2204), .I1(n2225), .CO(n28742));
    SB_CARRY mod_5_add_2009_19 (.CI(n28511), .I0(n2893), .I1(n2918), .CO(n28512));
    SB_LUT4 mod_5_add_1540_7_lut (.I0(n2205), .I1(n2205), .I2(n2225), 
            .I3(n28740), .O(n2304)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_7_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_2009_18_lut (.I0(n2894), .I1(n2894), .I2(n2918), 
            .I3(n28510), .O(n2993)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_18_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2009_18 (.CI(n28510), .I0(n2894), .I1(n2918), .CO(n28511));
    SB_CARRY mod_5_add_1540_7 (.CI(n28740), .I0(n2205), .I1(n2225), .CO(n28741));
    SB_LUT4 mod_5_add_2009_17_lut (.I0(n2895), .I1(n2895), .I2(n2918), 
            .I3(n28509), .O(n2994)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_17_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2009_17 (.CI(n28509), .I0(n2895), .I1(n2918), .CO(n28510));
    SB_LUT4 mod_5_add_2009_16_lut (.I0(n2896), .I1(n2896), .I2(n2918), 
            .I3(n28508), .O(n2995)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_16_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i2_2_lut (.I0(n1998), .I1(n2004), .I2(GND_net), .I3(GND_net), 
            .O(n18_adj_4769));
    defparam i2_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i12_4_lut_adj_1541 (.I0(n2003), .I1(n1999), .I2(n1996), .I3(n2007), 
            .O(n28_adj_4770));
    defparam i12_4_lut_adj_1541.LUT_INIT = 16'hfffe;
    SB_LUT4 i10_4_lut_adj_1542 (.I0(n1997), .I1(n2005), .I2(n2000), .I3(n2002), 
            .O(n26_adj_4771));
    defparam i10_4_lut_adj_1542.LUT_INIT = 16'hfffe;
    SB_LUT4 i11_4_lut_adj_1543 (.I0(n2001), .I1(n2008), .I2(n1994), .I3(n1995), 
            .O(n27_adj_4772));
    defparam i11_4_lut_adj_1543.LUT_INIT = 16'hfffe;
    SB_LUT4 mod_5_add_1540_6_lut (.I0(n2206), .I1(n2206), .I2(n2225), 
            .I3(n28739), .O(n2305)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_6_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2009_16 (.CI(n28508), .I0(n2896), .I1(n2918), .CO(n28509));
    SB_LUT4 mod_5_add_2009_15_lut (.I0(n2897), .I1(n2897), .I2(n2918), 
            .I3(n28507), .O(n2996)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_15_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY add_21_2 (.CI(VCC_net), .I0(bit_ctr[0]), .I1(GND_net), .CO(n27764));
    SB_CARRY mod_5_add_1540_6 (.CI(n28739), .I0(n2206), .I1(n2225), .CO(n28740));
    SB_LUT4 mod_5_add_1540_5_lut (.I0(n2207), .I1(n2207), .I2(n2225), 
            .I3(n28738), .O(n2306)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_5_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1540_5 (.CI(n28738), .I0(n2207), .I1(n2225), .CO(n28739));
    SB_LUT4 mod_5_add_1540_4_lut (.I0(n2208), .I1(n2208), .I2(n2225), 
            .I3(n28737), .O(n2307)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_4_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1540_4 (.CI(n28737), .I0(n2208), .I1(n2225), .CO(n28738));
    SB_LUT4 i9_4_lut_adj_1544 (.I0(bit_ctr[15]), .I1(n18_adj_4769), .I2(n2006), 
            .I3(n2009), .O(n25_adj_4773));
    defparam i9_4_lut_adj_1544.LUT_INIT = 16'hfefc;
    SB_LUT4 i15_4_lut_adj_1545 (.I0(n25_adj_4773), .I1(n27_adj_4772), .I2(n26_adj_4771), 
            .I3(n28_adj_4770), .O(n2027));
    defparam i15_4_lut_adj_1545.LUT_INIT = 16'hfffe;
    SB_LUT4 mod_5_add_1540_3_lut (.I0(n2209), .I1(n2209), .I2(n37630), 
            .I3(n28736), .O(n2308)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_3_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 i3_2_lut (.I0(n2491), .I1(n2504), .I2(GND_net), .I3(GND_net), 
            .O(n24_adj_4774));
    defparam i3_2_lut.LUT_INIT = 16'heeee;
    SB_CARRY mod_5_add_1540_3 (.CI(n28736), .I0(n2209), .I1(n37630), .CO(n28737));
    SB_LUT4 i13_4_lut_adj_1546 (.I0(n2496), .I1(n2505), .I2(n2500), .I3(n2499), 
            .O(n34_adj_4775));
    defparam i13_4_lut_adj_1546.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_3_lut_adj_1547 (.I0(bit_ctr[10]), .I1(n2497), .I2(n2509), 
            .I3(GND_net), .O(n22_adj_4776));
    defparam i1_3_lut_adj_1547.LUT_INIT = 16'hecec;
    SB_LUT4 i17_4_lut_adj_1548 (.I0(n2490), .I1(n34_adj_4775), .I2(n24_adj_4774), 
            .I3(n2494), .O(n38_adj_4777));
    defparam i17_4_lut_adj_1548.LUT_INIT = 16'hfffe;
    SB_LUT4 i15_4_lut_adj_1549 (.I0(n2501), .I1(n2502), .I2(n2506), .I3(n2492), 
            .O(n36_adj_4778));
    defparam i15_4_lut_adj_1549.LUT_INIT = 16'hfffe;
    SB_LUT4 i16_4_lut_adj_1550 (.I0(n2495), .I1(n2498), .I2(n2493), .I3(n22_adj_4776), 
            .O(n37_adj_4779));
    defparam i16_4_lut_adj_1550.LUT_INIT = 16'hfffe;
    SB_LUT4 i14_4_lut_adj_1551 (.I0(n2507), .I1(n2508), .I2(n2503), .I3(n2489), 
            .O(n35));
    defparam i14_4_lut_adj_1551.LUT_INIT = 16'hfffe;
    SB_LUT4 i20_4_lut (.I0(n35), .I1(n37_adj_4779), .I2(n36_adj_4778), 
            .I3(n38_adj_4777), .O(n2522));
    defparam i20_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i30870_1_lut (.I0(n2423), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n37623));
    defparam i30870_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mod_5_add_1540_2_lut (.I0(bit_ctr[13]), .I1(bit_ctr[13]), .I2(n37630), 
            .I3(VCC_net), .O(n2309)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_2_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_2009_15 (.CI(n28507), .I0(n2897), .I1(n2918), .CO(n28508));
    SB_LUT4 mod_5_add_2009_14_lut (.I0(n2898), .I1(n2898), .I2(n2918), 
            .I3(n28506), .O(n2997)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_14_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1540_2 (.CI(VCC_net), .I0(bit_ctr[13]), .I1(n37630), 
            .CO(n28736));
    SB_LUT4 mod_5_add_1607_21_lut (.I0(n2291), .I1(n2291), .I2(n2324), 
            .I3(n28735), .O(n2390)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_21_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2009_14 (.CI(n28506), .I0(n2898), .I1(n2918), .CO(n28507));
    SB_LUT4 mod_5_add_2009_13_lut (.I0(n2899), .I1(n2899), .I2(n2918), 
            .I3(n28505), .O(n2998)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_13_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2009_13 (.CI(n28505), .I0(n2899), .I1(n2918), .CO(n28506));
    SB_LUT4 mod_5_add_1607_20_lut (.I0(n2292), .I1(n2292), .I2(n2324), 
            .I3(n28734), .O(n2391)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_20_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_2009_12_lut (.I0(n2900), .I1(n2900), .I2(n2918), 
            .I3(n28504), .O(n2999)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_12_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1607_20 (.CI(n28734), .I0(n2292), .I1(n2324), .CO(n28735));
    SB_LUT4 add_21_14_lut (.I0(GND_net), .I1(bit_ctr[12]), .I2(GND_net), 
            .I3(n27775), .O(n255[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_2009_12 (.CI(n28504), .I0(n2900), .I1(n2918), .CO(n28505));
    SB_LUT4 mod_5_add_2009_11_lut (.I0(n2901), .I1(n2901), .I2(n2918), 
            .I3(n28503), .O(n3000)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_11_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1607_19_lut (.I0(n2293), .I1(n2293), .I2(n2324), 
            .I3(n28733), .O(n2392)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_19_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2009_11 (.CI(n28503), .I0(n2901), .I1(n2918), .CO(n28504));
    SB_CARRY mod_5_add_1607_19 (.CI(n28733), .I0(n2293), .I1(n2324), .CO(n28734));
    SB_LUT4 mod_5_add_2009_10_lut (.I0(n2902), .I1(n2902), .I2(n2918), 
            .I3(n28502), .O(n3001)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_10_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2009_10 (.CI(n28502), .I0(n2902), .I1(n2918), .CO(n28503));
    SB_LUT4 mod_5_add_1607_18_lut (.I0(n2294), .I1(n2294), .I2(n2324), 
            .I3(n28732), .O(n2393)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_18_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_2009_9_lut (.I0(n2903), .I1(n2903), .I2(n2918), 
            .I3(n28501), .O(n3002)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_9_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2009_9 (.CI(n28501), .I0(n2903), .I1(n2918), .CO(n28502));
    SB_CARRY mod_5_add_1607_18 (.CI(n28732), .I0(n2294), .I1(n2324), .CO(n28733));
    SB_LUT4 mod_5_add_2009_8_lut (.I0(n2904), .I1(n2904), .I2(n2918), 
            .I3(n28500), .O(n3003)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_8_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1607_17_lut (.I0(n2295), .I1(n2295), .I2(n2324), 
            .I3(n28731), .O(n2394)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_17_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY add_21_14 (.CI(n27775), .I0(bit_ctr[12]), .I1(GND_net), .CO(n27776));
    SB_CARRY mod_5_add_1607_17 (.CI(n28731), .I0(n2295), .I1(n2324), .CO(n28732));
    SB_LUT4 add_21_13_lut (.I0(GND_net), .I1(bit_ctr[11]), .I2(GND_net), 
            .I3(n27774), .O(n255[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_1607_16_lut (.I0(n2296), .I1(n2296), .I2(n2324), 
            .I3(n28730), .O(n2395)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_16_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1607_16 (.CI(n28730), .I0(n2296), .I1(n2324), .CO(n28731));
    SB_CARRY mod_5_add_2009_8 (.CI(n28500), .I0(n2904), .I1(n2918), .CO(n28501));
    SB_LUT4 mod_5_add_2009_7_lut (.I0(n2905), .I1(n2905), .I2(n2918), 
            .I3(n28499), .O(n3004)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_7_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1607_15_lut (.I0(n2297), .I1(n2297), .I2(n2324), 
            .I3(n28729), .O(n2396)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_15_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2009_7 (.CI(n28499), .I0(n2905), .I1(n2918), .CO(n28500));
    SB_LUT4 mod_5_add_2009_6_lut (.I0(n2906), .I1(n2906), .I2(n2918), 
            .I3(n28498), .O(n3005)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_6_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2009_6 (.CI(n28498), .I0(n2906), .I1(n2918), .CO(n28499));
    SB_LUT4 mod_5_add_2009_5_lut (.I0(n2907), .I1(n2907), .I2(n2918), 
            .I3(n28497), .O(n3006)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_5_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1607_15 (.CI(n28729), .I0(n2297), .I1(n2324), .CO(n28730));
    SB_LUT4 mod_5_add_1607_14_lut (.I0(n2298), .I1(n2298), .I2(n2324), 
            .I3(n28728), .O(n2397)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_14_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2009_5 (.CI(n28497), .I0(n2907), .I1(n2918), .CO(n28498));
    SB_LUT4 mod_5_add_2009_4_lut (.I0(n2908), .I1(n2908), .I2(n2918), 
            .I3(n28496), .O(n3007)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_4_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2009_4 (.CI(n28496), .I0(n2908), .I1(n2918), .CO(n28497));
    SB_LUT4 mod_5_add_2009_3_lut (.I0(n2909), .I1(n2909), .I2(n37632), 
            .I3(n28495), .O(n3008)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_3_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_2009_3 (.CI(n28495), .I0(n2909), .I1(n37632), .CO(n28496));
    SB_LUT4 i19470_2_lut (.I0(\neo_pixel_transmitter.done ), .I1(start), 
            .I2(GND_net), .I3(GND_net), .O(n24613));
    defparam i19470_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 mod_5_add_2009_2_lut (.I0(bit_ctr[6]), .I1(bit_ctr[6]), .I2(n37632), 
            .I3(VCC_net), .O(n3009)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_2_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1607_14 (.CI(n28728), .I0(n2298), .I1(n2324), .CO(n28729));
    SB_CARRY mod_5_add_2009_2 (.CI(VCC_net), .I0(bit_ctr[6]), .I1(n37632), 
            .CO(n28495));
    SB_LUT4 timer_1579_add_4_33_lut (.I0(GND_net), .I1(GND_net), .I2(timer[31]), 
            .I3(n28494), .O(n133[31])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1579_add_4_33_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 timer_1579_add_4_32_lut (.I0(GND_net), .I1(GND_net), .I2(timer[30]), 
            .I3(n28493), .O(n133[30])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1579_add_4_32_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1579_add_4_32 (.CI(n28493), .I0(GND_net), .I1(timer[30]), 
            .CO(n28494));
    SB_CARRY add_21_13 (.CI(n27774), .I0(bit_ctr[11]), .I1(GND_net), .CO(n27775));
    SB_LUT4 timer_1579_add_4_31_lut (.I0(GND_net), .I1(GND_net), .I2(timer[29]), 
            .I3(n28492), .O(n133[29])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1579_add_4_31_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1579_add_4_31 (.CI(n28492), .I0(GND_net), .I1(timer[29]), 
            .CO(n28493));
    SB_LUT4 timer_1579_add_4_30_lut (.I0(GND_net), .I1(GND_net), .I2(timer[28]), 
            .I3(n28491), .O(n133[28])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1579_add_4_30_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1579_add_4_30 (.CI(n28491), .I0(GND_net), .I1(timer[28]), 
            .CO(n28492));
    SB_LUT4 timer_1579_add_4_29_lut (.I0(GND_net), .I1(GND_net), .I2(timer[27]), 
            .I3(n28490), .O(n133[27])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1579_add_4_29_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1579_add_4_29 (.CI(n28490), .I0(GND_net), .I1(timer[27]), 
            .CO(n28491));
    SB_LUT4 timer_1579_add_4_28_lut (.I0(GND_net), .I1(GND_net), .I2(timer[26]), 
            .I3(n28489), .O(n133[26])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1579_add_4_28_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1579_add_4_28 (.CI(n28489), .I0(GND_net), .I1(timer[26]), 
            .CO(n28490));
    SB_LUT4 i1_2_lut_3_lut (.I0(n14), .I1(start), .I2(\neo_pixel_transmitter.done ), 
            .I3(GND_net), .O(n33365));
    defparam i1_2_lut_3_lut.LUT_INIT = 16'h2020;
    SB_LUT4 i29557_2_lut_3_lut (.I0(n24759), .I1(\neo_pixel_transmitter.done ), 
            .I2(\state[0] ), .I3(GND_net), .O(n36222));   // verilog/neopixel.v(35[12] 117[6])
    defparam i29557_2_lut_3_lut.LUT_INIT = 16'hfdfd;
    SB_LUT4 i30869_1_lut (.I0(n1928), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n37622));
    defparam i30869_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i7_3_lut_adj_1552 (.I0(bit_ctr[11]), .I1(n2403), .I2(n2409), 
            .I3(GND_net), .O(n27_adj_4781));
    defparam i7_3_lut_adj_1552.LUT_INIT = 16'hecec;
    SB_LUT4 i13_4_lut_adj_1553 (.I0(n2390), .I1(n2391), .I2(n2397), .I3(n2394), 
            .O(n33));
    defparam i13_4_lut_adj_1553.LUT_INIT = 16'hfffe;
    SB_LUT4 i12_4_lut_adj_1554 (.I0(n2392), .I1(n2405), .I2(n2400), .I3(n2398), 
            .O(n32));
    defparam i12_4_lut_adj_1554.LUT_INIT = 16'hfffe;
    SB_LUT4 i11_4_lut_adj_1555 (.I0(n2396), .I1(n2402), .I2(n2408), .I3(n2399), 
            .O(n31));
    defparam i11_4_lut_adj_1555.LUT_INIT = 16'hfffe;
    SB_LUT4 i15_4_lut_adj_1556 (.I0(n2393), .I1(n2406), .I2(n2395), .I3(n2407), 
            .O(n35_adj_4782));
    defparam i15_4_lut_adj_1556.LUT_INIT = 16'hfffe;
    SB_LUT4 i17_4_lut_adj_1557 (.I0(n33), .I1(n27_adj_4781), .I2(n2404), 
            .I3(n2401), .O(n37_adj_4783));
    defparam i17_4_lut_adj_1557.LUT_INIT = 16'hfffe;
    SB_LUT4 i19_4_lut_adj_1558 (.I0(n37_adj_4783), .I1(n35_adj_4782), .I2(n31), 
            .I3(n32), .O(n2423));
    defparam i19_4_lut_adj_1558.LUT_INIT = 16'hfffe;
    SB_LUT4 i19616_2_lut_4_lut (.I0(one_wire_N_553[9]), .I1(one_wire_N_553[11]), 
            .I2(one_wire_N_553[10]), .I3(n17526), .O(n24759));
    defparam i19616_2_lut_4_lut.LUT_INIT = 16'hffc8;
    SB_LUT4 mod_5_add_1607_13_lut (.I0(n2299), .I1(n2299), .I2(n2324), 
            .I3(n28727), .O(n2398)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_13_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 timer_1579_add_4_27_lut (.I0(GND_net), .I1(GND_net), .I2(timer[25]), 
            .I3(n28488), .O(n133[25])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1579_add_4_27_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1607_13 (.CI(n28727), .I0(n2299), .I1(n2324), .CO(n28728));
    SB_LUT4 mod_5_add_1607_12_lut (.I0(n2300), .I1(n2300), .I2(n2324), 
            .I3(n28726), .O(n2399)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_12_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY timer_1579_add_4_27 (.CI(n28488), .I0(GND_net), .I1(timer[25]), 
            .CO(n28489));
    SB_CARRY mod_5_add_1607_12 (.CI(n28726), .I0(n2300), .I1(n2324), .CO(n28727));
    SB_LUT4 mod_5_add_1607_11_lut (.I0(n2301), .I1(n2301), .I2(n2324), 
            .I3(n28725), .O(n2400)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_11_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 timer_1579_add_4_26_lut (.I0(GND_net), .I1(GND_net), .I2(timer[24]), 
            .I3(n28487), .O(n133[24])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1579_add_4_26_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1579_add_4_26 (.CI(n28487), .I0(GND_net), .I1(timer[24]), 
            .CO(n28488));
    SB_LUT4 timer_1579_add_4_25_lut (.I0(GND_net), .I1(GND_net), .I2(timer[23]), 
            .I3(n28486), .O(n133[23])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1579_add_4_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_21_12_lut (.I0(GND_net), .I1(bit_ctr[10]), .I2(GND_net), 
            .I3(n27773), .O(n255[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1579_add_4_25 (.CI(n28486), .I0(GND_net), .I1(timer[23]), 
            .CO(n28487));
    SB_LUT4 i2_3_lut_4_lut (.I0(n14), .I1(start), .I2(\neo_pixel_transmitter.done ), 
            .I3(\state[1] ), .O(n35064));
    defparam i2_3_lut_4_lut.LUT_INIT = 16'hffdf;
    SB_LUT4 timer_1579_add_4_24_lut (.I0(GND_net), .I1(GND_net), .I2(timer[22]), 
            .I3(n28485), .O(n133[22])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1579_add_4_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1579_add_4_24 (.CI(n28485), .I0(GND_net), .I1(timer[22]), 
            .CO(n28486));
    SB_LUT4 timer_1579_add_4_23_lut (.I0(GND_net), .I1(GND_net), .I2(timer[21]), 
            .I3(n28484), .O(n133[21])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1579_add_4_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1579_add_4_23 (.CI(n28484), .I0(GND_net), .I1(timer[21]), 
            .CO(n28485));
    SB_LUT4 sub_14_add_2_33_lut (.I0(one_wire_N_553[25]), .I1(timer[31]), 
            .I2(n1[31]), .I3(n27975), .O(n22_adj_4784)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_33_lut.LUT_INIT = 16'hebbe;
    SB_LUT4 timer_1579_add_4_22_lut (.I0(GND_net), .I1(GND_net), .I2(timer[20]), 
            .I3(n28483), .O(n133[20])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1579_add_4_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1579_add_4_22 (.CI(n28483), .I0(GND_net), .I1(timer[20]), 
            .CO(n28484));
    SB_LUT4 timer_1579_add_4_21_lut (.I0(GND_net), .I1(GND_net), .I2(timer[19]), 
            .I3(n28482), .O(n133[19])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1579_add_4_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1579_add_4_21 (.CI(n28482), .I0(GND_net), .I1(timer[19]), 
            .CO(n28483));
    SB_LUT4 timer_1579_add_4_20_lut (.I0(GND_net), .I1(GND_net), .I2(timer[18]), 
            .I3(n28481), .O(n133[18])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1579_add_4_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1579_add_4_20 (.CI(n28481), .I0(GND_net), .I1(timer[18]), 
            .CO(n28482));
    SB_LUT4 timer_1579_add_4_19_lut (.I0(GND_net), .I1(GND_net), .I2(timer[17]), 
            .I3(n28480), .O(n133[17])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1579_add_4_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1579_add_4_19 (.CI(n28480), .I0(GND_net), .I1(timer[17]), 
            .CO(n28481));
    SB_CARRY mod_5_add_1607_11 (.CI(n28725), .I0(n2301), .I1(n2324), .CO(n28726));
    SB_LUT4 timer_1579_add_4_18_lut (.I0(GND_net), .I1(GND_net), .I2(timer[16]), 
            .I3(n28479), .O(n133[16])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1579_add_4_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1579_add_4_18 (.CI(n28479), .I0(GND_net), .I1(timer[16]), 
            .CO(n28480));
    SB_LUT4 timer_1579_add_4_17_lut (.I0(GND_net), .I1(GND_net), .I2(timer[15]), 
            .I3(n28478), .O(n133[15])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1579_add_4_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i19_4_lut_adj_1559 (.I0(bit_ctr[26]), .I1(bit_ctr[16]), .I2(bit_ctr[20]), 
            .I3(bit_ctr[7]), .O(n46_adj_4785));
    defparam i19_4_lut_adj_1559.LUT_INIT = 16'hfffe;
    SB_LUT4 i17_4_lut_adj_1560 (.I0(bit_ctr[14]), .I1(bit_ctr[9]), .I2(bit_ctr[23]), 
            .I3(bit_ctr[10]), .O(n44_adj_4786));
    defparam i17_4_lut_adj_1560.LUT_INIT = 16'hfffe;
    SB_LUT4 i18_4_lut_adj_1561 (.I0(bit_ctr[27]), .I1(bit_ctr[12]), .I2(bit_ctr[15]), 
            .I3(bit_ctr[29]), .O(n45_adj_4787));
    defparam i18_4_lut_adj_1561.LUT_INIT = 16'hfffe;
    SB_LUT4 i16_4_lut_adj_1562 (.I0(bit_ctr[6]), .I1(bit_ctr[31]), .I2(bit_ctr[19]), 
            .I3(bit_ctr[21]), .O(n43_adj_4788));
    defparam i16_4_lut_adj_1562.LUT_INIT = 16'hfffe;
    SB_LUT4 i15_4_lut_adj_1563 (.I0(bit_ctr[17]), .I1(bit_ctr[28]), .I2(bit_ctr[11]), 
            .I3(bit_ctr[5]), .O(n42_adj_4789));
    defparam i15_4_lut_adj_1563.LUT_INIT = 16'hfffe;
    SB_LUT4 i13_2_lut (.I0(bit_ctr[18]), .I1(bit_ctr[8]), .I2(GND_net), 
            .I3(GND_net), .O(n40_adj_4790));
    defparam i13_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i21_4_lut_adj_1564 (.I0(bit_ctr[24]), .I1(n42_adj_4789), .I2(bit_ctr[13]), 
            .I3(bit_ctr[22]), .O(n48_adj_4791));
    defparam i21_4_lut_adj_1564.LUT_INIT = 16'hfffe;
    SB_LUT4 i25_4_lut_adj_1565 (.I0(n43_adj_4788), .I1(n45_adj_4787), .I2(n44_adj_4786), 
            .I3(n46_adj_4785), .O(n52_adj_4792));
    defparam i25_4_lut_adj_1565.LUT_INIT = 16'hfffe;
    SB_LUT4 i24_4_lut (.I0(bit_ctr[30]), .I1(n48_adj_4791), .I2(n40_adj_4790), 
            .I3(bit_ctr[25]), .O(n51));
    defparam i24_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut (.I0(bit_ctr[3]), .I1(n51), .I2(bit_ctr[4]), .I3(n52_adj_4792), 
            .O(\state_3__N_402[1] ));
    defparam i1_4_lut.LUT_INIT = 16'hffec;
    SB_CARRY timer_1579_add_4_17 (.CI(n28478), .I0(GND_net), .I1(timer[15]), 
            .CO(n28479));
    SB_LUT4 i2_3_lut (.I0(one_wire_N_553[3]), .I1(one_wire_N_553[4]), .I2(one_wire_N_553[2]), 
            .I3(GND_net), .O(n29522));
    defparam i2_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 i26764_2_lut (.I0(one_wire_N_553[4]), .I1(n24675), .I2(GND_net), 
            .I3(GND_net), .O(n33371));
    defparam i26764_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i6_4_lut_adj_1566 (.I0(one_wire_N_553[5]), .I1(one_wire_N_553[11]), 
            .I2(one_wire_N_553[7]), .I3(n17526), .O(n14_adj_4793));   // verilog/neopixel.v(104[14:39])
    defparam i6_4_lut_adj_1566.LUT_INIT = 16'hfffe;
    SB_LUT4 timer_1579_add_4_16_lut (.I0(GND_net), .I1(GND_net), .I2(timer[14]), 
            .I3(n28477), .O(n133[14])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1579_add_4_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1579_add_4_16 (.CI(n28477), .I0(GND_net), .I1(timer[14]), 
            .CO(n28478));
    SB_LUT4 timer_1579_add_4_15_lut (.I0(GND_net), .I1(GND_net), .I2(timer[13]), 
            .I3(n28476), .O(n133[13])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1579_add_4_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1579_add_4_15 (.CI(n28476), .I0(GND_net), .I1(timer[13]), 
            .CO(n28477));
    SB_LUT4 timer_1579_add_4_14_lut (.I0(GND_net), .I1(GND_net), .I2(timer[12]), 
            .I3(n28475), .O(n133[12])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1579_add_4_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1579_add_4_14 (.CI(n28475), .I0(GND_net), .I1(timer[12]), 
            .CO(n28476));
    SB_LUT4 mod_5_add_1607_10_lut (.I0(n2302), .I1(n2302), .I2(n2324), 
            .I3(n28724), .O(n2401)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_10_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 sub_14_add_2_32_lut (.I0(one_wire_N_553[24]), .I1(timer[30]), 
            .I2(n1[30]), .I3(n27974), .O(n23_adj_4794)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_32_lut.LUT_INIT = 16'hebbe;
    SB_LUT4 timer_1579_add_4_13_lut (.I0(GND_net), .I1(GND_net), .I2(timer[11]), 
            .I3(n28474), .O(n133[11])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1579_add_4_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1579_add_4_13 (.CI(n28474), .I0(GND_net), .I1(timer[11]), 
            .CO(n28475));
    SB_LUT4 timer_1579_add_4_12_lut (.I0(GND_net), .I1(GND_net), .I2(timer[10]), 
            .I3(n28473), .O(n133[10])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1579_add_4_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1607_10 (.CI(n28724), .I0(n2302), .I1(n2324), .CO(n28725));
    SB_CARRY timer_1579_add_4_12 (.CI(n28473), .I0(GND_net), .I1(timer[10]), 
            .CO(n28474));
    SB_LUT4 timer_1579_add_4_11_lut (.I0(GND_net), .I1(GND_net), .I2(timer[9]), 
            .I3(n28472), .O(n133[9])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1579_add_4_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1579_add_4_11 (.CI(n28472), .I0(GND_net), .I1(timer[9]), 
            .CO(n28473));
    SB_LUT4 timer_1579_add_4_10_lut (.I0(GND_net), .I1(GND_net), .I2(timer[8]), 
            .I3(n28471), .O(n133[8])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1579_add_4_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i7_4_lut_adj_1567 (.I0(one_wire_N_553[9]), .I1(n14_adj_4793), 
            .I2(n10_adj_4795), .I3(one_wire_N_553[6]), .O(n17393));   // verilog/neopixel.v(104[14:39])
    defparam i7_4_lut_adj_1567.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_adj_1568 (.I0(start), .I1(\neo_pixel_transmitter.done ), 
            .I2(GND_net), .I3(GND_net), .O(n17509));   // verilog/neopixel.v(79[18] 99[12])
    defparam i1_2_lut_adj_1568.LUT_INIT = 16'hbbbb;
    SB_LUT4 i270_2_lut (.I0(LED_c), .I1(\state_3__N_402[1] ), .I2(GND_net), 
            .I3(GND_net), .O(n1251));   // verilog/neopixel.v(40[18] 45[12])
    defparam i270_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i3439_4_lut (.I0(n24735), .I1(n1251), .I2(\state[1] ), .I3(n17509), 
            .O(n5449));
    defparam i3439_4_lut.LUT_INIT = 16'h3f35;
    SB_CARRY timer_1579_add_4_10 (.CI(n28471), .I0(GND_net), .I1(timer[8]), 
            .CO(n28472));
    SB_LUT4 i30865_4_lut (.I0(\state[1] ), .I1(n36280), .I2(\state[0] ), 
            .I3(n5449), .O(n18566));
    defparam i30865_4_lut.LUT_INIT = 16'h01f1;
    SB_LUT4 timer_1579_add_4_9_lut (.I0(GND_net), .I1(GND_net), .I2(timer[7]), 
            .I3(n28470), .O(n133[7])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1579_add_4_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i23_3_lut_4_lut (.I0(one_wire_N_553[4]), .I1(n24675), .I2(n29522), 
            .I3(\state[0] ), .O(n33377));
    defparam i23_3_lut_4_lut.LUT_INIT = 16'hf0ee;
    SB_LUT4 mod_5_add_1607_9_lut (.I0(n2303), .I1(n2303), .I2(n2324), 
            .I3(n28723), .O(n2402)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_9_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY timer_1579_add_4_9 (.CI(n28470), .I0(GND_net), .I1(timer[7]), 
            .CO(n28471));
    SB_LUT4 timer_1579_add_4_8_lut (.I0(GND_net), .I1(GND_net), .I2(timer[6]), 
            .I3(n28469), .O(n133[6])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1579_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1579_add_4_8 (.CI(n28469), .I0(GND_net), .I1(timer[6]), 
            .CO(n28470));
    SB_LUT4 timer_1579_add_4_7_lut (.I0(GND_net), .I1(GND_net), .I2(timer[5]), 
            .I3(n28468), .O(n133[5])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1579_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1579_add_4_7 (.CI(n28468), .I0(GND_net), .I1(timer[5]), 
            .CO(n28469));
    SB_CARRY mod_5_add_1607_9 (.CI(n28723), .I0(n2303), .I1(n2324), .CO(n28724));
    SB_LUT4 timer_1579_add_4_6_lut (.I0(GND_net), .I1(GND_net), .I2(timer[4]), 
            .I3(n28467), .O(n133[4])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1579_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1579_add_4_6 (.CI(n28467), .I0(GND_net), .I1(timer[4]), 
            .CO(n28468));
    SB_LUT4 timer_1579_add_4_5_lut (.I0(GND_net), .I1(GND_net), .I2(timer[3]), 
            .I3(n28466), .O(n133[3])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1579_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_14_add_2_32 (.CI(n27974), .I0(timer[30]), .I1(n1[30]), 
            .CO(n27975));
    SB_CARRY timer_1579_add_4_5 (.CI(n28466), .I0(GND_net), .I1(timer[3]), 
            .CO(n28467));
    SB_LUT4 timer_1579_add_4_4_lut (.I0(GND_net), .I1(GND_net), .I2(timer[2]), 
            .I3(n28465), .O(n133[2])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1579_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_1607_8_lut (.I0(n2304), .I1(n2304), .I2(n2324), 
            .I3(n28722), .O(n2403)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_8_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1607_8 (.CI(n28722), .I0(n2304), .I1(n2324), .CO(n28723));
    SB_CARRY timer_1579_add_4_4 (.CI(n28465), .I0(GND_net), .I1(timer[2]), 
            .CO(n28466));
    SB_LUT4 timer_1579_add_4_3_lut (.I0(GND_net), .I1(GND_net), .I2(timer[1]), 
            .I3(n28464), .O(n133[1])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1579_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1579_add_4_3 (.CI(n28464), .I0(GND_net), .I1(timer[1]), 
            .CO(n28465));
    SB_LUT4 timer_1579_add_4_2_lut (.I0(GND_net), .I1(GND_net), .I2(timer[0]), 
            .I3(VCC_net), .O(n133[0])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1579_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1579_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(timer[0]), 
            .CO(n28464));
    SB_LUT4 mod_5_add_2076_28_lut (.I0(n2984), .I1(n2984), .I2(n3017), 
            .I3(n28463), .O(n3083)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_28_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_2076_27_lut (.I0(n2985), .I1(n2985), .I2(n3017), 
            .I3(n28462), .O(n3084)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_27_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2076_27 (.CI(n28462), .I0(n2985), .I1(n3017), .CO(n28463));
    SB_LUT4 mod_5_add_2076_26_lut (.I0(n2986), .I1(n2986), .I2(n3017), 
            .I3(n28461), .O(n3085)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_26_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2076_26 (.CI(n28461), .I0(n2986), .I1(n3017), .CO(n28462));
    SB_LUT4 mod_5_add_2076_25_lut (.I0(n2987), .I1(n2987), .I2(n3017), 
            .I3(n28460), .O(n3086)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_25_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2076_25 (.CI(n28460), .I0(n2987), .I1(n3017), .CO(n28461));
    SB_LUT4 sub_14_add_2_31_lut (.I0(one_wire_N_553[19]), .I1(timer[29]), 
            .I2(n1[29]), .I3(n27973), .O(n28_adj_4796)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_31_lut.LUT_INIT = 16'hebbe;
    SB_LUT4 mod_5_add_2076_24_lut (.I0(n2988), .I1(n2988), .I2(n3017), 
            .I3(n28459), .O(n3087)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_24_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1607_7_lut (.I0(n2305), .I1(n2305), .I2(n2324), 
            .I3(n28721), .O(n2404)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_7_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2076_24 (.CI(n28459), .I0(n2988), .I1(n3017), .CO(n28460));
    SB_LUT4 mod_5_add_2076_23_lut (.I0(n2989), .I1(n2989), .I2(n3017), 
            .I3(n28458), .O(n3088)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_23_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1607_7 (.CI(n28721), .I0(n2305), .I1(n2324), .CO(n28722));
    SB_CARRY add_21_12 (.CI(n27773), .I0(bit_ctr[10]), .I1(GND_net), .CO(n27774));
    SB_LUT4 mod_5_add_1607_6_lut (.I0(n2306), .I1(n2306), .I2(n2324), 
            .I3(n28720), .O(n2405)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_6_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1607_6 (.CI(n28720), .I0(n2306), .I1(n2324), .CO(n28721));
    SB_CARRY mod_5_add_2076_23 (.CI(n28458), .I0(n2989), .I1(n3017), .CO(n28459));
    SB_CARRY sub_14_add_2_31 (.CI(n27973), .I0(timer[29]), .I1(n1[29]), 
            .CO(n27974));
    SB_LUT4 mod_5_add_2076_22_lut (.I0(n2990), .I1(n2990), .I2(n3017), 
            .I3(n28457), .O(n3089)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_22_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2076_22 (.CI(n28457), .I0(n2990), .I1(n3017), .CO(n28458));
    SB_LUT4 mod_5_add_2076_21_lut (.I0(n2991), .I1(n2991), .I2(n3017), 
            .I3(n28456), .O(n3090)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_21_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1607_5_lut (.I0(n2307), .I1(n2307), .I2(n2324), 
            .I3(n28719), .O(n2406)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_5_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1607_5 (.CI(n28719), .I0(n2307), .I1(n2324), .CO(n28720));
    SB_CARRY mod_5_add_2076_21 (.CI(n28456), .I0(n2991), .I1(n3017), .CO(n28457));
    SB_LUT4 mod_5_add_2076_20_lut (.I0(n2992), .I1(n2992), .I2(n3017), 
            .I3(n28455), .O(n3091)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_20_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2076_20 (.CI(n28455), .I0(n2992), .I1(n3017), .CO(n28456));
    SB_LUT4 mod_5_add_2076_19_lut (.I0(n2993), .I1(n2993), .I2(n3017), 
            .I3(n28454), .O(n3092)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_19_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 sub_14_add_2_30_lut (.I0(one_wire_N_553[26]), .I1(timer[28]), 
            .I2(n1[28]), .I3(n27972), .O(n26_adj_4797)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_30_lut.LUT_INIT = 16'hebbe;
    SB_CARRY mod_5_add_2076_19 (.CI(n28454), .I0(n2993), .I1(n3017), .CO(n28455));
    SB_LUT4 mod_5_add_2076_18_lut (.I0(n2994), .I1(n2994), .I2(n3017), 
            .I3(n28453), .O(n3093)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_18_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2076_18 (.CI(n28453), .I0(n2994), .I1(n3017), .CO(n28454));
    SB_LUT4 mod_5_add_2076_17_lut (.I0(n2995), .I1(n2995), .I2(n3017), 
            .I3(n28452), .O(n3094)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_17_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2076_17 (.CI(n28452), .I0(n2995), .I1(n3017), .CO(n28453));
    SB_LUT4 mod_5_add_2076_16_lut (.I0(n2996), .I1(n2996), .I2(n3017), 
            .I3(n28451), .O(n3095)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_16_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2076_16 (.CI(n28451), .I0(n2996), .I1(n3017), .CO(n28452));
    SB_LUT4 mod_5_add_2076_15_lut (.I0(n2997), .I1(n2997), .I2(n3017), 
            .I3(n28450), .O(n3096)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_15_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY sub_14_add_2_30 (.CI(n27972), .I0(timer[28]), .I1(n1[28]), 
            .CO(n27973));
    SB_CARRY mod_5_add_2076_15 (.CI(n28450), .I0(n2997), .I1(n3017), .CO(n28451));
    SB_LUT4 mod_5_add_2076_14_lut (.I0(n2998), .I1(n2998), .I2(n3017), 
            .I3(n28449), .O(n3097)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_14_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i1_2_lut_3_lut_4_lut (.I0(n8799), .I1(bit_ctr[30]), .I2(bit_ctr[31]), 
            .I3(bit_ctr[29]), .O(n29995));   // verilog/neopixel.v(22[26:36])
    defparam i1_2_lut_3_lut_4_lut.LUT_INIT = 16'h45ba;
    SB_LUT4 i1_2_lut_adj_1569 (.I0(\state[0] ), .I1(\neo_pixel_transmitter.done ), 
            .I2(GND_net), .I3(GND_net), .O(n78));
    defparam i1_2_lut_adj_1569.LUT_INIT = 16'h2222;
    SB_CARRY mod_5_add_2076_14 (.CI(n28449), .I0(n2998), .I1(n3017), .CO(n28450));
    SB_LUT4 mod_5_add_2076_13_lut (.I0(n2999), .I1(n2999), .I2(n3017), 
            .I3(n28448), .O(n3098)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_13_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2076_13 (.CI(n28448), .I0(n2999), .I1(n3017), .CO(n28449));
    SB_LUT4 mod_5_add_2076_12_lut (.I0(n3000), .I1(n3000), .I2(n3017), 
            .I3(n28447), .O(n3099)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_12_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2076_12 (.CI(n28447), .I0(n3000), .I1(n3017), .CO(n28448));
    SB_LUT4 mod_5_add_2076_11_lut (.I0(n3001), .I1(n3001), .I2(n3017), 
            .I3(n28446), .O(n3100)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_11_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 add_21_11_lut (.I0(GND_net), .I1(bit_ctr[9]), .I2(GND_net), 
            .I3(n27772), .O(n255[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_2076_11 (.CI(n28446), .I0(n3001), .I1(n3017), .CO(n28447));
    SB_LUT4 mod_5_add_2076_10_lut (.I0(n3002), .I1(n3002), .I2(n3017), 
            .I3(n28445), .O(n3101)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_10_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2076_10 (.CI(n28445), .I0(n3002), .I1(n3017), .CO(n28446));
    SB_LUT4 mod_5_add_2076_9_lut (.I0(n3003), .I1(n3003), .I2(n3017), 
            .I3(n28444), .O(n3102)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_9_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2076_9 (.CI(n28444), .I0(n3003), .I1(n3017), .CO(n28445));
    SB_LUT4 mod_5_add_2076_8_lut (.I0(n3004), .I1(n3004), .I2(n3017), 
            .I3(n28443), .O(n3103)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_8_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2076_8 (.CI(n28443), .I0(n3004), .I1(n3017), .CO(n28444));
    SB_LUT4 mod_5_add_2076_7_lut (.I0(n3005), .I1(n3005), .I2(n3017), 
            .I3(n28442), .O(n3104)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_7_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2076_7 (.CI(n28442), .I0(n3005), .I1(n3017), .CO(n28443));
    SB_LUT4 mod_5_add_2076_6_lut (.I0(n3006), .I1(n3006), .I2(n3017), 
            .I3(n28441), .O(n3105)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_6_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2076_6 (.CI(n28441), .I0(n3006), .I1(n3017), .CO(n28442));
    SB_LUT4 mod_5_add_2076_5_lut (.I0(n3007), .I1(n3007), .I2(n3017), 
            .I3(n28440), .O(n3106)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_5_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1607_4_lut (.I0(n2308), .I1(n2308), .I2(n2324), 
            .I3(n28718), .O(n2407)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_4_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1607_4 (.CI(n28718), .I0(n2308), .I1(n2324), .CO(n28719));
    SB_LUT4 sub_14_add_2_29_lut (.I0(one_wire_N_553[18]), .I1(timer[27]), 
            .I2(n1[27]), .I3(n27971), .O(n21_adj_4798)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_29_lut.LUT_INIT = 16'hebbe;
    SB_CARRY mod_5_add_2076_5 (.CI(n28440), .I0(n3007), .I1(n3017), .CO(n28441));
    SB_LUT4 mod_5_add_1607_3_lut (.I0(n2309), .I1(n2309), .I2(n37634), 
            .I3(n28717), .O(n2408)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_3_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY sub_14_add_2_29 (.CI(n27971), .I0(timer[27]), .I1(n1[27]), 
            .CO(n27972));
    SB_LUT4 mod_5_add_2076_4_lut (.I0(n3008), .I1(n3008), .I2(n3017), 
            .I3(n28439), .O(n3107)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_4_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2076_4 (.CI(n28439), .I0(n3008), .I1(n3017), .CO(n28440));
    SB_LUT4 mod_5_add_2076_3_lut (.I0(n3009), .I1(n3009), .I2(n37635), 
            .I3(n28438), .O(n3108)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_3_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1607_3 (.CI(n28717), .I0(n2309), .I1(n37634), .CO(n28718));
    SB_LUT4 mod_5_add_1607_2_lut (.I0(bit_ctr[12]), .I1(bit_ctr[12]), .I2(n37634), 
            .I3(VCC_net), .O(n2409)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_2_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1607_2 (.CI(VCC_net), .I0(bit_ctr[12]), .I1(n37634), 
            .CO(n28717));
    SB_LUT4 sub_14_add_2_28_lut (.I0(GND_net), .I1(timer[26]), .I2(n1[26]), 
            .I3(n27970), .O(one_wire_N_553[26])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_28_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_2076_3 (.CI(n28438), .I0(n3009), .I1(n37635), .CO(n28439));
    SB_LUT4 i26703_2_lut (.I0(one_wire_N_553[3]), .I1(one_wire_N_553[2]), 
            .I2(GND_net), .I3(GND_net), .O(n33451));
    defparam i26703_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i19532_2_lut (.I0(n29671), .I1(one_wire_N_553[3]), .I2(GND_net), 
            .I3(GND_net), .O(n24675));
    defparam i19532_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i16_4_lut_adj_1570 (.I0(n21_adj_4798), .I1(n23_adj_4794), .I2(n22_adj_4784), 
            .I3(n24_adj_4799), .O(n36_adj_4800));   // verilog/neopixel.v(104[14:39])
    defparam i16_4_lut_adj_1570.LUT_INIT = 16'hfffe;
    SB_LUT4 i17_4_lut_adj_1571 (.I0(n25_adj_4801), .I1(n27_adj_4802), .I2(n26_adj_4797), 
            .I3(n28_adj_4796), .O(n37_adj_4803));   // verilog/neopixel.v(104[14:39])
    defparam i17_4_lut_adj_1571.LUT_INIT = 16'hfffe;
    SB_LUT4 mod_5_add_2076_2_lut (.I0(bit_ctr[5]), .I1(bit_ctr[5]), .I2(n37635), 
            .I3(VCC_net), .O(n3109)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_2_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_2076_2 (.CI(VCC_net), .I0(bit_ctr[5]), .I1(n37635), 
            .CO(n28438));
    SB_LUT4 mod_5_add_2143_29_lut (.I0(n3083), .I1(n3083), .I2(n3116), 
            .I3(n28437), .O(n63)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_29_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_2143_28_lut (.I0(n3084), .I1(n3084), .I2(n3116), 
            .I3(n28436), .O(n61)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_28_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2143_28 (.CI(n28436), .I0(n3084), .I1(n3116), .CO(n28437));
    SB_LUT4 mod_5_add_2143_27_lut (.I0(n3085), .I1(n3085), .I2(n3116), 
            .I3(n28435), .O(n59)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_27_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2143_27 (.CI(n28435), .I0(n3085), .I1(n3116), .CO(n28436));
    SB_LUT4 mod_5_add_2143_26_lut (.I0(n3086), .I1(n3086), .I2(n3116), 
            .I3(n28434), .O(n57)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_26_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2143_26 (.CI(n28434), .I0(n3086), .I1(n3116), .CO(n28435));
    SB_LUT4 mod_5_i471_3_lut_3_lut_4_lut_4_lut (.I0(n8799), .I1(bit_ctr[30]), 
            .I2(bit_ctr[31]), .I3(bit_ctr[29]), .O(n708));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i471_3_lut_3_lut_4_lut_4_lut.LUT_INIT = 16'hb60c;
    SB_LUT4 mod_5_add_2143_25_lut (.I0(n3087), .I1(n3087), .I2(n3116), 
            .I3(n28433), .O(n55)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_25_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2143_25 (.CI(n28433), .I0(n3087), .I1(n3116), .CO(n28434));
    SB_LUT4 mod_5_add_2143_24_lut (.I0(n3088), .I1(n3088), .I2(n3116), 
            .I3(n28432), .O(n53)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_24_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2143_24 (.CI(n28432), .I0(n3088), .I1(n3116), .CO(n28433));
    SB_LUT4 mod_5_add_2143_23_lut (.I0(n3089), .I1(n3089), .I2(n3116), 
            .I3(n28431), .O(n51_adj_4804)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_23_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2143_23 (.CI(n28431), .I0(n3089), .I1(n3116), .CO(n28432));
    SB_LUT4 mod_5_add_2143_22_lut (.I0(n3090), .I1(n3090), .I2(n3116), 
            .I3(n28430), .O(n49_adj_4805)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_22_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY add_21_9 (.CI(n27770), .I0(bit_ctr[7]), .I1(GND_net), .CO(n27771));
    SB_CARRY mod_5_add_2143_22 (.CI(n28430), .I0(n3090), .I1(n3116), .CO(n28431));
    SB_LUT4 mod_5_add_2143_21_lut (.I0(n3091), .I1(n3091), .I2(n3116), 
            .I3(n28429), .O(n47_adj_4806)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_21_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2143_21 (.CI(n28429), .I0(n3091), .I1(n3116), .CO(n28430));
    SB_LUT4 mod_5_add_2143_20_lut (.I0(n3092), .I1(n3092), .I2(n3116), 
            .I3(n28428), .O(n45_adj_4807)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_20_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2143_20 (.CI(n28428), .I0(n3092), .I1(n3116), .CO(n28429));
    SB_LUT4 mod_5_add_2143_19_lut (.I0(n3093), .I1(n3093), .I2(n3116), 
            .I3(n28427), .O(n43_adj_4808)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_19_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2143_19 (.CI(n28427), .I0(n3093), .I1(n3116), .CO(n28428));
    SB_LUT4 i19_4_lut_adj_1572 (.I0(n37_adj_4803), .I1(n29_adj_4809), .I2(n36_adj_4800), 
            .I3(n30_adj_4810), .O(n17526));   // verilog/neopixel.v(104[14:39])
    defparam i19_4_lut_adj_1572.LUT_INIT = 16'hfffe;
    SB_LUT4 bit_ctr_0__bdd_4_lut (.I0(bit_ctr[0]), .I1(neopxl_color[18]), 
            .I2(neopxl_color[19]), .I3(bit_ctr[1]), .O(n37880));
    defparam bit_ctr_0__bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_LUT4 n37880_bdd_4_lut (.I0(n37880), .I1(neopxl_color[17]), .I2(neopxl_color[16]), 
            .I3(bit_ctr[1]), .O(n37883));
    defparam n37880_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_2_lut_adj_1573 (.I0(one_wire_N_553[9]), .I1(start), .I2(GND_net), 
            .I3(GND_net), .O(n10_adj_4811));
    defparam i1_2_lut_adj_1573.LUT_INIT = 16'heeee;
    SB_LUT4 i7_4_lut_adj_1574 (.I0(one_wire_N_553[11]), .I1(one_wire_N_553[5]), 
            .I2(one_wire_N_553[7]), .I3(n10_adj_4811), .O(n16_adj_4812));
    defparam i7_4_lut_adj_1574.LUT_INIT = 16'hfffe;
    SB_LUT4 i8_4_lut_adj_1575 (.I0(\state[1] ), .I1(n16_adj_4812), .I2(n10_adj_4795), 
            .I3(one_wire_N_553[6]), .O(n33545));
    defparam i8_4_lut_adj_1575.LUT_INIT = 16'hfffe;
    SB_LUT4 mod_5_add_2143_18_lut (.I0(n3094), .I1(n3094), .I2(n3116), 
            .I3(n28426), .O(n41)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_18_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2143_18 (.CI(n28426), .I0(n3094), .I1(n3116), .CO(n28427));
    SB_LUT4 i1_4_lut_adj_1576 (.I0(one_wire_N_553[4]), .I1(n32651), .I2(n24675), 
            .I3(n33451), .O(n116));
    defparam i1_4_lut_adj_1576.LUT_INIT = 16'h45cd;
    SB_LUT4 mod_5_add_2143_17_lut (.I0(n3095), .I1(n3095), .I2(n3116), 
            .I3(n28425), .O(n39_adj_4813)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_17_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2143_17 (.CI(n28425), .I0(n3095), .I1(n3116), .CO(n28426));
    SB_LUT4 i30388_3_lut (.I0(n33545), .I1(n116), .I2(n17526), .I3(GND_net), 
            .O(n35264));
    defparam i30388_3_lut.LUT_INIT = 16'hfbfb;
    SB_LUT4 mod_5_add_2143_16_lut (.I0(n3096), .I1(n3096), .I2(n3116), 
            .I3(n28424), .O(n37_adj_4814)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_16_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2143_16 (.CI(n28424), .I0(n3096), .I1(n3116), .CO(n28425));
    SB_LUT4 mod_5_add_2143_15_lut (.I0(n3097), .I1(n3097), .I2(n3116), 
            .I3(n28423), .O(n35_adj_4815)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_15_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2143_15 (.CI(n28423), .I0(n3097), .I1(n3116), .CO(n28424));
    SB_LUT4 mod_5_add_2143_14_lut (.I0(n3098), .I1(n3098), .I2(n3116), 
            .I3(n28422), .O(n33_adj_4816)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_14_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2143_14 (.CI(n28422), .I0(n3098), .I1(n3116), .CO(n28423));
    SB_LUT4 mod_5_add_2143_13_lut (.I0(n3099), .I1(n3099), .I2(n3116), 
            .I3(n28421), .O(n31_adj_4817)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_13_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2143_13 (.CI(n28421), .I0(n3099), .I1(n3116), .CO(n28422));
    SB_LUT4 mod_5_add_2143_12_lut (.I0(n3100), .I1(n3100), .I2(n3116), 
            .I3(n28420), .O(n29_adj_4818)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_12_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2143_12 (.CI(n28420), .I0(n3100), .I1(n3116), .CO(n28421));
    SB_LUT4 mod_5_add_2143_11_lut (.I0(n3101), .I1(n3101), .I2(n3116), 
            .I3(n28419), .O(n27_adj_4819)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_11_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2143_11 (.CI(n28419), .I0(n3101), .I1(n3116), .CO(n28420));
    SB_LUT4 mod_5_add_2143_10_lut (.I0(n3102), .I1(n3102), .I2(n3116), 
            .I3(n28418), .O(n25_adj_4820)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_10_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2143_10 (.CI(n28418), .I0(n3102), .I1(n3116), .CO(n28419));
    SB_LUT4 mod_5_add_2143_9_lut (.I0(n3103), .I1(n3103), .I2(n3116), 
            .I3(n28417), .O(n23_adj_4821)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_9_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2143_9 (.CI(n28417), .I0(n3103), .I1(n3116), .CO(n28418));
    SB_LUT4 mod_5_add_2143_8_lut (.I0(n3104), .I1(n3104), .I2(n3116), 
            .I3(n28416), .O(n21_adj_4822)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_8_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2143_8 (.CI(n28416), .I0(n3104), .I1(n3116), .CO(n28417));
    SB_CARRY sub_14_add_2_28 (.CI(n27970), .I0(timer[26]), .I1(n1[26]), 
            .CO(n27971));
    SB_LUT4 sub_14_add_2_27_lut (.I0(GND_net), .I1(timer[25]), .I2(n1[25]), 
            .I3(n27969), .O(one_wire_N_553[25])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_27_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_2143_7_lut (.I0(n3105), .I1(n3105), .I2(n3116), 
            .I3(n28415), .O(n19_adj_4823)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_7_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2143_7 (.CI(n28415), .I0(n3105), .I1(n3116), .CO(n28416));
    SB_CARRY sub_14_add_2_27 (.CI(n27969), .I0(timer[25]), .I1(n1[25]), 
            .CO(n27970));
    SB_LUT4 mod_5_add_2143_6_lut (.I0(n3106), .I1(n3106), .I2(n3116), 
            .I3(n28414), .O(n17_adj_4824)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_6_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2143_6 (.CI(n28414), .I0(n3106), .I1(n3116), .CO(n28415));
    SB_LUT4 mod_5_add_2143_5_lut (.I0(n3107), .I1(n3107), .I2(n3116), 
            .I3(n28413), .O(n15_adj_4825)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_5_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2143_5 (.CI(n28413), .I0(n3107), .I1(n3116), .CO(n28414));
    SB_LUT4 mod_5_add_2143_4_lut (.I0(n3108), .I1(n3108), .I2(n3116), 
            .I3(n28412), .O(n13_adj_4826)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_4_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2143_4 (.CI(n28412), .I0(n3108), .I1(n3116), .CO(n28413));
    SB_LUT4 bit_ctr_0__bdd_4_lut_31085 (.I0(bit_ctr[0]), .I1(neopxl_color[10]), 
            .I2(neopxl_color[11]), .I3(bit_ctr[1]), .O(n37826));
    defparam bit_ctr_0__bdd_4_lut_31085.LUT_INIT = 16'he4aa;
    SB_LUT4 n37826_bdd_4_lut (.I0(n37826), .I1(neopxl_color[9]), .I2(neopxl_color[8]), 
            .I3(bit_ctr[1]), .O(n35482));
    defparam n37826_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 mod_5_add_2143_3_lut (.I0(n3109), .I1(n3109), .I2(n37636), 
            .I3(n28411), .O(n11_adj_4827)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_3_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_2143_3 (.CI(n28411), .I0(n3109), .I1(n37636), .CO(n28412));
    SB_LUT4 mod_5_add_2143_2_lut (.I0(bit_ctr[4]), .I1(bit_ctr[4]), .I2(n37636), 
            .I3(VCC_net), .O(n3209)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_2_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 add_21_10_lut (.I0(GND_net), .I1(bit_ctr[8]), .I2(GND_net), 
            .I3(n27771), .O(n255[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_14_add_2_26_lut (.I0(GND_net), .I1(timer[24]), .I2(n1[24]), 
            .I3(n27968), .O(one_wire_N_553[24])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_26_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_2143_2 (.CI(VCC_net), .I0(bit_ctr[4]), .I1(n37636), 
            .CO(n28411));
    SB_LUT4 mod_5_add_803_9_lut (.I0(n1103), .I1(n1103), .I2(n1136), .I3(n28410), 
            .O(n1202)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_803_9_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_803_8_lut (.I0(n1104), .I1(n1104), .I2(n1136), .I3(n28409), 
            .O(n1203)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_803_8_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_803_8 (.CI(n28409), .I0(n1104), .I1(n1136), .CO(n28410));
    SB_LUT4 mod_5_add_803_7_lut (.I0(n1105), .I1(n1105), .I2(n1136), .I3(n28408), 
            .O(n1204)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_803_7_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_803_7 (.CI(n28408), .I0(n1105), .I1(n1136), .CO(n28409));
    SB_LUT4 mod_5_add_803_6_lut (.I0(n1106), .I1(n1106), .I2(n1136), .I3(n28407), 
            .O(n1205)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_803_6_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_803_6 (.CI(n28407), .I0(n1106), .I1(n1136), .CO(n28408));
    SB_LUT4 mod_5_add_803_5_lut (.I0(n1107), .I1(n1107), .I2(n1136), .I3(n28406), 
            .O(n1206)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_803_5_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_803_5 (.CI(n28406), .I0(n1107), .I1(n1136), .CO(n28407));
    SB_LUT4 mod_5_add_803_4_lut (.I0(n1108), .I1(n1108), .I2(n1136), .I3(n28405), 
            .O(n1207)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_803_4_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_803_4 (.CI(n28405), .I0(n1108), .I1(n1136), .CO(n28406));
    SB_CARRY sub_14_add_2_26 (.CI(n27968), .I0(timer[24]), .I1(n1[24]), 
            .CO(n27969));
    SB_LUT4 mod_5_add_803_3_lut (.I0(n1109), .I1(n1109), .I2(n37637), 
            .I3(n28404), .O(n1208)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_803_3_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_803_3 (.CI(n28404), .I0(n1109), .I1(n37637), .CO(n28405));
    SB_LUT4 sub_14_add_2_25_lut (.I0(one_wire_N_553[16]), .I1(timer[23]), 
            .I2(n1[23]), .I3(n27967), .O(n30_adj_4810)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_25_lut.LUT_INIT = 16'hebbe;
    SB_LUT4 mod_5_add_803_2_lut (.I0(bit_ctr[24]), .I1(bit_ctr[24]), .I2(n37637), 
            .I3(VCC_net), .O(n1209)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_803_2_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_803_2 (.CI(VCC_net), .I0(bit_ctr[24]), .I1(n37637), 
            .CO(n28404));
    SB_CARRY sub_14_add_2_25 (.CI(n27967), .I0(timer[23]), .I1(n1[23]), 
            .CO(n27968));
    SB_CARRY add_21_10 (.CI(n27771), .I0(bit_ctr[8]), .I1(GND_net), .CO(n27772));
    SB_LUT4 bit_ctr_0__bdd_4_lut_31040 (.I0(bit_ctr[0]), .I1(neopxl_color[14]), 
            .I2(neopxl_color[15]), .I3(bit_ctr[1]), .O(n37820));
    defparam bit_ctr_0__bdd_4_lut_31040.LUT_INIT = 16'he4aa;
    SB_LUT4 n37820_bdd_4_lut (.I0(n37820), .I1(neopxl_color[13]), .I2(neopxl_color[12]), 
            .I3(bit_ctr[1]), .O(n35485));
    defparam n37820_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 bit_ctr_0__bdd_4_lut_31035 (.I0(bit_ctr[0]), .I1(neopxl_color[2]), 
            .I2(neopxl_color[3]), .I3(bit_ctr[1]), .O(n37808));
    defparam bit_ctr_0__bdd_4_lut_31035.LUT_INIT = 16'he4aa;
    SB_LUT4 n37808_bdd_4_lut (.I0(n37808), .I1(neopxl_color[1]), .I2(neopxl_color[0]), 
            .I3(bit_ctr[1]), .O(n35491));
    defparam n37808_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 sub_14_add_2_24_lut (.I0(one_wire_N_553[13]), .I1(timer[22]), 
            .I2(n1[22]), .I3(n27966), .O(n24_adj_4799)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_24_lut.LUT_INIT = 16'hebbe;
    SB_CARRY sub_14_add_2_24 (.CI(n27966), .I0(timer[22]), .I1(n1[22]), 
            .CO(n27967));
    SB_LUT4 sub_14_add_2_23_lut (.I0(one_wire_N_553[14]), .I1(timer[21]), 
            .I2(n1[21]), .I3(n27965), .O(n25_adj_4801)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_23_lut.LUT_INIT = 16'hebbe;
    SB_CARRY sub_14_add_2_23 (.CI(n27965), .I0(timer[21]), .I1(n1[21]), 
            .CO(n27966));
    SB_LUT4 sub_14_add_2_22_lut (.I0(one_wire_N_553[15]), .I1(timer[20]), 
            .I2(n1[20]), .I3(n27964), .O(n29_adj_4809)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_22_lut.LUT_INIT = 16'hebbe;
    SB_LUT4 i4574_2_lut_3_lut_4_lut (.I0(bit_ctr[28]), .I1(n739), .I2(bit_ctr[27]), 
            .I3(n33419), .O(n60));   // verilog/neopixel.v(22[26:36])
    defparam i4574_2_lut_3_lut_4_lut.LUT_INIT = 16'hff90;
    SB_CARRY sub_14_add_2_22 (.CI(n27964), .I0(timer[20]), .I1(n1[20]), 
            .CO(n27965));
    SB_LUT4 sub_14_add_2_21_lut (.I0(GND_net), .I1(timer[19]), .I2(n1[19]), 
            .I3(n27963), .O(one_wire_N_553[19])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 bit_ctr_0__bdd_4_lut_31025 (.I0(bit_ctr[0]), .I1(neopxl_color[22]), 
            .I2(neopxl_color[23]), .I3(bit_ctr[1]), .O(n37742));
    defparam bit_ctr_0__bdd_4_lut_31025.LUT_INIT = 16'he4aa;
    SB_LUT4 n37742_bdd_4_lut (.I0(n37742), .I1(neopxl_color[21]), .I2(neopxl_color[20]), 
            .I3(bit_ctr[1]), .O(n37745));
    defparam n37742_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 bit_ctr_0__bdd_4_lut_30971 (.I0(bit_ctr[0]), .I1(neopxl_color[6]), 
            .I2(neopxl_color[7]), .I3(bit_ctr[1]), .O(n37730));
    defparam bit_ctr_0__bdd_4_lut_30971.LUT_INIT = 16'he4aa;
    SB_LUT4 n37730_bdd_4_lut (.I0(n37730), .I1(neopxl_color[5]), .I2(neopxl_color[4]), 
            .I3(bit_ctr[1]), .O(n36892));
    defparam n37730_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_CARRY sub_14_add_2_21 (.CI(n27963), .I0(timer[19]), .I1(n1[19]), 
            .CO(n27964));
    SB_LUT4 add_21_9_lut (.I0(GND_net), .I1(bit_ctr[7]), .I2(GND_net), 
            .I3(n27770), .O(n255[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_14_add_2_20_lut (.I0(GND_net), .I1(timer[18]), .I2(n1[18]), 
            .I3(n27962), .O(one_wire_N_553[18])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_14_add_2_20 (.CI(n27962), .I0(timer[18]), .I1(n1[18]), 
            .CO(n27963));
    SB_LUT4 sub_14_add_2_19_lut (.I0(one_wire_N_553[12]), .I1(timer[17]), 
            .I2(n1[17]), .I3(n27961), .O(n27_adj_4802)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_19_lut.LUT_INIT = 16'hebbe;
    SB_CARRY sub_14_add_2_19 (.CI(n27961), .I0(timer[17]), .I1(n1[17]), 
            .CO(n27962));
    SB_LUT4 sub_14_add_2_18_lut (.I0(GND_net), .I1(timer[16]), .I2(n1[16]), 
            .I3(n27960), .O(one_wire_N_553[16])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_14_add_2_18 (.CI(n27960), .I0(timer[16]), .I1(n1[16]), 
            .CO(n27961));
    SB_LUT4 sub_14_add_2_17_lut (.I0(GND_net), .I1(timer[15]), .I2(n1[15]), 
            .I3(n27959), .O(one_wire_N_553[15])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_14_add_2_17 (.CI(n27959), .I0(timer[15]), .I1(n1[15]), 
            .CO(n27960));
    SB_CARRY add_21_11 (.CI(n27772), .I0(bit_ctr[9]), .I1(GND_net), .CO(n27773));
    SB_LUT4 i26697_2_lut_4_lut (.I0(bit_ctr[28]), .I1(n8799), .I2(n608), 
            .I3(bit_ctr[29]), .O(n33444));
    defparam i26697_2_lut_4_lut.LUT_INIT = 16'h02a8;
    SB_LUT4 sub_14_add_2_16_lut (.I0(GND_net), .I1(timer[14]), .I2(n1[14]), 
            .I3(n27958), .O(one_wire_N_553[14])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_14_add_2_16 (.CI(n27958), .I0(timer[14]), .I1(n1[14]), 
            .CO(n27959));
    SB_LUT4 sub_14_add_2_15_lut (.I0(GND_net), .I1(timer[13]), .I2(n1[13]), 
            .I3(n27957), .O(one_wire_N_553[13])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_14_add_2_15 (.CI(n27957), .I0(timer[13]), .I1(n1[13]), 
            .CO(n27958));
    SB_LUT4 i26783_2_lut (.I0(one_wire_N_553[4]), .I1(n33451), .I2(GND_net), 
            .I3(GND_net), .O(n33533));
    defparam i26783_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i130_4_lut (.I0(n24659), .I1(n33551), .I2(\neo_pixel_transmitter.done ), 
            .I3(\state[1] ), .O(n103));
    defparam i130_4_lut.LUT_INIT = 16'h3530;
    SB_LUT4 i1_4_lut_adj_1577 (.I0(n33545), .I1(n33533), .I2(n33371), 
            .I3(n78), .O(n32559));
    defparam i1_4_lut_adj_1577.LUT_INIT = 16'h1505;
    SB_LUT4 i1_4_lut_adj_1578 (.I0(n17526), .I1(\state[0] ), .I2(n32559), 
            .I3(n103), .O(n18588));
    defparam i1_4_lut_adj_1578.LUT_INIT = 16'h5150;
    SB_LUT4 i3_1_lut (.I0(\neo_pixel_transmitter.done ), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(\neo_pixel_transmitter.done_N_616 ));   // verilog/neopixel.v(35[12] 117[6])
    defparam i3_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i30885_1_lut (.I0(n1235), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n37638));
    defparam i30885_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i1_1_lut (.I0(\neo_pixel_transmitter.t0 [0]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[0]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i1_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i6_4_lut_adj_1579 (.I0(n1205), .I1(n1206), .I2(n1204), .I3(n1207), 
            .O(n14_adj_4829));
    defparam i6_4_lut_adj_1579.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_3_lut_adj_1580 (.I0(bit_ctr[23]), .I1(n1203), .I2(n1209), 
            .I3(GND_net), .O(n9_adj_4830));
    defparam i1_3_lut_adj_1580.LUT_INIT = 16'hecec;
    SB_LUT4 i7_4_lut_adj_1581 (.I0(n9_adj_4830), .I1(n14_adj_4829), .I2(n1202), 
            .I3(n1208), .O(n1235));
    defparam i7_4_lut_adj_1581.LUT_INIT = 16'hfffe;
    SB_LUT4 sub_14_add_2_14_lut (.I0(GND_net), .I1(timer[12]), .I2(n1[12]), 
            .I3(n27956), .O(one_wire_N_553[12])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_14_add_2_14 (.CI(n27956), .I0(timer[12]), .I1(n1[12]), 
            .CO(n27957));
    SB_LUT4 sub_14_add_2_13_lut (.I0(GND_net), .I1(timer[11]), .I2(n1[11]), 
            .I3(n27955), .O(one_wire_N_553[11])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_14_inv_0_i2_1_lut (.I0(\neo_pixel_transmitter.t0 [1]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[1]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_DFFESS state_i0 (.Q(\state[0] ), .C(clk32MHz), .E(n18685), .D(state_3__N_402[0]), 
            .S(n33425));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF timer_1579__i1 (.Q(timer[1]), .C(clk32MHz), .D(n133[1]));   // verilog/neopixel.v(12[12:21])
    SB_CARRY sub_14_add_2_13 (.CI(n27955), .I0(timer[11]), .I1(n1[11]), 
            .CO(n27956));
    SB_LUT4 sub_14_add_2_12_lut (.I0(GND_net), .I1(timer[10]), .I2(n1[10]), 
            .I3(n27954), .O(one_wire_N_553[10])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_14_inv_0_i3_1_lut (.I0(\neo_pixel_transmitter.t0 [2]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[2]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1_2_lut_adj_1582 (.I0(bit_ctr[27]), .I1(n838), .I2(GND_net), 
            .I3(GND_net), .O(n16024));
    defparam i1_2_lut_adj_1582.LUT_INIT = 16'h9999;
    SB_LUT4 sub_14_inv_0_i4_1_lut (.I0(\neo_pixel_transmitter.t0 [3]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[3]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i5_1_lut (.I0(\neo_pixel_transmitter.t0 [4]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[4]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i6_1_lut (.I0(\neo_pixel_transmitter.t0 [5]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[5]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i7_1_lut (.I0(\neo_pixel_transmitter.t0 [6]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[6]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i8_1_lut (.I0(\neo_pixel_transmitter.t0 [7]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[7]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i8_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i3_2_lut_adj_1583 (.I0(n2302), .I1(n2292), .I2(GND_net), .I3(GND_net), 
            .O(n22_adj_4840));
    defparam i3_2_lut_adj_1583.LUT_INIT = 16'heeee;
    SB_LUT4 i11_4_lut_adj_1584 (.I0(bit_ctr[12]), .I1(n22_adj_4840), .I2(n2299), 
            .I3(n2309), .O(n30_adj_4841));
    defparam i11_4_lut_adj_1584.LUT_INIT = 16'hfefc;
    SB_LUT4 i15_4_lut_adj_1585 (.I0(n2294), .I1(n30_adj_4841), .I2(n2306), 
            .I3(n2297), .O(n34_adj_4842));
    defparam i15_4_lut_adj_1585.LUT_INIT = 16'hfffe;
    SB_LUT4 i13_4_lut_adj_1586 (.I0(n2301), .I1(n2307), .I2(n2291), .I3(n2305), 
            .O(n32_adj_4843));
    defparam i13_4_lut_adj_1586.LUT_INIT = 16'hfffe;
    SB_LUT4 i14_4_lut_adj_1587 (.I0(n2298), .I1(n2295), .I2(n2304), .I3(n2300), 
            .O(n33_adj_4844));
    defparam i14_4_lut_adj_1587.LUT_INIT = 16'hfffe;
    SB_LUT4 i12_4_lut_adj_1588 (.I0(n2308), .I1(n2296), .I2(n2303), .I3(n2293), 
            .O(n31_adj_4845));
    defparam i12_4_lut_adj_1588.LUT_INIT = 16'hfffe;
    SB_LUT4 i18_4_lut_adj_1589 (.I0(n31_adj_4845), .I1(n33_adj_4844), .I2(n32_adj_4843), 
            .I3(n34_adj_4842), .O(n2324));
    defparam i18_4_lut_adj_1589.LUT_INIT = 16'hfffe;
    SB_LUT4 i30877_1_lut (.I0(n2225), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n37630));
    defparam i30877_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_21_33_lut (.I0(GND_net), .I1(bit_ctr[31]), .I2(GND_net), 
            .I3(n27794), .O(n255[31])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_33_lut.LUT_INIT = 16'hC33C;
    SB_DFFE state_i1 (.Q(\state[1] ), .C(clk32MHz), .E(VCC_net), .D(n19040));   // verilog/neopixel.v(35[12] 117[6])
    SB_LUT4 i4298_2_lut_3_lut (.I0(bit_ctr[30]), .I1(bit_ctr[31]), .I2(bit_ctr[29]), 
            .I3(GND_net), .O(n8799));   // verilog/neopixel.v(22[26:36])
    defparam i4298_2_lut_3_lut.LUT_INIT = 16'h2020;
    SB_DFF \neo_pixel_transmitter.t0_i0_i1  (.Q(\neo_pixel_transmitter.t0 [1]), 
           .C(clk32MHz), .D(n19557));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i2  (.Q(\neo_pixel_transmitter.t0 [2]), 
           .C(clk32MHz), .D(n19556));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i3  (.Q(\neo_pixel_transmitter.t0 [3]), 
           .C(clk32MHz), .D(n19555));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i4  (.Q(\neo_pixel_transmitter.t0 [4]), 
           .C(clk32MHz), .D(n19554));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i5  (.Q(\neo_pixel_transmitter.t0 [5]), 
           .C(clk32MHz), .D(n19553));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i6  (.Q(\neo_pixel_transmitter.t0 [6]), 
           .C(clk32MHz), .D(n19552));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i7  (.Q(\neo_pixel_transmitter.t0 [7]), 
           .C(clk32MHz), .D(n19551));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i8  (.Q(\neo_pixel_transmitter.t0 [8]), 
           .C(clk32MHz), .D(n19550));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i9  (.Q(\neo_pixel_transmitter.t0 [9]), 
           .C(clk32MHz), .D(n19549));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i10  (.Q(\neo_pixel_transmitter.t0 [10]), 
           .C(clk32MHz), .D(n19548));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i11  (.Q(\neo_pixel_transmitter.t0 [11]), 
           .C(clk32MHz), .D(n19547));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i12  (.Q(\neo_pixel_transmitter.t0 [12]), 
           .C(clk32MHz), .D(n19546));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i13  (.Q(\neo_pixel_transmitter.t0 [13]), 
           .C(clk32MHz), .D(n19545));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i14  (.Q(\neo_pixel_transmitter.t0 [14]), 
           .C(clk32MHz), .D(n19544));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i15  (.Q(\neo_pixel_transmitter.t0 [15]), 
           .C(clk32MHz), .D(n19543));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i16  (.Q(\neo_pixel_transmitter.t0 [16]), 
           .C(clk32MHz), .D(n19542));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i17  (.Q(\neo_pixel_transmitter.t0 [17]), 
           .C(clk32MHz), .D(n19541));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i18  (.Q(\neo_pixel_transmitter.t0 [18]), 
           .C(clk32MHz), .D(n19540));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i19  (.Q(\neo_pixel_transmitter.t0 [19]), 
           .C(clk32MHz), .D(n19539));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i20  (.Q(\neo_pixel_transmitter.t0 [20]), 
           .C(clk32MHz), .D(n19538));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i21  (.Q(\neo_pixel_transmitter.t0 [21]), 
           .C(clk32MHz), .D(n19537));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i22  (.Q(\neo_pixel_transmitter.t0 [22]), 
           .C(clk32MHz), .D(n19536));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i23  (.Q(\neo_pixel_transmitter.t0 [23]), 
           .C(clk32MHz), .D(n19535));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i24  (.Q(\neo_pixel_transmitter.t0 [24]), 
           .C(clk32MHz), .D(n19534));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i25  (.Q(\neo_pixel_transmitter.t0 [25]), 
           .C(clk32MHz), .D(n19533));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i26  (.Q(\neo_pixel_transmitter.t0 [26]), 
           .C(clk32MHz), .D(n19529));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i27  (.Q(\neo_pixel_transmitter.t0 [27]), 
           .C(clk32MHz), .D(n19528));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i28  (.Q(\neo_pixel_transmitter.t0 [28]), 
           .C(clk32MHz), .D(n19527));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i29  (.Q(\neo_pixel_transmitter.t0 [29]), 
           .C(clk32MHz), .D(n19526));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i30  (.Q(\neo_pixel_transmitter.t0 [30]), 
           .C(clk32MHz), .D(n19525));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i31  (.Q(\neo_pixel_transmitter.t0 [31]), 
           .C(clk32MHz), .D(n19521));   // verilog/neopixel.v(35[12] 117[6])
    SB_CARRY sub_14_add_2_12 (.CI(n27954), .I0(timer[10]), .I1(n1[10]), 
            .CO(n27955));
    SB_LUT4 add_21_32_lut (.I0(GND_net), .I1(bit_ctr[30]), .I2(GND_net), 
            .I3(n27793), .O(n255[30])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_32_lut.LUT_INIT = 16'hC33C;
    SB_DFFESR bit_ctr_i0_i0 (.Q(bit_ctr[0]), .C(clk32MHz), .E(n18566), 
            .D(n255[0]), .R(n18886));   // verilog/neopixel.v(35[12] 117[6])
    SB_LUT4 i29756_3_lut_4_lut (.I0(bit_ctr[28]), .I1(n739), .I2(bit_ctr[27]), 
            .I3(n838), .O(n18794));
    defparam i29756_3_lut_4_lut.LUT_INIT = 16'h9969;
    SB_CARRY add_21_32 (.CI(n27793), .I0(bit_ctr[30]), .I1(GND_net), .CO(n27794));
    SB_LUT4 add_21_8_lut (.I0(GND_net), .I1(bit_ctr[6]), .I2(GND_net), 
            .I3(n27769), .O(n255[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i8_3_lut (.I0(bit_ctr[6]), .I1(n2907), .I2(n2909), .I3(GND_net), 
            .O(n33_adj_4846));
    defparam i8_3_lut.LUT_INIT = 16'hecec;
    SB_LUT4 mod_5_add_669_7_lut (.I0(GND_net), .I1(n905), .I2(VCC_net), 
            .I3(n27882), .O(n971[31])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_669_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i16_4_lut_adj_1590 (.I0(n2900), .I1(n2891), .I2(n2897), .I3(n2888), 
            .O(n41_adj_4847));
    defparam i16_4_lut_adj_1590.LUT_INIT = 16'hfffe;
    SB_LUT4 mod_5_add_669_6_lut (.I0(GND_net), .I1(n906), .I2(VCC_net), 
            .I3(n27881), .O(n971[30])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_669_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_14_add_2_11_lut (.I0(GND_net), .I1(timer[9]), .I2(n1[9]), 
            .I3(n27953), .O(one_wire_N_553[9])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_14_add_2_11 (.CI(n27953), .I0(timer[9]), .I1(n1[9]), 
            .CO(n27954));
    SB_LUT4 sub_14_inv_0_i9_1_lut (.I0(\neo_pixel_transmitter.t0 [8]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[8]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i9_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i13_3_lut_adj_1591 (.I0(n2906), .I1(n2887), .I2(n2892), .I3(GND_net), 
            .O(n38_adj_4850));
    defparam i13_3_lut_adj_1591.LUT_INIT = 16'hfefe;
    SB_LUT4 sub_14_add_2_10_lut (.I0(one_wire_N_553[10]), .I1(timer[8]), 
            .I2(n1[8]), .I3(n27952), .O(n10_adj_4795)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_10_lut.LUT_INIT = 16'hebbe;
    SB_LUT4 i18_4_lut_adj_1592 (.I0(n2896), .I1(n2885), .I2(n2905), .I3(n2902), 
            .O(n43_adj_4851));
    defparam i18_4_lut_adj_1592.LUT_INIT = 16'hfffe;
    SB_LUT4 i15_4_lut_adj_1593 (.I0(n2899), .I1(n2890), .I2(n2898), .I3(n2908), 
            .O(n40_adj_4852));
    defparam i15_4_lut_adj_1593.LUT_INIT = 16'hfffe;
    SB_LUT4 sub_14_inv_0_i10_1_lut (.I0(\neo_pixel_transmitter.t0 [9]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[9]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i10_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i21_4_lut_adj_1594 (.I0(n41_adj_4847), .I1(n33_adj_4846), .I2(n2889), 
            .I3(n2901), .O(n46_adj_4853));
    defparam i21_4_lut_adj_1594.LUT_INIT = 16'hfffe;
    SB_LUT4 add_21_31_lut (.I0(GND_net), .I1(bit_ctr[29]), .I2(GND_net), 
            .I3(n27792), .O(n255[29])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_31_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_669_6 (.CI(n27881), .I0(n906), .I1(VCC_net), .CO(n27882));
    SB_LUT4 i14_4_lut_adj_1595 (.I0(n2886), .I1(n2894), .I2(n2895), .I3(n2903), 
            .O(n39_adj_4854));
    defparam i14_4_lut_adj_1595.LUT_INIT = 16'hfffe;
    SB_LUT4 mod_5_add_669_5_lut (.I0(GND_net), .I1(n907), .I2(VCC_net), 
            .I3(n27880), .O(n971[29])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_669_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_14_add_2_10 (.CI(n27952), .I0(timer[8]), .I1(n1[8]), 
            .CO(n27953));
    SB_LUT4 sub_14_add_2_9_lut (.I0(GND_net), .I1(timer[7]), .I2(n1[7]), 
            .I3(n27951), .O(one_wire_N_553[7])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_669_5 (.CI(n27880), .I0(n907), .I1(VCC_net), .CO(n27881));
    SB_LUT4 i22_4_lut (.I0(n43_adj_4851), .I1(n2904), .I2(n38_adj_4850), 
            .I3(n2893), .O(n47_adj_4855));
    defparam i22_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 mod_5_i605_3_lut (.I0(n807), .I1(n60), .I2(n838), .I3(GND_net), 
            .O(n906));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i605_3_lut.LUT_INIT = 16'ha9a9;
    SB_CARRY sub_14_add_2_9 (.CI(n27951), .I0(timer[7]), .I1(n1[7]), .CO(n27952));
    SB_LUT4 i24_4_lut_adj_1596 (.I0(n47_adj_4855), .I1(n39_adj_4854), .I2(n46_adj_4853), 
            .I3(n40_adj_4852), .O(n2918));
    defparam i24_4_lut_adj_1596.LUT_INIT = 16'hfffe;
    SB_LUT4 sub_14_add_2_8_lut (.I0(GND_net), .I1(timer[6]), .I2(n1[6]), 
            .I3(n27950), .O(one_wire_N_553[6])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_669_4_lut (.I0(GND_net), .I1(n18794), .I2(VCC_net), 
            .I3(n27879), .O(n971[28])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_669_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i30878_1_lut (.I0(n2819), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n37631));
    defparam i30878_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i26801_2_lut_3_lut (.I0(n33545), .I1(one_wire_N_553[4]), .I2(n33451), 
            .I3(GND_net), .O(n33551));
    defparam i26801_2_lut_3_lut.LUT_INIT = 16'heaea;
    SB_CARRY sub_14_add_2_8 (.CI(n27950), .I0(timer[6]), .I1(n1[6]), .CO(n27951));
    SB_LUT4 sub_14_add_2_7_lut (.I0(GND_net), .I1(timer[5]), .I2(n1[5]), 
            .I3(n27949), .O(one_wire_N_553[5])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mux_788_Mux_0_i3_3_lut_3_lut (.I0(\neo_pixel_transmitter.done ), 
            .I1(start), .I2(\state[1] ), .I3(GND_net), .O(\neo_pixel_transmitter.done_N_610 ));   // verilog/neopixel.v(36[4] 116[11])
    defparam mux_788_Mux_0_i3_3_lut_3_lut.LUT_INIT = 16'ha1a1;
    SB_CARRY sub_14_add_2_7 (.CI(n27949), .I0(timer[5]), .I1(n1[5]), .CO(n27950));
    SB_LUT4 sub_14_add_2_6_lut (.I0(GND_net), .I1(timer[4]), .I2(n1[4]), 
            .I3(n27948), .O(one_wire_N_553[4])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_21_31 (.CI(n27792), .I0(bit_ctr[29]), .I1(GND_net), .CO(n27793));
    SB_CARRY mod_5_add_669_4 (.CI(n27879), .I0(n18794), .I1(VCC_net), 
            .CO(n27880));
    SB_LUT4 i18779_2_lut (.I0(bit_ctr[30]), .I1(bit_ctr[31]), .I2(GND_net), 
            .I3(GND_net), .O(n608));   // verilog/neopixel.v(22[26:36])
    defparam i18779_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i2_4_lut (.I0(n708), .I1(n608), .I2(n33444), .I3(n8799), 
            .O(n739));
    defparam i2_4_lut.LUT_INIT = 16'h0105;
    SB_CARRY sub_14_add_2_6 (.CI(n27948), .I0(timer[4]), .I1(n1[4]), .CO(n27949));
    SB_LUT4 sub_14_add_2_5_lut (.I0(GND_net), .I1(timer[3]), .I2(n1[3]), 
            .I3(n27947), .O(one_wire_N_553[3])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_2_lut_adj_1597 (.I0(bit_ctr[28]), .I1(n739), .I2(GND_net), 
            .I3(GND_net), .O(n16028));
    defparam i1_2_lut_adj_1597.LUT_INIT = 16'h6666;
    SB_LUT4 mod_5_add_669_3_lut (.I0(GND_net), .I1(n16024), .I2(GND_net), 
            .I3(n27878), .O(n971[27])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_669_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_14_add_2_5 (.CI(n27947), .I0(timer[3]), .I1(n1[3]), .CO(n27948));
    SB_LUT4 sub_14_add_2_4_lut (.I0(GND_net), .I1(timer[2]), .I2(n1[2]), 
            .I3(n27946), .O(one_wire_N_553[2])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_3_lut_2_lut (.I0(\state[0] ), .I1(\neo_pixel_transmitter.done ), 
            .I2(GND_net), .I3(GND_net), .O(n32651));
    defparam i1_3_lut_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY mod_5_add_669_3 (.CI(n27878), .I0(n16024), .I1(GND_net), 
            .CO(n27879));
    SB_CARRY sub_14_add_2_4 (.CI(n27946), .I0(timer[2]), .I1(n1[2]), .CO(n27947));
    SB_LUT4 i29826_3_lut_4_lut (.I0(n29522), .I1(start), .I2(\neo_pixel_transmitter.done ), 
            .I3(n17393), .O(n36280));
    defparam i29826_3_lut_4_lut.LUT_INIT = 16'hcfdf;
    SB_LUT4 i29726_3_lut (.I0(n29995), .I1(bit_ctr[28]), .I2(n739), .I3(GND_net), 
            .O(n33419));
    defparam i29726_3_lut.LUT_INIT = 16'ha6a6;
    SB_LUT4 sub_14_add_2_3_lut (.I0(n4_adj_4856), .I1(timer[1]), .I2(n1[1]), 
            .I3(n27945), .O(n29671)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_3_lut.LUT_INIT = 16'hebbe;
    SB_LUT4 i2_2_lut_3_lut (.I0(n17393), .I1(one_wire_N_553[4]), .I2(n24675), 
            .I3(GND_net), .O(n24735));
    defparam i2_2_lut_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i2_3_lut_4_lut_adj_1598 (.I0(\state[0] ), .I1(\state[1] ), .I2(LED_c), 
            .I3(\state_3__N_402[1] ), .O(n18886));   // verilog/neopixel.v(35[12] 117[6])
    defparam i2_3_lut_4_lut_adj_1598.LUT_INIT = 16'h8000;
    SB_LUT4 mod_5_add_669_2_lut (.I0(GND_net), .I1(bit_ctr[26]), .I2(GND_net), 
            .I3(VCC_net), .O(n971[26])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_669_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_14_add_2_3 (.CI(n27945), .I0(timer[1]), .I1(n1[1]), .CO(n27946));
    SB_LUT4 mod_5_i538_3_lut (.I0(n708), .I1(n33444), .I2(n739), .I3(GND_net), 
            .O(n807));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i538_3_lut.LUT_INIT = 16'ha9a9;
    SB_LUT4 mod_5_add_870_10_lut (.I0(n1202), .I1(n1202), .I2(n1235), 
            .I3(n28196), .O(n1301)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_870_10_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_870_9_lut (.I0(n1203), .I1(n1203), .I2(n1235), .I3(n28195), 
            .O(n1302)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_870_9_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_870_9 (.CI(n28195), .I0(n1203), .I1(n1235), .CO(n28196));
    SB_LUT4 mod_5_add_870_8_lut (.I0(n1204), .I1(n1204), .I2(n1235), .I3(n28194), 
            .O(n1303)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_870_8_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_870_8 (.CI(n28194), .I0(n1204), .I1(n1235), .CO(n28195));
    SB_LUT4 mod_5_add_870_7_lut (.I0(n1205), .I1(n1205), .I2(n1235), .I3(n28193), 
            .O(n1304)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_870_7_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_i604_4_lut (.I0(n807), .I1(n838), .I2(n60), .I3(GND_net), 
            .O(n905));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i604_4_lut.LUT_INIT = 16'h0101;
    SB_CARRY mod_5_add_870_7 (.CI(n28193), .I0(n1205), .I1(n1235), .CO(n28194));
    SB_LUT4 mod_5_add_870_6_lut (.I0(n1206), .I1(n1206), .I2(n1235), .I3(n28192), 
            .O(n1305)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_870_6_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_870_6 (.CI(n28192), .I0(n1206), .I1(n1235), .CO(n28193));
    SB_LUT4 mod_5_add_870_5_lut (.I0(n1207), .I1(n1207), .I2(n1235), .I3(n28191), 
            .O(n1306)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_870_5_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_870_5 (.CI(n28191), .I0(n1207), .I1(n1235), .CO(n28192));
    SB_LUT4 mod_5_add_870_4_lut (.I0(n1208), .I1(n1208), .I2(n1235), .I3(n28190), 
            .O(n1307)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_870_4_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_870_4 (.CI(n28190), .I0(n1208), .I1(n1235), .CO(n28191));
    SB_LUT4 sub_14_add_2_2_lut (.I0(one_wire_N_553[2]), .I1(timer[0]), .I2(n1[0]), 
            .I3(VCC_net), .O(n4_adj_4856)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_2_lut.LUT_INIT = 16'hebbe;
    SB_LUT4 mod_5_add_870_3_lut (.I0(n1209), .I1(n1209), .I2(n37638), 
            .I3(n28189), .O(n1308)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_870_3_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_870_3 (.CI(n28189), .I0(n1209), .I1(n37638), .CO(n28190));
    SB_LUT4 mod_5_add_870_2_lut (.I0(bit_ctr[23]), .I1(bit_ctr[23]), .I2(n37638), 
            .I3(VCC_net), .O(n1309)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_870_2_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_870_2 (.CI(VCC_net), .I0(bit_ctr[23]), .I1(n37638), 
            .CO(n28189));
    SB_LUT4 add_21_30_lut (.I0(GND_net), .I1(bit_ctr[28]), .I2(GND_net), 
            .I3(n27791), .O(n255[28])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_30_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_14_add_2_2 (.CI(VCC_net), .I0(timer[0]), .I1(n1[0]), 
            .CO(n27945));
    SB_DFF timer_1579__i2 (.Q(timer[2]), .C(clk32MHz), .D(n133[2]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1579__i3 (.Q(timer[3]), .C(clk32MHz), .D(n133[3]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1579__i4 (.Q(timer[4]), .C(clk32MHz), .D(n133[4]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1579__i5 (.Q(timer[5]), .C(clk32MHz), .D(n133[5]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1579__i6 (.Q(timer[6]), .C(clk32MHz), .D(n133[6]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1579__i7 (.Q(timer[7]), .C(clk32MHz), .D(n133[7]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1579__i8 (.Q(timer[8]), .C(clk32MHz), .D(n133[8]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1579__i9 (.Q(timer[9]), .C(clk32MHz), .D(n133[9]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1579__i10 (.Q(timer[10]), .C(clk32MHz), .D(n133[10]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1579__i11 (.Q(timer[11]), .C(clk32MHz), .D(n133[11]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1579__i12 (.Q(timer[12]), .C(clk32MHz), .D(n133[12]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1579__i13 (.Q(timer[13]), .C(clk32MHz), .D(n133[13]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1579__i14 (.Q(timer[14]), .C(clk32MHz), .D(n133[14]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1579__i15 (.Q(timer[15]), .C(clk32MHz), .D(n133[15]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1579__i16 (.Q(timer[16]), .C(clk32MHz), .D(n133[16]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1579__i17 (.Q(timer[17]), .C(clk32MHz), .D(n133[17]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1579__i18 (.Q(timer[18]), .C(clk32MHz), .D(n133[18]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1579__i19 (.Q(timer[19]), .C(clk32MHz), .D(n133[19]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1579__i20 (.Q(timer[20]), .C(clk32MHz), .D(n133[20]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1579__i21 (.Q(timer[21]), .C(clk32MHz), .D(n133[21]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1579__i22 (.Q(timer[22]), .C(clk32MHz), .D(n133[22]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1579__i23 (.Q(timer[23]), .C(clk32MHz), .D(n133[23]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1579__i24 (.Q(timer[24]), .C(clk32MHz), .D(n133[24]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1579__i25 (.Q(timer[25]), .C(clk32MHz), .D(n133[25]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1579__i26 (.Q(timer[26]), .C(clk32MHz), .D(n133[26]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1579__i27 (.Q(timer[27]), .C(clk32MHz), .D(n133[27]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1579__i28 (.Q(timer[28]), .C(clk32MHz), .D(n133[28]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1579__i29 (.Q(timer[29]), .C(clk32MHz), .D(n133[29]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1579__i30 (.Q(timer[30]), .C(clk32MHz), .D(n133[30]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1579__i31 (.Q(timer[31]), .C(clk32MHz), .D(n133[31]));   // verilog/neopixel.v(12[12:21])
    SB_DFFESR one_wire_108 (.Q(NEOPXL_c), .C(clk32MHz), .E(n18588), .D(\neo_pixel_transmitter.done_N_616 ), 
            .R(n33926));   // verilog/neopixel.v(35[12] 117[6])
    SB_CARRY add_21_30 (.CI(n27791), .I0(bit_ctr[28]), .I1(GND_net), .CO(n27792));
    SB_DFF start_103 (.Q(start), .C(clk32MHz), .D(n31453));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i0  (.Q(\neo_pixel_transmitter.t0 [0]), 
           .C(clk32MHz), .D(n19022));   // verilog/neopixel.v(35[12] 117[6])
    SB_CARRY mod_5_add_669_2 (.CI(VCC_net), .I0(bit_ctr[26]), .I1(GND_net), 
            .CO(n27878));
    SB_LUT4 i3_4_lut_4_lut (.I0(n33419), .I1(n16028), .I2(n807), .I3(bit_ctr[27]), 
            .O(n838));
    defparam i3_4_lut_4_lut.LUT_INIT = 16'h0405;
    SB_LUT4 i30379_3_lut_4_lut (.I0(n16028), .I1(bit_ctr[27]), .I2(n838), 
            .I3(n33419), .O(n907));   // verilog/neopixel.v(22[26:36])
    defparam i30379_3_lut_4_lut.LUT_INIT = 16'hf40b;
    SB_LUT4 i16_4_lut_adj_1599 (.I0(n2798), .I1(n2804), .I2(n2791), .I3(n2795), 
            .O(n40_adj_4857));
    defparam i16_4_lut_adj_1599.LUT_INIT = 16'hfffe;
    SB_LUT4 i14_4_lut_adj_1600 (.I0(n2796), .I1(n2793), .I2(n2788), .I3(n2808), 
            .O(n38_adj_4858));
    defparam i14_4_lut_adj_1600.LUT_INIT = 16'hfffe;
    SB_LUT4 mod_5_add_736_8_lut (.I0(n4), .I1(n4), .I2(n1037), .I3(n28867), 
            .O(n1103)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_736_8_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 add_21_29_lut (.I0(GND_net), .I1(bit_ctr[27]), .I2(GND_net), 
            .I3(n27790), .O(n255[27])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_29_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_736_7_lut (.I0(n1005), .I1(n1005), .I2(n1037), .I3(n28866), 
            .O(n1104)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_736_7_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_736_7 (.CI(n28866), .I0(n1005), .I1(n1037), .CO(n28867));
    SB_LUT4 mod_5_add_736_6_lut (.I0(n1006), .I1(n1006), .I2(n1037), .I3(n28865), 
            .O(n1105)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_736_6_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_736_6 (.CI(n28865), .I0(n1006), .I1(n1037), .CO(n28866));
    SB_LUT4 mod_5_add_736_5_lut (.I0(n1007), .I1(n1007), .I2(n1037), .I3(n28864), 
            .O(n1106)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_736_5_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_736_5 (.CI(n28864), .I0(n1007), .I1(n1037), .CO(n28865));
    SB_LUT4 mod_5_add_736_4_lut (.I0(n1008), .I1(n1008), .I2(n1037), .I3(n28863), 
            .O(n1107)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_736_4_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_736_4 (.CI(n28863), .I0(n1008), .I1(n1037), .CO(n28864));
    SB_LUT4 mod_5_add_736_3_lut (.I0(n1009), .I1(n1009), .I2(n37639), 
            .I3(n28862), .O(n1108)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_736_3_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_736_3 (.CI(n28862), .I0(n1009), .I1(n37639), .CO(n28863));
    SB_LUT4 mod_5_add_736_2_lut (.I0(bit_ctr[25]), .I1(bit_ctr[25]), .I2(n37639), 
            .I3(VCC_net), .O(n1109)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_736_2_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_736_2 (.CI(VCC_net), .I0(bit_ctr[25]), .I1(n37639), 
            .CO(n28862));
    SB_LUT4 mod_5_add_1004_12_lut (.I0(n1400), .I1(n1400), .I2(n1433), 
            .I3(n28861), .O(n1499)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1004_12_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i15_4_lut_adj_1601 (.I0(n2789), .I1(n2800), .I2(n2803), .I3(n2805), 
            .O(n39_adj_4859));
    defparam i15_4_lut_adj_1601.LUT_INIT = 16'hfffe;
    SB_LUT4 mod_5_add_1004_11_lut (.I0(n1401), .I1(n1401), .I2(n1433), 
            .I3(n28860), .O(n1500)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1004_11_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1004_11 (.CI(n28860), .I0(n1401), .I1(n1433), .CO(n28861));
    SB_LUT4 mod_5_add_1004_10_lut (.I0(n1402), .I1(n1402), .I2(n1433), 
            .I3(n28859), .O(n1501)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1004_10_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1004_10 (.CI(n28859), .I0(n1402), .I1(n1433), .CO(n28860));
    SB_LUT4 mod_5_add_1004_9_lut (.I0(n1403), .I1(n1403), .I2(n1433), 
            .I3(n28858), .O(n1502)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1004_9_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1004_9 (.CI(n28858), .I0(n1403), .I1(n1433), .CO(n28859));
    SB_LUT4 i13_4_lut_adj_1602 (.I0(n2792), .I1(n2787), .I2(n2801), .I3(n2799), 
            .O(n37_adj_4860));
    defparam i13_4_lut_adj_1602.LUT_INIT = 16'hfffe;
    SB_LUT4 mod_5_add_1004_8_lut (.I0(n1404), .I1(n1404), .I2(n1433), 
            .I3(n28857), .O(n1503)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1004_8_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1004_8 (.CI(n28857), .I0(n1404), .I1(n1433), .CO(n28858));
    SB_LUT4 mod_5_add_1004_7_lut (.I0(n1405), .I1(n1405), .I2(n1433), 
            .I3(n28856), .O(n1504)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1004_7_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1004_7 (.CI(n28856), .I0(n1405), .I1(n1433), .CO(n28857));
    SB_LUT4 mod_5_add_1004_6_lut (.I0(n1406), .I1(n1406), .I2(n1433), 
            .I3(n28855), .O(n1505)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1004_6_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1004_6 (.CI(n28855), .I0(n1406), .I1(n1433), .CO(n28856));
    SB_LUT4 mod_5_add_1004_5_lut (.I0(n1407), .I1(n1407), .I2(n1433), 
            .I3(n28854), .O(n1506)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1004_5_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1004_5 (.CI(n28854), .I0(n1407), .I1(n1433), .CO(n28855));
    SB_LUT4 mod_5_add_1004_4_lut (.I0(n1408), .I1(n1408), .I2(n1433), 
            .I3(n28853), .O(n1507)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1004_4_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1004_4 (.CI(n28853), .I0(n1408), .I1(n1433), .CO(n28854));
    SB_LUT4 mod_5_add_1004_3_lut (.I0(n1409), .I1(n1409), .I2(n37640), 
            .I3(n28852), .O(n1508)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1004_3_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1004_3 (.CI(n28852), .I0(n1409), .I1(n37640), .CO(n28853));
    SB_LUT4 mod_5_add_1004_2_lut (.I0(bit_ctr[21]), .I1(bit_ctr[21]), .I2(n37640), 
            .I3(VCC_net), .O(n1509)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1004_2_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1004_2 (.CI(VCC_net), .I0(bit_ctr[21]), .I1(n37640), 
            .CO(n28852));
    SB_LUT4 mod_5_add_1071_13_lut (.I0(n1499), .I1(n1499), .I2(n1532), 
            .I3(n28851), .O(n1598)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1071_13_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1071_12_lut (.I0(n1500), .I1(n1500), .I2(n1532), 
            .I3(n28850), .O(n1599)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1071_12_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1071_12 (.CI(n28850), .I0(n1500), .I1(n1532), .CO(n28851));
    SB_LUT4 mod_5_add_1071_11_lut (.I0(n1501), .I1(n1501), .I2(n1532), 
            .I3(n28849), .O(n1600)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1071_11_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1071_11 (.CI(n28849), .I0(n1501), .I1(n1532), .CO(n28850));
    SB_LUT4 mod_5_add_1071_10_lut (.I0(n1502), .I1(n1502), .I2(n1532), 
            .I3(n28848), .O(n1601)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1071_10_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1071_10 (.CI(n28848), .I0(n1502), .I1(n1532), .CO(n28849));
    SB_LUT4 mod_5_add_1071_9_lut (.I0(n1503), .I1(n1503), .I2(n1532), 
            .I3(n28847), .O(n1602)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1071_9_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1071_9 (.CI(n28847), .I0(n1503), .I1(n1532), .CO(n28848));
    SB_LUT4 mod_5_add_1071_8_lut (.I0(n1504), .I1(n1504), .I2(n1532), 
            .I3(n28846), .O(n1603)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1071_8_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1071_8 (.CI(n28846), .I0(n1504), .I1(n1532), .CO(n28847));
    SB_LUT4 mod_5_add_1071_7_lut (.I0(n1505), .I1(n1505), .I2(n1532), 
            .I3(n28845), .O(n1604)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1071_7_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1071_7 (.CI(n28845), .I0(n1505), .I1(n1532), .CO(n28846));
    SB_LUT4 mod_5_add_1071_6_lut (.I0(n1506), .I1(n1506), .I2(n1532), 
            .I3(n28844), .O(n1605)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1071_6_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1071_6 (.CI(n28844), .I0(n1506), .I1(n1532), .CO(n28845));
    SB_LUT4 mod_5_add_1071_5_lut (.I0(n1507), .I1(n1507), .I2(n1532), 
            .I3(n28843), .O(n1606)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1071_5_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1071_5 (.CI(n28843), .I0(n1507), .I1(n1532), .CO(n28844));
    SB_LUT4 mod_5_add_1071_4_lut (.I0(n1508), .I1(n1508), .I2(n1532), 
            .I3(n28842), .O(n1607)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1071_4_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1071_4 (.CI(n28842), .I0(n1508), .I1(n1532), .CO(n28843));
    SB_LUT4 mod_5_add_1071_3_lut (.I0(n1509), .I1(n1509), .I2(n37641), 
            .I3(n28841), .O(n1608)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1071_3_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1071_3 (.CI(n28841), .I0(n1509), .I1(n37641), .CO(n28842));
    SB_CARRY add_21_29 (.CI(n27790), .I0(bit_ctr[27]), .I1(GND_net), .CO(n27791));
    SB_LUT4 mod_5_add_1071_2_lut (.I0(bit_ctr[20]), .I1(bit_ctr[20]), .I2(n37641), 
            .I3(VCC_net), .O(n1609)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1071_2_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1071_2 (.CI(VCC_net), .I0(bit_ctr[20]), .I1(n37641), 
            .CO(n28841));
    SB_LUT4 mod_5_add_1138_14_lut (.I0(n1598), .I1(n1598), .I2(n1631), 
            .I3(n28840), .O(n1697)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1138_14_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1138_13_lut (.I0(n1599), .I1(n1599), .I2(n1631), 
            .I3(n28839), .O(n1698)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1138_13_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1138_13 (.CI(n28839), .I0(n1599), .I1(n1631), .CO(n28840));
    SB_LUT4 i10_2_lut (.I0(n2786), .I1(n2797), .I2(GND_net), .I3(GND_net), 
            .O(n34_adj_4861));
    defparam i10_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i18_4_lut_adj_1603 (.I0(n2794), .I1(n2806), .I2(n2807), .I3(n2790), 
            .O(n42_adj_4862));
    defparam i18_4_lut_adj_1603.LUT_INIT = 16'hfffe;
    SB_LUT4 mod_5_add_1138_12_lut (.I0(n1600), .I1(n1600), .I2(n1631), 
            .I3(n28838), .O(n1699)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1138_12_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i22_4_lut_adj_1604 (.I0(n37_adj_4860), .I1(n39_adj_4859), .I2(n38_adj_4858), 
            .I3(n40_adj_4857), .O(n46_adj_4863));
    defparam i22_4_lut_adj_1604.LUT_INIT = 16'hfffe;
    SB_CARRY mod_5_add_1138_12 (.CI(n28838), .I0(n1600), .I1(n1631), .CO(n28839));
    SB_LUT4 mod_5_add_1138_11_lut (.I0(n1601), .I1(n1601), .I2(n1631), 
            .I3(n28837), .O(n1700)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1138_11_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i9_3_lut (.I0(bit_ctr[7]), .I1(n2802), .I2(n2809), .I3(GND_net), 
            .O(n33_adj_4864));
    defparam i9_3_lut.LUT_INIT = 16'hecec;
    SB_LUT4 i23_4_lut_adj_1605 (.I0(n33_adj_4864), .I1(n46_adj_4863), .I2(n42_adj_4862), 
            .I3(n34_adj_4861), .O(n2819));
    defparam i23_4_lut_adj_1605.LUT_INIT = 16'hfffe;
    SB_CARRY mod_5_add_1138_11 (.CI(n28837), .I0(n1601), .I1(n1631), .CO(n28838));
    SB_LUT4 mod_5_add_1138_10_lut (.I0(n1602), .I1(n1602), .I2(n1631), 
            .I3(n28836), .O(n1701)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1138_10_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1138_10 (.CI(n28836), .I0(n1602), .I1(n1631), .CO(n28837));
    SB_LUT4 mod_5_add_1138_9_lut (.I0(n1603), .I1(n1603), .I2(n1631), 
            .I3(n28835), .O(n1702)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1138_9_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1138_9 (.CI(n28835), .I0(n1603), .I1(n1631), .CO(n28836));
    SB_LUT4 mod_5_add_1138_8_lut (.I0(n1604), .I1(n1604), .I2(n1631), 
            .I3(n28834), .O(n1703)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1138_8_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1138_8 (.CI(n28834), .I0(n1604), .I1(n1631), .CO(n28835));
    SB_LUT4 mod_5_add_1138_7_lut (.I0(n1605), .I1(n1605), .I2(n1631), 
            .I3(n28833), .O(n1704)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1138_7_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1138_7 (.CI(n28833), .I0(n1605), .I1(n1631), .CO(n28834));
    SB_LUT4 mod_5_add_1138_6_lut (.I0(n1606), .I1(n1606), .I2(n1631), 
            .I3(n28832), .O(n1705)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1138_6_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1138_6 (.CI(n28832), .I0(n1606), .I1(n1631), .CO(n28833));
    SB_LUT4 mod_5_add_1138_5_lut (.I0(n1607), .I1(n1607), .I2(n1631), 
            .I3(n28831), .O(n1706)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1138_5_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1138_5 (.CI(n28831), .I0(n1607), .I1(n1631), .CO(n28832));
    SB_LUT4 mod_5_add_1138_4_lut (.I0(n1608), .I1(n1608), .I2(n1631), 
            .I3(n28830), .O(n1707)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1138_4_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1138_4 (.CI(n28830), .I0(n1608), .I1(n1631), .CO(n28831));
    SB_LUT4 add_21_28_lut (.I0(GND_net), .I1(bit_ctr[26]), .I2(GND_net), 
            .I3(n27789), .O(n255[26])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_28_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_1138_3_lut (.I0(n1609), .I1(n1609), .I2(n37642), 
            .I3(n28829), .O(n1708)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1138_3_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1138_3 (.CI(n28829), .I0(n1609), .I1(n37642), .CO(n28830));
    SB_LUT4 mod_5_add_1138_2_lut (.I0(bit_ctr[19]), .I1(bit_ctr[19]), .I2(n37642), 
            .I3(VCC_net), .O(n1709)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1138_2_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1138_2 (.CI(VCC_net), .I0(bit_ctr[19]), .I1(n37642), 
            .CO(n28829));
    SB_LUT4 mod_5_add_1205_15_lut (.I0(n1697), .I1(n1697), .I2(n1730), 
            .I3(n28828), .O(n1796)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1205_15_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1205_14_lut (.I0(n1698), .I1(n1698), .I2(n1730), 
            .I3(n28827), .O(n1797)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1205_14_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1205_14 (.CI(n28827), .I0(n1698), .I1(n1730), .CO(n28828));
    SB_CARRY add_21_28 (.CI(n27789), .I0(bit_ctr[26]), .I1(GND_net), .CO(n27790));
    SB_LUT4 mod_5_add_1205_13_lut (.I0(n1699), .I1(n1699), .I2(n1730), 
            .I3(n28826), .O(n1798)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1205_13_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1205_13 (.CI(n28826), .I0(n1699), .I1(n1730), .CO(n28827));
    SB_LUT4 mod_5_add_1205_12_lut (.I0(n1700), .I1(n1700), .I2(n1730), 
            .I3(n28825), .O(n1799)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1205_12_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1205_12 (.CI(n28825), .I0(n1700), .I1(n1730), .CO(n28826));
    SB_LUT4 mod_5_add_1205_11_lut (.I0(n1701), .I1(n1701), .I2(n1730), 
            .I3(n28824), .O(n1800)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1205_11_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1205_11 (.CI(n28824), .I0(n1701), .I1(n1730), .CO(n28825));
    SB_LUT4 mod_5_add_1205_10_lut (.I0(n1702), .I1(n1702), .I2(n1730), 
            .I3(n28823), .O(n1801)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1205_10_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1205_10 (.CI(n28823), .I0(n1702), .I1(n1730), .CO(n28824));
    SB_LUT4 mod_5_add_1205_9_lut (.I0(n1703), .I1(n1703), .I2(n1730), 
            .I3(n28822), .O(n1802)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1205_9_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1205_9 (.CI(n28822), .I0(n1703), .I1(n1730), .CO(n28823));
    SB_LUT4 mod_5_add_1205_8_lut (.I0(n1704), .I1(n1704), .I2(n1730), 
            .I3(n28821), .O(n1803)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1205_8_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1205_8 (.CI(n28821), .I0(n1704), .I1(n1730), .CO(n28822));
    SB_LUT4 mod_5_add_1205_7_lut (.I0(n1705), .I1(n1705), .I2(n1730), 
            .I3(n28820), .O(n1804)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1205_7_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1205_7 (.CI(n28820), .I0(n1705), .I1(n1730), .CO(n28821));
    SB_LUT4 mod_5_add_1205_6_lut (.I0(n1706), .I1(n1706), .I2(n1730), 
            .I3(n28819), .O(n1805)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1205_6_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1205_6 (.CI(n28819), .I0(n1706), .I1(n1730), .CO(n28820));
    SB_LUT4 mod_5_add_1205_5_lut (.I0(n1707), .I1(n1707), .I2(n1730), 
            .I3(n28818), .O(n1806)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1205_5_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 add_21_27_lut (.I0(GND_net), .I1(bit_ctr[25]), .I2(GND_net), 
            .I3(n27788), .O(n255[25])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_27_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1205_5 (.CI(n28818), .I0(n1707), .I1(n1730), .CO(n28819));
    SB_LUT4 mod_5_add_1205_4_lut (.I0(n1708), .I1(n1708), .I2(n1730), 
            .I3(n28817), .O(n1807)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1205_4_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1205_4 (.CI(n28817), .I0(n1708), .I1(n1730), .CO(n28818));
    SB_LUT4 mod_5_add_1205_3_lut (.I0(n1709), .I1(n1709), .I2(n37643), 
            .I3(n28816), .O(n1808)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1205_3_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1205_3 (.CI(n28816), .I0(n1709), .I1(n37643), .CO(n28817));
    SB_LUT4 mod_5_add_1205_2_lut (.I0(bit_ctr[18]), .I1(bit_ctr[18]), .I2(n37643), 
            .I3(VCC_net), .O(n1809)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1205_2_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1205_2 (.CI(VCC_net), .I0(bit_ctr[18]), .I1(n37643), 
            .CO(n28816));
    SB_LUT4 mod_5_add_1272_16_lut (.I0(n1796), .I1(n1796), .I2(n1829), 
            .I3(n28815), .O(n1895)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_16_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1272_15_lut (.I0(n1797), .I1(n1797), .I2(n1829), 
            .I3(n28814), .O(n1896)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_15_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1272_15 (.CI(n28814), .I0(n1797), .I1(n1829), .CO(n28815));
    SB_LUT4 mod_5_add_1272_14_lut (.I0(n1798), .I1(n1798), .I2(n1829), 
            .I3(n28813), .O(n1897)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_14_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY add_21_27 (.CI(n27788), .I0(bit_ctr[25]), .I1(GND_net), .CO(n27789));
    SB_CARRY mod_5_add_1272_14 (.CI(n28813), .I0(n1798), .I1(n1829), .CO(n28814));
    SB_LUT4 mod_5_add_1272_13_lut (.I0(n1799), .I1(n1799), .I2(n1829), 
            .I3(n28812), .O(n1898)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_13_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1272_13 (.CI(n28812), .I0(n1799), .I1(n1829), .CO(n28813));
    SB_LUT4 mod_5_add_1272_12_lut (.I0(n1800), .I1(n1800), .I2(n1829), 
            .I3(n28811), .O(n1899)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_12_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1272_12 (.CI(n28811), .I0(n1800), .I1(n1829), .CO(n28812));
    SB_LUT4 mod_5_add_1272_11_lut (.I0(n1801), .I1(n1801), .I2(n1829), 
            .I3(n28810), .O(n1900)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_11_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1272_11 (.CI(n28810), .I0(n1801), .I1(n1829), .CO(n28811));
    SB_LUT4 mod_5_add_1272_10_lut (.I0(n1802), .I1(n1802), .I2(n1829), 
            .I3(n28809), .O(n1901)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_10_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1272_10 (.CI(n28809), .I0(n1802), .I1(n1829), .CO(n28810));
    SB_LUT4 mod_5_add_1272_9_lut (.I0(n1803), .I1(n1803), .I2(n1829), 
            .I3(n28808), .O(n1902)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_9_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1272_9 (.CI(n28808), .I0(n1803), .I1(n1829), .CO(n28809));
    SB_LUT4 mod_5_add_1272_8_lut (.I0(n1804), .I1(n1804), .I2(n1829), 
            .I3(n28807), .O(n1903)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_8_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1272_8 (.CI(n28807), .I0(n1804), .I1(n1829), .CO(n28808));
    SB_LUT4 mod_5_add_1272_7_lut (.I0(n1805), .I1(n1805), .I2(n1829), 
            .I3(n28806), .O(n1904)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_7_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1272_7 (.CI(n28806), .I0(n1805), .I1(n1829), .CO(n28807));
    SB_LUT4 mod_5_add_1272_6_lut (.I0(n1806), .I1(n1806), .I2(n1829), 
            .I3(n28805), .O(n1905)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_6_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1272_6 (.CI(n28805), .I0(n1806), .I1(n1829), .CO(n28806));
    SB_LUT4 mod_5_add_1272_5_lut (.I0(n1807), .I1(n1807), .I2(n1829), 
            .I3(n28804), .O(n1906)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_5_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1272_5 (.CI(n28804), .I0(n1807), .I1(n1829), .CO(n28805));
    SB_LUT4 add_21_26_lut (.I0(GND_net), .I1(bit_ctr[24]), .I2(GND_net), 
            .I3(n27787), .O(n255[24])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_26_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_1272_4_lut (.I0(n1808), .I1(n1808), .I2(n1829), 
            .I3(n28803), .O(n1907)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_4_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1272_4 (.CI(n28803), .I0(n1808), .I1(n1829), .CO(n28804));
    SB_LUT4 mod_5_add_1272_3_lut (.I0(n1809), .I1(n1809), .I2(n37644), 
            .I3(n28802), .O(n1908)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_3_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1272_3 (.CI(n28802), .I0(n1809), .I1(n37644), .CO(n28803));
    SB_LUT4 mod_5_add_1272_2_lut (.I0(bit_ctr[17]), .I1(bit_ctr[17]), .I2(n37644), 
            .I3(VCC_net), .O(n1909)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_2_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1272_2 (.CI(VCC_net), .I0(bit_ctr[17]), .I1(n37644), 
            .CO(n28802));
    SB_LUT4 i10_4_lut_adj_1606 (.I0(n2193), .I1(n2194), .I2(n2206), .I3(n2204), 
            .O(n28_adj_4865));
    defparam i10_4_lut_adj_1606.LUT_INIT = 16'hfffe;
    SB_LUT4 i14_4_lut_adj_1607 (.I0(n2203), .I1(n28_adj_4865), .I2(bit_ctr[13]), 
            .I3(n2209), .O(n32_adj_4866));
    defparam i14_4_lut_adj_1607.LUT_INIT = 16'hfeee;
    SB_LUT4 i12_4_lut_adj_1608 (.I0(n2208), .I1(n2201), .I2(n2192), .I3(n2196), 
            .O(n30_adj_4867));
    defparam i12_4_lut_adj_1608.LUT_INIT = 16'hfffe;
    SB_LUT4 i13_4_lut_adj_1609 (.I0(n2195), .I1(n2207), .I2(n2205), .I3(n2199), 
            .O(n31_adj_4868));
    defparam i13_4_lut_adj_1609.LUT_INIT = 16'hfffe;
    SB_LUT4 i11_4_lut_adj_1610 (.I0(n2202), .I1(n2197), .I2(n2198), .I3(n2200), 
            .O(n29_adj_4869));
    defparam i11_4_lut_adj_1610.LUT_INIT = 16'hfffe;
    SB_LUT4 i17_4_lut_adj_1611 (.I0(n29_adj_4869), .I1(n31_adj_4868), .I2(n30_adj_4867), 
            .I3(n32_adj_4866), .O(n2225));
    defparam i17_4_lut_adj_1611.LUT_INIT = 16'hfffe;
    SB_LUT4 mod_5_add_1339_17_lut (.I0(n1895), .I1(n1895), .I2(n1928), 
            .I3(n28801), .O(n1994)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_17_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i30876_1_lut (.I0(n2720), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n37629));
    defparam i30876_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mod_5_add_1339_16_lut (.I0(n1896), .I1(n1896), .I2(n1928), 
            .I3(n28800), .O(n1995)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_16_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1339_16 (.CI(n28800), .I0(n1896), .I1(n1928), .CO(n28801));
    SB_CARRY add_21_26 (.CI(n27787), .I0(bit_ctr[24]), .I1(GND_net), .CO(n27788));
    SB_LUT4 mod_5_add_1339_15_lut (.I0(n1897), .I1(n1897), .I2(n1928), 
            .I3(n28799), .O(n1996)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_15_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1339_15 (.CI(n28799), .I0(n1897), .I1(n1928), .CO(n28800));
    SB_LUT4 mod_5_add_1339_14_lut (.I0(n1898), .I1(n1898), .I2(n1928), 
            .I3(n28798), .O(n1997)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_14_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i30875_1_lut (.I0(n2126), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n37628));
    defparam i30875_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY mod_5_add_1339_14 (.CI(n28798), .I0(n1898), .I1(n1928), .CO(n28799));
    SB_LUT4 mod_5_add_1339_13_lut (.I0(n1899), .I1(n1899), .I2(n1928), 
            .I3(n28797), .O(n1998)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_13_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1339_13 (.CI(n28797), .I0(n1899), .I1(n1928), .CO(n28798));
    SB_LUT4 mod_5_add_1339_12_lut (.I0(n1900), .I1(n1900), .I2(n1928), 
            .I3(n28796), .O(n1999)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_12_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1339_12 (.CI(n28796), .I0(n1900), .I1(n1928), .CO(n28797));
    SB_LUT4 mod_5_add_1339_11_lut (.I0(n1901), .I1(n1901), .I2(n1928), 
            .I3(n28795), .O(n2000)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_11_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1339_11 (.CI(n28795), .I0(n1901), .I1(n1928), .CO(n28796));
    SB_LUT4 mod_5_add_1339_10_lut (.I0(n1902), .I1(n1902), .I2(n1928), 
            .I3(n28794), .O(n2001)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_10_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1339_10 (.CI(n28794), .I0(n1902), .I1(n1928), .CO(n28795));
    SB_LUT4 mod_5_add_1339_9_lut (.I0(n1903), .I1(n1903), .I2(n1928), 
            .I3(n28793), .O(n2002)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_9_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i5_2_lut (.I0(n2693), .I1(n2704), .I2(GND_net), .I3(GND_net), 
            .O(n28_adj_4870));
    defparam i5_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i15_4_lut_adj_1612 (.I0(n2699), .I1(n2706), .I2(n2694), .I3(n2691), 
            .O(n38_adj_4871));
    defparam i15_4_lut_adj_1612.LUT_INIT = 16'hfffe;
    SB_LUT4 i19494_2_lut (.I0(bit_ctr[8]), .I1(n2709), .I2(GND_net), .I3(GND_net), 
            .O(n24637));
    defparam i19494_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i13_4_lut_adj_1613 (.I0(n2701), .I1(n2696), .I2(n2697), .I3(n24637), 
            .O(n36_adj_4872));
    defparam i13_4_lut_adj_1613.LUT_INIT = 16'hfffe;
    SB_LUT4 i19_4_lut_adj_1614 (.I0(n2700), .I1(n38_adj_4871), .I2(n28_adj_4870), 
            .I3(n2705), .O(n42_adj_4873));
    defparam i19_4_lut_adj_1614.LUT_INIT = 16'hfffe;
    SB_LUT4 i17_4_lut_adj_1615 (.I0(n2702), .I1(n2690), .I2(n2689), .I3(n2708), 
            .O(n40_adj_4874));
    defparam i17_4_lut_adj_1615.LUT_INIT = 16'hfffe;
    SB_LUT4 i18_4_lut_adj_1616 (.I0(n2687), .I1(n36_adj_4872), .I2(n2703), 
            .I3(n2695), .O(n41_adj_4875));
    defparam i18_4_lut_adj_1616.LUT_INIT = 16'hfffe;
    SB_LUT4 i16_4_lut_adj_1617 (.I0(n2688), .I1(n2698), .I2(n2692), .I3(n2707), 
            .O(n39_adj_4876));
    defparam i16_4_lut_adj_1617.LUT_INIT = 16'hfffe;
    SB_LUT4 i22_4_lut_adj_1618 (.I0(n39_adj_4876), .I1(n41_adj_4875), .I2(n40_adj_4874), 
            .I3(n42_adj_4873), .O(n2720));
    defparam i22_4_lut_adj_1618.LUT_INIT = 16'hfffe;
    SB_LUT4 i30874_1_lut (.I0(n1334), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n37627));
    defparam i30874_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i3_4_lut (.I0(n24613), .I1(\state[1] ), .I2(n17393), .I3(n33377), 
            .O(n34121));
    defparam i3_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i2_4_lut_adj_1619 (.I0(\state[1] ), .I1(n34121), .I2(start), 
            .I3(n35064), .O(n34265));
    defparam i2_4_lut_adj_1619.LUT_INIT = 16'h8c00;
    SB_LUT4 bit_ctr_2__bdd_4_lut (.I0(bit_ctr[2]), .I1(n35482), .I2(n35485), 
            .I3(n30003), .O(n37664));
    defparam bit_ctr_2__bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_LUT4 n37664_bdd_4_lut (.I0(n37664), .I1(n36892), .I2(n35491), .I3(n30003), 
            .O(n37667));
    defparam n37664_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 sub_14_inv_0_i11_1_lut (.I0(\neo_pixel_transmitter.t0 [10]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[10]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i11_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i3_4_lut_adj_1620 (.I0(n31_adj_4817), .I1(n23_adj_4821), .I2(n55), 
            .I3(n39_adj_4813), .O(n34867));
    defparam i3_4_lut_adj_1620.LUT_INIT = 16'hfffe;
    SB_LUT4 i12_4_lut_adj_1621 (.I0(n25_adj_4820), .I1(n63), .I2(n27_adj_4819), 
            .I3(n11_adj_4827), .O(n28_adj_4877));
    defparam i12_4_lut_adj_1621.LUT_INIT = 16'hfffe;
    SB_LUT4 i10_4_lut_adj_1622 (.I0(n29_adj_4818), .I1(n61), .I2(n35_adj_4815), 
            .I3(n51_adj_4804), .O(n26_adj_4878));
    defparam i10_4_lut_adj_1622.LUT_INIT = 16'hfffe;
    SB_LUT4 i11_4_lut_adj_1623 (.I0(n59), .I1(n43_adj_4808), .I2(n47_adj_4806), 
            .I3(n57), .O(n27_adj_4879));
    defparam i11_4_lut_adj_1623.LUT_INIT = 16'hfffe;
    SB_LUT4 i9_4_lut_adj_1624 (.I0(n49_adj_4805), .I1(n15_adj_4825), .I2(n41), 
            .I3(n33_adj_4816), .O(n25_adj_4880));
    defparam i9_4_lut_adj_1624.LUT_INIT = 16'hfffe;
    SB_LUT4 i5_4_lut_adj_1625 (.I0(n45_adj_4807), .I1(n34867), .I2(bit_ctr[3]), 
            .I3(n3209), .O(n14_adj_4881));
    defparam i5_4_lut_adj_1625.LUT_INIT = 16'hfeee;
    SB_LUT4 i4_2_lut (.I0(n13_adj_4826), .I1(n19_adj_4823), .I2(GND_net), 
            .I3(GND_net), .O(n13_adj_4882));
    defparam i4_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i15_4_lut_adj_1626 (.I0(n25_adj_4880), .I1(n27_adj_4879), .I2(n26_adj_4878), 
            .I3(n28_adj_4877), .O(n35175));
    defparam i15_4_lut_adj_1626.LUT_INIT = 16'hfffe;
    SB_LUT4 i6_4_lut_adj_1627 (.I0(n17_adj_4824), .I1(n53), .I2(n37_adj_4814), 
            .I3(n21_adj_4822), .O(n15_adj_4883));
    defparam i6_4_lut_adj_1627.LUT_INIT = 16'hfffe;
    SB_LUT4 i27_4_lut (.I0(n15_adj_4883), .I1(n35175), .I2(n13_adj_4882), 
            .I3(n14_adj_4881), .O(n29627));
    defparam i27_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i19516_3_lut (.I0(one_wire_N_553[9]), .I1(one_wire_N_553[11]), 
            .I2(one_wire_N_553[10]), .I3(GND_net), .O(n24659));
    defparam i19516_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i284_2_lut (.I0(n24759), .I1(\neo_pixel_transmitter.done ), 
            .I2(GND_net), .I3(GND_net), .O(n1265));   // verilog/neopixel.v(103[9] 111[12])
    defparam i284_2_lut.LUT_INIT = 16'hdddd;
    SB_LUT4 i26638_4_lut (.I0(n17393), .I1(n29522), .I2(n33371), .I3(\state[0] ), 
            .O(n14));   // verilog/neopixel.v(35[12] 117[6])
    defparam i26638_4_lut.LUT_INIT = 16'hfaee;
    SB_LUT4 i15_4_lut_adj_1628 (.I0(n14), .I1(n36222), .I2(\state[1] ), 
            .I3(n17509), .O(n33425));   // verilog/neopixel.v(35[12] 117[6])
    defparam i15_4_lut_adj_1628.LUT_INIT = 16'h303a;
    SB_LUT4 i1_4_lut_adj_1629 (.I0(\state[0] ), .I1(n33365), .I2(n1265), 
            .I3(\state[1] ), .O(n18685));
    defparam i1_4_lut_adj_1629.LUT_INIT = 16'hafcc;
    SB_LUT4 mod_5_i2239_3_lut (.I0(n3209), .I1(bit_ctr[3]), .I2(n29627), 
            .I3(GND_net), .O(color_bit_N_596[4]));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i2239_3_lut.LUT_INIT = 16'h6a6a;
    SB_LUT4 i30040_4_lut (.I0(n37883), .I1(n30003), .I2(n37745), .I3(bit_ctr[2]), 
            .O(n36249));
    defparam i30040_4_lut.LUT_INIT = 16'h3022;
    SB_LUT4 i18599_4_lut (.I0(n37667), .I1(\state_3__N_402[1] ), .I2(n36249), 
            .I3(color_bit_N_596[4]), .O(state_3__N_402[0]));   // verilog/neopixel.v(40[18] 45[12])
    defparam i18599_4_lut.LUT_INIT = 16'h3022;
    SB_LUT4 sub_14_inv_0_i12_1_lut (.I0(\neo_pixel_transmitter.t0 [11]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[11]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i12_1_lut.LUT_INIT = 16'h5555;
    
endmodule
//
// Verilog Description of module pll32MHz
//

module pll32MHz (GND_net, CLK_c, VCC_net, clk32MHz) /* synthesis syn_module_defined=1 */ ;
    input GND_net;
    input CLK_c;
    input VCC_net;
    output clk32MHz;
    
    wire CLK_c /* synthesis SET_AS_NETWORK=CLK_c, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(3[9:12])
    wire clk32MHz /* synthesis SET_AS_NETWORK=clk32MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(33[6:14])
    
    SB_PLL40_CORE pll32MHz_inst (.REFERENCECLK(CLK_c), .PLLOUTGLOBAL(clk32MHz), 
            .BYPASS(GND_net), .RESETB(VCC_net)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=51, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=34, LSE_RLINE=37 */ ;   // verilog/TinyFPGA_B.v(34[10] 37[2])
    defparam pll32MHz_inst.FEEDBACK_PATH = "PHASE_AND_DELAY";
    defparam pll32MHz_inst.DELAY_ADJUSTMENT_MODE_FEEDBACK = "FIXED";
    defparam pll32MHz_inst.DELAY_ADJUSTMENT_MODE_RELATIVE = "FIXED";
    defparam pll32MHz_inst.SHIFTREG_DIV_MODE = 2'b00;
    defparam pll32MHz_inst.FDA_FEEDBACK = 4'b0000;
    defparam pll32MHz_inst.FDA_RELATIVE = 4'b0000;
    defparam pll32MHz_inst.PLLOUT_SELECT = "SHIFTREG_0deg";
    defparam pll32MHz_inst.DIVR = 4'b0000;
    defparam pll32MHz_inst.DIVF = 7'b0000001;
    defparam pll32MHz_inst.DIVQ = 3'b011;
    defparam pll32MHz_inst.FILTER_RANGE = 3'b001;
    defparam pll32MHz_inst.ENABLE_ICEGATE = 1'b0;
    defparam pll32MHz_inst.TEST_MODE = 1'b0;
    defparam pll32MHz_inst.EXTERNAL_DIVIDE_FACTOR = 1;
    
endmodule
//
// Verilog Description of module motorControl
//

module motorControl (GND_net, \Kp[2] , \Kp[3] , \Ki[0] , \Kp[0] , 
            \Kp[4] , \Kp[5] , \Kp[6] , \Kp[7] , \Kp[8] , \Kp[9] , 
            \Kp[10] , \Kp[11] , \Kp[12] , \Kp[13] , \Kp[14] , \Kp[15] , 
            \Kp[1] , PWMLimit, IntegralLimit, \Ki[1] , \Ki[2] , \Ki[3] , 
            \Ki[4] , \Ki[5] , \Ki[6] , \Ki[7] , \Ki[8] , \Ki[9] , 
            \Ki[10] , \Ki[11] , duty, clk32MHz, \Ki[12] , \Ki[13] , 
            \Ki[14] , \Ki[15] , VCC_net, setpoint, motor_state, n37633) /* synthesis syn_module_defined=1 */ ;
    input GND_net;
    input \Kp[2] ;
    input \Kp[3] ;
    input \Ki[0] ;
    input \Kp[0] ;
    input \Kp[4] ;
    input \Kp[5] ;
    input \Kp[6] ;
    input \Kp[7] ;
    input \Kp[8] ;
    input \Kp[9] ;
    input \Kp[10] ;
    input \Kp[11] ;
    input \Kp[12] ;
    input \Kp[13] ;
    input \Kp[14] ;
    input \Kp[15] ;
    input \Kp[1] ;
    input [23:0]PWMLimit;
    input [23:0]IntegralLimit;
    input \Ki[1] ;
    input \Ki[2] ;
    input \Ki[3] ;
    input \Ki[4] ;
    input \Ki[5] ;
    input \Ki[6] ;
    input \Ki[7] ;
    input \Ki[8] ;
    input \Ki[9] ;
    input \Ki[10] ;
    input \Ki[11] ;
    output [23:0]duty;
    input clk32MHz;
    input \Ki[12] ;
    input \Ki[13] ;
    input \Ki[14] ;
    input \Ki[15] ;
    input VCC_net;
    input [23:0]setpoint;
    input [23:0]motor_state;
    output n37633;
    
    wire clk32MHz /* synthesis SET_AS_NETWORK=clk32MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(33[6:14])
    
    wire n45;
    wire [23:0]n1;
    
    wire n28025;
    wire [23:0]\PID_CONTROLLER.integral ;   // verilog/motorControl.v(23[23:31])
    wire [23:0]duty_23__N_3646;
    wire [47:0]n106;
    wire [47:0]n155;
    
    wire n27868, n28026, n27869, n43, n28024;
    wire [23:0]n28;
    
    wire n162, n235;
    wire [23:0]\PID_CONTROLLER.integral_23__N_3546 ;
    
    wire \PID_CONTROLLER.integral_23__N_3594 ;
    wire [23:0]n3302;
    
    wire n308, n381, n454, n527, n600, n673, n746, n819, n892, 
        n965, n1038, n1111, n92, n23, n165, n238, n311, n384, 
        n457, n530, n603, n676, n749, n822, n895, n968, n1041, 
        n1114, n95, n26_adj_4313, n168, n241, n314, n387, n460, 
        n533, n606, n679, n752, n825, n898, n971, n1044, n1117, 
        n98, n29, n41, n28023;
    wire [23:0]n257;
    
    wire n256;
    wire [23:0]duty_23__N_3621;
    
    wire duty_23__N_3645;
    wire [23:0]duty_23__N_3522;
    
    wire n27867, n171, n244, n317, n390, n463, n536, n609, n682, 
        n755, n828, n901, n974, n1047, n1120, n101, n32, n174, 
        n247, n320, n393, n466, n539, n612, n685, n758, n17_adj_4317, 
        n9, n11, n831, n36526, n904, n36523, n977, n38414, n36890, 
        n1050, n36771, n38396, n36769, n104, n36767, n38390, n27, 
        n15, n13, n11_adj_4318, n36463, n21_adj_4319, n19_adj_4320, 
        n17_adj_4321, n9_adj_4322, n36469, n35, n16_adj_4324, n177, 
        n250, n323, n36444, n396, n8, n24_adj_4325, n469, n7_adj_4326, 
        n5_adj_4327, n36479, n36738, n36734, n25_adj_4328, n23_adj_4329, 
        n37006, n542, n615, n688, n761, n834, n31, n29_adj_4330, 
        n36858, n907, n37, n35_adj_4331, n33, n37065, n36773, 
        n38383, n36761, n980, n38378, n12, n36498, n38401, n10, 
        n30, n36956, n107, n38, n36506, n180, n38381, n36884, 
        n38407, n37042, n38372, n37097, n38369, n16_adj_4332, n36482, 
        n253, n24_adj_4333, n326, n6_adj_4334, n36898, n36899, n36484, 
        n399, n8_adj_4335, n38367, n36868, n36749;
    wire [23:0]\PID_CONTROLLER.integral_23__N_3597 ;
    
    wire n3_adj_4336, n4_adj_4337, n37000, n472, n37001, n12_adj_4338, 
        n36457, n10_adj_4339, n30_adj_4340, n36459, n545, n37071, 
        n36927, n618, n37120, n37121, n39, n37106, n6_adj_4341, 
        n37008, n37009, n691, n36446, n36872, n764, n36925, n36449, 
        n37022, n40, n37024, n4_adj_4342, n36896, n36897, n837, 
        n36500, n37069, n910, n36751, n37107, n37108, n110, n41_adj_4344, 
        n37080, n36487, n183, n37016, n37015, \PID_CONTROLLER.integral_23__N_3596 , 
        n37018, n256_adj_4345, n329, n402, n475, n548, n621, n694, 
        n767, n840, n113, n44, n186, n259_adj_4347, n332, n405, 
        n478, n551, n624, n697, n770, n116, n47, n189_adj_4349, 
        n262_adj_4350, n335, n408, n481, n554, n627, n700, n119, 
        n50, n192, n265_adj_4357, n338, n411, n484, n557, n630, 
        n122, n53, n195, n268_adj_4361, n341, n414, n487, n560, 
        n125, n56, n198, n271_adj_4371, n344, n417, n6_adj_4372;
    wire [3:0]n10026;
    wire [4:0]n10019;
    wire [1:0]n10037;
    
    wire n4_adj_4374;
    wire [2:0]n10032;
    
    wire n490, n12_adj_4375, n8_adj_4376, n11_adj_4377, n6_adj_4378, 
        n27573, n18_adj_4379, n13_adj_4380, n4_adj_4381, n34086, n77, 
        n8_adj_4382, n150, n223, n296, n369, n442, n515, n588, 
        n661, n734, n807, n880, n953, n1026, n1099;
    wire [23:0]n1_adj_4735;
    
    wire n28022, n74, n5_adj_4388, n147, n220, n293, n366, n439, 
        n512, n585, n658, n731, n804, n877, n950, n1023, n1096, 
        n80, n11_adj_4390, n153, n226, n299, n372, n445, n518, 
        n591, n664, n737, n810, n883, n956, n1029, n1102, n27866, 
        n28021, n83, n27865, n14_adj_4396, n156, n229, n302, n375, 
        n28020, n448, n521, n594, n667, n740, n813, n886, n959, 
        n1032, n1105, n86, n17_adj_4400, n77_adj_4402, n8_adj_4404, 
        n150_adj_4405, n223_adj_4407, n296_adj_4408, n159, n232, n305, 
        n378, n451, n524, n369_adj_4409, n597, n670, n442_adj_4410, 
        n743, n515_adj_4411, n816, n889, n962, n588_adj_4412, n1035, 
        n1108, n661_adj_4413, n734_adj_4414, n89, n20_adj_4415, n162_adj_4416, 
        n807_adj_4417, n235_adj_4418, n308_adj_4419, n381_adj_4420, 
        n454_adj_4421, n527_adj_4422, n880_adj_4423, n27864, n600_adj_4424, 
        n673_adj_4425, n953_adj_4426, n746_adj_4427, n27548, n819_adj_4428, 
        n892_adj_4429, n28019, n965_adj_4430, n1038_adj_4431, n1111_adj_4432, 
        n1026_adj_4433, n92_adj_4434, n23_adj_4435, n165_adj_4436, n238_adj_4437, 
        n1099_adj_4438, n27863, n28018, n28017, n311_adj_4439, n28016, 
        n28015, n27862, n27861, n28014, n384_adj_4442, n27514, n457_adj_4443, 
        n28013, n27860, n28012, n27859, n28011, n28010, n27858, 
        n28009, n28008, n4_adj_4446, n530_adj_4447, n27857, n603_adj_4448, 
        n28007, n676_adj_4449, n749_adj_4450, n28006, n27920, n28005, 
        n822_adj_4451, n895_adj_4452, n968_adj_4453, n1041_adj_4454, 
        n1114_adj_4455, n95_adj_4456, n26_adj_4457, n74_adj_4458, n168_adj_4459, 
        n27856, n5_adj_4460, n241_adj_4461, n27919, n314_adj_4462, 
        n28004, n387_adj_4463, n27471, n460_adj_4464, n533_adj_4465, 
        n606_adj_4466, n27855, n679_adj_4468, n147_adj_4469, n752_adj_4470, 
        n825_adj_4471, n27918, n220_adj_4472, n898_adj_4473, n971_adj_4474, 
        n27917, n293_adj_4475, n1044_adj_4476, n1117_adj_4477, n366_adj_4478, 
        n98_adj_4479, n29_adj_4480, n171_adj_4481, n244_adj_4482, n439_adj_4483, 
        n317_adj_4484, n390_adj_4485, n463_adj_4486, n536_adj_4487, 
        n609_adj_4488, n512_adj_4489, n585_adj_4490, n658_adj_4491, 
        n27916, n682_adj_4492, n731_adj_4493, n755_adj_4494, n828_adj_4495, 
        n901_adj_4496, n974_adj_4497, n1047_adj_4498, n804_adj_4499, 
        n877_adj_4500, n1120_adj_4501, n101_adj_4502, n950_adj_4503, 
        n32_adj_4504, n174_adj_4505, n247_adj_4506, n320_adj_4507, n393_adj_4508, 
        n466_adj_4509, n539_adj_4510, n612_adj_4511, n685_adj_4512, 
        n27998, n1023_adj_4513, n27997, n758_adj_4514, n831_adj_4515, 
        n904_adj_4516, n977_adj_4517, n1096_adj_4518, n1050_adj_4519, 
        n104_adj_4520, n35_adj_4521, n27915, n27914, n177_adj_4522, 
        n27996, n27995, n27913, n27994, n250_adj_4523, n323_adj_4524, 
        n27993, n27992, n27912, n27991, n396_adj_4525, n469_adj_4526, 
        n542_adj_4527, n615_adj_4528, n688_adj_4529, n27990, n761_adj_4531, 
        n27911, n834_adj_4532, n27989, n27910, n27909, n27988, n27908, 
        n27987, n27986, n27985, n80_adj_4533, n11_adj_4535;
    wire [5:0]n10308;
    
    wire n34185, n490_adj_4536, n29353;
    wire [4:0]n10316;
    
    wire n417_adj_4537, n29352, n344_adj_4538, n29351, n271_adj_4539, 
        n29350, n198_adj_4540, n29349, n56_adj_4541, n125_adj_4542;
    wire [6:0]n10299;
    
    wire n560_adj_4543, n29348, n487_adj_4544, n29347, n414_adj_4545, 
        n29346, n341_adj_4546, n29345, n268_adj_4547, n29344, n195_adj_4548, 
        n29343, n53_adj_4549, n122_adj_4550;
    wire [7:0]n10289;
    
    wire n630_adj_4551, n29342, n557_adj_4552, n29341, n484_adj_4553, 
        n29340, n411_adj_4554, n29339, n153_adj_4555, n338_adj_4556, 
        n29338, n27907, n265_adj_4557, n29337, n192_adj_4558, n29336, 
        n27984, n50_adj_4559, n119_adj_4560;
    wire [8:0]n10278;
    
    wire n700_adj_4561, n29335, n27906, n627_adj_4562, n29334, n554_adj_4563, 
        n29333, n481_adj_4564, n29332, n27983, n27982, n226_adj_4565, 
        n408_adj_4566, n29331, n299_adj_4567, n335_adj_4568, n29330, 
        n262_adj_4569, n29329, n372_adj_4570, n445_adj_4571, n189_adj_4572, 
        n29328, n518_adj_4573, n591_adj_4574, n27905, n664_adj_4575, 
        n47_adj_4576, n116_adj_4577, n27904, n737_adj_4578, n810_adj_4579, 
        n27981;
    wire [9:0]n10266;
    
    wire n770_adj_4580, n29327, n697_adj_4581, n29326, n624_adj_4582, 
        n29325, n883_adj_4583, n551_adj_4584, n29324, n478_adj_4585, 
        n29323, n405_adj_4586, n29322, n332_adj_4587, n29321, n259_adj_4588, 
        n29320, n186_adj_4589, n29319, n956_adj_4590, n44_adj_4591, 
        n113_adj_4592;
    wire [10:0]n10253;
    
    wire n840_adj_4593, n29318, n767_adj_4594, n29317, n694_adj_4595, 
        n29316, n621_adj_4596, n29315, n548_adj_4597, n29314, n475_adj_4598, 
        n29313, n402_adj_4599, n29312, n329_adj_4600, n29311, n256_adj_4601, 
        n29310, n183_adj_4602, n29309, n41_adj_4603, n110_adj_4604;
    wire [11:0]n10239;
    
    wire n910_adj_4605, n29308, n837_adj_4606, n29307, n764_adj_4607, 
        n29306, n691_adj_4608, n29305, n618_adj_4609, n29304, n1029_adj_4610, 
        n545_adj_4611, n29303, n472_adj_4612, n29302, n27903, n1102_adj_4613, 
        n27980, n399_adj_4614, n29301, n326_adj_4615, n29300, n27979, 
        n27902, n27978, n253_adj_4617, n29299, n27977, n27901, n180_adj_4618, 
        n29298, n38_adj_4619, n107_adj_4620;
    wire [12:0]n10224;
    
    wire n980_adj_4621, n29297, n907_adj_4622, n29296, n27976, n27900, 
        n39_adj_4623, n41_adj_4624, n45_adj_4625, n37_adj_4626, n29_adj_4627, 
        n31_adj_4628, n43_adj_4629, n23_adj_4630, n25_adj_4631, n35_adj_4632, 
        n11_adj_4633, n13_adj_4634, n15_adj_4635, n27_adj_4636, n33_adj_4637, 
        n9_adj_4638, n17_adj_4639, n19_adj_4640, n21_adj_4641, n36432, 
        n36426, n12_adj_4642, n10_adj_4643, n30_adj_4644, n29295, 
        n36442, n36706, n36702, n36998, n29294, n36842, n37063, 
        n16_adj_4645, n29293, n6_adj_4646, n36984, n36985, n8_adj_4647, 
        n29292, n24_adj_4648, n36412, n36410, n36874, n36931, n29291, 
        n4_adj_4649, n36976, n36977, n36422, n29290, n36420, n37073, 
        n36933, n37122, n37123, n29289, n37104, n36414, n37028, 
        n40_adj_4650, n29288, n37030, n29287, n41_adj_4651, n39_adj_4652, 
        n29286, n45_adj_4653, n43_adj_4654, n37_adj_4655;
    wire [13:0]n10208;
    
    wire n29285, n29284, n29_adj_4656, n31_adj_4657, n29283, n23_adj_4658, 
        n25_adj_4659, n29282, n35_adj_4660, n29281, n33_adj_4661, 
        n11_adj_4662, n29280, n13_adj_4663, n29279, n15_adj_4664, 
        n27_adj_4665, n9_adj_4666, n17_adj_4667, n19_adj_4668, n21_adj_4669, 
        n36398, n36392, n12_adj_4670, n10_adj_4671, n29278, n30_adj_4672, 
        n36408, n36674, n36670, n36990, n36826, n37061, n16_adj_4673, 
        n6_adj_4674, n36972, n36973, n29277, n8_adj_4675, n24_adj_4676, 
        n36375, n29276, n29275, n29274, n29273, n36373, n36876, 
        n36937, n4_adj_4677, n36970, n36971, n36387, n36385, n37075, 
        n36939, n37124, n37125, n37102, n36377, n37034, n40_adj_4678, 
        n37036;
    wire [14:0]n10191;
    
    wire n29272, n29271, n29270, n29269, n29268, n29267, n29266, 
        n29265, n29264, n29263, n29262, n29261, n27899, n29260, 
        n27898, n29259;
    wire [15:0]n10173;
    
    wire n29258, n29257, n29256, n29255, n29254, n29253, n29252, 
        n29251, n29250, n29249, n29248, n29247, n29246, n29245, 
        n29244;
    wire [16:0]n10154;
    
    wire n29243, n29242, n29241, n29240, n29239, n29238, n29237, 
        n29236, n29235, n29234, n29233, n29232, n29231, n29230, 
        n29229, n29228;
    wire [17:0]n10134;
    
    wire n29227, n29226, n29225, n29224, n29223, n29222, n29221, 
        n29220, n29219, n29218, n29217, n29216, n29215, n29214, 
        n29213, n29212, n29211;
    wire [18:0]n10113;
    
    wire n29210, n29209, n29208, n29207, n83_adj_4679, n29206, n29205, 
        n14_adj_4680, n29204, n29203, n29202, n156_adj_4681, n29201, 
        n29200, n29199, n29198, n29197, n229_adj_4682, n29196, n29195, 
        n29194, n29193, n302_adj_4684;
    wire [19:0]n10091;
    
    wire n29192, n29191, n29190, n29189, n375_adj_4685, n29188, 
        n29187, n29186, n29185, n29184, n29183, n29182, n29181, 
        n29180, n29179, n29178, n29177, n29176, n29175, n29174;
    wire [20:0]n10068;
    
    wire n29173, n29172, n29171, n29170, n29169, n29168, n29167, 
        n29166, n29165, n29164, n29163, n29162, n29161, n29160, 
        n29159, n29158, n29157, n29156, n29155, n29154;
    wire [0:0]n8179;
    wire [21:0]n10044;
    
    wire n29153, n29152, n29151, n29150, n29149, n29148, n29147, 
        n29146, n29145, n29144, n29143, n29142, n29141, n29140, 
        n29139, n29138, n29137, n29136, n29135, n29134, n29133, 
        n29132, n29131, n29130, n29129, n29128, n29127, n29126, 
        n29125, n29124, n29123, n29122, n29121, n29120, n29119, 
        n29118, n29117, n29116, n29115, n29114, n29113, n29112, 
        n29111;
    wire [5:0]n10011;
    
    wire n29110, n29109, n29108, n29107, n29106;
    wire [6:0]n10002;
    
    wire n29105, n29104, n29103, n29102, n29101, n29100;
    wire [7:0]n9992;
    
    wire n29099, n29098, n29097, n29096, n29095, n29094, n29093;
    wire [8:0]n9981;
    
    wire n29092, n29091, n29090, n29089, n29088, n29087, n29086, 
        n29085;
    wire [9:0]n9969;
    
    wire n29084, n29083, n29082, n29081, n29080, n29079, n29078, 
        n29077, n29076;
    wire [10:0]n9956;
    
    wire n29075, n29074, n29073, n29072, n29071, n29070, n29069, 
        n29068, n29067, n29066;
    wire [11:0]n9942;
    
    wire n29065, n29064, n29063, n29062, n29061, n29060, n29059, 
        n29058, n29057, n29056, n29055;
    wire [12:0]n9927;
    
    wire n29054, n29053, n29052, n29051, n29050, n29049, n29048, 
        n29047, n29046, n29045, n29044, n29043;
    wire [13:0]n9911;
    
    wire n29042, n29041, n29040, n29039, n29038, n29037, n29036, 
        n29035, n29034, n29033, n29032, n29031, n29030;
    wire [14:0]n9894;
    
    wire n29029, n29028, n29027, n29026, n29025, n29024, n29023, 
        n29022, n29021, n29020, n29019, n29018, n448_adj_4688, n29017, 
        n29016, n521_adj_4689;
    wire [15:0]n9876;
    
    wire n29015, n29014, n29013, n29012, n29011, n29010, n594_adj_4690, 
        n29009, n29008, n29007, n667_adj_4691, n29006, n29005, n29004, 
        n29003, n29002, n29001;
    wire [16:0]n9857;
    
    wire n29000, n28999, n28998, n28997, n28996, n28995, n28994, 
        n28993, n28992, n28991, n28990, n28989, n28988, n28987, 
        n28986, n28985;
    wire [17:0]n9837;
    
    wire n28984, n28983, n28982, n28981, n28980, n28979, n28978, 
        n28977, n28976, n28975, n28974, n28973, n28972, n28971, 
        n28970, n740_adj_4692, n813_adj_4693, n886_adj_4695, n959_adj_4696, 
        n1032_adj_4698, n1105_adj_4699, n86_adj_4700, n17_adj_4701, 
        n159_adj_4703, n28969, n28968, n20_adj_4707, n89_adj_4708;
    wire [18:0]n9816;
    
    wire n28967, n28966, n28965, n28964, n1108_adj_4709, n28963, 
        n1035_adj_4710, n28962, n962_adj_4711, n28961, n889_adj_4712, 
        n28960, n816_adj_4713, n28959, n743_adj_4714, n28958, n670_adj_4715, 
        n28957, n597_adj_4716, n28956, n232_adj_4717, n305_adj_4721, 
        n27680;
    wire [1:0]n10334;
    
    wire n4_adj_4722;
    wire [2:0]n10329;
    
    wire n524_adj_4723, n28955, n451_adj_4724, n28954, n27646, n4_adj_4725;
    wire [3:0]n10323;
    
    wire n378_adj_4726, n28953, n4_adj_4727, n6_adj_4728, n28952, 
        n27603, n28049, n28048, n28047, n28951, n28046, n28045, 
        n28044, n28950, n28043;
    wire [19:0]n9794;
    
    wire n28949, n28948, n28947, n28946, n28945, n28944, n28943, 
        n28042, n28942, n28941, n28041, n28940, n28939, n28938, 
        n28937, n28936, n28935, n28934, n28933, n28040, n28932, 
        n28931;
    wire [20:0]n9771;
    
    wire n28930, n28929, n28928, n28927, n28926, n28925, n28924, 
        n28923, n28922, n28921, n28920, n28919, n28918, n28917, 
        n28916, n28915, n28914, n28913, n28912, n28911;
    wire [0:0]n8175;
    wire [21:0]n9747;
    
    wire n28910, n28909, n28908, n28907, n28906, n28905, n28904, 
        n28039, n28903, n28902, n28901, n28900, n28899, n28898, 
        n28897, n28896, n28895, n28894, n28893, n28892, n28891, 
        n28890, n28889, n28888, n28887, n28886, n28885, n28884, 
        n28883, n28882, n28881, n28880, n28879, n28878, n28877, 
        n28876, n28875, n28874, n28873, n28872, n28871, n28870, 
        n27877, n28869, n28038, n28868, n28037, n27876, n28036, 
        n28035, n28034, n27875, n28033, n28032, n27874, n28031, 
        n28030, n27873, n27872, n27871, n28029, n28028, n27870, 
        n28027, n12_adj_4729, n8_adj_4730, n11_adj_4731, n6_adj_4732, 
        n27705, n18_adj_4733, n13_adj_4734;
    
    SB_LUT4 unary_minus_5_add_3_24_lut (.I0(\PID_CONTROLLER.integral [22]), 
            .I1(GND_net), .I2(n1[22]), .I3(n28025), .O(n45)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_24_lut.LUT_INIT = 16'h6996;
    SB_LUT4 add_12_16_lut (.I0(GND_net), .I1(n106[14]), .I2(n155[14]), 
            .I3(n27868), .O(duty_23__N_3646[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_5_add_3_24 (.CI(n28025), .I0(GND_net), .I1(n1[22]), 
            .CO(n28026));
    SB_CARRY add_12_16 (.CI(n27868), .I0(n106[14]), .I1(n155[14]), .CO(n27869));
    SB_LUT4 unary_minus_5_add_3_23_lut (.I0(\PID_CONTROLLER.integral [21]), 
            .I1(GND_net), .I2(n1[21]), .I3(n28024), .O(n43)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_23_lut.LUT_INIT = 16'h6996;
    SB_LUT4 mult_10_i110_2_lut (.I0(\Kp[2] ), .I1(n28[5]), .I2(GND_net), 
            .I3(GND_net), .O(n162));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i110_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i159_2_lut (.I0(\Kp[3] ), .I1(n28[5]), .I2(GND_net), 
            .I3(GND_net), .O(n235));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i159_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i2_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3546 [0]), 
            .I2(GND_net), .I3(GND_net), .O(n155[0]));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i2_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i2_2_lut (.I0(\Kp[0] ), .I1(n28[0]), .I2(GND_net), 
            .I3(GND_net), .O(n106[0]));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i2_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i19147_2_lut (.I0(n28[19]), .I1(\PID_CONTROLLER.integral_23__N_3594 ), 
            .I2(GND_net), .I3(GND_net), .O(n3302[19]));   // verilog/motorControl.v(31[7] 33[10])
    defparam i19147_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i19148_2_lut (.I0(n28[20]), .I1(\PID_CONTROLLER.integral_23__N_3594 ), 
            .I2(GND_net), .I3(GND_net), .O(n3302[20]));   // verilog/motorControl.v(31[7] 33[10])
    defparam i19148_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i19149_2_lut (.I0(n28[21]), .I1(\PID_CONTROLLER.integral_23__N_3594 ), 
            .I2(GND_net), .I3(GND_net), .O(n3302[21]));   // verilog/motorControl.v(31[7] 33[10])
    defparam i19149_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i208_2_lut (.I0(\Kp[4] ), .I1(n28[5]), .I2(GND_net), 
            .I3(GND_net), .O(n308));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i208_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i257_2_lut (.I0(\Kp[5] ), .I1(n28[5]), .I2(GND_net), 
            .I3(GND_net), .O(n381));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i257_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i306_2_lut (.I0(\Kp[6] ), .I1(n28[5]), .I2(GND_net), 
            .I3(GND_net), .O(n454));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i306_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i355_2_lut (.I0(\Kp[7] ), .I1(n28[5]), .I2(GND_net), 
            .I3(GND_net), .O(n527));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i355_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i404_2_lut (.I0(\Kp[8] ), .I1(n28[5]), .I2(GND_net), 
            .I3(GND_net), .O(n600));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i404_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i453_2_lut (.I0(\Kp[9] ), .I1(n28[5]), .I2(GND_net), 
            .I3(GND_net), .O(n673));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i453_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i502_2_lut (.I0(\Kp[10] ), .I1(n28[5]), .I2(GND_net), 
            .I3(GND_net), .O(n746));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i502_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i551_2_lut (.I0(\Kp[11] ), .I1(n28[5]), .I2(GND_net), 
            .I3(GND_net), .O(n819));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i551_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i600_2_lut (.I0(\Kp[12] ), .I1(n28[5]), .I2(GND_net), 
            .I3(GND_net), .O(n892));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i600_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i649_2_lut (.I0(\Kp[13] ), .I1(n28[5]), .I2(GND_net), 
            .I3(GND_net), .O(n965));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i649_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i698_2_lut (.I0(\Kp[14] ), .I1(n28[5]), .I2(GND_net), 
            .I3(GND_net), .O(n1038));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i698_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i747_2_lut (.I0(\Kp[15] ), .I1(n28[5]), .I2(GND_net), 
            .I3(GND_net), .O(n1111));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i747_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i63_2_lut (.I0(\Kp[1] ), .I1(n28[6]), .I2(GND_net), 
            .I3(GND_net), .O(n92));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i63_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i16_2_lut (.I0(\Kp[0] ), .I1(n28[7]), .I2(GND_net), 
            .I3(GND_net), .O(n23));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i16_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i112_2_lut (.I0(\Kp[2] ), .I1(n28[6]), .I2(GND_net), 
            .I3(GND_net), .O(n165));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i112_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i161_2_lut (.I0(\Kp[3] ), .I1(n28[6]), .I2(GND_net), 
            .I3(GND_net), .O(n238));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i161_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i210_2_lut (.I0(\Kp[4] ), .I1(n28[6]), .I2(GND_net), 
            .I3(GND_net), .O(n311));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i210_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i259_2_lut (.I0(\Kp[5] ), .I1(n28[6]), .I2(GND_net), 
            .I3(GND_net), .O(n384));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i259_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i308_2_lut (.I0(\Kp[6] ), .I1(n28[6]), .I2(GND_net), 
            .I3(GND_net), .O(n457));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i308_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i357_2_lut (.I0(\Kp[7] ), .I1(n28[6]), .I2(GND_net), 
            .I3(GND_net), .O(n530));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i357_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i406_2_lut (.I0(\Kp[8] ), .I1(n28[6]), .I2(GND_net), 
            .I3(GND_net), .O(n603));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i406_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i455_2_lut (.I0(\Kp[9] ), .I1(n28[6]), .I2(GND_net), 
            .I3(GND_net), .O(n676));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i455_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i504_2_lut (.I0(\Kp[10] ), .I1(n28[6]), .I2(GND_net), 
            .I3(GND_net), .O(n749));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i504_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i553_2_lut (.I0(\Kp[11] ), .I1(n28[6]), .I2(GND_net), 
            .I3(GND_net), .O(n822));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i553_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i602_2_lut (.I0(\Kp[12] ), .I1(n28[6]), .I2(GND_net), 
            .I3(GND_net), .O(n895));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i602_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i651_2_lut (.I0(\Kp[13] ), .I1(n28[6]), .I2(GND_net), 
            .I3(GND_net), .O(n968));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i651_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i700_2_lut (.I0(\Kp[14] ), .I1(n28[6]), .I2(GND_net), 
            .I3(GND_net), .O(n1041));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i700_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i749_2_lut (.I0(\Kp[15] ), .I1(n28[6]), .I2(GND_net), 
            .I3(GND_net), .O(n1114));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i749_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i65_2_lut (.I0(\Kp[1] ), .I1(n28[7]), .I2(GND_net), 
            .I3(GND_net), .O(n95));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i65_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i18_2_lut (.I0(\Kp[0] ), .I1(n28[8]), .I2(GND_net), 
            .I3(GND_net), .O(n26_adj_4313));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i18_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i114_2_lut (.I0(\Kp[2] ), .I1(n28[7]), .I2(GND_net), 
            .I3(GND_net), .O(n168));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i114_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i163_2_lut (.I0(\Kp[3] ), .I1(n28[7]), .I2(GND_net), 
            .I3(GND_net), .O(n241));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i163_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i212_2_lut (.I0(\Kp[4] ), .I1(n28[7]), .I2(GND_net), 
            .I3(GND_net), .O(n314));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i212_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i261_2_lut (.I0(\Kp[5] ), .I1(n28[7]), .I2(GND_net), 
            .I3(GND_net), .O(n387));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i261_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i310_2_lut (.I0(\Kp[6] ), .I1(n28[7]), .I2(GND_net), 
            .I3(GND_net), .O(n460));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i310_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i359_2_lut (.I0(\Kp[7] ), .I1(n28[7]), .I2(GND_net), 
            .I3(GND_net), .O(n533));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i359_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i408_2_lut (.I0(\Kp[8] ), .I1(n28[7]), .I2(GND_net), 
            .I3(GND_net), .O(n606));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i408_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i457_2_lut (.I0(\Kp[9] ), .I1(n28[7]), .I2(GND_net), 
            .I3(GND_net), .O(n679));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i457_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i506_2_lut (.I0(\Kp[10] ), .I1(n28[7]), .I2(GND_net), 
            .I3(GND_net), .O(n752));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i506_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i555_2_lut (.I0(\Kp[11] ), .I1(n28[7]), .I2(GND_net), 
            .I3(GND_net), .O(n825));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i555_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i604_2_lut (.I0(\Kp[12] ), .I1(n28[7]), .I2(GND_net), 
            .I3(GND_net), .O(n898));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i604_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i653_2_lut (.I0(\Kp[13] ), .I1(n28[7]), .I2(GND_net), 
            .I3(GND_net), .O(n971));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i653_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i702_2_lut (.I0(\Kp[14] ), .I1(n28[7]), .I2(GND_net), 
            .I3(GND_net), .O(n1044));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i702_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i751_2_lut (.I0(\Kp[15] ), .I1(n28[7]), .I2(GND_net), 
            .I3(GND_net), .O(n1117));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i751_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i67_2_lut (.I0(\Kp[1] ), .I1(n28[8]), .I2(GND_net), 
            .I3(GND_net), .O(n98));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i67_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i20_2_lut (.I0(\Kp[0] ), .I1(n28[9]), .I2(GND_net), 
            .I3(GND_net), .O(n29));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i20_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY unary_minus_5_add_3_23 (.CI(n28024), .I0(GND_net), .I1(n1[21]), 
            .CO(n28025));
    SB_LUT4 unary_minus_5_add_3_22_lut (.I0(\PID_CONTROLLER.integral [20]), 
            .I1(GND_net), .I2(n1[20]), .I3(n28023), .O(n41)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_22_lut.LUT_INIT = 16'h6996;
    SB_LUT4 mux_17_i24_3_lut (.I0(duty_23__N_3646[23]), .I1(n257[23]), .I2(n256), 
            .I3(GND_net), .O(duty_23__N_3621[23]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_17_i24_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_i24_3_lut (.I0(duty_23__N_3621[23]), .I1(PWMLimit[23]), 
            .I2(duty_23__N_3645), .I3(GND_net), .O(duty_23__N_3522[23]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_i24_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_17_i23_3_lut (.I0(duty_23__N_3646[22]), .I1(n257[22]), .I2(n256), 
            .I3(GND_net), .O(duty_23__N_3621[22]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_17_i23_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_i23_3_lut (.I0(duty_23__N_3621[22]), .I1(PWMLimit[22]), 
            .I2(duty_23__N_3645), .I3(GND_net), .O(duty_23__N_3522[22]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_i23_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_17_i22_3_lut (.I0(duty_23__N_3646[21]), .I1(n257[21]), .I2(n256), 
            .I3(GND_net), .O(duty_23__N_3621[21]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_17_i22_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_12_15_lut (.I0(GND_net), .I1(n106[13]), .I2(n155[13]), 
            .I3(n27867), .O(duty_23__N_3646[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 duty_23__I_0_i22_3_lut (.I0(duty_23__N_3621[21]), .I1(PWMLimit[21]), 
            .I2(duty_23__N_3645), .I3(GND_net), .O(duty_23__N_3522[21]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_i22_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_17_i21_3_lut (.I0(duty_23__N_3646[20]), .I1(n257[20]), .I2(n256), 
            .I3(GND_net), .O(duty_23__N_3621[20]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_17_i21_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_i21_3_lut (.I0(duty_23__N_3621[20]), .I1(PWMLimit[20]), 
            .I2(duty_23__N_3645), .I3(GND_net), .O(duty_23__N_3522[20]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_i21_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_17_i20_3_lut (.I0(duty_23__N_3646[19]), .I1(n257[19]), .I2(n256), 
            .I3(GND_net), .O(duty_23__N_3621[19]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_17_i20_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_i20_3_lut (.I0(duty_23__N_3621[19]), .I1(PWMLimit[19]), 
            .I2(duty_23__N_3645), .I3(GND_net), .O(duty_23__N_3522[19]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_i20_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_17_i19_3_lut (.I0(duty_23__N_3646[18]), .I1(n257[18]), .I2(n256), 
            .I3(GND_net), .O(duty_23__N_3621[18]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_17_i19_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_i19_3_lut (.I0(duty_23__N_3621[18]), .I1(PWMLimit[18]), 
            .I2(duty_23__N_3645), .I3(GND_net), .O(duty_23__N_3522[18]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_i19_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_17_i18_3_lut (.I0(duty_23__N_3646[17]), .I1(n257[17]), .I2(n256), 
            .I3(GND_net), .O(duty_23__N_3621[17]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_17_i18_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_i18_3_lut (.I0(duty_23__N_3621[17]), .I1(PWMLimit[17]), 
            .I2(duty_23__N_3645), .I3(GND_net), .O(duty_23__N_3522[17]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_i18_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_17_i17_3_lut (.I0(duty_23__N_3646[16]), .I1(n257[16]), .I2(n256), 
            .I3(GND_net), .O(duty_23__N_3621[16]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_17_i17_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_i17_3_lut (.I0(duty_23__N_3621[16]), .I1(PWMLimit[16]), 
            .I2(duty_23__N_3645), .I3(GND_net), .O(duty_23__N_3522[16]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_i17_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_17_i16_3_lut (.I0(duty_23__N_3646[15]), .I1(n257[15]), .I2(n256), 
            .I3(GND_net), .O(duty_23__N_3621[15]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_17_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_i16_3_lut (.I0(duty_23__N_3621[15]), .I1(PWMLimit[15]), 
            .I2(duty_23__N_3645), .I3(GND_net), .O(duty_23__N_3522[15]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_17_i15_3_lut (.I0(duty_23__N_3646[14]), .I1(n257[14]), .I2(n256), 
            .I3(GND_net), .O(duty_23__N_3621[14]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_17_i15_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_i15_3_lut (.I0(duty_23__N_3621[14]), .I1(PWMLimit[14]), 
            .I2(duty_23__N_3645), .I3(GND_net), .O(duty_23__N_3522[14]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_i15_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_17_i14_3_lut (.I0(duty_23__N_3646[13]), .I1(n257[13]), .I2(n256), 
            .I3(GND_net), .O(duty_23__N_3621[13]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_17_i14_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_i14_3_lut (.I0(duty_23__N_3621[13]), .I1(PWMLimit[13]), 
            .I2(duty_23__N_3645), .I3(GND_net), .O(duty_23__N_3522[13]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_i14_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_17_i13_3_lut (.I0(duty_23__N_3646[12]), .I1(n257[12]), .I2(n256), 
            .I3(GND_net), .O(duty_23__N_3621[12]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_17_i13_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_i13_3_lut (.I0(duty_23__N_3621[12]), .I1(PWMLimit[12]), 
            .I2(duty_23__N_3645), .I3(GND_net), .O(duty_23__N_3522[12]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_i13_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 unary_minus_5_inv_0_i1_1_lut (.I0(IntegralLimit[0]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[0]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i1_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mux_17_i12_3_lut (.I0(duty_23__N_3646[11]), .I1(n257[11]), .I2(n256), 
            .I3(GND_net), .O(duty_23__N_3621[11]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_17_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_i12_3_lut (.I0(duty_23__N_3621[11]), .I1(PWMLimit[11]), 
            .I2(duty_23__N_3645), .I3(GND_net), .O(duty_23__N_3522[11]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_17_i11_3_lut (.I0(duty_23__N_3646[10]), .I1(n257[10]), .I2(n256), 
            .I3(GND_net), .O(duty_23__N_3621[10]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_17_i11_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_i11_3_lut (.I0(duty_23__N_3621[10]), .I1(PWMLimit[10]), 
            .I2(duty_23__N_3645), .I3(GND_net), .O(duty_23__N_3522[10]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_i11_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_17_i10_3_lut (.I0(duty_23__N_3646[9]), .I1(n257[9]), .I2(n256), 
            .I3(GND_net), .O(duty_23__N_3621[9]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_17_i10_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_i10_3_lut (.I0(duty_23__N_3621[9]), .I1(PWMLimit[9]), 
            .I2(duty_23__N_3645), .I3(GND_net), .O(duty_23__N_3522[9]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_i10_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_17_i9_3_lut (.I0(duty_23__N_3646[8]), .I1(n257[8]), .I2(n256), 
            .I3(GND_net), .O(duty_23__N_3621[8]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_17_i9_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_i9_3_lut (.I0(duty_23__N_3621[8]), .I1(PWMLimit[8]), 
            .I2(duty_23__N_3645), .I3(GND_net), .O(duty_23__N_3522[8]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_i9_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_17_i8_3_lut (.I0(duty_23__N_3646[7]), .I1(n257[7]), .I2(n256), 
            .I3(GND_net), .O(duty_23__N_3621[7]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_17_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_i8_3_lut (.I0(duty_23__N_3621[7]), .I1(PWMLimit[7]), 
            .I2(duty_23__N_3645), .I3(GND_net), .O(duty_23__N_3522[7]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_17_i7_3_lut (.I0(duty_23__N_3646[6]), .I1(n257[6]), .I2(n256), 
            .I3(GND_net), .O(duty_23__N_3621[6]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_17_i7_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_i7_3_lut (.I0(duty_23__N_3621[6]), .I1(PWMLimit[6]), 
            .I2(duty_23__N_3645), .I3(GND_net), .O(duty_23__N_3522[6]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_i7_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_17_i6_3_lut (.I0(duty_23__N_3646[5]), .I1(n257[5]), .I2(n256), 
            .I3(GND_net), .O(duty_23__N_3621[5]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_17_i6_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_i6_3_lut (.I0(duty_23__N_3621[5]), .I1(PWMLimit[5]), 
            .I2(duty_23__N_3645), .I3(GND_net), .O(duty_23__N_3522[5]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_i6_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_17_i5_3_lut (.I0(duty_23__N_3646[4]), .I1(n257[4]), .I2(n256), 
            .I3(GND_net), .O(duty_23__N_3621[4]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_17_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_i5_3_lut (.I0(duty_23__N_3621[4]), .I1(PWMLimit[4]), 
            .I2(duty_23__N_3645), .I3(GND_net), .O(duty_23__N_3522[4]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_17_i4_3_lut (.I0(duty_23__N_3646[3]), .I1(n257[3]), .I2(n256), 
            .I3(GND_net), .O(duty_23__N_3621[3]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_17_i4_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_i4_3_lut (.I0(duty_23__N_3621[3]), .I1(PWMLimit[3]), 
            .I2(duty_23__N_3645), .I3(GND_net), .O(duty_23__N_3522[3]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_i4_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_10_i116_2_lut (.I0(\Kp[2] ), .I1(n28[8]), .I2(GND_net), 
            .I3(GND_net), .O(n171));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i116_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i165_2_lut (.I0(\Kp[3] ), .I1(n28[8]), .I2(GND_net), 
            .I3(GND_net), .O(n244));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i165_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i214_2_lut (.I0(\Kp[4] ), .I1(n28[8]), .I2(GND_net), 
            .I3(GND_net), .O(n317));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i214_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i263_2_lut (.I0(\Kp[5] ), .I1(n28[8]), .I2(GND_net), 
            .I3(GND_net), .O(n390));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i263_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i312_2_lut (.I0(\Kp[6] ), .I1(n28[8]), .I2(GND_net), 
            .I3(GND_net), .O(n463));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i312_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_17_i3_3_lut (.I0(duty_23__N_3646[2]), .I1(n257[2]), .I2(n256), 
            .I3(GND_net), .O(duty_23__N_3621[2]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_17_i3_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_i3_3_lut (.I0(duty_23__N_3621[2]), .I1(PWMLimit[2]), 
            .I2(duty_23__N_3645), .I3(GND_net), .O(duty_23__N_3522[2]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_i3_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_10_i361_2_lut (.I0(\Kp[7] ), .I1(n28[8]), .I2(GND_net), 
            .I3(GND_net), .O(n536));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i361_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i410_2_lut (.I0(\Kp[8] ), .I1(n28[8]), .I2(GND_net), 
            .I3(GND_net), .O(n609));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i410_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i459_2_lut (.I0(\Kp[9] ), .I1(n28[8]), .I2(GND_net), 
            .I3(GND_net), .O(n682));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i459_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i508_2_lut (.I0(\Kp[10] ), .I1(n28[8]), .I2(GND_net), 
            .I3(GND_net), .O(n755));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i508_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i557_2_lut (.I0(\Kp[11] ), .I1(n28[8]), .I2(GND_net), 
            .I3(GND_net), .O(n828));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i557_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i606_2_lut (.I0(\Kp[12] ), .I1(n28[8]), .I2(GND_net), 
            .I3(GND_net), .O(n901));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i606_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i655_2_lut (.I0(\Kp[13] ), .I1(n28[8]), .I2(GND_net), 
            .I3(GND_net), .O(n974));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i655_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i704_2_lut (.I0(\Kp[14] ), .I1(n28[8]), .I2(GND_net), 
            .I3(GND_net), .O(n1047));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i704_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i753_2_lut (.I0(\Kp[15] ), .I1(n28[8]), .I2(GND_net), 
            .I3(GND_net), .O(n1120));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i753_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i69_2_lut (.I0(\Kp[1] ), .I1(n28[9]), .I2(GND_net), 
            .I3(GND_net), .O(n101));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i69_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i22_2_lut (.I0(\Kp[0] ), .I1(n28[10]), .I2(GND_net), 
            .I3(GND_net), .O(n32));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i22_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i118_2_lut (.I0(\Kp[2] ), .I1(n28[9]), .I2(GND_net), 
            .I3(GND_net), .O(n174));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i118_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i167_2_lut (.I0(\Kp[3] ), .I1(n28[9]), .I2(GND_net), 
            .I3(GND_net), .O(n247));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i167_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i216_2_lut (.I0(\Kp[4] ), .I1(n28[9]), .I2(GND_net), 
            .I3(GND_net), .O(n320));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i216_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i265_2_lut (.I0(\Kp[5] ), .I1(n28[9]), .I2(GND_net), 
            .I3(GND_net), .O(n393));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i265_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i314_2_lut (.I0(\Kp[6] ), .I1(n28[9]), .I2(GND_net), 
            .I3(GND_net), .O(n466));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i314_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_inv_0_i2_1_lut (.I0(IntegralLimit[1]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[1]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i363_2_lut (.I0(\Kp[7] ), .I1(n28[9]), .I2(GND_net), 
            .I3(GND_net), .O(n539));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i363_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i412_2_lut (.I0(\Kp[8] ), .I1(n28[9]), .I2(GND_net), 
            .I3(GND_net), .O(n612));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i412_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i19150_2_lut (.I0(n28[22]), .I1(\PID_CONTROLLER.integral_23__N_3594 ), 
            .I2(GND_net), .I3(GND_net), .O(n3302[22]));   // verilog/motorControl.v(31[7] 33[10])
    defparam i19150_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i461_2_lut (.I0(\Kp[9] ), .I1(n28[9]), .I2(GND_net), 
            .I3(GND_net), .O(n685));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i461_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_inv_0_i3_1_lut (.I0(IntegralLimit[2]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[2]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i510_2_lut (.I0(\Kp[10] ), .I1(n28[9]), .I2(GND_net), 
            .I3(GND_net), .O(n758));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i510_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 IntegralLimit_23__I_0_i17_2_lut (.I0(\PID_CONTROLLER.integral [8]), 
            .I1(IntegralLimit[8]), .I2(GND_net), .I3(GND_net), .O(n17_adj_4317));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i17_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 IntegralLimit_23__I_0_i9_2_lut (.I0(\PID_CONTROLLER.integral [4]), 
            .I1(IntegralLimit[4]), .I2(GND_net), .I3(GND_net), .O(n9));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i9_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 IntegralLimit_23__I_0_i11_2_lut (.I0(\PID_CONTROLLER.integral [5]), 
            .I1(IntegralLimit[5]), .I2(GND_net), .I3(GND_net), .O(n11));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i11_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_10_i559_2_lut (.I0(\Kp[11] ), .I1(n28[9]), .I2(GND_net), 
            .I3(GND_net), .O(n831));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i559_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i29771_4_lut (.I0(\PID_CONTROLLER.integral [3]), .I1(\PID_CONTROLLER.integral [2]), 
            .I2(IntegralLimit[3]), .I3(IntegralLimit[2]), .O(n36526));
    defparam i29771_4_lut.LUT_INIT = 16'h7bde;
    SB_LUT4 mult_10_i608_2_lut (.I0(\Kp[12] ), .I1(n28[9]), .I2(GND_net), 
            .I3(GND_net), .O(n904));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i608_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i29768_3_lut (.I0(n11), .I1(n9), .I2(n36526), .I3(GND_net), 
            .O(n36523));
    defparam i29768_3_lut.LUT_INIT = 16'habab;
    SB_LUT4 mult_10_i657_2_lut (.I0(\Kp[13] ), .I1(n28[9]), .I2(GND_net), 
            .I3(GND_net), .O(n977));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i657_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 IntegralLimit_23__I_0_i13_rep_132_2_lut (.I0(\PID_CONTROLLER.integral [6]), 
            .I1(IntegralLimit[6]), .I2(GND_net), .I3(GND_net), .O(n38414));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i13_rep_132_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i30135_4_lut (.I0(\PID_CONTROLLER.integral [7]), .I1(n38414), 
            .I2(IntegralLimit[7]), .I3(n36523), .O(n36890));
    defparam i30135_4_lut.LUT_INIT = 16'hffde;
    SB_LUT4 mult_10_i706_2_lut (.I0(\Kp[14] ), .I1(n28[9]), .I2(GND_net), 
            .I3(GND_net), .O(n1050));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i706_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i30016_4_lut (.I0(\PID_CONTROLLER.integral [9]), .I1(n17_adj_4317), 
            .I2(IntegralLimit[9]), .I3(n36890), .O(n36771));
    defparam i30016_4_lut.LUT_INIT = 16'hdeff;
    SB_LUT4 IntegralLimit_23__I_0_i21_rep_114_2_lut (.I0(\PID_CONTROLLER.integral [10]), 
            .I1(IntegralLimit[10]), .I2(GND_net), .I3(GND_net), .O(n38396));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i21_rep_114_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i30014_4_lut (.I0(\PID_CONTROLLER.integral [9]), .I1(n17_adj_4317), 
            .I2(IntegralLimit[9]), .I3(n9), .O(n36769));
    defparam i30014_4_lut.LUT_INIT = 16'hffde;
    SB_LUT4 mult_10_i71_2_lut (.I0(\Kp[1] ), .I1(n28[10]), .I2(GND_net), 
            .I3(GND_net), .O(n104));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i71_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i30012_4_lut (.I0(\PID_CONTROLLER.integral [11]), .I1(n38396), 
            .I2(IntegralLimit[11]), .I3(n36769), .O(n36767));
    defparam i30012_4_lut.LUT_INIT = 16'hdeff;
    SB_LUT4 IntegralLimit_23__I_0_i25_rep_108_2_lut (.I0(\PID_CONTROLLER.integral [12]), 
            .I1(IntegralLimit[12]), .I2(GND_net), .I3(GND_net), .O(n38390));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i25_rep_108_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i29708_4_lut (.I0(n27), .I1(n15), .I2(n13), .I3(n11_adj_4318), 
            .O(n36463));
    defparam i29708_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i29714_4_lut (.I0(n21_adj_4319), .I1(n19_adj_4320), .I2(n17_adj_4321), 
            .I3(n9_adj_4322), .O(n36469));
    defparam i29714_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 mult_10_i24_2_lut (.I0(\Kp[0] ), .I1(n28[11]), .I2(GND_net), 
            .I3(GND_net), .O(n35));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i24_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 \PID_CONTROLLER.integral_23__I_0_i16_3_lut  (.I0(\PID_CONTROLLER.integral [9]), 
            .I1(\PID_CONTROLLER.integral [21]), .I2(n43), .I3(GND_net), 
            .O(n16_adj_4324));   // verilog/motorControl.v(31[38:63])
    defparam \PID_CONTROLLER.integral_23__I_0_i16_3_lut .LUT_INIT = 16'hcaca;
    SB_LUT4 mult_10_i120_2_lut (.I0(\Kp[2] ), .I1(n28[10]), .I2(GND_net), 
            .I3(GND_net), .O(n177));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i120_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i169_2_lut (.I0(\Kp[3] ), .I1(n28[10]), .I2(GND_net), 
            .I3(GND_net), .O(n250));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i169_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i218_2_lut (.I0(\Kp[4] ), .I1(n28[10]), .I2(GND_net), 
            .I3(GND_net), .O(n323));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i218_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i29689_2_lut (.I0(n43), .I1(n19_adj_4320), .I2(GND_net), .I3(GND_net), 
            .O(n36444));
    defparam i29689_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 mult_10_i267_2_lut (.I0(\Kp[5] ), .I1(n28[10]), .I2(GND_net), 
            .I3(GND_net), .O(n396));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i267_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 \PID_CONTROLLER.integral_23__I_0_i8_3_lut  (.I0(\PID_CONTROLLER.integral [4]), 
            .I1(\PID_CONTROLLER.integral [8]), .I2(n17_adj_4321), .I3(GND_net), 
            .O(n8));   // verilog/motorControl.v(31[38:63])
    defparam \PID_CONTROLLER.integral_23__I_0_i8_3_lut .LUT_INIT = 16'hcaca;
    SB_LUT4 \PID_CONTROLLER.integral_23__I_0_i24_3_lut  (.I0(n16_adj_4324), 
            .I1(\PID_CONTROLLER.integral [22]), .I2(n45), .I3(GND_net), 
            .O(n24_adj_4325));   // verilog/motorControl.v(31[38:63])
    defparam \PID_CONTROLLER.integral_23__I_0_i24_3_lut .LUT_INIT = 16'hcaca;
    SB_LUT4 mult_10_i316_2_lut (.I0(\Kp[6] ), .I1(n28[10]), .I2(GND_net), 
            .I3(GND_net), .O(n469));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i316_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i29724_2_lut (.I0(n7_adj_4326), .I1(n5_adj_4327), .I2(GND_net), 
            .I3(GND_net), .O(n36479));
    defparam i29724_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i29983_4_lut (.I0(n13), .I1(n11_adj_4318), .I2(n9_adj_4322), 
            .I3(n36479), .O(n36738));
    defparam i29983_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i29979_4_lut (.I0(n19_adj_4320), .I1(n17_adj_4321), .I2(n15), 
            .I3(n36738), .O(n36734));
    defparam i29979_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i30251_4_lut (.I0(n25_adj_4328), .I1(n23_adj_4329), .I2(n21_adj_4319), 
            .I3(n36734), .O(n37006));
    defparam i30251_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 mult_10_i365_2_lut (.I0(\Kp[7] ), .I1(n28[10]), .I2(GND_net), 
            .I3(GND_net), .O(n542));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i365_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i414_2_lut (.I0(\Kp[8] ), .I1(n28[10]), .I2(GND_net), 
            .I3(GND_net), .O(n615));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i414_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i463_2_lut (.I0(\Kp[9] ), .I1(n28[10]), .I2(GND_net), 
            .I3(GND_net), .O(n688));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i463_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i512_2_lut (.I0(\Kp[10] ), .I1(n28[10]), .I2(GND_net), 
            .I3(GND_net), .O(n761));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i512_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i561_2_lut (.I0(\Kp[11] ), .I1(n28[10]), .I2(GND_net), 
            .I3(GND_net), .O(n834));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i561_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i30103_4_lut (.I0(n31), .I1(n29_adj_4330), .I2(n27), .I3(n37006), 
            .O(n36858));
    defparam i30103_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 mult_10_i610_2_lut (.I0(\Kp[12] ), .I1(n28[10]), .I2(GND_net), 
            .I3(GND_net), .O(n907));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i610_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i30310_4_lut (.I0(n37), .I1(n35_adj_4331), .I2(n33), .I3(n36858), 
            .O(n37065));
    defparam i30310_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i30018_4_lut (.I0(\PID_CONTROLLER.integral [7]), .I1(n38414), 
            .I2(IntegralLimit[7]), .I3(n11), .O(n36773));
    defparam i30018_4_lut.LUT_INIT = 16'hffde;
    SB_LUT4 IntegralLimit_23__I_0_i27_rep_101_2_lut (.I0(\PID_CONTROLLER.integral [13]), 
            .I1(IntegralLimit[13]), .I2(GND_net), .I3(GND_net), .O(n38383));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i27_rep_101_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i30006_4_lut (.I0(\PID_CONTROLLER.integral [14]), .I1(n38383), 
            .I2(IntegralLimit[14]), .I3(n36773), .O(n36761));
    defparam i30006_4_lut.LUT_INIT = 16'hdeff;
    SB_LUT4 mult_10_i659_2_lut (.I0(\Kp[13] ), .I1(n28[10]), .I2(GND_net), 
            .I3(GND_net), .O(n980));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i659_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 IntegralLimit_23__I_0_i31_rep_96_2_lut (.I0(\PID_CONTROLLER.integral [15]), 
            .I1(IntegralLimit[15]), .I2(GND_net), .I3(GND_net), .O(n38378));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i31_rep_96_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 IntegralLimit_23__I_0_i12_3_lut (.I0(IntegralLimit[7]), .I1(IntegralLimit[16]), 
            .I2(\PID_CONTROLLER.integral [16]), .I3(GND_net), .O(n12));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i12_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i29743_4_lut (.I0(\PID_CONTROLLER.integral [16]), .I1(\PID_CONTROLLER.integral [7]), 
            .I2(IntegralLimit[16]), .I3(IntegralLimit[7]), .O(n36498));
    defparam i29743_4_lut.LUT_INIT = 16'h7bde;
    SB_LUT4 IntegralLimit_23__I_0_i35_rep_119_2_lut (.I0(\PID_CONTROLLER.integral [17]), 
            .I1(IntegralLimit[17]), .I2(GND_net), .I3(GND_net), .O(n38401));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i35_rep_119_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 IntegralLimit_23__I_0_i10_3_lut (.I0(IntegralLimit[5]), .I1(IntegralLimit[6]), 
            .I2(\PID_CONTROLLER.integral [6]), .I3(GND_net), .O(n10));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i10_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 IntegralLimit_23__I_0_i30_3_lut (.I0(n12), .I1(IntegralLimit[17]), 
            .I2(\PID_CONTROLLER.integral [17]), .I3(GND_net), .O(n30));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i30_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i30201_4_lut (.I0(\PID_CONTROLLER.integral [11]), .I1(n38396), 
            .I2(IntegralLimit[11]), .I3(n36771), .O(n36956));
    defparam i30201_4_lut.LUT_INIT = 16'hffde;
    SB_LUT4 mult_10_i73_2_lut (.I0(\Kp[1] ), .I1(n28[11]), .I2(GND_net), 
            .I3(GND_net), .O(n107));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i73_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i26_2_lut (.I0(\Kp[0] ), .I1(n28[12]), .I2(GND_net), 
            .I3(GND_net), .O(n38));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i26_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i29751_4_lut (.I0(\PID_CONTROLLER.integral [13]), .I1(n38390), 
            .I2(IntegralLimit[13]), .I3(n36956), .O(n36506));
    defparam i29751_4_lut.LUT_INIT = 16'h5a7b;
    SB_LUT4 mult_10_i122_2_lut (.I0(\Kp[2] ), .I1(n28[11]), .I2(GND_net), 
            .I3(GND_net), .O(n180));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i122_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 IntegralLimit_23__I_0_i29_rep_99_2_lut (.I0(\PID_CONTROLLER.integral [14]), 
            .I1(IntegralLimit[14]), .I2(GND_net), .I3(GND_net), .O(n38381));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i29_rep_99_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i30129_4_lut (.I0(\PID_CONTROLLER.integral [15]), .I1(n38381), 
            .I2(IntegralLimit[15]), .I3(n36506), .O(n36884));
    defparam i30129_4_lut.LUT_INIT = 16'hffde;
    SB_LUT4 IntegralLimit_23__I_0_i33_rep_125_2_lut (.I0(\PID_CONTROLLER.integral [16]), 
            .I1(IntegralLimit[16]), .I2(GND_net), .I3(GND_net), .O(n38407));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i33_rep_125_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i30287_4_lut (.I0(\PID_CONTROLLER.integral [17]), .I1(n38407), 
            .I2(IntegralLimit[17]), .I3(n36884), .O(n37042));
    defparam i30287_4_lut.LUT_INIT = 16'hffde;
    SB_LUT4 IntegralLimit_23__I_0_i37_rep_90_2_lut (.I0(\PID_CONTROLLER.integral [18]), 
            .I1(IntegralLimit[18]), .I2(GND_net), .I3(GND_net), .O(n38372));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i37_rep_90_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i30342_4_lut (.I0(\PID_CONTROLLER.integral [19]), .I1(n38372), 
            .I2(IntegralLimit[19]), .I3(n37042), .O(n37097));
    defparam i30342_4_lut.LUT_INIT = 16'hffde;
    SB_LUT4 IntegralLimit_23__I_0_i41_rep_87_2_lut (.I0(\PID_CONTROLLER.integral [20]), 
            .I1(IntegralLimit[20]), .I2(GND_net), .I3(GND_net), .O(n38369));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i41_rep_87_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 IntegralLimit_23__I_0_i16_3_lut (.I0(IntegralLimit[9]), .I1(IntegralLimit[21]), 
            .I2(\PID_CONTROLLER.integral [21]), .I3(GND_net), .O(n16_adj_4332));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i16_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i29727_4_lut (.I0(\PID_CONTROLLER.integral [21]), .I1(\PID_CONTROLLER.integral [9]), 
            .I2(IntegralLimit[21]), .I3(IntegralLimit[9]), .O(n36482));
    defparam i29727_4_lut.LUT_INIT = 16'h7bde;
    SB_LUT4 mult_10_i171_2_lut (.I0(\Kp[3] ), .I1(n28[11]), .I2(GND_net), 
            .I3(GND_net), .O(n253));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i171_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 IntegralLimit_23__I_0_i24_3_lut (.I0(n16_adj_4332), .I1(IntegralLimit[22]), 
            .I2(\PID_CONTROLLER.integral [22]), .I3(GND_net), .O(n24_adj_4333));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i24_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 mult_10_i220_2_lut (.I0(\Kp[4] ), .I1(n28[11]), .I2(GND_net), 
            .I3(GND_net), .O(n326));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i220_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 IntegralLimit_23__I_0_i6_3_lut (.I0(IntegralLimit[2]), .I1(IntegralLimit[3]), 
            .I2(\PID_CONTROLLER.integral [3]), .I3(GND_net), .O(n6_adj_4334));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i6_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i30143_3_lut (.I0(n6_adj_4334), .I1(IntegralLimit[10]), .I2(\PID_CONTROLLER.integral [10]), 
            .I3(GND_net), .O(n36898));   // verilog/motorControl.v(31[10:34])
    defparam i30143_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i30144_3_lut (.I0(n36898), .I1(IntegralLimit[11]), .I2(\PID_CONTROLLER.integral [11]), 
            .I3(GND_net), .O(n36899));   // verilog/motorControl.v(31[10:34])
    defparam i30144_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i29729_4_lut (.I0(\PID_CONTROLLER.integral [21]), .I1(n38390), 
            .I2(IntegralLimit[21]), .I3(n36767), .O(n36484));
    defparam i29729_4_lut.LUT_INIT = 16'h5a7b;
    SB_LUT4 mult_10_i269_2_lut (.I0(\Kp[5] ), .I1(n28[11]), .I2(GND_net), 
            .I3(GND_net), .O(n399));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i269_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i30113_4_lut (.I0(n24_adj_4333), .I1(n8_adj_4335), .I2(n38367), 
            .I3(n36482), .O(n36868));   // verilog/motorControl.v(31[10:34])
    defparam i30113_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i29994_3_lut (.I0(n36899), .I1(IntegralLimit[12]), .I2(\PID_CONTROLLER.integral [12]), 
            .I3(GND_net), .O(n36749));   // verilog/motorControl.v(31[10:34])
    defparam i29994_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 \PID_CONTROLLER.integral_23__I_0_i4_4_lut  (.I0(\PID_CONTROLLER.integral_23__N_3597 [0]), 
            .I1(\PID_CONTROLLER.integral [1]), .I2(n3_adj_4336), .I3(\PID_CONTROLLER.integral [0]), 
            .O(n4_adj_4337));   // verilog/motorControl.v(31[38:63])
    defparam \PID_CONTROLLER.integral_23__I_0_i4_4_lut .LUT_INIT = 16'hc5c0;
    SB_LUT4 i30245_3_lut (.I0(n4_adj_4337), .I1(\PID_CONTROLLER.integral [13]), 
            .I2(n27), .I3(GND_net), .O(n37000));   // verilog/motorControl.v(31[38:63])
    defparam i30245_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_10_i318_2_lut (.I0(\Kp[6] ), .I1(n28[11]), .I2(GND_net), 
            .I3(GND_net), .O(n472));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i318_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i30246_3_lut (.I0(n37000), .I1(\PID_CONTROLLER.integral [14]), 
            .I2(n29_adj_4330), .I3(GND_net), .O(n37001));   // verilog/motorControl.v(31[38:63])
    defparam i30246_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 \PID_CONTROLLER.integral_23__I_0_i12_3_lut  (.I0(\PID_CONTROLLER.integral [7]), 
            .I1(\PID_CONTROLLER.integral [16]), .I2(n33), .I3(GND_net), 
            .O(n12_adj_4338));   // verilog/motorControl.v(31[38:63])
    defparam \PID_CONTROLLER.integral_23__I_0_i12_3_lut .LUT_INIT = 16'hcaca;
    SB_LUT4 i29702_2_lut (.I0(n33), .I1(n15), .I2(GND_net), .I3(GND_net), 
            .O(n36457));
    defparam i29702_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 \PID_CONTROLLER.integral_23__I_0_i10_3_lut  (.I0(\PID_CONTROLLER.integral [5]), 
            .I1(\PID_CONTROLLER.integral [6]), .I2(n13), .I3(GND_net), 
            .O(n10_adj_4339));   // verilog/motorControl.v(31[38:63])
    defparam \PID_CONTROLLER.integral_23__I_0_i10_3_lut .LUT_INIT = 16'hcaca;
    SB_LUT4 \PID_CONTROLLER.integral_23__I_0_i30_3_lut  (.I0(n12_adj_4338), 
            .I1(\PID_CONTROLLER.integral [17]), .I2(n35_adj_4331), .I3(GND_net), 
            .O(n30_adj_4340));   // verilog/motorControl.v(31[38:63])
    defparam \PID_CONTROLLER.integral_23__I_0_i30_3_lut .LUT_INIT = 16'hcaca;
    SB_LUT4 i29704_4_lut (.I0(n33), .I1(n31), .I2(n29_adj_4330), .I3(n36463), 
            .O(n36459));
    defparam i29704_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 mult_10_i367_2_lut (.I0(\Kp[7] ), .I1(n28[11]), .I2(GND_net), 
            .I3(GND_net), .O(n545));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i367_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i30316_4_lut (.I0(n30_adj_4340), .I1(n10_adj_4339), .I2(n35_adj_4331), 
            .I3(n36457), .O(n37071));   // verilog/motorControl.v(31[38:63])
    defparam i30316_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i30172_3_lut (.I0(n37001), .I1(\PID_CONTROLLER.integral [15]), 
            .I2(n31), .I3(GND_net), .O(n36927));   // verilog/motorControl.v(31[38:63])
    defparam i30172_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_10_i416_2_lut (.I0(\Kp[8] ), .I1(n28[11]), .I2(GND_net), 
            .I3(GND_net), .O(n618));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i416_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i30365_4_lut (.I0(n36927), .I1(n37071), .I2(n35_adj_4331), 
            .I3(n36459), .O(n37120));   // verilog/motorControl.v(31[38:63])
    defparam i30365_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i30366_3_lut (.I0(n37120), .I1(\PID_CONTROLLER.integral [18]), 
            .I2(n37), .I3(GND_net), .O(n37121));   // verilog/motorControl.v(31[38:63])
    defparam i30366_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i30351_3_lut (.I0(n37121), .I1(\PID_CONTROLLER.integral [19]), 
            .I2(n39), .I3(GND_net), .O(n37106));   // verilog/motorControl.v(31[38:63])
    defparam i30351_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 \PID_CONTROLLER.integral_23__I_0_i6_3_lut  (.I0(\PID_CONTROLLER.integral [2]), 
            .I1(\PID_CONTROLLER.integral [3]), .I2(n7_adj_4326), .I3(GND_net), 
            .O(n6_adj_4341));   // verilog/motorControl.v(31[38:63])
    defparam \PID_CONTROLLER.integral_23__I_0_i6_3_lut .LUT_INIT = 16'hcaca;
    SB_LUT4 i30253_3_lut (.I0(n6_adj_4341), .I1(\PID_CONTROLLER.integral [10]), 
            .I2(n21_adj_4319), .I3(GND_net), .O(n37008));   // verilog/motorControl.v(31[38:63])
    defparam i30253_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i30254_3_lut (.I0(n37008), .I1(\PID_CONTROLLER.integral [11]), 
            .I2(n23_adj_4329), .I3(GND_net), .O(n37009));   // verilog/motorControl.v(31[38:63])
    defparam i30254_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_10_i465_2_lut (.I0(\Kp[9] ), .I1(n28[11]), .I2(GND_net), 
            .I3(GND_net), .O(n691));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i465_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i29691_4_lut (.I0(n43), .I1(n25_adj_4328), .I2(n23_adj_4329), 
            .I3(n36469), .O(n36446));
    defparam i29691_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i30117_4_lut (.I0(n24_adj_4325), .I1(n8), .I2(n45), .I3(n36444), 
            .O(n36872));   // verilog/motorControl.v(31[38:63])
    defparam i30117_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 mult_10_i514_2_lut (.I0(\Kp[10] ), .I1(n28[11]), .I2(GND_net), 
            .I3(GND_net), .O(n764));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i514_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i30170_3_lut (.I0(n37009), .I1(\PID_CONTROLLER.integral [12]), 
            .I2(n25_adj_4328), .I3(GND_net), .O(n36925));   // verilog/motorControl.v(31[38:63])
    defparam i30170_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i29694_4_lut (.I0(n43), .I1(n41), .I2(n39), .I3(n37065), 
            .O(n36449));
    defparam i29694_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i30267_4_lut (.I0(n36925), .I1(n36872), .I2(n45), .I3(n36446), 
            .O(n37022));   // verilog/motorControl.v(31[38:63])
    defparam i30267_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i30335_3_lut (.I0(n37106), .I1(\PID_CONTROLLER.integral [20]), 
            .I2(n41), .I3(GND_net), .O(n40));   // verilog/motorControl.v(31[38:63])
    defparam i30335_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i30269_4_lut (.I0(n40), .I1(n37022), .I2(n45), .I3(n36449), 
            .O(n37024));   // verilog/motorControl.v(31[38:63])
    defparam i30269_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 IntegralLimit_23__I_0_i4_4_lut (.I0(\PID_CONTROLLER.integral [0]), 
            .I1(IntegralLimit[1]), .I2(\PID_CONTROLLER.integral [1]), .I3(IntegralLimit[0]), 
            .O(n4_adj_4342));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i4_4_lut.LUT_INIT = 16'h4d0c;
    SB_LUT4 i30141_3_lut (.I0(n4_adj_4342), .I1(IntegralLimit[13]), .I2(\PID_CONTROLLER.integral [13]), 
            .I3(GND_net), .O(n36896));   // verilog/motorControl.v(31[10:34])
    defparam i30141_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i30142_3_lut (.I0(n36896), .I1(IntegralLimit[14]), .I2(\PID_CONTROLLER.integral [14]), 
            .I3(GND_net), .O(n36897));   // verilog/motorControl.v(31[10:34])
    defparam i30142_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 mult_10_i563_2_lut (.I0(\Kp[11] ), .I1(n28[11]), .I2(GND_net), 
            .I3(GND_net), .O(n837));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i563_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i29745_4_lut (.I0(\PID_CONTROLLER.integral [16]), .I1(n38378), 
            .I2(IntegralLimit[16]), .I3(n36761), .O(n36500));
    defparam i29745_4_lut.LUT_INIT = 16'h5a7b;
    SB_LUT4 i30314_4_lut (.I0(n30), .I1(n10), .I2(n38401), .I3(n36498), 
            .O(n37069));   // verilog/motorControl.v(31[10:34])
    defparam i30314_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 mult_10_i612_2_lut (.I0(\Kp[12] ), .I1(n28[11]), .I2(GND_net), 
            .I3(GND_net), .O(n910));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i612_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i29996_3_lut (.I0(n36897), .I1(IntegralLimit[15]), .I2(\PID_CONTROLLER.integral [15]), 
            .I3(GND_net), .O(n36751));   // verilog/motorControl.v(31[10:34])
    defparam i29996_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i30352_4_lut (.I0(n36751), .I1(n37069), .I2(n38401), .I3(n36500), 
            .O(n37107));   // verilog/motorControl.v(31[10:34])
    defparam i30352_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i30353_3_lut (.I0(n37107), .I1(IntegralLimit[18]), .I2(\PID_CONTROLLER.integral [18]), 
            .I3(GND_net), .O(n37108));   // verilog/motorControl.v(31[10:34])
    defparam i30353_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 mult_10_i75_2_lut (.I0(\Kp[1] ), .I1(n28[12]), .I2(GND_net), 
            .I3(GND_net), .O(n110));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i75_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i28_2_lut (.I0(\Kp[0] ), .I1(n28[13]), .I2(GND_net), 
            .I3(GND_net), .O(n41_adj_4344));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i28_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i30325_3_lut (.I0(n37108), .I1(IntegralLimit[19]), .I2(\PID_CONTROLLER.integral [19]), 
            .I3(GND_net), .O(n37080));   // verilog/motorControl.v(31[10:34])
    defparam i30325_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i29732_4_lut (.I0(\PID_CONTROLLER.integral [21]), .I1(n38369), 
            .I2(IntegralLimit[21]), .I3(n37097), .O(n36487));
    defparam i29732_4_lut.LUT_INIT = 16'h5a7b;
    SB_LUT4 IntegralLimit_23__I_0_i45_rep_85_2_lut (.I0(\PID_CONTROLLER.integral [22]), 
            .I1(IntegralLimit[22]), .I2(GND_net), .I3(GND_net), .O(n38367));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i45_rep_85_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_10_i124_2_lut (.I0(\Kp[2] ), .I1(n28[12]), .I2(GND_net), 
            .I3(GND_net), .O(n183));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i124_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i30261_4_lut (.I0(n36749), .I1(n36868), .I2(n38367), .I3(n36484), 
            .O(n37016));   // verilog/motorControl.v(31[10:34])
    defparam i30261_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i30260_3_lut (.I0(n37080), .I1(IntegralLimit[20]), .I2(\PID_CONTROLLER.integral [20]), 
            .I3(GND_net), .O(n37015));   // verilog/motorControl.v(31[10:34])
    defparam i30260_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i30270_3_lut (.I0(n37024), .I1(\PID_CONTROLLER.integral_23__N_3597 [23]), 
            .I2(\PID_CONTROLLER.integral [23]), .I3(GND_net), .O(\PID_CONTROLLER.integral_23__N_3596 ));   // verilog/motorControl.v(31[38:63])
    defparam i30270_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i30263_4_lut (.I0(n37015), .I1(n37016), .I2(n38367), .I3(n36487), 
            .O(n37018));   // verilog/motorControl.v(31[10:34])
    defparam i30263_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 mult_10_i173_2_lut (.I0(\Kp[3] ), .I1(n28[12]), .I2(GND_net), 
            .I3(GND_net), .O(n256_adj_4345));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i173_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i222_2_lut (.I0(\Kp[4] ), .I1(n28[12]), .I2(GND_net), 
            .I3(GND_net), .O(n329));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i222_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 \PID_CONTROLLER.integral_23__I_830_4_lut  (.I0(n37018), .I1(\PID_CONTROLLER.integral_23__N_3596 ), 
            .I2(\PID_CONTROLLER.integral [23]), .I3(IntegralLimit[23]), 
            .O(\PID_CONTROLLER.integral_23__N_3594 ));   // verilog/motorControl.v(31[10:63])
    defparam \PID_CONTROLLER.integral_23__I_830_4_lut .LUT_INIT = 16'h80c8;
    SB_LUT4 mult_10_i271_2_lut (.I0(\Kp[5] ), .I1(n28[12]), .I2(GND_net), 
            .I3(GND_net), .O(n402));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i271_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i320_2_lut (.I0(\Kp[6] ), .I1(n28[12]), .I2(GND_net), 
            .I3(GND_net), .O(n475));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i320_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i369_2_lut (.I0(\Kp[7] ), .I1(n28[12]), .I2(GND_net), 
            .I3(GND_net), .O(n548));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i369_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i418_2_lut (.I0(\Kp[8] ), .I1(n28[12]), .I2(GND_net), 
            .I3(GND_net), .O(n621));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i418_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i467_2_lut (.I0(\Kp[9] ), .I1(n28[12]), .I2(GND_net), 
            .I3(GND_net), .O(n694));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i467_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i516_2_lut (.I0(\Kp[10] ), .I1(n28[12]), .I2(GND_net), 
            .I3(GND_net), .O(n767));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i516_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i565_2_lut (.I0(\Kp[11] ), .I1(n28[12]), .I2(GND_net), 
            .I3(GND_net), .O(n840));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i565_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i77_2_lut (.I0(\Kp[1] ), .I1(n28[13]), .I2(GND_net), 
            .I3(GND_net), .O(n113));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i77_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i30_2_lut (.I0(\Kp[0] ), .I1(n28[14]), .I2(GND_net), 
            .I3(GND_net), .O(n44));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i30_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i126_2_lut (.I0(\Kp[2] ), .I1(n28[13]), .I2(GND_net), 
            .I3(GND_net), .O(n186));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i126_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i175_2_lut (.I0(\Kp[3] ), .I1(n28[13]), .I2(GND_net), 
            .I3(GND_net), .O(n259_adj_4347));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i175_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i224_2_lut (.I0(\Kp[4] ), .I1(n28[13]), .I2(GND_net), 
            .I3(GND_net), .O(n332));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i224_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i273_2_lut (.I0(\Kp[5] ), .I1(n28[13]), .I2(GND_net), 
            .I3(GND_net), .O(n405));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i273_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i322_2_lut (.I0(\Kp[6] ), .I1(n28[13]), .I2(GND_net), 
            .I3(GND_net), .O(n478));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i322_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i371_2_lut (.I0(\Kp[7] ), .I1(n28[13]), .I2(GND_net), 
            .I3(GND_net), .O(n551));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i371_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i420_2_lut (.I0(\Kp[8] ), .I1(n28[13]), .I2(GND_net), 
            .I3(GND_net), .O(n624));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i420_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i469_2_lut (.I0(\Kp[9] ), .I1(n28[13]), .I2(GND_net), 
            .I3(GND_net), .O(n697));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i469_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i518_2_lut (.I0(\Kp[10] ), .I1(n28[13]), .I2(GND_net), 
            .I3(GND_net), .O(n770));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i518_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i79_2_lut (.I0(\Kp[1] ), .I1(n28[14]), .I2(GND_net), 
            .I3(GND_net), .O(n116));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i79_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i32_2_lut (.I0(\Kp[0] ), .I1(n28[15]), .I2(GND_net), 
            .I3(GND_net), .O(n47));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i32_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i128_2_lut (.I0(\Kp[2] ), .I1(n28[14]), .I2(GND_net), 
            .I3(GND_net), .O(n189_adj_4349));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i128_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i177_2_lut (.I0(\Kp[3] ), .I1(n28[14]), .I2(GND_net), 
            .I3(GND_net), .O(n262_adj_4350));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i177_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i226_2_lut (.I0(\Kp[4] ), .I1(n28[14]), .I2(GND_net), 
            .I3(GND_net), .O(n335));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i226_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i275_2_lut (.I0(\Kp[5] ), .I1(n28[14]), .I2(GND_net), 
            .I3(GND_net), .O(n408));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i275_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i324_2_lut (.I0(\Kp[6] ), .I1(n28[14]), .I2(GND_net), 
            .I3(GND_net), .O(n481));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i324_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i373_2_lut (.I0(\Kp[7] ), .I1(n28[14]), .I2(GND_net), 
            .I3(GND_net), .O(n554));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i373_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i422_2_lut (.I0(\Kp[8] ), .I1(n28[14]), .I2(GND_net), 
            .I3(GND_net), .O(n627));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i422_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i471_2_lut (.I0(\Kp[9] ), .I1(n28[14]), .I2(GND_net), 
            .I3(GND_net), .O(n700));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i471_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i19151_2_lut (.I0(n28[23]), .I1(\PID_CONTROLLER.integral_23__N_3594 ), 
            .I2(GND_net), .I3(GND_net), .O(n3302[23]));   // verilog/motorControl.v(31[7] 33[10])
    defparam i19151_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_inv_0_i4_1_lut (.I0(IntegralLimit[3]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[3]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_5_inv_0_i5_1_lut (.I0(IntegralLimit[4]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[4]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_5_inv_0_i6_1_lut (.I0(IntegralLimit[5]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[5]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_5_inv_0_i7_1_lut (.I0(IntegralLimit[6]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[6]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_5_inv_0_i8_1_lut (.I0(IntegralLimit[7]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[7]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i8_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i81_2_lut (.I0(\Kp[1] ), .I1(n28[15]), .I2(GND_net), 
            .I3(GND_net), .O(n119));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i81_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i34_2_lut (.I0(\Kp[0] ), .I1(n28[16]), .I2(GND_net), 
            .I3(GND_net), .O(n50));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i34_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i130_2_lut (.I0(\Kp[2] ), .I1(n28[15]), .I2(GND_net), 
            .I3(GND_net), .O(n192));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i130_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i179_2_lut (.I0(\Kp[3] ), .I1(n28[15]), .I2(GND_net), 
            .I3(GND_net), .O(n265_adj_4357));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i179_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i228_2_lut (.I0(\Kp[4] ), .I1(n28[15]), .I2(GND_net), 
            .I3(GND_net), .O(n338));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i228_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i277_2_lut (.I0(\Kp[5] ), .I1(n28[15]), .I2(GND_net), 
            .I3(GND_net), .O(n411));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i277_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i326_2_lut (.I0(\Kp[6] ), .I1(n28[15]), .I2(GND_net), 
            .I3(GND_net), .O(n484));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i326_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i375_2_lut (.I0(\Kp[7] ), .I1(n28[15]), .I2(GND_net), 
            .I3(GND_net), .O(n557));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i375_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i424_2_lut (.I0(\Kp[8] ), .I1(n28[15]), .I2(GND_net), 
            .I3(GND_net), .O(n630));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i424_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_inv_0_i9_1_lut (.I0(IntegralLimit[8]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[8]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i9_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_5_inv_0_i10_1_lut (.I0(IntegralLimit[9]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[9]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i10_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i83_2_lut (.I0(\Kp[1] ), .I1(n28[16]), .I2(GND_net), 
            .I3(GND_net), .O(n122));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i83_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i36_2_lut (.I0(\Kp[0] ), .I1(n28[17]), .I2(GND_net), 
            .I3(GND_net), .O(n53));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i36_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i132_2_lut (.I0(\Kp[2] ), .I1(n28[16]), .I2(GND_net), 
            .I3(GND_net), .O(n195));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i132_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i181_2_lut (.I0(\Kp[3] ), .I1(n28[16]), .I2(GND_net), 
            .I3(GND_net), .O(n268_adj_4361));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i181_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_inv_0_i11_1_lut (.I0(IntegralLimit[10]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[10]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i11_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i230_2_lut (.I0(\Kp[4] ), .I1(n28[16]), .I2(GND_net), 
            .I3(GND_net), .O(n341));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i230_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i279_2_lut (.I0(\Kp[5] ), .I1(n28[16]), .I2(GND_net), 
            .I3(GND_net), .O(n414));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i279_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i328_2_lut (.I0(\Kp[6] ), .I1(n28[16]), .I2(GND_net), 
            .I3(GND_net), .O(n487));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i328_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i377_2_lut (.I0(\Kp[7] ), .I1(n28[16]), .I2(GND_net), 
            .I3(GND_net), .O(n560));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i377_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i85_2_lut (.I0(\Kp[1] ), .I1(n28[17]), .I2(GND_net), 
            .I3(GND_net), .O(n125));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i85_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i38_2_lut (.I0(\Kp[0] ), .I1(n28[18]), .I2(GND_net), 
            .I3(GND_net), .O(n56));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i38_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_inv_0_i12_1_lut (.I0(IntegralLimit[11]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[11]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i12_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_5_inv_0_i13_1_lut (.I0(IntegralLimit[12]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[12]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i13_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_5_inv_0_i14_1_lut (.I0(IntegralLimit[13]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[13]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i14_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i134_2_lut (.I0(\Kp[2] ), .I1(n28[17]), .I2(GND_net), 
            .I3(GND_net), .O(n198));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i134_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_inv_0_i15_1_lut (.I0(IntegralLimit[14]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[14]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i15_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_5_inv_0_i16_1_lut (.I0(IntegralLimit[15]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[15]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i16_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_5_inv_0_i17_1_lut (.I0(IntegralLimit[16]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[16]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i17_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_5_inv_0_i18_1_lut (.I0(IntegralLimit[17]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[17]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i18_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i183_2_lut (.I0(\Kp[3] ), .I1(n28[17]), .I2(GND_net), 
            .I3(GND_net), .O(n271_adj_4371));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i183_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i232_2_lut (.I0(\Kp[4] ), .I1(n28[17]), .I2(GND_net), 
            .I3(GND_net), .O(n344));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i232_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i281_2_lut (.I0(\Kp[5] ), .I1(n28[17]), .I2(GND_net), 
            .I3(GND_net), .O(n417));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i281_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i2_4_lut (.I0(n6_adj_4372), .I1(\Kp[4] ), .I2(n10026[2]), 
            .I3(n28[18]), .O(n10019[3]));   // verilog/motorControl.v(34[16:22])
    defparam i2_4_lut.LUT_INIT = 16'h965a;
    SB_LUT4 unary_minus_5_inv_0_i19_1_lut (.I0(IntegralLimit[18]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[18]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i19_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i22463_4_lut (.I0(\Kp[0] ), .I1(\Kp[1] ), .I2(n28[22]), .I3(n28[21]), 
            .O(n10037[0]));   // verilog/motorControl.v(34[16:22])
    defparam i22463_4_lut.LUT_INIT = 16'h6ca0;
    SB_LUT4 i2_4_lut_adj_1485 (.I0(n4_adj_4374), .I1(\Kp[3] ), .I2(n10032[1]), 
            .I3(n28[19]), .O(n10026[2]));   // verilog/motorControl.v(34[16:22])
    defparam i2_4_lut_adj_1485.LUT_INIT = 16'h965a;
    SB_LUT4 mult_10_i330_2_lut (.I0(\Kp[6] ), .I1(n28[17]), .I2(GND_net), 
            .I3(GND_net), .O(n490));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i330_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i2_4_lut_adj_1486 (.I0(\Kp[0] ), .I1(\Kp[3] ), .I2(n28[23]), 
            .I3(n28[20]), .O(n12_adj_4375));   // verilog/motorControl.v(34[16:22])
    defparam i2_4_lut_adj_1486.LUT_INIT = 16'h9c50;
    SB_LUT4 i22399_4_lut (.I0(n10026[2]), .I1(\Kp[4] ), .I2(n6_adj_4372), 
            .I3(n28[18]), .O(n8_adj_4376));   // verilog/motorControl.v(34[16:22])
    defparam i22399_4_lut.LUT_INIT = 16'he8a0;
    SB_LUT4 i1_4_lut (.I0(\Kp[4] ), .I1(\Kp[2] ), .I2(n28[19]), .I3(n28[21]), 
            .O(n11_adj_4377));   // verilog/motorControl.v(34[16:22])
    defparam i1_4_lut.LUT_INIT = 16'h6ca0;
    SB_LUT4 i22430_4_lut (.I0(n10032[1]), .I1(\Kp[3] ), .I2(n4_adj_4374), 
            .I3(n28[19]), .O(n6_adj_4378));   // verilog/motorControl.v(34[16:22])
    defparam i22430_4_lut.LUT_INIT = 16'he8a0;
    SB_LUT4 i22465_4_lut (.I0(\Kp[0] ), .I1(\Kp[1] ), .I2(n28[22]), .I3(n28[21]), 
            .O(n27573));   // verilog/motorControl.v(34[16:22])
    defparam i22465_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i8_4_lut (.I0(n6_adj_4378), .I1(n11_adj_4377), .I2(n8_adj_4376), 
            .I3(n12_adj_4375), .O(n18_adj_4379));   // verilog/motorControl.v(34[16:22])
    defparam i8_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut (.I0(\Kp[5] ), .I1(\Kp[1] ), .I2(n28[18]), .I3(n28[22]), 
            .O(n13_adj_4380));   // verilog/motorControl.v(34[16:22])
    defparam i3_4_lut.LUT_INIT = 16'h6ca0;
    SB_LUT4 i9_4_lut (.I0(n13_adj_4380), .I1(n18_adj_4379), .I2(n27573), 
            .I3(n4_adj_4381), .O(n34086));   // verilog/motorControl.v(34[16:22])
    defparam i9_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 mult_11_i53_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3546 [1]), 
            .I2(GND_net), .I3(GND_net), .O(n77));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i53_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i6_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3546 [2]), 
            .I2(GND_net), .I3(GND_net), .O(n8_adj_4382));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i6_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i102_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3546 [1]), 
            .I2(GND_net), .I3(GND_net), .O(n150));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i102_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i151_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3546 [1]), 
            .I2(GND_net), .I3(GND_net), .O(n223));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i151_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i200_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3546 [1]), 
            .I2(GND_net), .I3(GND_net), .O(n296));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i200_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i249_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3546 [1]), 
            .I2(GND_net), .I3(GND_net), .O(n369));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i249_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i298_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3546 [1]), 
            .I2(GND_net), .I3(GND_net), .O(n442));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i298_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i347_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3546 [1]), 
            .I2(GND_net), .I3(GND_net), .O(n515));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i347_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i396_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3546 [1]), 
            .I2(GND_net), .I3(GND_net), .O(n588));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i396_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i445_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral_23__N_3546 [1]), 
            .I2(GND_net), .I3(GND_net), .O(n661));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i445_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i494_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral_23__N_3546 [1]), 
            .I2(GND_net), .I3(GND_net), .O(n734));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i494_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i543_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral_23__N_3546 [1]), 
            .I2(GND_net), .I3(GND_net), .O(n807));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i543_2_lut.LUT_INIT = 16'h8888;
    SB_DFF result_i0 (.Q(duty[0]), .C(clk32MHz), .D(duty_23__N_3522[0]));   // verilog/motorControl.v(29[14] 48[8])
    SB_LUT4 mult_11_i592_2_lut (.I0(\Ki[12] ), .I1(\PID_CONTROLLER.integral_23__N_3546 [1]), 
            .I2(GND_net), .I3(GND_net), .O(n880));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i592_2_lut.LUT_INIT = 16'h8888;
    SB_DFF \PID_CONTROLLER.integral_i0  (.Q(\PID_CONTROLLER.integral [0]), 
           .C(clk32MHz), .D(\PID_CONTROLLER.integral_23__N_3546 [0]));   // verilog/motorControl.v(29[14] 48[8])
    SB_LUT4 mult_11_i641_2_lut (.I0(\Ki[13] ), .I1(\PID_CONTROLLER.integral_23__N_3546 [1]), 
            .I2(GND_net), .I3(GND_net), .O(n953));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i641_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i690_2_lut (.I0(\Ki[14] ), .I1(\PID_CONTROLLER.integral_23__N_3546 [1]), 
            .I2(GND_net), .I3(GND_net), .O(n1026));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i690_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i739_2_lut (.I0(\Ki[15] ), .I1(\PID_CONTROLLER.integral_23__N_3546 [1]), 
            .I2(GND_net), .I3(GND_net), .O(n1099));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i739_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_inv_0_i24_1_lut (.I0(IntegralLimit[23]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[23]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i24_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_16_inv_0_i1_1_lut (.I0(PWMLimit[0]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4735[0]));   // verilog/motorControl.v(39[18:27])
    defparam unary_minus_16_inv_0_i1_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_16_inv_0_i2_1_lut (.I0(PWMLimit[1]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4735[1]));   // verilog/motorControl.v(39[18:27])
    defparam unary_minus_16_inv_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY unary_minus_5_add_3_22 (.CI(n28023), .I0(GND_net), .I1(n1[20]), 
            .CO(n28024));
    SB_LUT4 unary_minus_16_inv_0_i3_1_lut (.I0(PWMLimit[2]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4735[2]));   // verilog/motorControl.v(39[18:27])
    defparam unary_minus_16_inv_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_16_inv_0_i4_1_lut (.I0(PWMLimit[3]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4735[3]));   // verilog/motorControl.v(39[18:27])
    defparam unary_minus_16_inv_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_5_add_3_21_lut (.I0(\PID_CONTROLLER.integral [19]), 
            .I1(GND_net), .I2(n1[19]), .I3(n28022), .O(n39)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_21_lut.LUT_INIT = 16'h6996;
    SB_LUT4 mult_11_i51_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3546 [0]), 
            .I2(GND_net), .I3(GND_net), .O(n74));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i51_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i4_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3546 [1]), 
            .I2(GND_net), .I3(GND_net), .O(n5_adj_4388));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i4_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i100_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3546 [0]), 
            .I2(GND_net), .I3(GND_net), .O(n147));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i100_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i149_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3546 [0]), 
            .I2(GND_net), .I3(GND_net), .O(n220));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i149_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i198_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3546 [0]), 
            .I2(GND_net), .I3(GND_net), .O(n293));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i198_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_16_inv_0_i5_1_lut (.I0(PWMLimit[4]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4735[4]));   // verilog/motorControl.v(39[18:27])
    defparam unary_minus_16_inv_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_11_i247_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3546 [0]), 
            .I2(GND_net), .I3(GND_net), .O(n366));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i247_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i296_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3546 [0]), 
            .I2(GND_net), .I3(GND_net), .O(n439));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i296_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i345_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3546 [0]), 
            .I2(GND_net), .I3(GND_net), .O(n512));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i345_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i394_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3546 [0]), 
            .I2(GND_net), .I3(GND_net), .O(n585));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i394_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i443_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral_23__N_3546 [0]), 
            .I2(GND_net), .I3(GND_net), .O(n658));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i443_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i492_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral_23__N_3546 [0]), 
            .I2(GND_net), .I3(GND_net), .O(n731));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i492_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i541_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral_23__N_3546 [0]), 
            .I2(GND_net), .I3(GND_net), .O(n804));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i541_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i590_2_lut (.I0(\Ki[12] ), .I1(\PID_CONTROLLER.integral_23__N_3546 [0]), 
            .I2(GND_net), .I3(GND_net), .O(n877));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i590_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i639_2_lut (.I0(\Ki[13] ), .I1(\PID_CONTROLLER.integral_23__N_3546 [0]), 
            .I2(GND_net), .I3(GND_net), .O(n950));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i639_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i688_2_lut (.I0(\Ki[14] ), .I1(\PID_CONTROLLER.integral_23__N_3546 [0]), 
            .I2(GND_net), .I3(GND_net), .O(n1023));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i688_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i737_2_lut (.I0(\Ki[15] ), .I1(\PID_CONTROLLER.integral_23__N_3546 [0]), 
            .I2(GND_net), .I3(GND_net), .O(n1096));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i737_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i55_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3546 [2]), 
            .I2(GND_net), .I3(GND_net), .O(n80));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i55_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i8_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3546 [3]), 
            .I2(GND_net), .I3(GND_net), .O(n11_adj_4390));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i8_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i104_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3546 [2]), 
            .I2(GND_net), .I3(GND_net), .O(n153));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i104_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i153_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3546 [2]), 
            .I2(GND_net), .I3(GND_net), .O(n226));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i153_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_16_inv_0_i6_1_lut (.I0(PWMLimit[5]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4735[5]));   // verilog/motorControl.v(39[18:27])
    defparam unary_minus_16_inv_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_12_15 (.CI(n27867), .I0(n106[13]), .I1(n155[13]), .CO(n27868));
    SB_LUT4 mult_11_i202_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3546 [2]), 
            .I2(GND_net), .I3(GND_net), .O(n299));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i202_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i251_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3546 [2]), 
            .I2(GND_net), .I3(GND_net), .O(n372));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i251_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i300_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3546 [2]), 
            .I2(GND_net), .I3(GND_net), .O(n445));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i300_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i349_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3546 [2]), 
            .I2(GND_net), .I3(GND_net), .O(n518));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i349_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i398_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3546 [2]), 
            .I2(GND_net), .I3(GND_net), .O(n591));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i398_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i447_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral_23__N_3546 [2]), 
            .I2(GND_net), .I3(GND_net), .O(n664));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i447_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i496_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral_23__N_3546 [2]), 
            .I2(GND_net), .I3(GND_net), .O(n737));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i496_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i545_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral_23__N_3546 [2]), 
            .I2(GND_net), .I3(GND_net), .O(n810));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i545_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i594_2_lut (.I0(\Ki[12] ), .I1(\PID_CONTROLLER.integral_23__N_3546 [2]), 
            .I2(GND_net), .I3(GND_net), .O(n883));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i594_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i643_2_lut (.I0(\Ki[13] ), .I1(\PID_CONTROLLER.integral_23__N_3546 [2]), 
            .I2(GND_net), .I3(GND_net), .O(n956));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i643_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i692_2_lut (.I0(\Ki[14] ), .I1(\PID_CONTROLLER.integral_23__N_3546 [2]), 
            .I2(GND_net), .I3(GND_net), .O(n1029));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i692_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i741_2_lut (.I0(\Ki[15] ), .I1(\PID_CONTROLLER.integral_23__N_3546 [2]), 
            .I2(GND_net), .I3(GND_net), .O(n1102));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i741_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_16_inv_0_i7_1_lut (.I0(PWMLimit[6]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4735[6]));   // verilog/motorControl.v(39[18:27])
    defparam unary_minus_16_inv_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY unary_minus_5_add_3_21 (.CI(n28022), .I0(GND_net), .I1(n1[19]), 
            .CO(n28023));
    SB_LUT4 add_12_14_lut (.I0(GND_net), .I1(n106[12]), .I2(n155[12]), 
            .I3(n27866), .O(duty_23__N_3646[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_12_14 (.CI(n27866), .I0(n106[12]), .I1(n155[12]), .CO(n27867));
    SB_LUT4 unary_minus_5_add_3_20_lut (.I0(\PID_CONTROLLER.integral [18]), 
            .I1(GND_net), .I2(n1[18]), .I3(n28021), .O(n37)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_20_lut.LUT_INIT = 16'h6996;
    SB_LUT4 unary_minus_16_inv_0_i8_1_lut (.I0(PWMLimit[7]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4735[7]));   // verilog/motorControl.v(39[18:27])
    defparam unary_minus_16_inv_0_i8_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_16_inv_0_i9_1_lut (.I0(PWMLimit[8]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4735[8]));   // verilog/motorControl.v(39[18:27])
    defparam unary_minus_16_inv_0_i9_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_11_i57_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3546 [3]), 
            .I2(GND_net), .I3(GND_net), .O(n83));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i57_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_12_13_lut (.I0(GND_net), .I1(n106[11]), .I2(n155[11]), 
            .I3(n27865), .O(duty_23__N_3646[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i10_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3546 [4]), 
            .I2(GND_net), .I3(GND_net), .O(n14_adj_4396));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i10_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i106_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3546 [3]), 
            .I2(GND_net), .I3(GND_net), .O(n156));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i106_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i155_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3546 [3]), 
            .I2(GND_net), .I3(GND_net), .O(n229));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i155_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i204_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3546 [3]), 
            .I2(GND_net), .I3(GND_net), .O(n302));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i204_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY unary_minus_5_add_3_20 (.CI(n28021), .I0(GND_net), .I1(n1[18]), 
            .CO(n28022));
    SB_LUT4 mult_11_i253_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3546 [3]), 
            .I2(GND_net), .I3(GND_net), .O(n375));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i253_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_add_3_19_lut (.I0(\PID_CONTROLLER.integral [17]), 
            .I1(GND_net), .I2(n1[17]), .I3(n28020), .O(n35_adj_4331)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_19_lut.LUT_INIT = 16'h6996;
    SB_LUT4 unary_minus_16_inv_0_i10_1_lut (.I0(PWMLimit[9]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4735[9]));   // verilog/motorControl.v(39[18:27])
    defparam unary_minus_16_inv_0_i10_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_11_i302_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3546 [3]), 
            .I2(GND_net), .I3(GND_net), .O(n448));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i302_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_16_inv_0_i11_1_lut (.I0(PWMLimit[10]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4735[10]));   // verilog/motorControl.v(39[18:27])
    defparam unary_minus_16_inv_0_i11_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_11_i351_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3546 [3]), 
            .I2(GND_net), .I3(GND_net), .O(n521));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i351_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i400_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3546 [3]), 
            .I2(GND_net), .I3(GND_net), .O(n594));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i400_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_12_13 (.CI(n27865), .I0(n106[11]), .I1(n155[11]), .CO(n27866));
    SB_LUT4 mult_11_i449_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral_23__N_3546 [3]), 
            .I2(GND_net), .I3(GND_net), .O(n667));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i449_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i498_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral_23__N_3546 [3]), 
            .I2(GND_net), .I3(GND_net), .O(n740));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i498_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i547_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral_23__N_3546 [3]), 
            .I2(GND_net), .I3(GND_net), .O(n813));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i547_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i596_2_lut (.I0(\Ki[12] ), .I1(\PID_CONTROLLER.integral_23__N_3546 [3]), 
            .I2(GND_net), .I3(GND_net), .O(n886));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i596_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i645_2_lut (.I0(\Ki[13] ), .I1(\PID_CONTROLLER.integral_23__N_3546 [3]), 
            .I2(GND_net), .I3(GND_net), .O(n959));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i645_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i694_2_lut (.I0(\Ki[14] ), .I1(\PID_CONTROLLER.integral_23__N_3546 [3]), 
            .I2(GND_net), .I3(GND_net), .O(n1032));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i694_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i743_2_lut (.I0(\Ki[15] ), .I1(\PID_CONTROLLER.integral_23__N_3546 [3]), 
            .I2(GND_net), .I3(GND_net), .O(n1105));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i743_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_16_inv_0_i12_1_lut (.I0(PWMLimit[11]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4735[11]));   // verilog/motorControl.v(39[18:27])
    defparam unary_minus_16_inv_0_i12_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_11_i59_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3546 [4]), 
            .I2(GND_net), .I3(GND_net), .O(n86));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i59_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i12_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3546 [5]), 
            .I2(GND_net), .I3(GND_net), .O(n17_adj_4400));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i12_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i53_2_lut (.I0(\Kp[1] ), .I1(n28[1]), .I2(GND_net), 
            .I3(GND_net), .O(n77_adj_4402));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i53_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i6_2_lut (.I0(\Kp[0] ), .I1(n28[2]), .I2(GND_net), 
            .I3(GND_net), .O(n8_adj_4404));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i6_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i102_2_lut (.I0(\Kp[2] ), .I1(n28[1]), .I2(GND_net), 
            .I3(GND_net), .O(n150_adj_4405));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i102_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_16_inv_0_i13_1_lut (.I0(PWMLimit[12]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4735[12]));   // verilog/motorControl.v(39[18:27])
    defparam unary_minus_16_inv_0_i13_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i151_2_lut (.I0(\Kp[3] ), .I1(n28[1]), .I2(GND_net), 
            .I3(GND_net), .O(n223_adj_4407));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i151_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i200_2_lut (.I0(\Kp[4] ), .I1(n28[1]), .I2(GND_net), 
            .I3(GND_net), .O(n296_adj_4408));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i200_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i108_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3546 [4]), 
            .I2(GND_net), .I3(GND_net), .O(n159));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i108_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i157_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3546 [4]), 
            .I2(GND_net), .I3(GND_net), .O(n232));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i157_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i206_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3546 [4]), 
            .I2(GND_net), .I3(GND_net), .O(n305));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i206_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i255_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3546 [4]), 
            .I2(GND_net), .I3(GND_net), .O(n378));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i255_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i304_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3546 [4]), 
            .I2(GND_net), .I3(GND_net), .O(n451));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i304_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i353_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3546 [4]), 
            .I2(GND_net), .I3(GND_net), .O(n524));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i353_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i249_2_lut (.I0(\Kp[5] ), .I1(n28[1]), .I2(GND_net), 
            .I3(GND_net), .O(n369_adj_4409));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i249_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i402_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3546 [4]), 
            .I2(GND_net), .I3(GND_net), .O(n597));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i402_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i451_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral_23__N_3546 [4]), 
            .I2(GND_net), .I3(GND_net), .O(n670));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i451_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i298_2_lut (.I0(\Kp[6] ), .I1(n28[1]), .I2(GND_net), 
            .I3(GND_net), .O(n442_adj_4410));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i298_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i500_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral_23__N_3546 [4]), 
            .I2(GND_net), .I3(GND_net), .O(n743));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i500_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i347_2_lut (.I0(\Kp[7] ), .I1(n28[1]), .I2(GND_net), 
            .I3(GND_net), .O(n515_adj_4411));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i347_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i549_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral_23__N_3546 [4]), 
            .I2(GND_net), .I3(GND_net), .O(n816));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i549_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i598_2_lut (.I0(\Ki[12] ), .I1(\PID_CONTROLLER.integral_23__N_3546 [4]), 
            .I2(GND_net), .I3(GND_net), .O(n889));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i598_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i647_2_lut (.I0(\Ki[13] ), .I1(\PID_CONTROLLER.integral_23__N_3546 [4]), 
            .I2(GND_net), .I3(GND_net), .O(n962));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i647_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i396_2_lut (.I0(\Kp[8] ), .I1(n28[1]), .I2(GND_net), 
            .I3(GND_net), .O(n588_adj_4412));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i396_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i696_2_lut (.I0(\Ki[14] ), .I1(\PID_CONTROLLER.integral_23__N_3546 [4]), 
            .I2(GND_net), .I3(GND_net), .O(n1035));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i696_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i745_2_lut (.I0(\Ki[15] ), .I1(\PID_CONTROLLER.integral_23__N_3546 [4]), 
            .I2(GND_net), .I3(GND_net), .O(n1108));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i745_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i445_2_lut (.I0(\Kp[9] ), .I1(n28[1]), .I2(GND_net), 
            .I3(GND_net), .O(n661_adj_4413));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i445_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i494_2_lut (.I0(\Kp[10] ), .I1(n28[1]), .I2(GND_net), 
            .I3(GND_net), .O(n734_adj_4414));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i494_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i61_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3546 [5]), 
            .I2(GND_net), .I3(GND_net), .O(n89));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i61_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i14_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3546 [6]), 
            .I2(GND_net), .I3(GND_net), .O(n20_adj_4415));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i14_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i110_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3546 [5]), 
            .I2(GND_net), .I3(GND_net), .O(n162_adj_4416));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i110_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY unary_minus_5_add_3_19 (.CI(n28020), .I0(GND_net), .I1(n1[17]), 
            .CO(n28021));
    SB_LUT4 mult_10_i543_2_lut (.I0(\Kp[11] ), .I1(n28[1]), .I2(GND_net), 
            .I3(GND_net), .O(n807_adj_4417));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i543_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i159_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3546 [5]), 
            .I2(GND_net), .I3(GND_net), .O(n235_adj_4418));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i159_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i208_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3546 [5]), 
            .I2(GND_net), .I3(GND_net), .O(n308_adj_4419));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i208_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i257_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3546 [5]), 
            .I2(GND_net), .I3(GND_net), .O(n381_adj_4420));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i257_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i306_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3546 [5]), 
            .I2(GND_net), .I3(GND_net), .O(n454_adj_4421));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i306_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i355_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3546 [5]), 
            .I2(GND_net), .I3(GND_net), .O(n527_adj_4422));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i355_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i592_2_lut (.I0(\Kp[12] ), .I1(n28[1]), .I2(GND_net), 
            .I3(GND_net), .O(n880_adj_4423));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i592_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_12_12_lut (.I0(GND_net), .I1(n106[10]), .I2(n155[10]), 
            .I3(n27864), .O(duty_23__N_3646[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i404_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3546 [5]), 
            .I2(GND_net), .I3(GND_net), .O(n600_adj_4424));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i404_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i453_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral_23__N_3546 [5]), 
            .I2(GND_net), .I3(GND_net), .O(n673_adj_4425));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i453_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i641_2_lut (.I0(\Kp[13] ), .I1(n28[1]), .I2(GND_net), 
            .I3(GND_net), .O(n953_adj_4426));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i641_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i502_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral_23__N_3546 [5]), 
            .I2(GND_net), .I3(GND_net), .O(n746_adj_4427));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i502_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i22453_3_lut_4_lut (.I0(\Kp[2] ), .I1(n28[20]), .I2(n27548), 
            .I3(n10037[0]), .O(n4_adj_4381));   // verilog/motorControl.v(34[16:22])
    defparam i22453_3_lut_4_lut.LUT_INIT = 16'hf880;
    SB_LUT4 mult_11_i551_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral_23__N_3546 [5]), 
            .I2(GND_net), .I3(GND_net), .O(n819_adj_4428));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i551_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i2_3_lut_4_lut (.I0(\Kp[2] ), .I1(n28[20]), .I2(n10037[0]), 
            .I3(n27548), .O(n10032[1]));   // verilog/motorControl.v(34[16:22])
    defparam i2_3_lut_4_lut.LUT_INIT = 16'h8778;
    SB_LUT4 mult_11_i600_2_lut (.I0(\Ki[12] ), .I1(\PID_CONTROLLER.integral_23__N_3546 [5]), 
            .I2(GND_net), .I3(GND_net), .O(n892_adj_4429));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i600_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_add_3_18_lut (.I0(\PID_CONTROLLER.integral [16]), 
            .I1(GND_net), .I2(n1[16]), .I3(n28019), .O(n33)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_18_lut.LUT_INIT = 16'h6996;
    SB_LUT4 mult_11_i649_2_lut (.I0(\Ki[13] ), .I1(\PID_CONTROLLER.integral_23__N_3546 [5]), 
            .I2(GND_net), .I3(GND_net), .O(n965_adj_4430));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i649_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i22440_2_lut_3_lut_4_lut (.I0(\Kp[0] ), .I1(n28[21]), .I2(n28[20]), 
            .I3(\Kp[1] ), .O(n10032[0]));   // verilog/motorControl.v(34[16:22])
    defparam i22440_2_lut_3_lut_4_lut.LUT_INIT = 16'h7888;
    SB_LUT4 mult_11_i698_2_lut (.I0(\Ki[14] ), .I1(\PID_CONTROLLER.integral_23__N_3546 [5]), 
            .I2(GND_net), .I3(GND_net), .O(n1038_adj_4431));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i698_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_12_12 (.CI(n27864), .I0(n106[10]), .I1(n155[10]), .CO(n27865));
    SB_LUT4 i22442_2_lut_3_lut_4_lut (.I0(\Kp[0] ), .I1(n28[21]), .I2(n28[20]), 
            .I3(\Kp[1] ), .O(n27548));   // verilog/motorControl.v(34[16:22])
    defparam i22442_2_lut_3_lut_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 mult_11_i747_2_lut (.I0(\Ki[15] ), .I1(\PID_CONTROLLER.integral_23__N_3546 [5]), 
            .I2(GND_net), .I3(GND_net), .O(n1111_adj_4432));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i747_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i690_2_lut (.I0(\Kp[14] ), .I1(n28[1]), .I2(GND_net), 
            .I3(GND_net), .O(n1026_adj_4433));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i690_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i63_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3546 [6]), 
            .I2(GND_net), .I3(GND_net), .O(n92_adj_4434));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i63_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i16_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3546 [7]), 
            .I2(GND_net), .I3(GND_net), .O(n23_adj_4435));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i16_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i112_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3546 [6]), 
            .I2(GND_net), .I3(GND_net), .O(n165_adj_4436));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i112_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i161_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3546 [6]), 
            .I2(GND_net), .I3(GND_net), .O(n238_adj_4437));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i161_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY unary_minus_5_add_3_18 (.CI(n28019), .I0(GND_net), .I1(n1[16]), 
            .CO(n28020));
    SB_LUT4 mult_10_i739_2_lut (.I0(\Kp[15] ), .I1(n28[1]), .I2(GND_net), 
            .I3(GND_net), .O(n1099_adj_4438));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i739_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_12_11_lut (.I0(GND_net), .I1(n106[9]), .I2(n155[9]), .I3(n27863), 
            .O(duty_23__N_3646[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_5_add_3_17_lut (.I0(\PID_CONTROLLER.integral [15]), 
            .I1(GND_net), .I2(n1[15]), .I3(n28018), .O(n31)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_17_lut.LUT_INIT = 16'h6996;
    SB_CARRY unary_minus_5_add_3_17 (.CI(n28018), .I0(GND_net), .I1(n1[15]), 
            .CO(n28019));
    SB_LUT4 unary_minus_5_add_3_16_lut (.I0(\PID_CONTROLLER.integral [14]), 
            .I1(GND_net), .I2(n1[14]), .I3(n28017), .O(n29_adj_4330)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_16_lut.LUT_INIT = 16'h6996;
    SB_CARRY unary_minus_5_add_3_16 (.CI(n28017), .I0(GND_net), .I1(n1[14]), 
            .CO(n28018));
    SB_LUT4 mult_11_i210_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3546 [6]), 
            .I2(GND_net), .I3(GND_net), .O(n311_adj_4439));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i210_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_12_11 (.CI(n27863), .I0(n106[9]), .I1(n155[9]), .CO(n27864));
    SB_LUT4 unary_minus_5_add_3_15_lut (.I0(\PID_CONTROLLER.integral [13]), 
            .I1(GND_net), .I2(n1[13]), .I3(n28016), .O(n27)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_15_lut.LUT_INIT = 16'h6996;
    SB_CARRY unary_minus_5_add_3_15 (.CI(n28016), .I0(GND_net), .I1(n1[13]), 
            .CO(n28017));
    SB_LUT4 unary_minus_5_add_3_14_lut (.I0(\PID_CONTROLLER.integral [12]), 
            .I1(GND_net), .I2(n1[12]), .I3(n28015), .O(n25_adj_4328)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_14_lut.LUT_INIT = 16'h6996;
    SB_LUT4 add_12_10_lut (.I0(GND_net), .I1(n106[8]), .I2(n155[8]), .I3(n27862), 
            .O(duty_23__N_3646[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_12_10 (.CI(n27862), .I0(n106[8]), .I1(n155[8]), .CO(n27863));
    SB_CARRY unary_minus_5_add_3_14 (.CI(n28015), .I0(GND_net), .I1(n1[12]), 
            .CO(n28016));
    SB_LUT4 add_12_9_lut (.I0(GND_net), .I1(n106[7]), .I2(n155[7]), .I3(n27861), 
            .O(duty_23__N_3646[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_5_add_3_13_lut (.I0(\PID_CONTROLLER.integral [11]), 
            .I1(GND_net), .I2(n1[11]), .I3(n28014), .O(n23_adj_4329)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_13_lut.LUT_INIT = 16'h6996;
    SB_CARRY add_12_9 (.CI(n27861), .I0(n106[7]), .I1(n155[7]), .CO(n27862));
    SB_LUT4 mult_11_i259_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3546 [6]), 
            .I2(GND_net), .I3(GND_net), .O(n384_adj_4442));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i259_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i2_3_lut_4_lut_adj_1487 (.I0(\Kp[2] ), .I1(n28[19]), .I2(n10032[0]), 
            .I3(n27514), .O(n10026[1]));   // verilog/motorControl.v(34[16:22])
    defparam i2_3_lut_4_lut_adj_1487.LUT_INIT = 16'h8778;
    SB_CARRY unary_minus_5_add_3_13 (.CI(n28014), .I0(GND_net), .I1(n1[11]), 
            .CO(n28015));
    SB_LUT4 mult_11_i308_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3546 [6]), 
            .I2(GND_net), .I3(GND_net), .O(n457_adj_4443));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i308_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_add_3_12_lut (.I0(\PID_CONTROLLER.integral [10]), 
            .I1(GND_net), .I2(n1[10]), .I3(n28013), .O(n21_adj_4319)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_12_lut.LUT_INIT = 16'h6996;
    SB_CARRY unary_minus_5_add_3_12 (.CI(n28013), .I0(GND_net), .I1(n1[10]), 
            .CO(n28014));
    SB_LUT4 add_12_8_lut (.I0(GND_net), .I1(n106[6]), .I2(n155[6]), .I3(n27860), 
            .O(duty_23__N_3646[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_5_add_3_11_lut (.I0(\PID_CONTROLLER.integral [9]), 
            .I1(GND_net), .I2(n1[9]), .I3(n28012), .O(n19_adj_4320)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_11_lut.LUT_INIT = 16'h6996;
    SB_CARRY add_12_8 (.CI(n27860), .I0(n106[6]), .I1(n155[6]), .CO(n27861));
    SB_LUT4 i22422_3_lut_4_lut (.I0(\Kp[2] ), .I1(n28[19]), .I2(n27514), 
            .I3(n10032[0]), .O(n4_adj_4374));   // verilog/motorControl.v(34[16:22])
    defparam i22422_3_lut_4_lut.LUT_INIT = 16'hf880;
    SB_CARRY unary_minus_5_add_3_11 (.CI(n28012), .I0(GND_net), .I1(n1[9]), 
            .CO(n28013));
    SB_LUT4 i22409_2_lut_3_lut_4_lut (.I0(\Kp[0] ), .I1(n28[20]), .I2(n28[19]), 
            .I3(\Kp[1] ), .O(n10026[0]));   // verilog/motorControl.v(34[16:22])
    defparam i22409_2_lut_3_lut_4_lut.LUT_INIT = 16'h7888;
    SB_LUT4 i22411_2_lut_3_lut_4_lut (.I0(\Kp[0] ), .I1(n28[20]), .I2(n28[19]), 
            .I3(\Kp[1] ), .O(n27514));   // verilog/motorControl.v(34[16:22])
    defparam i22411_2_lut_3_lut_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 add_12_7_lut (.I0(GND_net), .I1(n106[5]), .I2(n155[5]), .I3(n27859), 
            .O(duty_23__N_3646[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_5_add_3_10_lut (.I0(\PID_CONTROLLER.integral [8]), 
            .I1(GND_net), .I2(n1[8]), .I3(n28011), .O(n17_adj_4321)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_10_lut.LUT_INIT = 16'h6996;
    SB_CARRY unary_minus_5_add_3_10 (.CI(n28011), .I0(GND_net), .I1(n1[8]), 
            .CO(n28012));
    SB_LUT4 unary_minus_5_add_3_9_lut (.I0(\PID_CONTROLLER.integral [7]), 
            .I1(GND_net), .I2(n1[7]), .I3(n28010), .O(n15)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_9_lut.LUT_INIT = 16'h6996;
    SB_CARRY unary_minus_5_add_3_9 (.CI(n28010), .I0(GND_net), .I1(n1[7]), 
            .CO(n28011));
    SB_CARRY add_12_7 (.CI(n27859), .I0(n106[5]), .I1(n155[5]), .CO(n27860));
    SB_LUT4 add_12_6_lut (.I0(GND_net), .I1(n106[4]), .I2(n155[4]), .I3(n27858), 
            .O(duty_23__N_3646[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_5_add_3_8_lut (.I0(\PID_CONTROLLER.integral [6]), 
            .I1(GND_net), .I2(n1[6]), .I3(n28009), .O(n13)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_8_lut.LUT_INIT = 16'h6996;
    SB_CARRY unary_minus_5_add_3_8 (.CI(n28009), .I0(GND_net), .I1(n1[6]), 
            .CO(n28010));
    SB_LUT4 unary_minus_5_add_3_7_lut (.I0(\PID_CONTROLLER.integral [5]), 
            .I1(GND_net), .I2(n1[5]), .I3(n28008), .O(n11_adj_4318)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_7_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i22391_3_lut_4_lut (.I0(\Kp[3] ), .I1(n28[18]), .I2(n4_adj_4446), 
            .I3(n10026[1]), .O(n6_adj_4372));   // verilog/motorControl.v(34[16:22])
    defparam i22391_3_lut_4_lut.LUT_INIT = 16'hf880;
    SB_LUT4 mult_11_i357_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3546 [6]), 
            .I2(GND_net), .I3(GND_net), .O(n530_adj_4447));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i357_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY unary_minus_5_add_3_7 (.CI(n28008), .I0(GND_net), .I1(n1[5]), 
            .CO(n28009));
    SB_CARRY add_12_6 (.CI(n27858), .I0(n106[4]), .I1(n155[4]), .CO(n27859));
    SB_LUT4 add_12_5_lut (.I0(GND_net), .I1(n106[3]), .I2(n155[3]), .I3(n27857), 
            .O(duty_23__N_3646[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i406_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3546 [6]), 
            .I2(GND_net), .I3(GND_net), .O(n603_adj_4448));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i406_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_add_3_6_lut (.I0(\PID_CONTROLLER.integral [4]), 
            .I1(GND_net), .I2(n1[4]), .I3(n28007), .O(n9_adj_4322)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_6_lut.LUT_INIT = 16'h6996;
    SB_LUT4 mult_11_i455_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral_23__N_3546 [6]), 
            .I2(GND_net), .I3(GND_net), .O(n676_adj_4449));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i455_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i504_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral_23__N_3546 [6]), 
            .I2(GND_net), .I3(GND_net), .O(n749_adj_4450));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i504_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY unary_minus_5_add_3_6 (.CI(n28007), .I0(GND_net), .I1(n1[4]), 
            .CO(n28008));
    SB_LUT4 unary_minus_5_add_3_5_lut (.I0(\PID_CONTROLLER.integral [3]), 
            .I1(GND_net), .I2(n1[3]), .I3(n28006), .O(n7_adj_4326)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_5_lut.LUT_INIT = 16'h6996;
    SB_LUT4 add_751_25_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [23]), 
            .I2(n3302[23]), .I3(n27920), .O(\PID_CONTROLLER.integral_23__N_3546 [23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_751_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_5_add_3_5 (.CI(n28006), .I0(GND_net), .I1(n1[3]), 
            .CO(n28007));
    SB_LUT4 unary_minus_5_add_3_4_lut (.I0(\PID_CONTROLLER.integral [2]), 
            .I1(GND_net), .I2(n1[2]), .I3(n28005), .O(n5_adj_4327)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_4_lut.LUT_INIT = 16'h6996;
    SB_CARRY add_12_5 (.CI(n27857), .I0(n106[3]), .I1(n155[3]), .CO(n27858));
    SB_CARRY unary_minus_5_add_3_4 (.CI(n28005), .I0(GND_net), .I1(n1[2]), 
            .CO(n28006));
    SB_LUT4 mult_11_i553_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral_23__N_3546 [6]), 
            .I2(GND_net), .I3(GND_net), .O(n822_adj_4451));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i553_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i602_2_lut (.I0(\Ki[12] ), .I1(\PID_CONTROLLER.integral_23__N_3546 [6]), 
            .I2(GND_net), .I3(GND_net), .O(n895_adj_4452));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i602_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i651_2_lut (.I0(\Ki[13] ), .I1(\PID_CONTROLLER.integral_23__N_3546 [6]), 
            .I2(GND_net), .I3(GND_net), .O(n968_adj_4453));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i651_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i700_2_lut (.I0(\Ki[14] ), .I1(\PID_CONTROLLER.integral_23__N_3546 [6]), 
            .I2(GND_net), .I3(GND_net), .O(n1041_adj_4454));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i700_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i749_2_lut (.I0(\Ki[15] ), .I1(\PID_CONTROLLER.integral_23__N_3546 [6]), 
            .I2(GND_net), .I3(GND_net), .O(n1114_adj_4455));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i749_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i65_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3546 [7]), 
            .I2(GND_net), .I3(GND_net), .O(n95_adj_4456));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i65_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i18_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3546 [8]), 
            .I2(GND_net), .I3(GND_net), .O(n26_adj_4457));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i18_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i51_2_lut (.I0(\Kp[1] ), .I1(n28[0]), .I2(GND_net), 
            .I3(GND_net), .O(n74_adj_4458));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i51_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i114_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3546 [7]), 
            .I2(GND_net), .I3(GND_net), .O(n168_adj_4459));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i114_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_12_4_lut (.I0(GND_net), .I1(n106[2]), .I2(n155[2]), .I3(n27856), 
            .O(duty_23__N_3646[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i4_2_lut (.I0(\Kp[0] ), .I1(n28[1]), .I2(GND_net), 
            .I3(GND_net), .O(n5_adj_4460));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i4_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i163_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3546 [7]), 
            .I2(GND_net), .I3(GND_net), .O(n241_adj_4461));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i163_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_751_24_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [22]), 
            .I2(n3302[22]), .I3(n27919), .O(\PID_CONTROLLER.integral_23__N_3546 [22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_751_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_12_4 (.CI(n27856), .I0(n106[2]), .I1(n155[2]), .CO(n27857));
    SB_LUT4 mult_11_i212_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3546 [7]), 
            .I2(GND_net), .I3(GND_net), .O(n314_adj_4462));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i212_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i2_3_lut_4_lut_adj_1488 (.I0(\Kp[3] ), .I1(n28[18]), .I2(n10026[1]), 
            .I3(n4_adj_4446), .O(n10019[2]));   // verilog/motorControl.v(34[16:22])
    defparam i2_3_lut_4_lut_adj_1488.LUT_INIT = 16'h8778;
    SB_LUT4 unary_minus_5_add_3_3_lut (.I0(\PID_CONTROLLER.integral [1]), 
            .I1(GND_net), .I2(n1[1]), .I3(n28004), .O(n3_adj_4336)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_3_lut.LUT_INIT = 16'h6996;
    SB_LUT4 mult_11_i261_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3546 [7]), 
            .I2(GND_net), .I3(GND_net), .O(n387_adj_4463));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i261_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i2_3_lut_4_lut_adj_1489 (.I0(\Kp[2] ), .I1(n28[18]), .I2(n10026[0]), 
            .I3(n27471), .O(n10019[1]));   // verilog/motorControl.v(34[16:22])
    defparam i2_3_lut_4_lut_adj_1489.LUT_INIT = 16'h8778;
    SB_LUT4 mult_11_i310_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3546 [7]), 
            .I2(GND_net), .I3(GND_net), .O(n460_adj_4464));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i310_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i359_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3546 [7]), 
            .I2(GND_net), .I3(GND_net), .O(n533_adj_4465));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i359_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i408_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3546 [7]), 
            .I2(GND_net), .I3(GND_net), .O(n606_adj_4466));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i408_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i18692_2_lut (.I0(n28[0]), .I1(\PID_CONTROLLER.integral_23__N_3594 ), 
            .I2(GND_net), .I3(GND_net), .O(n3302[0]));   // verilog/motorControl.v(31[7] 33[10])
    defparam i18692_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_751_24 (.CI(n27919), .I0(\PID_CONTROLLER.integral [22]), 
            .I1(n3302[22]), .CO(n27920));
    SB_CARRY unary_minus_5_add_3_3 (.CI(n28004), .I0(GND_net), .I1(n1[1]), 
            .CO(n28005));
    SB_LUT4 unary_minus_5_add_3_2_lut (.I0(GND_net), .I1(GND_net), .I2(n1[0]), 
            .I3(VCC_net), .O(\PID_CONTROLLER.integral_23__N_3597 [0])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_12_3_lut (.I0(GND_net), .I1(n106[1]), .I2(n155[1]), .I3(n27855), 
            .O(duty_23__N_3646[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_5_add_3_2 (.CI(VCC_net), .I0(GND_net), .I1(n1[0]), 
            .CO(n28004));
    SB_LUT4 mult_11_i457_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral_23__N_3546 [7]), 
            .I2(GND_net), .I3(GND_net), .O(n679_adj_4468));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i457_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i22383_3_lut_4_lut (.I0(\Kp[2] ), .I1(n28[18]), .I2(n27471), 
            .I3(n10026[0]), .O(n4_adj_4446));   // verilog/motorControl.v(34[16:22])
    defparam i22383_3_lut_4_lut.LUT_INIT = 16'hf880;
    SB_LUT4 mult_10_i100_2_lut (.I0(\Kp[2] ), .I1(n28[0]), .I2(GND_net), 
            .I3(GND_net), .O(n147_adj_4469));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i100_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i506_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral_23__N_3546 [7]), 
            .I2(GND_net), .I3(GND_net), .O(n752_adj_4470));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i506_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i555_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral_23__N_3546 [7]), 
            .I2(GND_net), .I3(GND_net), .O(n825_adj_4471));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i555_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_751_23_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [21]), 
            .I2(n3302[21]), .I3(n27918), .O(\PID_CONTROLLER.integral_23__N_3546 [21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_751_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_751_23 (.CI(n27918), .I0(\PID_CONTROLLER.integral [21]), 
            .I1(n3302[21]), .CO(n27919));
    SB_LUT4 mult_10_i149_2_lut (.I0(\Kp[3] ), .I1(n28[0]), .I2(GND_net), 
            .I3(GND_net), .O(n220_adj_4472));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i149_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_12_3 (.CI(n27855), .I0(n106[1]), .I1(n155[1]), .CO(n27856));
    SB_LUT4 mult_11_i604_2_lut (.I0(\Ki[12] ), .I1(\PID_CONTROLLER.integral_23__N_3546 [7]), 
            .I2(GND_net), .I3(GND_net), .O(n898_adj_4473));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i604_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i653_2_lut (.I0(\Ki[13] ), .I1(\PID_CONTROLLER.integral_23__N_3546 [7]), 
            .I2(GND_net), .I3(GND_net), .O(n971_adj_4474));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i653_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_751_22_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [20]), 
            .I2(n3302[20]), .I3(n27917), .O(\PID_CONTROLLER.integral_23__N_3546 [20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_751_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i198_2_lut (.I0(\Kp[4] ), .I1(n28[0]), .I2(GND_net), 
            .I3(GND_net), .O(n293_adj_4475));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i198_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i702_2_lut (.I0(\Ki[14] ), .I1(\PID_CONTROLLER.integral_23__N_3546 [7]), 
            .I2(GND_net), .I3(GND_net), .O(n1044_adj_4476));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i702_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i751_2_lut (.I0(\Ki[15] ), .I1(\PID_CONTROLLER.integral_23__N_3546 [7]), 
            .I2(GND_net), .I3(GND_net), .O(n1117_adj_4477));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i751_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i247_2_lut (.I0(\Kp[5] ), .I1(n28[0]), .I2(GND_net), 
            .I3(GND_net), .O(n366_adj_4478));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i247_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i67_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3546 [8]), 
            .I2(GND_net), .I3(GND_net), .O(n98_adj_4479));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i67_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i20_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3546 [9]), 
            .I2(GND_net), .I3(GND_net), .O(n29_adj_4480));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i20_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i116_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3546 [8]), 
            .I2(GND_net), .I3(GND_net), .O(n171_adj_4481));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i116_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i19129_2_lut (.I0(n28[1]), .I1(\PID_CONTROLLER.integral_23__N_3594 ), 
            .I2(GND_net), .I3(GND_net), .O(n3302[1]));   // verilog/motorControl.v(31[7] 33[10])
    defparam i19129_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i165_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3546 [8]), 
            .I2(GND_net), .I3(GND_net), .O(n244_adj_4482));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i165_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i19130_2_lut (.I0(n28[2]), .I1(\PID_CONTROLLER.integral_23__N_3594 ), 
            .I2(GND_net), .I3(GND_net), .O(n3302[2]));   // verilog/motorControl.v(31[7] 33[10])
    defparam i19130_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i296_2_lut (.I0(\Kp[6] ), .I1(n28[0]), .I2(GND_net), 
            .I3(GND_net), .O(n439_adj_4483));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i296_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i214_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3546 [8]), 
            .I2(GND_net), .I3(GND_net), .O(n317_adj_4484));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i214_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i263_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3546 [8]), 
            .I2(GND_net), .I3(GND_net), .O(n390_adj_4485));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i263_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i312_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3546 [8]), 
            .I2(GND_net), .I3(GND_net), .O(n463_adj_4486));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i312_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i361_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3546 [8]), 
            .I2(GND_net), .I3(GND_net), .O(n536_adj_4487));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i361_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i410_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3546 [8]), 
            .I2(GND_net), .I3(GND_net), .O(n609_adj_4488));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i410_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_17_i2_3_lut (.I0(duty_23__N_3646[1]), .I1(n257[1]), .I2(n256), 
            .I3(GND_net), .O(duty_23__N_3621[1]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_17_i2_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_i2_3_lut (.I0(duty_23__N_3621[1]), .I1(PWMLimit[1]), 
            .I2(duty_23__N_3645), .I3(GND_net), .O(duty_23__N_3522[1]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_i2_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_10_i345_2_lut (.I0(\Kp[7] ), .I1(n28[0]), .I2(GND_net), 
            .I3(GND_net), .O(n512_adj_4489));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i345_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i394_2_lut (.I0(\Kp[8] ), .I1(n28[0]), .I2(GND_net), 
            .I3(GND_net), .O(n585_adj_4490));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i394_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_751_22 (.CI(n27917), .I0(\PID_CONTROLLER.integral [20]), 
            .I1(n3302[20]), .CO(n27918));
    SB_LUT4 mult_10_i443_2_lut (.I0(\Kp[9] ), .I1(n28[0]), .I2(GND_net), 
            .I3(GND_net), .O(n658_adj_4491));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i443_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_751_21_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [19]), 
            .I2(n3302[19]), .I3(n27916), .O(\PID_CONTROLLER.integral_23__N_3546 [19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_751_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i459_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral_23__N_3546 [8]), 
            .I2(GND_net), .I3(GND_net), .O(n682_adj_4492));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i459_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_12_2_lut (.I0(GND_net), .I1(n106[0]), .I2(n155[0]), .I3(GND_net), 
            .O(duty_23__N_3646[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_12_2 (.CI(GND_net), .I0(n106[0]), .I1(n155[0]), .CO(n27855));
    SB_CARRY add_751_21 (.CI(n27916), .I0(\PID_CONTROLLER.integral [19]), 
            .I1(n3302[19]), .CO(n27917));
    SB_LUT4 mult_10_i492_2_lut (.I0(\Kp[10] ), .I1(n28[0]), .I2(GND_net), 
            .I3(GND_net), .O(n731_adj_4493));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i492_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i508_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral_23__N_3546 [8]), 
            .I2(GND_net), .I3(GND_net), .O(n755_adj_4494));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i508_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i557_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral_23__N_3546 [8]), 
            .I2(GND_net), .I3(GND_net), .O(n828_adj_4495));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i557_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i606_2_lut (.I0(\Ki[12] ), .I1(\PID_CONTROLLER.integral_23__N_3546 [8]), 
            .I2(GND_net), .I3(GND_net), .O(n901_adj_4496));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i606_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i655_2_lut (.I0(\Ki[13] ), .I1(\PID_CONTROLLER.integral_23__N_3546 [8]), 
            .I2(GND_net), .I3(GND_net), .O(n974_adj_4497));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i655_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i704_2_lut (.I0(\Ki[14] ), .I1(\PID_CONTROLLER.integral_23__N_3546 [8]), 
            .I2(GND_net), .I3(GND_net), .O(n1047_adj_4498));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i704_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i541_2_lut (.I0(\Kp[11] ), .I1(n28[0]), .I2(GND_net), 
            .I3(GND_net), .O(n804_adj_4499));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i541_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i590_2_lut (.I0(\Kp[12] ), .I1(n28[0]), .I2(GND_net), 
            .I3(GND_net), .O(n877_adj_4500));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i590_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i753_2_lut (.I0(\Ki[15] ), .I1(\PID_CONTROLLER.integral_23__N_3546 [8]), 
            .I2(GND_net), .I3(GND_net), .O(n1120_adj_4501));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i753_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i69_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3546 [9]), 
            .I2(GND_net), .I3(GND_net), .O(n101_adj_4502));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i69_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i639_2_lut (.I0(\Kp[13] ), .I1(n28[0]), .I2(GND_net), 
            .I3(GND_net), .O(n950_adj_4503));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i639_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i22_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3546 [10]), 
            .I2(GND_net), .I3(GND_net), .O(n32_adj_4504));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i22_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i118_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3546 [9]), 
            .I2(GND_net), .I3(GND_net), .O(n174_adj_4505));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i118_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i167_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3546 [9]), 
            .I2(GND_net), .I3(GND_net), .O(n247_adj_4506));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i167_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i216_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3546 [9]), 
            .I2(GND_net), .I3(GND_net), .O(n320_adj_4507));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i216_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i265_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3546 [9]), 
            .I2(GND_net), .I3(GND_net), .O(n393_adj_4508));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i265_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i314_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3546 [9]), 
            .I2(GND_net), .I3(GND_net), .O(n466_adj_4509));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i314_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i363_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3546 [9]), 
            .I2(GND_net), .I3(GND_net), .O(n539_adj_4510));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i363_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i22370_2_lut_3_lut_4_lut (.I0(\Kp[0] ), .I1(n28[19]), .I2(n28[18]), 
            .I3(\Kp[1] ), .O(n10019[0]));   // verilog/motorControl.v(34[16:22])
    defparam i22370_2_lut_3_lut_4_lut.LUT_INIT = 16'h7888;
    SB_LUT4 mult_11_i412_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3546 [9]), 
            .I2(GND_net), .I3(GND_net), .O(n612_adj_4511));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i412_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i461_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral_23__N_3546 [9]), 
            .I2(GND_net), .I3(GND_net), .O(n685_adj_4512));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i461_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 sub_3_add_2_25_lut (.I0(GND_net), .I1(setpoint[23]), .I2(motor_state[23]), 
            .I3(n27998), .O(n28[23])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_3_add_2_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i688_2_lut (.I0(\Kp[14] ), .I1(n28[0]), .I2(GND_net), 
            .I3(GND_net), .O(n1023_adj_4513));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i688_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 sub_3_add_2_24_lut (.I0(GND_net), .I1(setpoint[22]), .I2(motor_state[22]), 
            .I3(n27997), .O(n28[22])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_3_add_2_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i510_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral_23__N_3546 [9]), 
            .I2(GND_net), .I3(GND_net), .O(n758_adj_4514));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i510_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i559_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral_23__N_3546 [9]), 
            .I2(GND_net), .I3(GND_net), .O(n831_adj_4515));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i559_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i608_2_lut (.I0(\Ki[12] ), .I1(\PID_CONTROLLER.integral_23__N_3546 [9]), 
            .I2(GND_net), .I3(GND_net), .O(n904_adj_4516));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i608_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i657_2_lut (.I0(\Ki[13] ), .I1(\PID_CONTROLLER.integral_23__N_3546 [9]), 
            .I2(GND_net), .I3(GND_net), .O(n977_adj_4517));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i657_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i737_2_lut (.I0(\Kp[15] ), .I1(n28[0]), .I2(GND_net), 
            .I3(GND_net), .O(n1096_adj_4518));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i737_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i706_2_lut (.I0(\Ki[14] ), .I1(\PID_CONTROLLER.integral_23__N_3546 [9]), 
            .I2(GND_net), .I3(GND_net), .O(n1050_adj_4519));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i706_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i71_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3546 [10]), 
            .I2(GND_net), .I3(GND_net), .O(n104_adj_4520));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i71_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i24_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3546 [11]), 
            .I2(GND_net), .I3(GND_net), .O(n35_adj_4521));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i24_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i22372_2_lut_3_lut_4_lut (.I0(\Kp[0] ), .I1(n28[19]), .I2(n28[18]), 
            .I3(\Kp[1] ), .O(n27471));   // verilog/motorControl.v(34[16:22])
    defparam i22372_2_lut_3_lut_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 add_751_20_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [18]), 
            .I2(n3302[18]), .I3(n27915), .O(\PID_CONTROLLER.integral_23__N_3546 [18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_751_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_751_20 (.CI(n27915), .I0(\PID_CONTROLLER.integral [18]), 
            .I1(n3302[18]), .CO(n27916));
    SB_LUT4 add_751_19_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [17]), 
            .I2(n3302[17]), .I3(n27914), .O(\PID_CONTROLLER.integral_23__N_3546 [17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_751_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i120_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3546 [10]), 
            .I2(GND_net), .I3(GND_net), .O(n177_adj_4522));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i120_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY sub_3_add_2_24 (.CI(n27997), .I0(setpoint[22]), .I1(motor_state[22]), 
            .CO(n27998));
    SB_LUT4 sub_3_add_2_23_lut (.I0(GND_net), .I1(setpoint[21]), .I2(motor_state[21]), 
            .I3(n27996), .O(n28[21])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_3_add_2_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_751_19 (.CI(n27914), .I0(\PID_CONTROLLER.integral [17]), 
            .I1(n3302[17]), .CO(n27915));
    SB_CARRY sub_3_add_2_23 (.CI(n27996), .I0(setpoint[21]), .I1(motor_state[21]), 
            .CO(n27997));
    SB_LUT4 sub_3_add_2_22_lut (.I0(GND_net), .I1(setpoint[20]), .I2(motor_state[20]), 
            .I3(n27995), .O(n28[20])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_3_add_2_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_3_add_2_22 (.CI(n27995), .I0(setpoint[20]), .I1(motor_state[20]), 
            .CO(n27996));
    SB_LUT4 add_751_18_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [16]), 
            .I2(n3302[16]), .I3(n27913), .O(\PID_CONTROLLER.integral_23__N_3546 [16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_751_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_3_add_2_21_lut (.I0(GND_net), .I1(setpoint[19]), .I2(motor_state[19]), 
            .I3(n27994), .O(n28[19])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_3_add_2_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_3_add_2_21 (.CI(n27994), .I0(setpoint[19]), .I1(motor_state[19]), 
            .CO(n27995));
    SB_CARRY add_751_18 (.CI(n27913), .I0(\PID_CONTROLLER.integral [16]), 
            .I1(n3302[16]), .CO(n27914));
    SB_LUT4 mult_11_i169_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3546 [10]), 
            .I2(GND_net), .I3(GND_net), .O(n250_adj_4523));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i169_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i218_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3546 [10]), 
            .I2(GND_net), .I3(GND_net), .O(n323_adj_4524));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i218_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 sub_3_add_2_20_lut (.I0(GND_net), .I1(setpoint[18]), .I2(motor_state[18]), 
            .I3(n27993), .O(n28[18])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_3_add_2_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_3_add_2_20 (.CI(n27993), .I0(setpoint[18]), .I1(motor_state[18]), 
            .CO(n27994));
    SB_LUT4 sub_3_add_2_19_lut (.I0(GND_net), .I1(setpoint[17]), .I2(motor_state[17]), 
            .I3(n27992), .O(n28[17])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_3_add_2_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_751_17_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [15]), 
            .I2(n3302[15]), .I3(n27912), .O(\PID_CONTROLLER.integral_23__N_3546 [15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_751_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_751_17 (.CI(n27912), .I0(\PID_CONTROLLER.integral [15]), 
            .I1(n3302[15]), .CO(n27913));
    SB_CARRY sub_3_add_2_19 (.CI(n27992), .I0(setpoint[17]), .I1(motor_state[17]), 
            .CO(n27993));
    SB_LUT4 sub_3_add_2_18_lut (.I0(GND_net), .I1(setpoint[16]), .I2(motor_state[16]), 
            .I3(n27991), .O(n28[16])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_3_add_2_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i267_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3546 [10]), 
            .I2(GND_net), .I3(GND_net), .O(n396_adj_4525));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i267_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i316_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3546 [10]), 
            .I2(GND_net), .I3(GND_net), .O(n469_adj_4526));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i316_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY sub_3_add_2_18 (.CI(n27991), .I0(setpoint[16]), .I1(motor_state[16]), 
            .CO(n27992));
    SB_LUT4 mult_11_i365_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3546 [10]), 
            .I2(GND_net), .I3(GND_net), .O(n542_adj_4527));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i365_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i414_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3546 [10]), 
            .I2(GND_net), .I3(GND_net), .O(n615_adj_4528));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i414_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i463_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral_23__N_3546 [10]), 
            .I2(GND_net), .I3(GND_net), .O(n688_adj_4529));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i463_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_16_inv_0_i14_1_lut (.I0(PWMLimit[13]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4735[13]));   // verilog/motorControl.v(39[18:27])
    defparam unary_minus_16_inv_0_i14_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_3_add_2_17_lut (.I0(GND_net), .I1(setpoint[15]), .I2(motor_state[15]), 
            .I3(n27990), .O(n28[15])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_3_add_2_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i512_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral_23__N_3546 [10]), 
            .I2(GND_net), .I3(GND_net), .O(n761_adj_4531));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i512_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_751_16_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [14]), 
            .I2(n3302[14]), .I3(n27911), .O(\PID_CONTROLLER.integral_23__N_3546 [14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_751_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i561_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral_23__N_3546 [10]), 
            .I2(GND_net), .I3(GND_net), .O(n834_adj_4532));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i561_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_751_16 (.CI(n27911), .I0(\PID_CONTROLLER.integral [14]), 
            .I1(n3302[14]), .CO(n27912));
    SB_CARRY sub_3_add_2_17 (.CI(n27990), .I0(setpoint[15]), .I1(motor_state[15]), 
            .CO(n27991));
    SB_LUT4 sub_3_add_2_16_lut (.I0(GND_net), .I1(setpoint[14]), .I2(motor_state[14]), 
            .I3(n27989), .O(n28[14])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_3_add_2_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_751_15_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [13]), 
            .I2(n3302[13]), .I3(n27910), .O(\PID_CONTROLLER.integral_23__N_3546 [13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_751_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_3_add_2_16 (.CI(n27989), .I0(setpoint[14]), .I1(motor_state[14]), 
            .CO(n27990));
    SB_CARRY add_751_15 (.CI(n27910), .I0(\PID_CONTROLLER.integral [13]), 
            .I1(n3302[13]), .CO(n27911));
    SB_LUT4 add_751_14_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [12]), 
            .I2(n3302[12]), .I3(n27909), .O(\PID_CONTROLLER.integral_23__N_3546 [12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_751_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_751_14 (.CI(n27909), .I0(\PID_CONTROLLER.integral [12]), 
            .I1(n3302[12]), .CO(n27910));
    SB_LUT4 sub_3_add_2_15_lut (.I0(GND_net), .I1(setpoint[13]), .I2(motor_state[13]), 
            .I3(n27988), .O(n28[13])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_3_add_2_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_3_add_2_15 (.CI(n27988), .I0(setpoint[13]), .I1(motor_state[13]), 
            .CO(n27989));
    SB_LUT4 add_751_13_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [11]), 
            .I2(n3302[11]), .I3(n27908), .O(\PID_CONTROLLER.integral_23__N_3546 [11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_751_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_3_add_2_14_lut (.I0(GND_net), .I1(setpoint[12]), .I2(motor_state[12]), 
            .I3(n27987), .O(n28[12])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_3_add_2_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_3_add_2_14 (.CI(n27987), .I0(setpoint[12]), .I1(motor_state[12]), 
            .CO(n27988));
    SB_LUT4 sub_3_add_2_13_lut (.I0(GND_net), .I1(setpoint[11]), .I2(motor_state[11]), 
            .I3(n27986), .O(n28[11])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_3_add_2_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_3_add_2_13 (.CI(n27986), .I0(setpoint[11]), .I1(motor_state[11]), 
            .CO(n27987));
    SB_LUT4 sub_3_add_2_12_lut (.I0(GND_net), .I1(setpoint[10]), .I2(motor_state[10]), 
            .I3(n27985), .O(n28[10])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_3_add_2_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i55_2_lut (.I0(\Kp[1] ), .I1(n28[2]), .I2(GND_net), 
            .I3(GND_net), .O(n80_adj_4533));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i55_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i8_2_lut (.I0(\Kp[0] ), .I1(n28[3]), .I2(GND_net), 
            .I3(GND_net), .O(n11_adj_4535));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i8_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5283_7_lut (.I0(GND_net), .I1(n34185), .I2(n490_adj_4536), 
            .I3(n29353), .O(n10308[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5283_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5283_6_lut (.I0(GND_net), .I1(n10316[3]), .I2(n417_adj_4537), 
            .I3(n29352), .O(n10308[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5283_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5283_6 (.CI(n29352), .I0(n10316[3]), .I1(n417_adj_4537), 
            .CO(n29353));
    SB_LUT4 add_5283_5_lut (.I0(GND_net), .I1(n10316[2]), .I2(n344_adj_4538), 
            .I3(n29351), .O(n10308[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5283_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5283_5 (.CI(n29351), .I0(n10316[2]), .I1(n344_adj_4538), 
            .CO(n29352));
    SB_LUT4 add_5283_4_lut (.I0(GND_net), .I1(n10316[1]), .I2(n271_adj_4539), 
            .I3(n29350), .O(n10308[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5283_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5283_4 (.CI(n29350), .I0(n10316[1]), .I1(n271_adj_4539), 
            .CO(n29351));
    SB_LUT4 add_5283_3_lut (.I0(GND_net), .I1(n10316[0]), .I2(n198_adj_4540), 
            .I3(n29349), .O(n10308[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5283_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5283_3 (.CI(n29349), .I0(n10316[0]), .I1(n198_adj_4540), 
            .CO(n29350));
    SB_LUT4 add_5283_2_lut (.I0(GND_net), .I1(n56_adj_4541), .I2(n125_adj_4542), 
            .I3(GND_net), .O(n10308[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5283_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5283_2 (.CI(GND_net), .I0(n56_adj_4541), .I1(n125_adj_4542), 
            .CO(n29349));
    SB_LUT4 add_5282_8_lut (.I0(GND_net), .I1(n10308[5]), .I2(n560_adj_4543), 
            .I3(n29348), .O(n10299[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5282_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5282_7_lut (.I0(GND_net), .I1(n10308[4]), .I2(n487_adj_4544), 
            .I3(n29347), .O(n10299[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5282_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5282_7 (.CI(n29347), .I0(n10308[4]), .I1(n487_adj_4544), 
            .CO(n29348));
    SB_LUT4 add_5282_6_lut (.I0(GND_net), .I1(n10308[3]), .I2(n414_adj_4545), 
            .I3(n29346), .O(n10299[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5282_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5282_6 (.CI(n29346), .I0(n10308[3]), .I1(n414_adj_4545), 
            .CO(n29347));
    SB_LUT4 add_5282_5_lut (.I0(GND_net), .I1(n10308[2]), .I2(n341_adj_4546), 
            .I3(n29345), .O(n10299[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5282_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5282_5 (.CI(n29345), .I0(n10308[2]), .I1(n341_adj_4546), 
            .CO(n29346));
    SB_LUT4 add_5282_4_lut (.I0(GND_net), .I1(n10308[1]), .I2(n268_adj_4547), 
            .I3(n29344), .O(n10299[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5282_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5282_4 (.CI(n29344), .I0(n10308[1]), .I1(n268_adj_4547), 
            .CO(n29345));
    SB_LUT4 add_5282_3_lut (.I0(GND_net), .I1(n10308[0]), .I2(n195_adj_4548), 
            .I3(n29343), .O(n10299[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5282_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5282_3 (.CI(n29343), .I0(n10308[0]), .I1(n195_adj_4548), 
            .CO(n29344));
    SB_LUT4 add_5282_2_lut (.I0(GND_net), .I1(n53_adj_4549), .I2(n122_adj_4550), 
            .I3(GND_net), .O(n10299[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5282_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5282_2 (.CI(GND_net), .I0(n53_adj_4549), .I1(n122_adj_4550), 
            .CO(n29343));
    SB_LUT4 add_5281_9_lut (.I0(GND_net), .I1(n10299[6]), .I2(n630_adj_4551), 
            .I3(n29342), .O(n10289[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5281_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5281_8_lut (.I0(GND_net), .I1(n10299[5]), .I2(n557_adj_4552), 
            .I3(n29341), .O(n10289[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5281_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5281_8 (.CI(n29341), .I0(n10299[5]), .I1(n557_adj_4552), 
            .CO(n29342));
    SB_LUT4 add_5281_7_lut (.I0(GND_net), .I1(n10299[4]), .I2(n484_adj_4553), 
            .I3(n29340), .O(n10289[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5281_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5281_7 (.CI(n29340), .I0(n10299[4]), .I1(n484_adj_4553), 
            .CO(n29341));
    SB_LUT4 add_5281_6_lut (.I0(GND_net), .I1(n10299[3]), .I2(n411_adj_4554), 
            .I3(n29339), .O(n10289[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5281_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5281_6 (.CI(n29339), .I0(n10299[3]), .I1(n411_adj_4554), 
            .CO(n29340));
    SB_CARRY add_751_13 (.CI(n27908), .I0(\PID_CONTROLLER.integral [11]), 
            .I1(n3302[11]), .CO(n27909));
    SB_LUT4 mult_10_i104_2_lut (.I0(\Kp[2] ), .I1(n28[2]), .I2(GND_net), 
            .I3(GND_net), .O(n153_adj_4555));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i104_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5281_5_lut (.I0(GND_net), .I1(n10299[2]), .I2(n338_adj_4556), 
            .I3(n29338), .O(n10289[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5281_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5281_5 (.CI(n29338), .I0(n10299[2]), .I1(n338_adj_4556), 
            .CO(n29339));
    SB_CARRY sub_3_add_2_12 (.CI(n27985), .I0(setpoint[10]), .I1(motor_state[10]), 
            .CO(n27986));
    SB_LUT4 add_751_12_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [10]), 
            .I2(n3302[10]), .I3(n27907), .O(\PID_CONTROLLER.integral_23__N_3546 [10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_751_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5281_4_lut (.I0(GND_net), .I1(n10299[1]), .I2(n265_adj_4557), 
            .I3(n29337), .O(n10289[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5281_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5281_4 (.CI(n29337), .I0(n10299[1]), .I1(n265_adj_4557), 
            .CO(n29338));
    SB_LUT4 add_5281_3_lut (.I0(GND_net), .I1(n10299[0]), .I2(n192_adj_4558), 
            .I3(n29336), .O(n10289[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5281_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_3_add_2_11_lut (.I0(GND_net), .I1(setpoint[9]), .I2(motor_state[9]), 
            .I3(n27984), .O(n28[9])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_3_add_2_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5281_3 (.CI(n29336), .I0(n10299[0]), .I1(n192_adj_4558), 
            .CO(n29337));
    SB_LUT4 add_5281_2_lut (.I0(GND_net), .I1(n50_adj_4559), .I2(n119_adj_4560), 
            .I3(GND_net), .O(n10289[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5281_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5281_2 (.CI(GND_net), .I0(n50_adj_4559), .I1(n119_adj_4560), 
            .CO(n29336));
    SB_CARRY add_751_12 (.CI(n27907), .I0(\PID_CONTROLLER.integral [10]), 
            .I1(n3302[10]), .CO(n27908));
    SB_LUT4 add_5280_10_lut (.I0(GND_net), .I1(n10289[7]), .I2(n700_adj_4561), 
            .I3(n29335), .O(n10278[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5280_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_751_11_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [9]), 
            .I2(n3302[9]), .I3(n27906), .O(\PID_CONTROLLER.integral_23__N_3546 [9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_751_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5280_9_lut (.I0(GND_net), .I1(n10289[6]), .I2(n627_adj_4562), 
            .I3(n29334), .O(n10278[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5280_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5280_9 (.CI(n29334), .I0(n10289[6]), .I1(n627_adj_4562), 
            .CO(n29335));
    SB_LUT4 add_5280_8_lut (.I0(GND_net), .I1(n10289[5]), .I2(n554_adj_4563), 
            .I3(n29333), .O(n10278[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5280_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5280_8 (.CI(n29333), .I0(n10289[5]), .I1(n554_adj_4563), 
            .CO(n29334));
    SB_LUT4 add_5280_7_lut (.I0(GND_net), .I1(n10289[4]), .I2(n481_adj_4564), 
            .I3(n29332), .O(n10278[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5280_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5280_7 (.CI(n29332), .I0(n10289[4]), .I1(n481_adj_4564), 
            .CO(n29333));
    SB_CARRY sub_3_add_2_11 (.CI(n27984), .I0(setpoint[9]), .I1(motor_state[9]), 
            .CO(n27985));
    SB_LUT4 sub_3_add_2_10_lut (.I0(GND_net), .I1(setpoint[8]), .I2(motor_state[8]), 
            .I3(n27983), .O(n28[8])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_3_add_2_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_3_add_2_10 (.CI(n27983), .I0(setpoint[8]), .I1(motor_state[8]), 
            .CO(n27984));
    SB_LUT4 sub_3_add_2_9_lut (.I0(GND_net), .I1(setpoint[7]), .I2(motor_state[7]), 
            .I3(n27982), .O(n28[7])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_3_add_2_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i153_2_lut (.I0(\Kp[3] ), .I1(n28[2]), .I2(GND_net), 
            .I3(GND_net), .O(n226_adj_4565));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i153_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5280_6_lut (.I0(GND_net), .I1(n10289[3]), .I2(n408_adj_4566), 
            .I3(n29331), .O(n10278[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5280_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i202_2_lut (.I0(\Kp[4] ), .I1(n28[2]), .I2(GND_net), 
            .I3(GND_net), .O(n299_adj_4567));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i202_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5280_6 (.CI(n29331), .I0(n10289[3]), .I1(n408_adj_4566), 
            .CO(n29332));
    SB_LUT4 add_5280_5_lut (.I0(GND_net), .I1(n10289[2]), .I2(n335_adj_4568), 
            .I3(n29330), .O(n10278[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5280_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5280_5 (.CI(n29330), .I0(n10289[2]), .I1(n335_adj_4568), 
            .CO(n29331));
    SB_CARRY add_751_11 (.CI(n27906), .I0(\PID_CONTROLLER.integral [9]), 
            .I1(n3302[9]), .CO(n27907));
    SB_LUT4 add_5280_4_lut (.I0(GND_net), .I1(n10289[1]), .I2(n262_adj_4569), 
            .I3(n29329), .O(n10278[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5280_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i251_2_lut (.I0(\Kp[5] ), .I1(n28[2]), .I2(GND_net), 
            .I3(GND_net), .O(n372_adj_4570));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i251_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5280_4 (.CI(n29329), .I0(n10289[1]), .I1(n262_adj_4569), 
            .CO(n29330));
    SB_LUT4 mult_10_i300_2_lut (.I0(\Kp[6] ), .I1(n28[2]), .I2(GND_net), 
            .I3(GND_net), .O(n445_adj_4571));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i300_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5280_3_lut (.I0(GND_net), .I1(n10289[0]), .I2(n189_adj_4572), 
            .I3(n29328), .O(n10278[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5280_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5280_3 (.CI(n29328), .I0(n10289[0]), .I1(n189_adj_4572), 
            .CO(n29329));
    SB_LUT4 mult_10_i349_2_lut (.I0(\Kp[7] ), .I1(n28[2]), .I2(GND_net), 
            .I3(GND_net), .O(n518_adj_4573));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i349_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i398_2_lut (.I0(\Kp[8] ), .I1(n28[2]), .I2(GND_net), 
            .I3(GND_net), .O(n591_adj_4574));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i398_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_751_10_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [8]), 
            .I2(n3302[8]), .I3(n27905), .O(\PID_CONTROLLER.integral_23__N_3546 [8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_751_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i447_2_lut (.I0(\Kp[9] ), .I1(n28[2]), .I2(GND_net), 
            .I3(GND_net), .O(n664_adj_4575));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i447_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5280_2_lut (.I0(GND_net), .I1(n47_adj_4576), .I2(n116_adj_4577), 
            .I3(GND_net), .O(n10278[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5280_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_751_10 (.CI(n27905), .I0(\PID_CONTROLLER.integral [8]), 
            .I1(n3302[8]), .CO(n27906));
    SB_LUT4 add_751_9_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [7]), 
            .I2(n3302[7]), .I3(n27904), .O(\PID_CONTROLLER.integral_23__N_3546 [7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_751_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i496_2_lut (.I0(\Kp[10] ), .I1(n28[2]), .I2(GND_net), 
            .I3(GND_net), .O(n737_adj_4578));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i496_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY sub_3_add_2_9 (.CI(n27982), .I0(setpoint[7]), .I1(motor_state[7]), 
            .CO(n27983));
    SB_CARRY add_5280_2 (.CI(GND_net), .I0(n47_adj_4576), .I1(n116_adj_4577), 
            .CO(n29328));
    SB_LUT4 mult_10_i545_2_lut (.I0(\Kp[11] ), .I1(n28[2]), .I2(GND_net), 
            .I3(GND_net), .O(n810_adj_4579));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i545_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 sub_3_add_2_8_lut (.I0(GND_net), .I1(setpoint[6]), .I2(motor_state[6]), 
            .I3(n27981), .O(n28[6])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_3_add_2_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5279_11_lut (.I0(GND_net), .I1(n10278[8]), .I2(n770_adj_4580), 
            .I3(n29327), .O(n10266[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5279_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_751_9 (.CI(n27904), .I0(\PID_CONTROLLER.integral [7]), 
            .I1(n3302[7]), .CO(n27905));
    SB_LUT4 add_5279_10_lut (.I0(GND_net), .I1(n10278[7]), .I2(n697_adj_4581), 
            .I3(n29326), .O(n10266[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5279_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5279_10 (.CI(n29326), .I0(n10278[7]), .I1(n697_adj_4581), 
            .CO(n29327));
    SB_LUT4 add_5279_9_lut (.I0(GND_net), .I1(n10278[6]), .I2(n624_adj_4582), 
            .I3(n29325), .O(n10266[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5279_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i594_2_lut (.I0(\Kp[12] ), .I1(n28[2]), .I2(GND_net), 
            .I3(GND_net), .O(n883_adj_4583));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i594_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5279_9 (.CI(n29325), .I0(n10278[6]), .I1(n624_adj_4582), 
            .CO(n29326));
    SB_LUT4 add_5279_8_lut (.I0(GND_net), .I1(n10278[5]), .I2(n551_adj_4584), 
            .I3(n29324), .O(n10266[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5279_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5279_8 (.CI(n29324), .I0(n10278[5]), .I1(n551_adj_4584), 
            .CO(n29325));
    SB_LUT4 add_5279_7_lut (.I0(GND_net), .I1(n10278[4]), .I2(n478_adj_4585), 
            .I3(n29323), .O(n10266[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5279_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5279_7 (.CI(n29323), .I0(n10278[4]), .I1(n478_adj_4585), 
            .CO(n29324));
    SB_LUT4 add_5279_6_lut (.I0(GND_net), .I1(n10278[3]), .I2(n405_adj_4586), 
            .I3(n29322), .O(n10266[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5279_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5279_6 (.CI(n29322), .I0(n10278[3]), .I1(n405_adj_4586), 
            .CO(n29323));
    SB_LUT4 add_5279_5_lut (.I0(GND_net), .I1(n10278[2]), .I2(n332_adj_4587), 
            .I3(n29321), .O(n10266[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5279_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5279_5 (.CI(n29321), .I0(n10278[2]), .I1(n332_adj_4587), 
            .CO(n29322));
    SB_LUT4 add_5279_4_lut (.I0(GND_net), .I1(n10278[1]), .I2(n259_adj_4588), 
            .I3(n29320), .O(n10266[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5279_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5279_4 (.CI(n29320), .I0(n10278[1]), .I1(n259_adj_4588), 
            .CO(n29321));
    SB_LUT4 add_5279_3_lut (.I0(GND_net), .I1(n10278[0]), .I2(n186_adj_4589), 
            .I3(n29319), .O(n10266[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5279_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i643_2_lut (.I0(\Kp[13] ), .I1(n28[2]), .I2(GND_net), 
            .I3(GND_net), .O(n956_adj_4590));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i643_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5279_3 (.CI(n29319), .I0(n10278[0]), .I1(n186_adj_4589), 
            .CO(n29320));
    SB_LUT4 add_5279_2_lut (.I0(GND_net), .I1(n44_adj_4591), .I2(n113_adj_4592), 
            .I3(GND_net), .O(n10266[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5279_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5279_2 (.CI(GND_net), .I0(n44_adj_4591), .I1(n113_adj_4592), 
            .CO(n29319));
    SB_LUT4 add_5278_12_lut (.I0(GND_net), .I1(n10266[9]), .I2(n840_adj_4593), 
            .I3(n29318), .O(n10253[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5278_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5278_11_lut (.I0(GND_net), .I1(n10266[8]), .I2(n767_adj_4594), 
            .I3(n29317), .O(n10253[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5278_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5278_11 (.CI(n29317), .I0(n10266[8]), .I1(n767_adj_4594), 
            .CO(n29318));
    SB_LUT4 add_5278_10_lut (.I0(GND_net), .I1(n10266[7]), .I2(n694_adj_4595), 
            .I3(n29316), .O(n10253[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5278_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5278_10 (.CI(n29316), .I0(n10266[7]), .I1(n694_adj_4595), 
            .CO(n29317));
    SB_LUT4 add_5278_9_lut (.I0(GND_net), .I1(n10266[6]), .I2(n621_adj_4596), 
            .I3(n29315), .O(n10253[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5278_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5278_9 (.CI(n29315), .I0(n10266[6]), .I1(n621_adj_4596), 
            .CO(n29316));
    SB_LUT4 add_5278_8_lut (.I0(GND_net), .I1(n10266[5]), .I2(n548_adj_4597), 
            .I3(n29314), .O(n10253[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5278_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5278_8 (.CI(n29314), .I0(n10266[5]), .I1(n548_adj_4597), 
            .CO(n29315));
    SB_LUT4 add_5278_7_lut (.I0(GND_net), .I1(n10266[4]), .I2(n475_adj_4598), 
            .I3(n29313), .O(n10253[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5278_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5278_7 (.CI(n29313), .I0(n10266[4]), .I1(n475_adj_4598), 
            .CO(n29314));
    SB_LUT4 add_5278_6_lut (.I0(GND_net), .I1(n10266[3]), .I2(n402_adj_4599), 
            .I3(n29312), .O(n10253[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5278_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5278_6 (.CI(n29312), .I0(n10266[3]), .I1(n402_adj_4599), 
            .CO(n29313));
    SB_LUT4 add_5278_5_lut (.I0(GND_net), .I1(n10266[2]), .I2(n329_adj_4600), 
            .I3(n29311), .O(n10253[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5278_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5278_5 (.CI(n29311), .I0(n10266[2]), .I1(n329_adj_4600), 
            .CO(n29312));
    SB_LUT4 add_5278_4_lut (.I0(GND_net), .I1(n10266[1]), .I2(n256_adj_4601), 
            .I3(n29310), .O(n10253[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5278_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5278_4 (.CI(n29310), .I0(n10266[1]), .I1(n256_adj_4601), 
            .CO(n29311));
    SB_LUT4 add_5278_3_lut (.I0(GND_net), .I1(n10266[0]), .I2(n183_adj_4602), 
            .I3(n29309), .O(n10253[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5278_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5278_3 (.CI(n29309), .I0(n10266[0]), .I1(n183_adj_4602), 
            .CO(n29310));
    SB_LUT4 add_5278_2_lut (.I0(GND_net), .I1(n41_adj_4603), .I2(n110_adj_4604), 
            .I3(GND_net), .O(n10253[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5278_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5278_2 (.CI(GND_net), .I0(n41_adj_4603), .I1(n110_adj_4604), 
            .CO(n29309));
    SB_LUT4 add_5277_13_lut (.I0(GND_net), .I1(n10253[10]), .I2(n910_adj_4605), 
            .I3(n29308), .O(n10239[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5277_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5277_12_lut (.I0(GND_net), .I1(n10253[9]), .I2(n837_adj_4606), 
            .I3(n29307), .O(n10239[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5277_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5277_12 (.CI(n29307), .I0(n10253[9]), .I1(n837_adj_4606), 
            .CO(n29308));
    SB_LUT4 add_5277_11_lut (.I0(GND_net), .I1(n10253[8]), .I2(n764_adj_4607), 
            .I3(n29306), .O(n10239[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5277_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5277_11 (.CI(n29306), .I0(n10253[8]), .I1(n764_adj_4607), 
            .CO(n29307));
    SB_LUT4 add_5277_10_lut (.I0(GND_net), .I1(n10253[7]), .I2(n691_adj_4608), 
            .I3(n29305), .O(n10239[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5277_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5277_10 (.CI(n29305), .I0(n10253[7]), .I1(n691_adj_4608), 
            .CO(n29306));
    SB_LUT4 add_5277_9_lut (.I0(GND_net), .I1(n10253[6]), .I2(n618_adj_4609), 
            .I3(n29304), .O(n10239[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5277_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i692_2_lut (.I0(\Kp[14] ), .I1(n28[2]), .I2(GND_net), 
            .I3(GND_net), .O(n1029_adj_4610));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i692_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5277_9 (.CI(n29304), .I0(n10253[6]), .I1(n618_adj_4609), 
            .CO(n29305));
    SB_CARRY sub_3_add_2_8 (.CI(n27981), .I0(setpoint[6]), .I1(motor_state[6]), 
            .CO(n27982));
    SB_LUT4 add_5277_8_lut (.I0(GND_net), .I1(n10253[5]), .I2(n545_adj_4611), 
            .I3(n29303), .O(n10239[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5277_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5277_8 (.CI(n29303), .I0(n10253[5]), .I1(n545_adj_4611), 
            .CO(n29304));
    SB_LUT4 add_5277_7_lut (.I0(GND_net), .I1(n10253[4]), .I2(n472_adj_4612), 
            .I3(n29302), .O(n10239[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5277_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5277_7 (.CI(n29302), .I0(n10253[4]), .I1(n472_adj_4612), 
            .CO(n29303));
    SB_LUT4 add_751_8_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [6]), 
            .I2(n3302[6]), .I3(n27903), .O(\PID_CONTROLLER.integral_23__N_3546 [6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_751_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_751_8 (.CI(n27903), .I0(\PID_CONTROLLER.integral [6]), 
            .I1(n3302[6]), .CO(n27904));
    SB_LUT4 mult_10_i741_2_lut (.I0(\Kp[15] ), .I1(n28[2]), .I2(GND_net), 
            .I3(GND_net), .O(n1102_adj_4613));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i741_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 sub_3_add_2_7_lut (.I0(GND_net), .I1(setpoint[5]), .I2(motor_state[5]), 
            .I3(n27980), .O(n28[5])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_3_add_2_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5277_6_lut (.I0(GND_net), .I1(n10253[3]), .I2(n399_adj_4614), 
            .I3(n29301), .O(n10239[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5277_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_3_add_2_7 (.CI(n27980), .I0(setpoint[5]), .I1(motor_state[5]), 
            .CO(n27981));
    SB_CARRY add_5277_6 (.CI(n29301), .I0(n10253[3]), .I1(n399_adj_4614), 
            .CO(n29302));
    SB_LUT4 add_5277_5_lut (.I0(GND_net), .I1(n10253[2]), .I2(n326_adj_4615), 
            .I3(n29300), .O(n10239[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5277_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_3_add_2_6_lut (.I0(GND_net), .I1(setpoint[4]), .I2(motor_state[4]), 
            .I3(n27979), .O(n28[4])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_3_add_2_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_3_add_2_6 (.CI(n27979), .I0(setpoint[4]), .I1(motor_state[4]), 
            .CO(n27980));
    SB_CARRY add_5277_5 (.CI(n29300), .I0(n10253[2]), .I1(n326_adj_4615), 
            .CO(n29301));
    SB_LUT4 add_751_7_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [5]), 
            .I2(n3302[5]), .I3(n27902), .O(\PID_CONTROLLER.integral_23__N_3546 [5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_751_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_3_add_2_5_lut (.I0(GND_net), .I1(setpoint[3]), .I2(motor_state[3]), 
            .I3(n27978), .O(n28[3])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_3_add_2_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_3_add_2_5 (.CI(n27978), .I0(setpoint[3]), .I1(motor_state[3]), 
            .CO(n27979));
    SB_LUT4 add_5277_4_lut (.I0(GND_net), .I1(n10253[1]), .I2(n253_adj_4617), 
            .I3(n29299), .O(n10239[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5277_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_3_add_2_4_lut (.I0(GND_net), .I1(setpoint[2]), .I2(motor_state[2]), 
            .I3(n27977), .O(n28[2])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_3_add_2_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_5_inv_0_i20_1_lut (.I0(IntegralLimit[19]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[19]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i20_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_5277_4 (.CI(n29299), .I0(n10253[1]), .I1(n253_adj_4617), 
            .CO(n29300));
    SB_CARRY add_751_7 (.CI(n27902), .I0(\PID_CONTROLLER.integral [5]), 
            .I1(n3302[5]), .CO(n27903));
    SB_LUT4 add_751_6_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [4]), 
            .I2(n3302[4]), .I3(n27901), .O(\PID_CONTROLLER.integral_23__N_3546 [4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_751_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_3_add_2_4 (.CI(n27977), .I0(setpoint[2]), .I1(motor_state[2]), 
            .CO(n27978));
    SB_LUT4 add_5277_3_lut (.I0(GND_net), .I1(n10253[0]), .I2(n180_adj_4618), 
            .I3(n29298), .O(n10239[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5277_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5277_3 (.CI(n29298), .I0(n10253[0]), .I1(n180_adj_4618), 
            .CO(n29299));
    SB_LUT4 add_5277_2_lut (.I0(GND_net), .I1(n38_adj_4619), .I2(n107_adj_4620), 
            .I3(GND_net), .O(n10239[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5277_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_751_6 (.CI(n27901), .I0(\PID_CONTROLLER.integral [4]), 
            .I1(n3302[4]), .CO(n27902));
    SB_CARRY add_5277_2 (.CI(GND_net), .I0(n38_adj_4619), .I1(n107_adj_4620), 
            .CO(n29298));
    SB_LUT4 add_5276_14_lut (.I0(GND_net), .I1(n10239[11]), .I2(n980_adj_4621), 
            .I3(n29297), .O(n10224[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5276_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5276_13_lut (.I0(GND_net), .I1(n10239[10]), .I2(n907_adj_4622), 
            .I3(n29296), .O(n10224[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5276_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_3_add_2_3_lut (.I0(GND_net), .I1(setpoint[1]), .I2(motor_state[1]), 
            .I3(n27976), .O(n28[1])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_3_add_2_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5276_13 (.CI(n29296), .I0(n10239[10]), .I1(n907_adj_4622), 
            .CO(n29297));
    SB_LUT4 add_751_5_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [3]), 
            .I2(n3302[3]), .I3(n27900), .O(\PID_CONTROLLER.integral_23__N_3546 [3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_751_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 duty_23__I_831_i39_2_lut (.I0(PWMLimit[19]), .I1(duty_23__N_3646[19]), 
            .I2(GND_net), .I3(GND_net), .O(n39_adj_4623));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_831_i39_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_831_i41_2_lut (.I0(PWMLimit[20]), .I1(duty_23__N_3646[20]), 
            .I2(GND_net), .I3(GND_net), .O(n41_adj_4624));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_831_i41_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 unary_minus_5_inv_0_i22_1_lut (.I0(IntegralLimit[21]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[21]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i22_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 duty_23__I_831_i45_2_lut (.I0(PWMLimit[22]), .I1(duty_23__N_3646[22]), 
            .I2(GND_net), .I3(GND_net), .O(n45_adj_4625));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_831_i45_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_831_i37_2_lut (.I0(PWMLimit[18]), .I1(duty_23__N_3646[18]), 
            .I2(GND_net), .I3(GND_net), .O(n37_adj_4626));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_831_i37_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_831_i29_2_lut (.I0(PWMLimit[14]), .I1(duty_23__N_3646[14]), 
            .I2(GND_net), .I3(GND_net), .O(n29_adj_4627));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_831_i29_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_831_i31_2_lut (.I0(PWMLimit[15]), .I1(duty_23__N_3646[15]), 
            .I2(GND_net), .I3(GND_net), .O(n31_adj_4628));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_831_i31_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_831_i43_2_lut (.I0(PWMLimit[21]), .I1(duty_23__N_3646[21]), 
            .I2(GND_net), .I3(GND_net), .O(n43_adj_4629));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_831_i43_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_831_i23_2_lut (.I0(PWMLimit[11]), .I1(duty_23__N_3646[11]), 
            .I2(GND_net), .I3(GND_net), .O(n23_adj_4630));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_831_i23_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_831_i25_2_lut (.I0(PWMLimit[12]), .I1(duty_23__N_3646[12]), 
            .I2(GND_net), .I3(GND_net), .O(n25_adj_4631));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_831_i25_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_831_i35_2_lut (.I0(PWMLimit[17]), .I1(duty_23__N_3646[17]), 
            .I2(GND_net), .I3(GND_net), .O(n35_adj_4632));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_831_i35_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_831_i11_2_lut (.I0(PWMLimit[5]), .I1(duty_23__N_3646[5]), 
            .I2(GND_net), .I3(GND_net), .O(n11_adj_4633));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_831_i11_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_831_i13_2_lut (.I0(PWMLimit[6]), .I1(duty_23__N_3646[6]), 
            .I2(GND_net), .I3(GND_net), .O(n13_adj_4634));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_831_i13_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_831_i15_2_lut (.I0(PWMLimit[7]), .I1(duty_23__N_3646[7]), 
            .I2(GND_net), .I3(GND_net), .O(n15_adj_4635));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_831_i15_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_831_i27_2_lut (.I0(PWMLimit[13]), .I1(duty_23__N_3646[13]), 
            .I2(GND_net), .I3(GND_net), .O(n27_adj_4636));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_831_i27_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_831_i33_2_lut (.I0(PWMLimit[16]), .I1(duty_23__N_3646[16]), 
            .I2(GND_net), .I3(GND_net), .O(n33_adj_4637));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_831_i33_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_831_i9_2_lut (.I0(PWMLimit[4]), .I1(duty_23__N_3646[4]), 
            .I2(GND_net), .I3(GND_net), .O(n9_adj_4638));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_831_i9_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_831_i17_2_lut (.I0(PWMLimit[8]), .I1(duty_23__N_3646[8]), 
            .I2(GND_net), .I3(GND_net), .O(n17_adj_4639));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_831_i17_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_831_i19_2_lut (.I0(PWMLimit[9]), .I1(duty_23__N_3646[9]), 
            .I2(GND_net), .I3(GND_net), .O(n19_adj_4640));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_831_i19_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_831_i21_2_lut (.I0(PWMLimit[10]), .I1(duty_23__N_3646[10]), 
            .I2(GND_net), .I3(GND_net), .O(n21_adj_4641));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_831_i21_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i29677_4_lut (.I0(n21_adj_4641), .I1(n19_adj_4640), .I2(n17_adj_4639), 
            .I3(n9_adj_4638), .O(n36432));
    defparam i29677_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i29671_4_lut (.I0(n27_adj_4636), .I1(n15_adj_4635), .I2(n13_adj_4634), 
            .I3(n11_adj_4633), .O(n36426));
    defparam i29671_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 duty_23__I_831_i12_3_lut (.I0(duty_23__N_3646[7]), .I1(duty_23__N_3646[16]), 
            .I2(n33_adj_4637), .I3(GND_net), .O(n12_adj_4642));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_831_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_831_i10_3_lut (.I0(duty_23__N_3646[5]), .I1(duty_23__N_3646[6]), 
            .I2(n13_adj_4634), .I3(GND_net), .O(n10_adj_4643));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_831_i10_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_831_i30_3_lut (.I0(n12_adj_4642), .I1(duty_23__N_3646[17]), 
            .I2(n35_adj_4632), .I3(GND_net), .O(n30_adj_4644));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_831_i30_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_5276_12_lut (.I0(GND_net), .I1(n10239[9]), .I2(n834_adj_4532), 
            .I3(n29295), .O(n10224[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5276_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i29951_4_lut (.I0(n13_adj_4634), .I1(n11_adj_4633), .I2(n9_adj_4638), 
            .I3(n36442), .O(n36706));
    defparam i29951_4_lut.LUT_INIT = 16'heeef;
    SB_CARRY add_5276_12 (.CI(n29295), .I0(n10239[9]), .I1(n834_adj_4532), 
            .CO(n29296));
    SB_LUT4 i29947_4_lut (.I0(n19_adj_4640), .I1(n17_adj_4639), .I2(n15_adj_4635), 
            .I3(n36706), .O(n36702));
    defparam i29947_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i30243_4_lut (.I0(n25_adj_4631), .I1(n23_adj_4630), .I2(n21_adj_4641), 
            .I3(n36702), .O(n36998));
    defparam i30243_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 add_5276_11_lut (.I0(GND_net), .I1(n10239[8]), .I2(n761_adj_4531), 
            .I3(n29294), .O(n10224[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5276_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i30087_4_lut (.I0(n31_adj_4628), .I1(n29_adj_4627), .I2(n27_adj_4636), 
            .I3(n36998), .O(n36842));
    defparam i30087_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i30308_4_lut (.I0(n37_adj_4626), .I1(n35_adj_4632), .I2(n33_adj_4637), 
            .I3(n36842), .O(n37063));
    defparam i30308_4_lut.LUT_INIT = 16'hfffe;
    SB_CARRY add_5276_11 (.CI(n29294), .I0(n10239[8]), .I1(n761_adj_4531), 
            .CO(n29295));
    SB_LUT4 duty_23__I_831_i16_3_lut (.I0(duty_23__N_3646[9]), .I1(duty_23__N_3646[21]), 
            .I2(n43_adj_4629), .I3(GND_net), .O(n16_adj_4645));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_831_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_5276_10_lut (.I0(GND_net), .I1(n10239[7]), .I2(n688_adj_4529), 
            .I3(n29293), .O(n10224[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5276_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i30229_3_lut (.I0(n6_adj_4646), .I1(duty_23__N_3646[10]), .I2(n21_adj_4641), 
            .I3(GND_net), .O(n36984));   // verilog/motorControl.v(36[10:25])
    defparam i30229_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i30230_3_lut (.I0(n36984), .I1(duty_23__N_3646[11]), .I2(n23_adj_4630), 
            .I3(GND_net), .O(n36985));   // verilog/motorControl.v(36[10:25])
    defparam i30230_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_5276_10 (.CI(n29293), .I0(n10239[7]), .I1(n688_adj_4529), 
            .CO(n29294));
    SB_LUT4 duty_23__I_831_i8_3_lut (.I0(duty_23__N_3646[4]), .I1(duty_23__N_3646[8]), 
            .I2(n17_adj_4639), .I3(GND_net), .O(n8_adj_4647));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_831_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_5276_9_lut (.I0(GND_net), .I1(n10239[6]), .I2(n615_adj_4528), 
            .I3(n29292), .O(n10224[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5276_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 duty_23__I_831_i24_3_lut (.I0(n16_adj_4645), .I1(duty_23__N_3646[22]), 
            .I2(n45_adj_4625), .I3(GND_net), .O(n24_adj_4648));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_831_i24_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i29657_4_lut (.I0(n43_adj_4629), .I1(n25_adj_4631), .I2(n23_adj_4630), 
            .I3(n36432), .O(n36412));
    defparam i29657_4_lut.LUT_INIT = 16'haaab;
    SB_CARRY add_5276_9 (.CI(n29292), .I0(n10239[6]), .I1(n615_adj_4528), 
            .CO(n29293));
    SB_LUT4 i30119_4_lut (.I0(n24_adj_4648), .I1(n8_adj_4647), .I2(n45_adj_4625), 
            .I3(n36410), .O(n36874));   // verilog/motorControl.v(36[10:25])
    defparam i30119_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i30176_3_lut (.I0(n36985), .I1(duty_23__N_3646[12]), .I2(n25_adj_4631), 
            .I3(GND_net), .O(n36931));   // verilog/motorControl.v(36[10:25])
    defparam i30176_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_5276_8_lut (.I0(GND_net), .I1(n10239[5]), .I2(n542_adj_4527), 
            .I3(n29291), .O(n10224[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5276_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 duty_23__I_831_i4_4_lut (.I0(duty_23__N_3646[0]), .I1(duty_23__N_3646[1]), 
            .I2(PWMLimit[1]), .I3(PWMLimit[0]), .O(n4_adj_4649));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_831_i4_4_lut.LUT_INIT = 16'h0c8e;
    SB_LUT4 i30221_3_lut (.I0(n4_adj_4649), .I1(duty_23__N_3646[13]), .I2(n27_adj_4636), 
            .I3(GND_net), .O(n36976));   // verilog/motorControl.v(36[10:25])
    defparam i30221_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_5276_8 (.CI(n29291), .I0(n10239[5]), .I1(n542_adj_4527), 
            .CO(n29292));
    SB_LUT4 i30222_3_lut (.I0(n36976), .I1(duty_23__N_3646[14]), .I2(n29_adj_4627), 
            .I3(GND_net), .O(n36977));   // verilog/motorControl.v(36[10:25])
    defparam i30222_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i29667_4_lut (.I0(n33_adj_4637), .I1(n31_adj_4628), .I2(n29_adj_4627), 
            .I3(n36426), .O(n36422));
    defparam i29667_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 add_5276_7_lut (.I0(GND_net), .I1(n10239[4]), .I2(n469_adj_4526), 
            .I3(n29290), .O(n10224[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5276_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i30318_4_lut (.I0(n30_adj_4644), .I1(n10_adj_4643), .I2(n35_adj_4632), 
            .I3(n36420), .O(n37073));   // verilog/motorControl.v(36[10:25])
    defparam i30318_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i30178_3_lut (.I0(n36977), .I1(duty_23__N_3646[15]), .I2(n31_adj_4628), 
            .I3(GND_net), .O(n36933));   // verilog/motorControl.v(36[10:25])
    defparam i30178_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_5276_7 (.CI(n29290), .I0(n10239[4]), .I1(n469_adj_4526), 
            .CO(n29291));
    SB_LUT4 i30367_4_lut (.I0(n36933), .I1(n37073), .I2(n35_adj_4632), 
            .I3(n36422), .O(n37122));   // verilog/motorControl.v(36[10:25])
    defparam i30367_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i30368_3_lut (.I0(n37122), .I1(duty_23__N_3646[18]), .I2(n37_adj_4626), 
            .I3(GND_net), .O(n37123));   // verilog/motorControl.v(36[10:25])
    defparam i30368_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_5276_6_lut (.I0(GND_net), .I1(n10239[3]), .I2(n396_adj_4525), 
            .I3(n29289), .O(n10224[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5276_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i30349_3_lut (.I0(n37123), .I1(duty_23__N_3646[19]), .I2(n39_adj_4623), 
            .I3(GND_net), .O(n37104));   // verilog/motorControl.v(36[10:25])
    defparam i30349_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i29659_4_lut (.I0(n43_adj_4629), .I1(n41_adj_4624), .I2(n39_adj_4623), 
            .I3(n37063), .O(n36414));
    defparam i29659_4_lut.LUT_INIT = 16'haaab;
    SB_CARRY add_5276_6 (.CI(n29289), .I0(n10239[3]), .I1(n396_adj_4525), 
            .CO(n29290));
    SB_LUT4 i30273_4_lut (.I0(n36931), .I1(n36874), .I2(n45_adj_4625), 
            .I3(n36412), .O(n37028));   // verilog/motorControl.v(36[10:25])
    defparam i30273_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i30337_3_lut (.I0(n37104), .I1(duty_23__N_3646[20]), .I2(n41_adj_4624), 
            .I3(GND_net), .O(n40_adj_4650));   // verilog/motorControl.v(36[10:25])
    defparam i30337_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_5276_5_lut (.I0(GND_net), .I1(n10239[2]), .I2(n323_adj_4524), 
            .I3(n29288), .O(n10224[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5276_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i30275_4_lut (.I0(n40_adj_4650), .I1(n37028), .I2(n45_adj_4625), 
            .I3(n36414), .O(n37030));   // verilog/motorControl.v(36[10:25])
    defparam i30275_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i30276_3_lut (.I0(n37030), .I1(PWMLimit[23]), .I2(duty_23__N_3646[23]), 
            .I3(GND_net), .O(duty_23__N_3645));   // verilog/motorControl.v(36[10:25])
    defparam i30276_3_lut.LUT_INIT = 16'h8e8e;
    SB_CARRY add_5276_5 (.CI(n29288), .I0(n10239[2]), .I1(n323_adj_4524), 
            .CO(n29289));
    SB_LUT4 add_5276_4_lut (.I0(GND_net), .I1(n10239[1]), .I2(n250_adj_4523), 
            .I3(n29287), .O(n10224[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5276_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_15_i41_2_lut (.I0(duty_23__N_3646[20]), .I1(n257[20]), 
            .I2(GND_net), .I3(GND_net), .O(n41_adj_4651));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i41_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_5276_4 (.CI(n29287), .I0(n10239[1]), .I1(n250_adj_4523), 
            .CO(n29288));
    SB_LUT4 LessThan_15_i39_2_lut (.I0(duty_23__N_3646[19]), .I1(n257[19]), 
            .I2(GND_net), .I3(GND_net), .O(n39_adj_4652));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i39_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_5276_3_lut (.I0(GND_net), .I1(n10239[0]), .I2(n177_adj_4522), 
            .I3(n29286), .O(n10224[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5276_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_15_i45_2_lut (.I0(duty_23__N_3646[22]), .I1(n257[22]), 
            .I2(GND_net), .I3(GND_net), .O(n45_adj_4653));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i45_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_5276_3 (.CI(n29286), .I0(n10239[0]), .I1(n177_adj_4522), 
            .CO(n29287));
    SB_LUT4 add_5276_2_lut (.I0(GND_net), .I1(n35_adj_4521), .I2(n104_adj_4520), 
            .I3(GND_net), .O(n10224[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5276_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_15_i43_2_lut (.I0(duty_23__N_3646[21]), .I1(n257[21]), 
            .I2(GND_net), .I3(GND_net), .O(n43_adj_4654));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i43_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_5276_2 (.CI(GND_net), .I0(n35_adj_4521), .I1(n104_adj_4520), 
            .CO(n29286));
    SB_LUT4 LessThan_15_i37_2_lut (.I0(duty_23__N_3646[18]), .I1(n257[18]), 
            .I2(GND_net), .I3(GND_net), .O(n37_adj_4655));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i37_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_5275_15_lut (.I0(GND_net), .I1(n10224[12]), .I2(n1050_adj_4519), 
            .I3(n29285), .O(n10208[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5275_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5275_14_lut (.I0(GND_net), .I1(n10224[11]), .I2(n977_adj_4517), 
            .I3(n29284), .O(n10208[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5275_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_15_i29_2_lut (.I0(duty_23__N_3646[14]), .I1(n257[14]), 
            .I2(GND_net), .I3(GND_net), .O(n29_adj_4656));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i29_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_5275_14 (.CI(n29284), .I0(n10224[11]), .I1(n977_adj_4517), 
            .CO(n29285));
    SB_LUT4 LessThan_15_i31_2_lut (.I0(duty_23__N_3646[15]), .I1(n257[15]), 
            .I2(GND_net), .I3(GND_net), .O(n31_adj_4657));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i31_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_5275_13_lut (.I0(GND_net), .I1(n10224[10]), .I2(n904_adj_4516), 
            .I3(n29283), .O(n10208[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5275_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_15_i23_2_lut (.I0(duty_23__N_3646[11]), .I1(n257[11]), 
            .I2(GND_net), .I3(GND_net), .O(n23_adj_4658));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i23_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_5275_13 (.CI(n29283), .I0(n10224[10]), .I1(n904_adj_4516), 
            .CO(n29284));
    SB_LUT4 LessThan_15_i25_2_lut (.I0(duty_23__N_3646[12]), .I1(n257[12]), 
            .I2(GND_net), .I3(GND_net), .O(n25_adj_4659));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i25_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_5275_12_lut (.I0(GND_net), .I1(n10224[9]), .I2(n831_adj_4515), 
            .I3(n29282), .O(n10208[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5275_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5275_12 (.CI(n29282), .I0(n10224[9]), .I1(n831_adj_4515), 
            .CO(n29283));
    SB_LUT4 LessThan_15_i35_2_lut (.I0(duty_23__N_3646[17]), .I1(n257[17]), 
            .I2(GND_net), .I3(GND_net), .O(n35_adj_4660));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i35_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_5275_11_lut (.I0(GND_net), .I1(n10224[8]), .I2(n758_adj_4514), 
            .I3(n29281), .O(n10208[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5275_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_15_i33_2_lut (.I0(duty_23__N_3646[16]), .I1(n257[16]), 
            .I2(GND_net), .I3(GND_net), .O(n33_adj_4661));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i33_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_5275_11 (.CI(n29281), .I0(n10224[8]), .I1(n758_adj_4514), 
            .CO(n29282));
    SB_LUT4 LessThan_15_i11_2_lut (.I0(duty_23__N_3646[5]), .I1(n257[5]), 
            .I2(GND_net), .I3(GND_net), .O(n11_adj_4662));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i11_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_5275_10_lut (.I0(GND_net), .I1(n10224[7]), .I2(n685_adj_4512), 
            .I3(n29280), .O(n10208[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5275_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_15_i13_2_lut (.I0(duty_23__N_3646[6]), .I1(n257[6]), 
            .I2(GND_net), .I3(GND_net), .O(n13_adj_4663));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i13_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_5275_10 (.CI(n29280), .I0(n10224[7]), .I1(n685_adj_4512), 
            .CO(n29281));
    SB_LUT4 add_5275_9_lut (.I0(GND_net), .I1(n10224[6]), .I2(n612_adj_4511), 
            .I3(n29279), .O(n10208[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5275_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5275_9 (.CI(n29279), .I0(n10224[6]), .I1(n612_adj_4511), 
            .CO(n29280));
    SB_LUT4 LessThan_15_i15_2_lut (.I0(duty_23__N_3646[7]), .I1(n257[7]), 
            .I2(GND_net), .I3(GND_net), .O(n15_adj_4664));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i15_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_15_i27_2_lut (.I0(duty_23__N_3646[13]), .I1(n257[13]), 
            .I2(GND_net), .I3(GND_net), .O(n27_adj_4665));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i27_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_15_i9_2_lut (.I0(duty_23__N_3646[4]), .I1(n257[4]), 
            .I2(GND_net), .I3(GND_net), .O(n9_adj_4666));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i9_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_15_i17_2_lut (.I0(duty_23__N_3646[8]), .I1(n257[8]), 
            .I2(GND_net), .I3(GND_net), .O(n17_adj_4667));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i17_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_15_i19_2_lut (.I0(duty_23__N_3646[9]), .I1(n257[9]), 
            .I2(GND_net), .I3(GND_net), .O(n19_adj_4668));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i19_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_15_i21_2_lut (.I0(duty_23__N_3646[10]), .I1(n257[10]), 
            .I2(GND_net), .I3(GND_net), .O(n21_adj_4669));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i21_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i29643_4_lut (.I0(n21_adj_4669), .I1(n19_adj_4668), .I2(n17_adj_4667), 
            .I3(n9_adj_4666), .O(n36398));
    defparam i29643_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i29637_4_lut (.I0(n27_adj_4665), .I1(n15_adj_4664), .I2(n13_adj_4663), 
            .I3(n11_adj_4662), .O(n36392));
    defparam i29637_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 LessThan_15_i12_3_lut (.I0(n257[7]), .I1(n257[16]), .I2(n33_adj_4661), 
            .I3(GND_net), .O(n12_adj_4670));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_15_i10_3_lut (.I0(n257[5]), .I1(n257[6]), .I2(n13_adj_4663), 
            .I3(GND_net), .O(n10_adj_4671));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i10_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_5275_8_lut (.I0(GND_net), .I1(n10224[5]), .I2(n539_adj_4510), 
            .I3(n29278), .O(n10208[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5275_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_15_i30_3_lut (.I0(n12_adj_4670), .I1(n257[17]), .I2(n35_adj_4660), 
            .I3(GND_net), .O(n30_adj_4672));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i30_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i29919_4_lut (.I0(n13_adj_4663), .I1(n11_adj_4662), .I2(n9_adj_4666), 
            .I3(n36408), .O(n36674));
    defparam i29919_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i29915_4_lut (.I0(n19_adj_4668), .I1(n17_adj_4667), .I2(n15_adj_4664), 
            .I3(n36674), .O(n36670));
    defparam i29915_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i30235_4_lut (.I0(n25_adj_4659), .I1(n23_adj_4658), .I2(n21_adj_4669), 
            .I3(n36670), .O(n36990));
    defparam i30235_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i30071_4_lut (.I0(n31_adj_4657), .I1(n29_adj_4656), .I2(n27_adj_4665), 
            .I3(n36990), .O(n36826));
    defparam i30071_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i30306_4_lut (.I0(n37_adj_4655), .I1(n35_adj_4660), .I2(n33_adj_4661), 
            .I3(n36826), .O(n37061));
    defparam i30306_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 LessThan_15_i16_3_lut (.I0(n257[9]), .I1(n257[21]), .I2(n43_adj_4654), 
            .I3(GND_net), .O(n16_adj_4673));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i30217_3_lut (.I0(n6_adj_4674), .I1(n257[10]), .I2(n21_adj_4669), 
            .I3(GND_net), .O(n36972));   // verilog/motorControl.v(38[19:35])
    defparam i30217_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i30218_3_lut (.I0(n36972), .I1(n257[11]), .I2(n23_adj_4658), 
            .I3(GND_net), .O(n36973));   // verilog/motorControl.v(38[19:35])
    defparam i30218_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_5275_8 (.CI(n29278), .I0(n10224[5]), .I1(n539_adj_4510), 
            .CO(n29279));
    SB_LUT4 add_5275_7_lut (.I0(GND_net), .I1(n10224[4]), .I2(n466_adj_4509), 
            .I3(n29277), .O(n10208[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5275_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_15_i8_3_lut (.I0(n257[4]), .I1(n257[8]), .I2(n17_adj_4667), 
            .I3(GND_net), .O(n8_adj_4675));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_15_i24_3_lut (.I0(n16_adj_4673), .I1(n257[22]), .I2(n45_adj_4653), 
            .I3(GND_net), .O(n24_adj_4676));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i24_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i29620_4_lut (.I0(n43_adj_4654), .I1(n25_adj_4659), .I2(n23_adj_4658), 
            .I3(n36398), .O(n36375));
    defparam i29620_4_lut.LUT_INIT = 16'haaab;
    SB_CARRY add_5275_7 (.CI(n29277), .I0(n10224[4]), .I1(n466_adj_4509), 
            .CO(n29278));
    SB_LUT4 add_5275_6_lut (.I0(GND_net), .I1(n10224[3]), .I2(n393_adj_4508), 
            .I3(n29276), .O(n10208[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5275_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_3_add_2_3 (.CI(n27976), .I0(setpoint[1]), .I1(motor_state[1]), 
            .CO(n27977));
    SB_CARRY add_5275_6 (.CI(n29276), .I0(n10224[3]), .I1(n393_adj_4508), 
            .CO(n29277));
    SB_LUT4 add_5275_5_lut (.I0(GND_net), .I1(n10224[2]), .I2(n320_adj_4507), 
            .I3(n29275), .O(n10208[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5275_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5275_5 (.CI(n29275), .I0(n10224[2]), .I1(n320_adj_4507), 
            .CO(n29276));
    SB_LUT4 add_5275_4_lut (.I0(GND_net), .I1(n10224[1]), .I2(n247_adj_4506), 
            .I3(n29274), .O(n10208[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5275_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_751_5 (.CI(n27900), .I0(\PID_CONTROLLER.integral [3]), 
            .I1(n3302[3]), .CO(n27901));
    SB_CARRY add_5275_4 (.CI(n29274), .I0(n10224[1]), .I1(n247_adj_4506), 
            .CO(n29275));
    SB_LUT4 add_5275_3_lut (.I0(GND_net), .I1(n10224[0]), .I2(n174_adj_4505), 
            .I3(n29273), .O(n10208[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5275_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5275_3 (.CI(n29273), .I0(n10224[0]), .I1(n174_adj_4505), 
            .CO(n29274));
    SB_LUT4 add_5275_2_lut (.I0(GND_net), .I1(n32_adj_4504), .I2(n101_adj_4502), 
            .I3(GND_net), .O(n10208[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5275_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5275_2 (.CI(GND_net), .I0(n32_adj_4504), .I1(n101_adj_4502), 
            .CO(n29273));
    SB_LUT4 i30121_4_lut (.I0(n24_adj_4676), .I1(n8_adj_4675), .I2(n45_adj_4653), 
            .I3(n36373), .O(n36876));   // verilog/motorControl.v(38[19:35])
    defparam i30121_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i30182_3_lut (.I0(n36973), .I1(n257[12]), .I2(n25_adj_4659), 
            .I3(GND_net), .O(n36937));   // verilog/motorControl.v(38[19:35])
    defparam i30182_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_15_i4_4_lut (.I0(duty_23__N_3646[0]), .I1(n257[1]), 
            .I2(duty_23__N_3646[1]), .I3(n257[0]), .O(n4_adj_4677));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i4_4_lut.LUT_INIT = 16'h4d0c;
    SB_LUT4 i30215_3_lut (.I0(n4_adj_4677), .I1(n257[13]), .I2(n27_adj_4665), 
            .I3(GND_net), .O(n36970));   // verilog/motorControl.v(38[19:35])
    defparam i30215_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i30216_3_lut (.I0(n36970), .I1(n257[14]), .I2(n29_adj_4656), 
            .I3(GND_net), .O(n36971));   // verilog/motorControl.v(38[19:35])
    defparam i30216_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i29632_4_lut (.I0(n33_adj_4661), .I1(n31_adj_4657), .I2(n29_adj_4656), 
            .I3(n36392), .O(n36387));
    defparam i29632_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i30320_4_lut (.I0(n30_adj_4672), .I1(n10_adj_4671), .I2(n35_adj_4660), 
            .I3(n36385), .O(n37075));   // verilog/motorControl.v(38[19:35])
    defparam i30320_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i30184_3_lut (.I0(n36971), .I1(n257[15]), .I2(n31_adj_4657), 
            .I3(GND_net), .O(n36939));   // verilog/motorControl.v(38[19:35])
    defparam i30184_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i30369_4_lut (.I0(n36939), .I1(n37075), .I2(n35_adj_4660), 
            .I3(n36387), .O(n37124));   // verilog/motorControl.v(38[19:35])
    defparam i30369_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i30370_3_lut (.I0(n37124), .I1(n257[18]), .I2(n37_adj_4655), 
            .I3(GND_net), .O(n37125));   // verilog/motorControl.v(38[19:35])
    defparam i30370_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i30347_3_lut (.I0(n37125), .I1(n257[19]), .I2(n39_adj_4652), 
            .I3(GND_net), .O(n37102));   // verilog/motorControl.v(38[19:35])
    defparam i30347_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i29622_4_lut (.I0(n43_adj_4654), .I1(n41_adj_4651), .I2(n39_adj_4652), 
            .I3(n37061), .O(n36377));
    defparam i29622_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i30279_4_lut (.I0(n36937), .I1(n36876), .I2(n45_adj_4653), 
            .I3(n36375), .O(n37034));   // verilog/motorControl.v(38[19:35])
    defparam i30279_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i30339_3_lut (.I0(n37102), .I1(n257[20]), .I2(n41_adj_4651), 
            .I3(GND_net), .O(n40_adj_4678));   // verilog/motorControl.v(38[19:35])
    defparam i30339_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i30281_4_lut (.I0(n40_adj_4678), .I1(n37034), .I2(n45_adj_4653), 
            .I3(n36377), .O(n37036));   // verilog/motorControl.v(38[19:35])
    defparam i30281_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i30282_3_lut (.I0(n37036), .I1(duty_23__N_3646[23]), .I2(n257[23]), 
            .I3(GND_net), .O(n256));   // verilog/motorControl.v(38[19:35])
    defparam i30282_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 mux_17_i1_3_lut (.I0(duty_23__N_3646[0]), .I1(n257[0]), .I2(n256), 
            .I3(GND_net), .O(duty_23__N_3621[0]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_17_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_i1_3_lut (.I0(duty_23__N_3621[0]), .I1(PWMLimit[0]), 
            .I2(duty_23__N_3645), .I3(GND_net), .O(duty_23__N_3522[0]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_5274_16_lut (.I0(GND_net), .I1(n10208[13]), .I2(n1120_adj_4501), 
            .I3(n29272), .O(n10191[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5274_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5274_15_lut (.I0(GND_net), .I1(n10208[12]), .I2(n1047_adj_4498), 
            .I3(n29271), .O(n10191[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5274_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5274_15 (.CI(n29271), .I0(n10208[12]), .I1(n1047_adj_4498), 
            .CO(n29272));
    SB_LUT4 add_5274_14_lut (.I0(GND_net), .I1(n10208[11]), .I2(n974_adj_4497), 
            .I3(n29270), .O(n10191[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5274_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5274_14 (.CI(n29270), .I0(n10208[11]), .I1(n974_adj_4497), 
            .CO(n29271));
    SB_LUT4 add_5274_13_lut (.I0(GND_net), .I1(n10208[10]), .I2(n901_adj_4496), 
            .I3(n29269), .O(n10191[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5274_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5274_13 (.CI(n29269), .I0(n10208[10]), .I1(n901_adj_4496), 
            .CO(n29270));
    SB_LUT4 add_5274_12_lut (.I0(GND_net), .I1(n10208[9]), .I2(n828_adj_4495), 
            .I3(n29268), .O(n10191[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5274_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5274_12 (.CI(n29268), .I0(n10208[9]), .I1(n828_adj_4495), 
            .CO(n29269));
    SB_LUT4 add_5274_11_lut (.I0(GND_net), .I1(n10208[8]), .I2(n755_adj_4494), 
            .I3(n29267), .O(n10191[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5274_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5274_11 (.CI(n29267), .I0(n10208[8]), .I1(n755_adj_4494), 
            .CO(n29268));
    SB_LUT4 add_5274_10_lut (.I0(GND_net), .I1(n10208[7]), .I2(n682_adj_4492), 
            .I3(n29266), .O(n10191[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5274_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5274_10 (.CI(n29266), .I0(n10208[7]), .I1(n682_adj_4492), 
            .CO(n29267));
    SB_DFF result_i1 (.Q(duty[1]), .C(clk32MHz), .D(duty_23__N_3522[1]));   // verilog/motorControl.v(29[14] 48[8])
    SB_LUT4 add_5274_9_lut (.I0(GND_net), .I1(n10208[6]), .I2(n609_adj_4488), 
            .I3(n29265), .O(n10191[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5274_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5274_9 (.CI(n29265), .I0(n10208[6]), .I1(n609_adj_4488), 
            .CO(n29266));
    SB_LUT4 add_5274_8_lut (.I0(GND_net), .I1(n10208[5]), .I2(n536_adj_4487), 
            .I3(n29264), .O(n10191[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5274_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5274_8 (.CI(n29264), .I0(n10208[5]), .I1(n536_adj_4487), 
            .CO(n29265));
    SB_LUT4 add_5274_7_lut (.I0(GND_net), .I1(n10208[4]), .I2(n463_adj_4486), 
            .I3(n29263), .O(n10191[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5274_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5274_7 (.CI(n29263), .I0(n10208[4]), .I1(n463_adj_4486), 
            .CO(n29264));
    SB_LUT4 add_5274_6_lut (.I0(GND_net), .I1(n10208[3]), .I2(n390_adj_4485), 
            .I3(n29262), .O(n10191[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5274_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5274_6 (.CI(n29262), .I0(n10208[3]), .I1(n390_adj_4485), 
            .CO(n29263));
    SB_LUT4 add_5274_5_lut (.I0(GND_net), .I1(n10208[2]), .I2(n317_adj_4484), 
            .I3(n29261), .O(n10191[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5274_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_751_4_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [2]), 
            .I2(n3302[2]), .I3(n27899), .O(\PID_CONTROLLER.integral_23__N_3546 [2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_751_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5274_5 (.CI(n29261), .I0(n10208[2]), .I1(n317_adj_4484), 
            .CO(n29262));
    SB_LUT4 add_5274_4_lut (.I0(GND_net), .I1(n10208[1]), .I2(n244_adj_4482), 
            .I3(n29260), .O(n10191[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5274_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5274_4 (.CI(n29260), .I0(n10208[1]), .I1(n244_adj_4482), 
            .CO(n29261));
    SB_LUT4 unary_minus_5_inv_0_i21_1_lut (.I0(IntegralLimit[20]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[20]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i21_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_3_add_2_2_lut (.I0(GND_net), .I1(setpoint[0]), .I2(motor_state[0]), 
            .I3(VCC_net), .O(n28[0])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_3_add_2_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_3_add_2_2 (.CI(VCC_net), .I0(setpoint[0]), .I1(motor_state[0]), 
            .CO(n27976));
    SB_CARRY add_751_4 (.CI(n27899), .I0(\PID_CONTROLLER.integral [2]), 
            .I1(n3302[2]), .CO(n27900));
    SB_LUT4 add_751_3_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [1]), 
            .I2(n3302[1]), .I3(n27898), .O(\PID_CONTROLLER.integral_23__N_3546 [1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_751_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5274_3_lut (.I0(GND_net), .I1(n10208[0]), .I2(n171_adj_4481), 
            .I3(n29259), .O(n10191[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5274_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5274_3 (.CI(n29259), .I0(n10208[0]), .I1(n171_adj_4481), 
            .CO(n29260));
    SB_LUT4 add_5274_2_lut (.I0(GND_net), .I1(n29_adj_4480), .I2(n98_adj_4479), 
            .I3(GND_net), .O(n10191[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5274_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5274_2 (.CI(GND_net), .I0(n29_adj_4480), .I1(n98_adj_4479), 
            .CO(n29259));
    SB_LUT4 add_5273_17_lut (.I0(GND_net), .I1(n10191[14]), .I2(GND_net), 
            .I3(n29258), .O(n10173[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5273_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5273_16_lut (.I0(GND_net), .I1(n10191[13]), .I2(n1117_adj_4477), 
            .I3(n29257), .O(n10173[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5273_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5273_16 (.CI(n29257), .I0(n10191[13]), .I1(n1117_adj_4477), 
            .CO(n29258));
    SB_LUT4 add_5273_15_lut (.I0(GND_net), .I1(n10191[12]), .I2(n1044_adj_4476), 
            .I3(n29256), .O(n10173[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5273_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5273_15 (.CI(n29256), .I0(n10191[12]), .I1(n1044_adj_4476), 
            .CO(n29257));
    SB_LUT4 add_5273_14_lut (.I0(GND_net), .I1(n10191[11]), .I2(n971_adj_4474), 
            .I3(n29255), .O(n10173[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5273_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5273_14 (.CI(n29255), .I0(n10191[11]), .I1(n971_adj_4474), 
            .CO(n29256));
    SB_LUT4 add_5273_13_lut (.I0(GND_net), .I1(n10191[10]), .I2(n898_adj_4473), 
            .I3(n29254), .O(n10173[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5273_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5273_13 (.CI(n29254), .I0(n10191[10]), .I1(n898_adj_4473), 
            .CO(n29255));
    SB_LUT4 add_5273_12_lut (.I0(GND_net), .I1(n10191[9]), .I2(n825_adj_4471), 
            .I3(n29253), .O(n10173[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5273_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5273_12 (.CI(n29253), .I0(n10191[9]), .I1(n825_adj_4471), 
            .CO(n29254));
    SB_LUT4 add_5273_11_lut (.I0(GND_net), .I1(n10191[8]), .I2(n752_adj_4470), 
            .I3(n29252), .O(n10173[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5273_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_751_3 (.CI(n27898), .I0(\PID_CONTROLLER.integral [1]), 
            .I1(n3302[1]), .CO(n27899));
    SB_CARRY add_5273_11 (.CI(n29252), .I0(n10191[8]), .I1(n752_adj_4470), 
            .CO(n29253));
    SB_LUT4 add_5273_10_lut (.I0(GND_net), .I1(n10191[7]), .I2(n679_adj_4468), 
            .I3(n29251), .O(n10173[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5273_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5273_10 (.CI(n29251), .I0(n10191[7]), .I1(n679_adj_4468), 
            .CO(n29252));
    SB_LUT4 add_751_2_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [0]), 
            .I2(n3302[0]), .I3(GND_net), .O(\PID_CONTROLLER.integral_23__N_3546 [0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_751_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5273_9_lut (.I0(GND_net), .I1(n10191[6]), .I2(n606_adj_4466), 
            .I3(n29250), .O(n10173[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5273_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5273_9 (.CI(n29250), .I0(n10191[6]), .I1(n606_adj_4466), 
            .CO(n29251));
    SB_LUT4 add_5273_8_lut (.I0(GND_net), .I1(n10191[5]), .I2(n533_adj_4465), 
            .I3(n29249), .O(n10173[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5273_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5273_8 (.CI(n29249), .I0(n10191[5]), .I1(n533_adj_4465), 
            .CO(n29250));
    SB_LUT4 add_5273_7_lut (.I0(GND_net), .I1(n10191[4]), .I2(n460_adj_4464), 
            .I3(n29248), .O(n10173[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5273_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5273_7 (.CI(n29248), .I0(n10191[4]), .I1(n460_adj_4464), 
            .CO(n29249));
    SB_LUT4 add_5273_6_lut (.I0(GND_net), .I1(n10191[3]), .I2(n387_adj_4463), 
            .I3(n29247), .O(n10173[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5273_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5273_6 (.CI(n29247), .I0(n10191[3]), .I1(n387_adj_4463), 
            .CO(n29248));
    SB_LUT4 add_5273_5_lut (.I0(GND_net), .I1(n10191[2]), .I2(n314_adj_4462), 
            .I3(n29246), .O(n10173[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5273_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5273_5 (.CI(n29246), .I0(n10191[2]), .I1(n314_adj_4462), 
            .CO(n29247));
    SB_LUT4 add_5273_4_lut (.I0(GND_net), .I1(n10191[1]), .I2(n241_adj_4461), 
            .I3(n29245), .O(n10173[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5273_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5273_4 (.CI(n29245), .I0(n10191[1]), .I1(n241_adj_4461), 
            .CO(n29246));
    SB_LUT4 add_5273_3_lut (.I0(GND_net), .I1(n10191[0]), .I2(n168_adj_4459), 
            .I3(n29244), .O(n10173[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5273_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5273_3 (.CI(n29244), .I0(n10191[0]), .I1(n168_adj_4459), 
            .CO(n29245));
    SB_LUT4 add_5273_2_lut (.I0(GND_net), .I1(n26_adj_4457), .I2(n95_adj_4456), 
            .I3(GND_net), .O(n10173[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5273_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5273_2 (.CI(GND_net), .I0(n26_adj_4457), .I1(n95_adj_4456), 
            .CO(n29244));
    SB_LUT4 add_5272_18_lut (.I0(GND_net), .I1(n10173[15]), .I2(GND_net), 
            .I3(n29243), .O(n10154[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5272_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5272_17_lut (.I0(GND_net), .I1(n10173[14]), .I2(GND_net), 
            .I3(n29242), .O(n10154[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5272_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5272_17 (.CI(n29242), .I0(n10173[14]), .I1(GND_net), 
            .CO(n29243));
    SB_LUT4 add_5272_16_lut (.I0(GND_net), .I1(n10173[13]), .I2(n1114_adj_4455), 
            .I3(n29241), .O(n10154[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5272_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5272_16 (.CI(n29241), .I0(n10173[13]), .I1(n1114_adj_4455), 
            .CO(n29242));
    SB_LUT4 add_5272_15_lut (.I0(GND_net), .I1(n10173[12]), .I2(n1041_adj_4454), 
            .I3(n29240), .O(n10154[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5272_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5272_15 (.CI(n29240), .I0(n10173[12]), .I1(n1041_adj_4454), 
            .CO(n29241));
    SB_LUT4 add_5272_14_lut (.I0(GND_net), .I1(n10173[11]), .I2(n968_adj_4453), 
            .I3(n29239), .O(n10154[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5272_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5272_14 (.CI(n29239), .I0(n10173[11]), .I1(n968_adj_4453), 
            .CO(n29240));
    SB_LUT4 add_5272_13_lut (.I0(GND_net), .I1(n10173[10]), .I2(n895_adj_4452), 
            .I3(n29238), .O(n10154[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5272_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5272_13 (.CI(n29238), .I0(n10173[10]), .I1(n895_adj_4452), 
            .CO(n29239));
    SB_LUT4 add_5272_12_lut (.I0(GND_net), .I1(n10173[9]), .I2(n822_adj_4451), 
            .I3(n29237), .O(n10154[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5272_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5272_12 (.CI(n29237), .I0(n10173[9]), .I1(n822_adj_4451), 
            .CO(n29238));
    SB_LUT4 add_5272_11_lut (.I0(GND_net), .I1(n10173[8]), .I2(n749_adj_4450), 
            .I3(n29236), .O(n10154[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5272_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5272_11 (.CI(n29236), .I0(n10173[8]), .I1(n749_adj_4450), 
            .CO(n29237));
    SB_LUT4 add_5272_10_lut (.I0(GND_net), .I1(n10173[7]), .I2(n676_adj_4449), 
            .I3(n29235), .O(n10154[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5272_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5272_10 (.CI(n29235), .I0(n10173[7]), .I1(n676_adj_4449), 
            .CO(n29236));
    SB_LUT4 add_5272_9_lut (.I0(GND_net), .I1(n10173[6]), .I2(n603_adj_4448), 
            .I3(n29234), .O(n10154[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5272_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5272_9 (.CI(n29234), .I0(n10173[6]), .I1(n603_adj_4448), 
            .CO(n29235));
    SB_LUT4 add_5272_8_lut (.I0(GND_net), .I1(n10173[5]), .I2(n530_adj_4447), 
            .I3(n29233), .O(n10154[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5272_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5272_8 (.CI(n29233), .I0(n10173[5]), .I1(n530_adj_4447), 
            .CO(n29234));
    SB_CARRY add_751_2 (.CI(GND_net), .I0(\PID_CONTROLLER.integral [0]), 
            .I1(n3302[0]), .CO(n27898));
    SB_LUT4 add_5272_7_lut (.I0(GND_net), .I1(n10173[4]), .I2(n457_adj_4443), 
            .I3(n29232), .O(n10154[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5272_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5272_7 (.CI(n29232), .I0(n10173[4]), .I1(n457_adj_4443), 
            .CO(n29233));
    SB_LUT4 add_5272_6_lut (.I0(GND_net), .I1(n10173[3]), .I2(n384_adj_4442), 
            .I3(n29231), .O(n10154[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5272_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5272_6 (.CI(n29231), .I0(n10173[3]), .I1(n384_adj_4442), 
            .CO(n29232));
    SB_LUT4 add_5272_5_lut (.I0(GND_net), .I1(n10173[2]), .I2(n311_adj_4439), 
            .I3(n29230), .O(n10154[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5272_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5272_5 (.CI(n29230), .I0(n10173[2]), .I1(n311_adj_4439), 
            .CO(n29231));
    SB_LUT4 add_5272_4_lut (.I0(GND_net), .I1(n10173[1]), .I2(n238_adj_4437), 
            .I3(n29229), .O(n10154[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5272_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5272_4 (.CI(n29229), .I0(n10173[1]), .I1(n238_adj_4437), 
            .CO(n29230));
    SB_LUT4 add_5272_3_lut (.I0(GND_net), .I1(n10173[0]), .I2(n165_adj_4436), 
            .I3(n29228), .O(n10154[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5272_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5272_3 (.CI(n29228), .I0(n10173[0]), .I1(n165_adj_4436), 
            .CO(n29229));
    SB_LUT4 add_5272_2_lut (.I0(GND_net), .I1(n23_adj_4435), .I2(n92_adj_4434), 
            .I3(GND_net), .O(n10154[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5272_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5272_2 (.CI(GND_net), .I0(n23_adj_4435), .I1(n92_adj_4434), 
            .CO(n29228));
    SB_LUT4 add_5271_19_lut (.I0(GND_net), .I1(n10154[16]), .I2(GND_net), 
            .I3(n29227), .O(n10134[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5271_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5271_18_lut (.I0(GND_net), .I1(n10154[15]), .I2(GND_net), 
            .I3(n29226), .O(n10134[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5271_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5271_18 (.CI(n29226), .I0(n10154[15]), .I1(GND_net), 
            .CO(n29227));
    SB_LUT4 add_5271_17_lut (.I0(GND_net), .I1(n10154[14]), .I2(GND_net), 
            .I3(n29225), .O(n10134[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5271_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5271_17 (.CI(n29225), .I0(n10154[14]), .I1(GND_net), 
            .CO(n29226));
    SB_LUT4 add_5271_16_lut (.I0(GND_net), .I1(n10154[13]), .I2(n1111_adj_4432), 
            .I3(n29224), .O(n10134[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5271_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5271_16 (.CI(n29224), .I0(n10154[13]), .I1(n1111_adj_4432), 
            .CO(n29225));
    SB_LUT4 add_5271_15_lut (.I0(GND_net), .I1(n10154[12]), .I2(n1038_adj_4431), 
            .I3(n29223), .O(n10134[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5271_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5271_15 (.CI(n29223), .I0(n10154[12]), .I1(n1038_adj_4431), 
            .CO(n29224));
    SB_LUT4 add_5271_14_lut (.I0(GND_net), .I1(n10154[11]), .I2(n965_adj_4430), 
            .I3(n29222), .O(n10134[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5271_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5271_14 (.CI(n29222), .I0(n10154[11]), .I1(n965_adj_4430), 
            .CO(n29223));
    SB_LUT4 add_5271_13_lut (.I0(GND_net), .I1(n10154[10]), .I2(n892_adj_4429), 
            .I3(n29221), .O(n10134[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5271_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5271_13 (.CI(n29221), .I0(n10154[10]), .I1(n892_adj_4429), 
            .CO(n29222));
    SB_LUT4 add_5271_12_lut (.I0(GND_net), .I1(n10154[9]), .I2(n819_adj_4428), 
            .I3(n29220), .O(n10134[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5271_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5271_12 (.CI(n29220), .I0(n10154[9]), .I1(n819_adj_4428), 
            .CO(n29221));
    SB_LUT4 add_5271_11_lut (.I0(GND_net), .I1(n10154[8]), .I2(n746_adj_4427), 
            .I3(n29219), .O(n10134[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5271_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5271_11 (.CI(n29219), .I0(n10154[8]), .I1(n746_adj_4427), 
            .CO(n29220));
    SB_LUT4 add_5271_10_lut (.I0(GND_net), .I1(n10154[7]), .I2(n673_adj_4425), 
            .I3(n29218), .O(n10134[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5271_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5271_10 (.CI(n29218), .I0(n10154[7]), .I1(n673_adj_4425), 
            .CO(n29219));
    SB_LUT4 add_5271_9_lut (.I0(GND_net), .I1(n10154[6]), .I2(n600_adj_4424), 
            .I3(n29217), .O(n10134[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5271_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5271_9 (.CI(n29217), .I0(n10154[6]), .I1(n600_adj_4424), 
            .CO(n29218));
    SB_LUT4 add_5271_8_lut (.I0(GND_net), .I1(n10154[5]), .I2(n527_adj_4422), 
            .I3(n29216), .O(n10134[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5271_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5271_8 (.CI(n29216), .I0(n10154[5]), .I1(n527_adj_4422), 
            .CO(n29217));
    SB_LUT4 add_5271_7_lut (.I0(GND_net), .I1(n10154[4]), .I2(n454_adj_4421), 
            .I3(n29215), .O(n10134[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5271_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5271_7 (.CI(n29215), .I0(n10154[4]), .I1(n454_adj_4421), 
            .CO(n29216));
    SB_LUT4 add_5271_6_lut (.I0(GND_net), .I1(n10154[3]), .I2(n381_adj_4420), 
            .I3(n29214), .O(n10134[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5271_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5271_6 (.CI(n29214), .I0(n10154[3]), .I1(n381_adj_4420), 
            .CO(n29215));
    SB_LUT4 add_5271_5_lut (.I0(GND_net), .I1(n10154[2]), .I2(n308_adj_4419), 
            .I3(n29213), .O(n10134[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5271_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5271_5 (.CI(n29213), .I0(n10154[2]), .I1(n308_adj_4419), 
            .CO(n29214));
    SB_LUT4 add_5271_4_lut (.I0(GND_net), .I1(n10154[1]), .I2(n235_adj_4418), 
            .I3(n29212), .O(n10134[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5271_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5271_4 (.CI(n29212), .I0(n10154[1]), .I1(n235_adj_4418), 
            .CO(n29213));
    SB_LUT4 add_5271_3_lut (.I0(GND_net), .I1(n10154[0]), .I2(n162_adj_4416), 
            .I3(n29211), .O(n10134[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5271_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5271_3 (.CI(n29211), .I0(n10154[0]), .I1(n162_adj_4416), 
            .CO(n29212));
    SB_LUT4 add_5271_2_lut (.I0(GND_net), .I1(n20_adj_4415), .I2(n89), 
            .I3(GND_net), .O(n10134[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5271_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5271_2 (.CI(GND_net), .I0(n20_adj_4415), .I1(n89), .CO(n29211));
    SB_LUT4 add_5270_20_lut (.I0(GND_net), .I1(n10134[17]), .I2(GND_net), 
            .I3(n29210), .O(n10113[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5270_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5270_19_lut (.I0(GND_net), .I1(n10134[16]), .I2(GND_net), 
            .I3(n29209), .O(n10113[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5270_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5270_19 (.CI(n29209), .I0(n10134[16]), .I1(GND_net), 
            .CO(n29210));
    SB_LUT4 add_5270_18_lut (.I0(GND_net), .I1(n10134[15]), .I2(GND_net), 
            .I3(n29208), .O(n10113[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5270_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5270_18 (.CI(n29208), .I0(n10134[15]), .I1(GND_net), 
            .CO(n29209));
    SB_LUT4 add_5270_17_lut (.I0(GND_net), .I1(n10134[14]), .I2(GND_net), 
            .I3(n29207), .O(n10113[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5270_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5270_17 (.CI(n29207), .I0(n10134[14]), .I1(GND_net), 
            .CO(n29208));
    SB_LUT4 mult_10_i57_2_lut (.I0(\Kp[1] ), .I1(n28[3]), .I2(GND_net), 
            .I3(GND_net), .O(n83_adj_4679));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i57_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5270_16_lut (.I0(GND_net), .I1(n10134[13]), .I2(n1108), 
            .I3(n29206), .O(n10113[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5270_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5270_16 (.CI(n29206), .I0(n10134[13]), .I1(n1108), .CO(n29207));
    SB_LUT4 add_5270_15_lut (.I0(GND_net), .I1(n10134[12]), .I2(n1035), 
            .I3(n29205), .O(n10113[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5270_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i10_2_lut (.I0(\Kp[0] ), .I1(n28[4]), .I2(GND_net), 
            .I3(GND_net), .O(n14_adj_4680));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i10_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5270_15 (.CI(n29205), .I0(n10134[12]), .I1(n1035), .CO(n29206));
    SB_LUT4 add_5270_14_lut (.I0(GND_net), .I1(n10134[11]), .I2(n962), 
            .I3(n29204), .O(n10113[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5270_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5270_14 (.CI(n29204), .I0(n10134[11]), .I1(n962), .CO(n29205));
    SB_LUT4 add_5270_13_lut (.I0(GND_net), .I1(n10134[10]), .I2(n889), 
            .I3(n29203), .O(n10113[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5270_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5270_13 (.CI(n29203), .I0(n10134[10]), .I1(n889), .CO(n29204));
    SB_LUT4 add_5270_12_lut (.I0(GND_net), .I1(n10134[9]), .I2(n816), 
            .I3(n29202), .O(n10113[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5270_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5270_12 (.CI(n29202), .I0(n10134[9]), .I1(n816), .CO(n29203));
    SB_LUT4 mult_10_i106_2_lut (.I0(\Kp[2] ), .I1(n28[3]), .I2(GND_net), 
            .I3(GND_net), .O(n156_adj_4681));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i106_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5270_11_lut (.I0(GND_net), .I1(n10134[8]), .I2(n743), 
            .I3(n29201), .O(n10113[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5270_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5270_11 (.CI(n29201), .I0(n10134[8]), .I1(n743), .CO(n29202));
    SB_LUT4 add_5270_10_lut (.I0(GND_net), .I1(n10134[7]), .I2(n670), 
            .I3(n29200), .O(n10113[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5270_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5270_10 (.CI(n29200), .I0(n10134[7]), .I1(n670), .CO(n29201));
    SB_LUT4 add_5270_9_lut (.I0(GND_net), .I1(n10134[6]), .I2(n597), .I3(n29199), 
            .O(n10113[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5270_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5270_9 (.CI(n29199), .I0(n10134[6]), .I1(n597), .CO(n29200));
    SB_LUT4 add_5270_8_lut (.I0(GND_net), .I1(n10134[5]), .I2(n524), .I3(n29198), 
            .O(n10113[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5270_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5270_8 (.CI(n29198), .I0(n10134[5]), .I1(n524), .CO(n29199));
    SB_LUT4 add_5270_7_lut (.I0(GND_net), .I1(n10134[4]), .I2(n451), .I3(n29197), 
            .O(n10113[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5270_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i155_2_lut (.I0(\Kp[3] ), .I1(n28[3]), .I2(GND_net), 
            .I3(GND_net), .O(n229_adj_4682));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i155_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5270_7 (.CI(n29197), .I0(n10134[4]), .I1(n451), .CO(n29198));
    SB_LUT4 add_5270_6_lut (.I0(GND_net), .I1(n10134[3]), .I2(n378), .I3(n29196), 
            .O(n10113[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5270_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5270_6 (.CI(n29196), .I0(n10134[3]), .I1(n378), .CO(n29197));
    SB_LUT4 add_5270_5_lut (.I0(GND_net), .I1(n10134[2]), .I2(n305), .I3(n29195), 
            .O(n10113[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5270_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5270_5 (.CI(n29195), .I0(n10134[2]), .I1(n305), .CO(n29196));
    SB_LUT4 add_5270_4_lut (.I0(GND_net), .I1(n10134[1]), .I2(n232), .I3(n29194), 
            .O(n10113[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5270_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_16_inv_0_i15_1_lut (.I0(PWMLimit[14]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4735[14]));   // verilog/motorControl.v(39[18:27])
    defparam unary_minus_16_inv_0_i15_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_5270_4 (.CI(n29194), .I0(n10134[1]), .I1(n232), .CO(n29195));
    SB_LUT4 add_5270_3_lut (.I0(GND_net), .I1(n10134[0]), .I2(n159), .I3(n29193), 
            .O(n10113[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5270_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i204_2_lut (.I0(\Kp[4] ), .I1(n28[3]), .I2(GND_net), 
            .I3(GND_net), .O(n302_adj_4684));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i204_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5270_3 (.CI(n29193), .I0(n10134[0]), .I1(n159), .CO(n29194));
    SB_LUT4 add_5270_2_lut (.I0(GND_net), .I1(n17_adj_4400), .I2(n86), 
            .I3(GND_net), .O(n10113[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5270_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5270_2 (.CI(GND_net), .I0(n17_adj_4400), .I1(n86), .CO(n29193));
    SB_LUT4 add_5269_21_lut (.I0(GND_net), .I1(n10113[18]), .I2(GND_net), 
            .I3(n29192), .O(n10091[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5269_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5269_20_lut (.I0(GND_net), .I1(n10113[17]), .I2(GND_net), 
            .I3(n29191), .O(n10091[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5269_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5269_20 (.CI(n29191), .I0(n10113[17]), .I1(GND_net), 
            .CO(n29192));
    SB_LUT4 add_5269_19_lut (.I0(GND_net), .I1(n10113[16]), .I2(GND_net), 
            .I3(n29190), .O(n10091[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5269_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5269_19 (.CI(n29190), .I0(n10113[16]), .I1(GND_net), 
            .CO(n29191));
    SB_LUT4 add_5269_18_lut (.I0(GND_net), .I1(n10113[15]), .I2(GND_net), 
            .I3(n29189), .O(n10091[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5269_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5269_18 (.CI(n29189), .I0(n10113[15]), .I1(GND_net), 
            .CO(n29190));
    SB_LUT4 mult_10_i253_2_lut (.I0(\Kp[5] ), .I1(n28[3]), .I2(GND_net), 
            .I3(GND_net), .O(n375_adj_4685));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i253_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5269_17_lut (.I0(GND_net), .I1(n10113[14]), .I2(GND_net), 
            .I3(n29188), .O(n10091[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5269_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5269_17 (.CI(n29188), .I0(n10113[14]), .I1(GND_net), 
            .CO(n29189));
    SB_LUT4 add_5269_16_lut (.I0(GND_net), .I1(n10113[13]), .I2(n1105), 
            .I3(n29187), .O(n10091[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5269_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5269_16 (.CI(n29187), .I0(n10113[13]), .I1(n1105), .CO(n29188));
    SB_LUT4 add_5269_15_lut (.I0(GND_net), .I1(n10113[12]), .I2(n1032), 
            .I3(n29186), .O(n10091[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5269_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5269_15 (.CI(n29186), .I0(n10113[12]), .I1(n1032), .CO(n29187));
    SB_LUT4 add_5269_14_lut (.I0(GND_net), .I1(n10113[11]), .I2(n959), 
            .I3(n29185), .O(n10091[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5269_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5269_14 (.CI(n29185), .I0(n10113[11]), .I1(n959), .CO(n29186));
    SB_LUT4 add_5269_13_lut (.I0(GND_net), .I1(n10113[10]), .I2(n886), 
            .I3(n29184), .O(n10091[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5269_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5269_13 (.CI(n29184), .I0(n10113[10]), .I1(n886), .CO(n29185));
    SB_LUT4 add_5269_12_lut (.I0(GND_net), .I1(n10113[9]), .I2(n813), 
            .I3(n29183), .O(n10091[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5269_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5269_12 (.CI(n29183), .I0(n10113[9]), .I1(n813), .CO(n29184));
    SB_LUT4 add_5269_11_lut (.I0(GND_net), .I1(n10113[8]), .I2(n740), 
            .I3(n29182), .O(n10091[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5269_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5269_11 (.CI(n29182), .I0(n10113[8]), .I1(n740), .CO(n29183));
    SB_LUT4 add_5269_10_lut (.I0(GND_net), .I1(n10113[7]), .I2(n667), 
            .I3(n29181), .O(n10091[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5269_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5269_10 (.CI(n29181), .I0(n10113[7]), .I1(n667), .CO(n29182));
    SB_LUT4 add_5269_9_lut (.I0(GND_net), .I1(n10113[6]), .I2(n594), .I3(n29180), 
            .O(n10091[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5269_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5269_9 (.CI(n29180), .I0(n10113[6]), .I1(n594), .CO(n29181));
    SB_LUT4 add_5269_8_lut (.I0(GND_net), .I1(n10113[5]), .I2(n521), .I3(n29179), 
            .O(n10091[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5269_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5269_8 (.CI(n29179), .I0(n10113[5]), .I1(n521), .CO(n29180));
    SB_LUT4 add_5269_7_lut (.I0(GND_net), .I1(n10113[4]), .I2(n448), .I3(n29178), 
            .O(n10091[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5269_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5269_7 (.CI(n29178), .I0(n10113[4]), .I1(n448), .CO(n29179));
    SB_LUT4 add_5269_6_lut (.I0(GND_net), .I1(n10113[3]), .I2(n375), .I3(n29177), 
            .O(n10091[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5269_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5269_6 (.CI(n29177), .I0(n10113[3]), .I1(n375), .CO(n29178));
    SB_LUT4 add_5269_5_lut (.I0(GND_net), .I1(n10113[2]), .I2(n302), .I3(n29176), 
            .O(n10091[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5269_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5269_5 (.CI(n29176), .I0(n10113[2]), .I1(n302), .CO(n29177));
    SB_LUT4 add_5269_4_lut (.I0(GND_net), .I1(n10113[1]), .I2(n229), .I3(n29175), 
            .O(n10091[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5269_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5269_4 (.CI(n29175), .I0(n10113[1]), .I1(n229), .CO(n29176));
    SB_LUT4 add_5269_3_lut (.I0(GND_net), .I1(n10113[0]), .I2(n156), .I3(n29174), 
            .O(n10091[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5269_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5269_3 (.CI(n29174), .I0(n10113[0]), .I1(n156), .CO(n29175));
    SB_LUT4 add_5269_2_lut (.I0(GND_net), .I1(n14_adj_4396), .I2(n83), 
            .I3(GND_net), .O(n10091[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5269_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5269_2 (.CI(GND_net), .I0(n14_adj_4396), .I1(n83), .CO(n29174));
    SB_LUT4 add_5268_22_lut (.I0(GND_net), .I1(n10091[19]), .I2(GND_net), 
            .I3(n29173), .O(n10068[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5268_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5268_21_lut (.I0(GND_net), .I1(n10091[18]), .I2(GND_net), 
            .I3(n29172), .O(n10068[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5268_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5268_21 (.CI(n29172), .I0(n10091[18]), .I1(GND_net), 
            .CO(n29173));
    SB_LUT4 add_5268_20_lut (.I0(GND_net), .I1(n10091[17]), .I2(GND_net), 
            .I3(n29171), .O(n10068[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5268_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5268_20 (.CI(n29171), .I0(n10091[17]), .I1(GND_net), 
            .CO(n29172));
    SB_LUT4 add_5268_19_lut (.I0(GND_net), .I1(n10091[16]), .I2(GND_net), 
            .I3(n29170), .O(n10068[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5268_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5268_19 (.CI(n29170), .I0(n10091[16]), .I1(GND_net), 
            .CO(n29171));
    SB_LUT4 add_5268_18_lut (.I0(GND_net), .I1(n10091[15]), .I2(GND_net), 
            .I3(n29169), .O(n10068[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5268_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5268_18 (.CI(n29169), .I0(n10091[15]), .I1(GND_net), 
            .CO(n29170));
    SB_LUT4 add_5268_17_lut (.I0(GND_net), .I1(n10091[14]), .I2(GND_net), 
            .I3(n29168), .O(n10068[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5268_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5268_17 (.CI(n29168), .I0(n10091[14]), .I1(GND_net), 
            .CO(n29169));
    SB_LUT4 add_5268_16_lut (.I0(GND_net), .I1(n10091[13]), .I2(n1102), 
            .I3(n29167), .O(n10068[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5268_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5268_16 (.CI(n29167), .I0(n10091[13]), .I1(n1102), .CO(n29168));
    SB_LUT4 add_5268_15_lut (.I0(GND_net), .I1(n10091[12]), .I2(n1029), 
            .I3(n29166), .O(n10068[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5268_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5268_15 (.CI(n29166), .I0(n10091[12]), .I1(n1029), .CO(n29167));
    SB_LUT4 add_5268_14_lut (.I0(GND_net), .I1(n10091[11]), .I2(n956), 
            .I3(n29165), .O(n10068[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5268_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5268_14 (.CI(n29165), .I0(n10091[11]), .I1(n956), .CO(n29166));
    SB_LUT4 add_5268_13_lut (.I0(GND_net), .I1(n10091[10]), .I2(n883), 
            .I3(n29164), .O(n10068[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5268_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5268_13 (.CI(n29164), .I0(n10091[10]), .I1(n883), .CO(n29165));
    SB_LUT4 add_5268_12_lut (.I0(GND_net), .I1(n10091[9]), .I2(n810), 
            .I3(n29163), .O(n10068[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5268_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5268_12 (.CI(n29163), .I0(n10091[9]), .I1(n810), .CO(n29164));
    SB_LUT4 add_5268_11_lut (.I0(GND_net), .I1(n10091[8]), .I2(n737), 
            .I3(n29162), .O(n10068[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5268_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5268_11 (.CI(n29162), .I0(n10091[8]), .I1(n737), .CO(n29163));
    SB_LUT4 add_5268_10_lut (.I0(GND_net), .I1(n10091[7]), .I2(n664), 
            .I3(n29161), .O(n10068[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5268_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5268_10 (.CI(n29161), .I0(n10091[7]), .I1(n664), .CO(n29162));
    SB_LUT4 add_5268_9_lut (.I0(GND_net), .I1(n10091[6]), .I2(n591), .I3(n29160), 
            .O(n10068[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5268_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5268_9 (.CI(n29160), .I0(n10091[6]), .I1(n591), .CO(n29161));
    SB_LUT4 add_5268_8_lut (.I0(GND_net), .I1(n10091[5]), .I2(n518), .I3(n29159), 
            .O(n10068[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5268_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5268_8 (.CI(n29159), .I0(n10091[5]), .I1(n518), .CO(n29160));
    SB_LUT4 add_5268_7_lut (.I0(GND_net), .I1(n10091[4]), .I2(n445), .I3(n29158), 
            .O(n10068[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5268_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5268_7 (.CI(n29158), .I0(n10091[4]), .I1(n445), .CO(n29159));
    SB_LUT4 add_5268_6_lut (.I0(GND_net), .I1(n10091[3]), .I2(n372), .I3(n29157), 
            .O(n10068[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5268_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5268_6 (.CI(n29157), .I0(n10091[3]), .I1(n372), .CO(n29158));
    SB_LUT4 add_5268_5_lut (.I0(GND_net), .I1(n10091[2]), .I2(n299), .I3(n29156), 
            .O(n10068[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5268_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5268_5 (.CI(n29156), .I0(n10091[2]), .I1(n299), .CO(n29157));
    SB_LUT4 add_5268_4_lut (.I0(GND_net), .I1(n10091[1]), .I2(n226), .I3(n29155), 
            .O(n10068[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5268_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5268_4 (.CI(n29155), .I0(n10091[1]), .I1(n226), .CO(n29156));
    SB_LUT4 add_5268_3_lut (.I0(GND_net), .I1(n10091[0]), .I2(n153), .I3(n29154), 
            .O(n10068[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5268_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5268_3 (.CI(n29154), .I0(n10091[0]), .I1(n153), .CO(n29155));
    SB_LUT4 add_5268_2_lut (.I0(GND_net), .I1(n11_adj_4390), .I2(n80), 
            .I3(GND_net), .O(n10068[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5268_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5268_2 (.CI(GND_net), .I0(n11_adj_4390), .I1(n80), .CO(n29154));
    SB_LUT4 mult_11_add_1225_24_lut (.I0(\PID_CONTROLLER.integral_23__N_3546 [23]), 
            .I1(n10044[21]), .I2(GND_net), .I3(n29153), .O(n8179[0])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_24_lut.LUT_INIT = 16'h6996;
    SB_LUT4 mult_11_add_1225_23_lut (.I0(GND_net), .I1(n10044[20]), .I2(GND_net), 
            .I3(n29152), .O(n155[22])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_23 (.CI(n29152), .I0(n10044[20]), .I1(GND_net), 
            .CO(n29153));
    SB_LUT4 mult_11_add_1225_22_lut (.I0(GND_net), .I1(n10044[19]), .I2(GND_net), 
            .I3(n29151), .O(n155[21])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_22 (.CI(n29151), .I0(n10044[19]), .I1(GND_net), 
            .CO(n29152));
    SB_LUT4 mult_11_add_1225_21_lut (.I0(GND_net), .I1(n10044[18]), .I2(GND_net), 
            .I3(n29150), .O(n155[20])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_21 (.CI(n29150), .I0(n10044[18]), .I1(GND_net), 
            .CO(n29151));
    SB_LUT4 mult_11_add_1225_20_lut (.I0(GND_net), .I1(n10044[17]), .I2(GND_net), 
            .I3(n29149), .O(n155[19])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_20 (.CI(n29149), .I0(n10044[17]), .I1(GND_net), 
            .CO(n29150));
    SB_LUT4 mult_11_add_1225_19_lut (.I0(GND_net), .I1(n10044[16]), .I2(GND_net), 
            .I3(n29148), .O(n155[18])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_19 (.CI(n29148), .I0(n10044[16]), .I1(GND_net), 
            .CO(n29149));
    SB_LUT4 mult_11_add_1225_18_lut (.I0(GND_net), .I1(n10044[15]), .I2(GND_net), 
            .I3(n29147), .O(n155[17])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_18 (.CI(n29147), .I0(n10044[15]), .I1(GND_net), 
            .CO(n29148));
    SB_LUT4 mult_11_add_1225_17_lut (.I0(GND_net), .I1(n10044[14]), .I2(GND_net), 
            .I3(n29146), .O(n155[16])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_17 (.CI(n29146), .I0(n10044[14]), .I1(GND_net), 
            .CO(n29147));
    SB_LUT4 mult_11_add_1225_16_lut (.I0(GND_net), .I1(n10044[13]), .I2(n1096), 
            .I3(n29145), .O(n155[15])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_16 (.CI(n29145), .I0(n10044[13]), .I1(n1096), 
            .CO(n29146));
    SB_LUT4 mult_11_add_1225_15_lut (.I0(GND_net), .I1(n10044[12]), .I2(n1023), 
            .I3(n29144), .O(n155[14])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_15 (.CI(n29144), .I0(n10044[12]), .I1(n1023), 
            .CO(n29145));
    SB_LUT4 mult_11_add_1225_14_lut (.I0(GND_net), .I1(n10044[11]), .I2(n950), 
            .I3(n29143), .O(n155[13])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_14 (.CI(n29143), .I0(n10044[11]), .I1(n950), 
            .CO(n29144));
    SB_LUT4 mult_11_add_1225_13_lut (.I0(GND_net), .I1(n10044[10]), .I2(n877), 
            .I3(n29142), .O(n155[12])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_13 (.CI(n29142), .I0(n10044[10]), .I1(n877), 
            .CO(n29143));
    SB_LUT4 mult_11_add_1225_12_lut (.I0(GND_net), .I1(n10044[9]), .I2(n804), 
            .I3(n29141), .O(n155[11])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_12 (.CI(n29141), .I0(n10044[9]), .I1(n804), 
            .CO(n29142));
    SB_LUT4 mult_11_add_1225_11_lut (.I0(GND_net), .I1(n10044[8]), .I2(n731), 
            .I3(n29140), .O(n155[10])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_11 (.CI(n29140), .I0(n10044[8]), .I1(n731), 
            .CO(n29141));
    SB_LUT4 mult_11_add_1225_10_lut (.I0(GND_net), .I1(n10044[7]), .I2(n658), 
            .I3(n29139), .O(n155[9])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_10 (.CI(n29139), .I0(n10044[7]), .I1(n658), 
            .CO(n29140));
    SB_LUT4 mult_11_add_1225_9_lut (.I0(GND_net), .I1(n10044[6]), .I2(n585), 
            .I3(n29138), .O(n155[8])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_9 (.CI(n29138), .I0(n10044[6]), .I1(n585), 
            .CO(n29139));
    SB_LUT4 mult_11_add_1225_8_lut (.I0(GND_net), .I1(n10044[5]), .I2(n512), 
            .I3(n29137), .O(n155[7])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_8 (.CI(n29137), .I0(n10044[5]), .I1(n512), 
            .CO(n29138));
    SB_LUT4 mult_11_add_1225_7_lut (.I0(GND_net), .I1(n10044[4]), .I2(n439), 
            .I3(n29136), .O(n155[6])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_7 (.CI(n29136), .I0(n10044[4]), .I1(n439), 
            .CO(n29137));
    SB_LUT4 mult_11_add_1225_6_lut (.I0(GND_net), .I1(n10044[3]), .I2(n366), 
            .I3(n29135), .O(n155[5])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_6 (.CI(n29135), .I0(n10044[3]), .I1(n366), 
            .CO(n29136));
    SB_LUT4 mult_11_add_1225_5_lut (.I0(GND_net), .I1(n10044[2]), .I2(n293), 
            .I3(n29134), .O(n155[4])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_5 (.CI(n29134), .I0(n10044[2]), .I1(n293), 
            .CO(n29135));
    SB_LUT4 mult_11_add_1225_4_lut (.I0(GND_net), .I1(n10044[1]), .I2(n220), 
            .I3(n29133), .O(n155[3])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_4 (.CI(n29133), .I0(n10044[1]), .I1(n220), 
            .CO(n29134));
    SB_LUT4 mult_11_add_1225_3_lut (.I0(GND_net), .I1(n10044[0]), .I2(n147), 
            .I3(n29132), .O(n155[2])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_3 (.CI(n29132), .I0(n10044[0]), .I1(n147), 
            .CO(n29133));
    SB_LUT4 mult_11_add_1225_2_lut (.I0(GND_net), .I1(n5_adj_4388), .I2(n74), 
            .I3(GND_net), .O(n155[1])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_2 (.CI(GND_net), .I0(n5_adj_4388), .I1(n74), 
            .CO(n29132));
    SB_LUT4 add_5267_23_lut (.I0(GND_net), .I1(n10068[20]), .I2(GND_net), 
            .I3(n29131), .O(n10044[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5267_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5267_22_lut (.I0(GND_net), .I1(n10068[19]), .I2(GND_net), 
            .I3(n29130), .O(n10044[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5267_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5267_22 (.CI(n29130), .I0(n10068[19]), .I1(GND_net), 
            .CO(n29131));
    SB_LUT4 add_5267_21_lut (.I0(GND_net), .I1(n10068[18]), .I2(GND_net), 
            .I3(n29129), .O(n10044[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5267_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5267_21 (.CI(n29129), .I0(n10068[18]), .I1(GND_net), 
            .CO(n29130));
    SB_LUT4 add_5267_20_lut (.I0(GND_net), .I1(n10068[17]), .I2(GND_net), 
            .I3(n29128), .O(n10044[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5267_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5267_20 (.CI(n29128), .I0(n10068[17]), .I1(GND_net), 
            .CO(n29129));
    SB_LUT4 add_5267_19_lut (.I0(GND_net), .I1(n10068[16]), .I2(GND_net), 
            .I3(n29127), .O(n10044[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5267_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5267_19 (.CI(n29127), .I0(n10068[16]), .I1(GND_net), 
            .CO(n29128));
    SB_LUT4 add_5267_18_lut (.I0(GND_net), .I1(n10068[15]), .I2(GND_net), 
            .I3(n29126), .O(n10044[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5267_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5267_18 (.CI(n29126), .I0(n10068[15]), .I1(GND_net), 
            .CO(n29127));
    SB_LUT4 add_5267_17_lut (.I0(GND_net), .I1(n10068[14]), .I2(GND_net), 
            .I3(n29125), .O(n10044[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5267_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5267_17 (.CI(n29125), .I0(n10068[14]), .I1(GND_net), 
            .CO(n29126));
    SB_LUT4 add_5267_16_lut (.I0(GND_net), .I1(n10068[13]), .I2(n1099), 
            .I3(n29124), .O(n10044[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5267_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5267_16 (.CI(n29124), .I0(n10068[13]), .I1(n1099), .CO(n29125));
    SB_LUT4 add_5267_15_lut (.I0(GND_net), .I1(n10068[12]), .I2(n1026), 
            .I3(n29123), .O(n10044[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5267_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5267_15 (.CI(n29123), .I0(n10068[12]), .I1(n1026), .CO(n29124));
    SB_LUT4 add_5267_14_lut (.I0(GND_net), .I1(n10068[11]), .I2(n953), 
            .I3(n29122), .O(n10044[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5267_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5267_14 (.CI(n29122), .I0(n10068[11]), .I1(n953), .CO(n29123));
    SB_LUT4 add_5267_13_lut (.I0(GND_net), .I1(n10068[10]), .I2(n880), 
            .I3(n29121), .O(n10044[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5267_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5267_13 (.CI(n29121), .I0(n10068[10]), .I1(n880), .CO(n29122));
    SB_LUT4 add_5267_12_lut (.I0(GND_net), .I1(n10068[9]), .I2(n807), 
            .I3(n29120), .O(n10044[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5267_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5267_12 (.CI(n29120), .I0(n10068[9]), .I1(n807), .CO(n29121));
    SB_LUT4 add_5267_11_lut (.I0(GND_net), .I1(n10068[8]), .I2(n734), 
            .I3(n29119), .O(n10044[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5267_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5267_11 (.CI(n29119), .I0(n10068[8]), .I1(n734), .CO(n29120));
    SB_LUT4 add_5267_10_lut (.I0(GND_net), .I1(n10068[7]), .I2(n661), 
            .I3(n29118), .O(n10044[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5267_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5267_10 (.CI(n29118), .I0(n10068[7]), .I1(n661), .CO(n29119));
    SB_LUT4 add_5267_9_lut (.I0(GND_net), .I1(n10068[6]), .I2(n588), .I3(n29117), 
            .O(n10044[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5267_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5267_9 (.CI(n29117), .I0(n10068[6]), .I1(n588), .CO(n29118));
    SB_LUT4 add_5267_8_lut (.I0(GND_net), .I1(n10068[5]), .I2(n515), .I3(n29116), 
            .O(n10044[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5267_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5267_8 (.CI(n29116), .I0(n10068[5]), .I1(n515), .CO(n29117));
    SB_LUT4 add_5267_7_lut (.I0(GND_net), .I1(n10068[4]), .I2(n442), .I3(n29115), 
            .O(n10044[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5267_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5267_7 (.CI(n29115), .I0(n10068[4]), .I1(n442), .CO(n29116));
    SB_LUT4 add_5267_6_lut (.I0(GND_net), .I1(n10068[3]), .I2(n369), .I3(n29114), 
            .O(n10044[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5267_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5267_6 (.CI(n29114), .I0(n10068[3]), .I1(n369), .CO(n29115));
    SB_LUT4 add_5267_5_lut (.I0(GND_net), .I1(n10068[2]), .I2(n296), .I3(n29113), 
            .O(n10044[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5267_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5267_5 (.CI(n29113), .I0(n10068[2]), .I1(n296), .CO(n29114));
    SB_LUT4 add_5267_4_lut (.I0(GND_net), .I1(n10068[1]), .I2(n223), .I3(n29112), 
            .O(n10044[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5267_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5267_4 (.CI(n29112), .I0(n10068[1]), .I1(n223), .CO(n29113));
    SB_LUT4 add_5267_3_lut (.I0(GND_net), .I1(n10068[0]), .I2(n150), .I3(n29111), 
            .O(n10044[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5267_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5267_3 (.CI(n29111), .I0(n10068[0]), .I1(n150), .CO(n29112));
    SB_LUT4 add_5267_2_lut (.I0(GND_net), .I1(n8_adj_4382), .I2(n77), 
            .I3(GND_net), .O(n10044[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5267_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5267_2 (.CI(GND_net), .I0(n8_adj_4382), .I1(n77), .CO(n29111));
    SB_LUT4 add_5261_7_lut (.I0(GND_net), .I1(n34086), .I2(n490), .I3(n29110), 
            .O(n10011[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5261_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5261_6_lut (.I0(GND_net), .I1(n10019[3]), .I2(n417), .I3(n29109), 
            .O(n10011[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5261_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5261_6 (.CI(n29109), .I0(n10019[3]), .I1(n417), .CO(n29110));
    SB_LUT4 add_5261_5_lut (.I0(GND_net), .I1(n10019[2]), .I2(n344), .I3(n29108), 
            .O(n10011[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5261_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5261_5 (.CI(n29108), .I0(n10019[2]), .I1(n344), .CO(n29109));
    SB_LUT4 add_5261_4_lut (.I0(GND_net), .I1(n10019[1]), .I2(n271_adj_4371), 
            .I3(n29107), .O(n10011[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5261_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5261_4 (.CI(n29107), .I0(n10019[1]), .I1(n271_adj_4371), 
            .CO(n29108));
    SB_LUT4 add_5261_3_lut (.I0(GND_net), .I1(n10019[0]), .I2(n198), .I3(n29106), 
            .O(n10011[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5261_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5261_3 (.CI(n29106), .I0(n10019[0]), .I1(n198), .CO(n29107));
    SB_LUT4 add_5261_2_lut (.I0(GND_net), .I1(n56), .I2(n125), .I3(GND_net), 
            .O(n10011[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5261_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5261_2 (.CI(GND_net), .I0(n56), .I1(n125), .CO(n29106));
    SB_LUT4 add_5260_8_lut (.I0(GND_net), .I1(n10011[5]), .I2(n560), .I3(n29105), 
            .O(n10002[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5260_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5260_7_lut (.I0(GND_net), .I1(n10011[4]), .I2(n487), .I3(n29104), 
            .O(n10002[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5260_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5260_7 (.CI(n29104), .I0(n10011[4]), .I1(n487), .CO(n29105));
    SB_LUT4 add_5260_6_lut (.I0(GND_net), .I1(n10011[3]), .I2(n414), .I3(n29103), 
            .O(n10002[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5260_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5260_6 (.CI(n29103), .I0(n10011[3]), .I1(n414), .CO(n29104));
    SB_LUT4 add_5260_5_lut (.I0(GND_net), .I1(n10011[2]), .I2(n341), .I3(n29102), 
            .O(n10002[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5260_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5260_5 (.CI(n29102), .I0(n10011[2]), .I1(n341), .CO(n29103));
    SB_LUT4 add_5260_4_lut (.I0(GND_net), .I1(n10011[1]), .I2(n268_adj_4361), 
            .I3(n29101), .O(n10002[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5260_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5260_4 (.CI(n29101), .I0(n10011[1]), .I1(n268_adj_4361), 
            .CO(n29102));
    SB_LUT4 add_5260_3_lut (.I0(GND_net), .I1(n10011[0]), .I2(n195), .I3(n29100), 
            .O(n10002[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5260_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5260_3 (.CI(n29100), .I0(n10011[0]), .I1(n195), .CO(n29101));
    SB_LUT4 add_5260_2_lut (.I0(GND_net), .I1(n53), .I2(n122), .I3(GND_net), 
            .O(n10002[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5260_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5260_2 (.CI(GND_net), .I0(n53), .I1(n122), .CO(n29100));
    SB_LUT4 add_5259_9_lut (.I0(GND_net), .I1(n10002[6]), .I2(n630), .I3(n29099), 
            .O(n9992[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5259_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5259_8_lut (.I0(GND_net), .I1(n10002[5]), .I2(n557), .I3(n29098), 
            .O(n9992[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5259_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5259_8 (.CI(n29098), .I0(n10002[5]), .I1(n557), .CO(n29099));
    SB_LUT4 add_5259_7_lut (.I0(GND_net), .I1(n10002[4]), .I2(n484), .I3(n29097), 
            .O(n9992[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5259_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5259_7 (.CI(n29097), .I0(n10002[4]), .I1(n484), .CO(n29098));
    SB_LUT4 add_5259_6_lut (.I0(GND_net), .I1(n10002[3]), .I2(n411), .I3(n29096), 
            .O(n9992[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5259_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5259_6 (.CI(n29096), .I0(n10002[3]), .I1(n411), .CO(n29097));
    SB_LUT4 add_5259_5_lut (.I0(GND_net), .I1(n10002[2]), .I2(n338), .I3(n29095), 
            .O(n9992[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5259_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5259_5 (.CI(n29095), .I0(n10002[2]), .I1(n338), .CO(n29096));
    SB_LUT4 add_5259_4_lut (.I0(GND_net), .I1(n10002[1]), .I2(n265_adj_4357), 
            .I3(n29094), .O(n9992[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5259_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5259_4 (.CI(n29094), .I0(n10002[1]), .I1(n265_adj_4357), 
            .CO(n29095));
    SB_LUT4 add_5259_3_lut (.I0(GND_net), .I1(n10002[0]), .I2(n192), .I3(n29093), 
            .O(n9992[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5259_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5259_3 (.CI(n29093), .I0(n10002[0]), .I1(n192), .CO(n29094));
    SB_LUT4 add_5259_2_lut (.I0(GND_net), .I1(n50), .I2(n119), .I3(GND_net), 
            .O(n9992[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5259_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5259_2 (.CI(GND_net), .I0(n50), .I1(n119), .CO(n29093));
    SB_LUT4 add_5258_10_lut (.I0(GND_net), .I1(n9992[7]), .I2(n700), .I3(n29092), 
            .O(n9981[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5258_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5258_9_lut (.I0(GND_net), .I1(n9992[6]), .I2(n627), .I3(n29091), 
            .O(n9981[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5258_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5258_9 (.CI(n29091), .I0(n9992[6]), .I1(n627), .CO(n29092));
    SB_LUT4 add_5258_8_lut (.I0(GND_net), .I1(n9992[5]), .I2(n554), .I3(n29090), 
            .O(n9981[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5258_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5258_8 (.CI(n29090), .I0(n9992[5]), .I1(n554), .CO(n29091));
    SB_LUT4 add_5258_7_lut (.I0(GND_net), .I1(n9992[4]), .I2(n481), .I3(n29089), 
            .O(n9981[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5258_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5258_7 (.CI(n29089), .I0(n9992[4]), .I1(n481), .CO(n29090));
    SB_LUT4 add_5258_6_lut (.I0(GND_net), .I1(n9992[3]), .I2(n408), .I3(n29088), 
            .O(n9981[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5258_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5258_6 (.CI(n29088), .I0(n9992[3]), .I1(n408), .CO(n29089));
    SB_LUT4 add_5258_5_lut (.I0(GND_net), .I1(n9992[2]), .I2(n335), .I3(n29087), 
            .O(n9981[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5258_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5258_5 (.CI(n29087), .I0(n9992[2]), .I1(n335), .CO(n29088));
    SB_LUT4 add_5258_4_lut (.I0(GND_net), .I1(n9992[1]), .I2(n262_adj_4350), 
            .I3(n29086), .O(n9981[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5258_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5258_4 (.CI(n29086), .I0(n9992[1]), .I1(n262_adj_4350), 
            .CO(n29087));
    SB_LUT4 add_5258_3_lut (.I0(GND_net), .I1(n9992[0]), .I2(n189_adj_4349), 
            .I3(n29085), .O(n9981[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5258_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5258_3 (.CI(n29085), .I0(n9992[0]), .I1(n189_adj_4349), 
            .CO(n29086));
    SB_LUT4 add_5258_2_lut (.I0(GND_net), .I1(n47), .I2(n116), .I3(GND_net), 
            .O(n9981[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5258_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5258_2 (.CI(GND_net), .I0(n47), .I1(n116), .CO(n29085));
    SB_LUT4 add_5257_11_lut (.I0(GND_net), .I1(n9981[8]), .I2(n770), .I3(n29084), 
            .O(n9969[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5257_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5257_10_lut (.I0(GND_net), .I1(n9981[7]), .I2(n697), .I3(n29083), 
            .O(n9969[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5257_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5257_10 (.CI(n29083), .I0(n9981[7]), .I1(n697), .CO(n29084));
    SB_LUT4 add_5257_9_lut (.I0(GND_net), .I1(n9981[6]), .I2(n624), .I3(n29082), 
            .O(n9969[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5257_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5257_9 (.CI(n29082), .I0(n9981[6]), .I1(n624), .CO(n29083));
    SB_LUT4 add_5257_8_lut (.I0(GND_net), .I1(n9981[5]), .I2(n551), .I3(n29081), 
            .O(n9969[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5257_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5257_8 (.CI(n29081), .I0(n9981[5]), .I1(n551), .CO(n29082));
    SB_LUT4 add_5257_7_lut (.I0(GND_net), .I1(n9981[4]), .I2(n478), .I3(n29080), 
            .O(n9969[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5257_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5257_7 (.CI(n29080), .I0(n9981[4]), .I1(n478), .CO(n29081));
    SB_LUT4 add_5257_6_lut (.I0(GND_net), .I1(n9981[3]), .I2(n405), .I3(n29079), 
            .O(n9969[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5257_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5257_6 (.CI(n29079), .I0(n9981[3]), .I1(n405), .CO(n29080));
    SB_LUT4 add_5257_5_lut (.I0(GND_net), .I1(n9981[2]), .I2(n332), .I3(n29078), 
            .O(n9969[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5257_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5257_5 (.CI(n29078), .I0(n9981[2]), .I1(n332), .CO(n29079));
    SB_LUT4 add_5257_4_lut (.I0(GND_net), .I1(n9981[1]), .I2(n259_adj_4347), 
            .I3(n29077), .O(n9969[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5257_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5257_4 (.CI(n29077), .I0(n9981[1]), .I1(n259_adj_4347), 
            .CO(n29078));
    SB_LUT4 add_5257_3_lut (.I0(GND_net), .I1(n9981[0]), .I2(n186), .I3(n29076), 
            .O(n9969[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5257_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5257_3 (.CI(n29076), .I0(n9981[0]), .I1(n186), .CO(n29077));
    SB_LUT4 add_5257_2_lut (.I0(GND_net), .I1(n44), .I2(n113), .I3(GND_net), 
            .O(n9969[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5257_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5257_2 (.CI(GND_net), .I0(n44), .I1(n113), .CO(n29076));
    SB_LUT4 add_5256_12_lut (.I0(GND_net), .I1(n9969[9]), .I2(n840), .I3(n29075), 
            .O(n9956[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5256_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5256_11_lut (.I0(GND_net), .I1(n9969[8]), .I2(n767), .I3(n29074), 
            .O(n9956[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5256_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5256_11 (.CI(n29074), .I0(n9969[8]), .I1(n767), .CO(n29075));
    SB_LUT4 add_5256_10_lut (.I0(GND_net), .I1(n9969[7]), .I2(n694), .I3(n29073), 
            .O(n9956[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5256_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5256_10 (.CI(n29073), .I0(n9969[7]), .I1(n694), .CO(n29074));
    SB_LUT4 add_5256_9_lut (.I0(GND_net), .I1(n9969[6]), .I2(n621), .I3(n29072), 
            .O(n9956[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5256_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5256_9 (.CI(n29072), .I0(n9969[6]), .I1(n621), .CO(n29073));
    SB_LUT4 add_5256_8_lut (.I0(GND_net), .I1(n9969[5]), .I2(n548), .I3(n29071), 
            .O(n9956[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5256_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5256_8 (.CI(n29071), .I0(n9969[5]), .I1(n548), .CO(n29072));
    SB_LUT4 add_5256_7_lut (.I0(GND_net), .I1(n9969[4]), .I2(n475), .I3(n29070), 
            .O(n9956[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5256_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5256_7 (.CI(n29070), .I0(n9969[4]), .I1(n475), .CO(n29071));
    SB_LUT4 add_5256_6_lut (.I0(GND_net), .I1(n9969[3]), .I2(n402), .I3(n29069), 
            .O(n9956[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5256_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5256_6 (.CI(n29069), .I0(n9969[3]), .I1(n402), .CO(n29070));
    SB_LUT4 add_5256_5_lut (.I0(GND_net), .I1(n9969[2]), .I2(n329), .I3(n29068), 
            .O(n9956[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5256_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5256_5 (.CI(n29068), .I0(n9969[2]), .I1(n329), .CO(n29069));
    SB_LUT4 add_5256_4_lut (.I0(GND_net), .I1(n9969[1]), .I2(n256_adj_4345), 
            .I3(n29067), .O(n9956[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5256_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5256_4 (.CI(n29067), .I0(n9969[1]), .I1(n256_adj_4345), 
            .CO(n29068));
    SB_LUT4 add_5256_3_lut (.I0(GND_net), .I1(n9969[0]), .I2(n183), .I3(n29066), 
            .O(n9956[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5256_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5256_3 (.CI(n29066), .I0(n9969[0]), .I1(n183), .CO(n29067));
    SB_LUT4 add_5256_2_lut (.I0(GND_net), .I1(n41_adj_4344), .I2(n110), 
            .I3(GND_net), .O(n9956[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5256_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5256_2 (.CI(GND_net), .I0(n41_adj_4344), .I1(n110), .CO(n29066));
    SB_LUT4 add_5255_13_lut (.I0(GND_net), .I1(n9956[10]), .I2(n910), 
            .I3(n29065), .O(n9942[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5255_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5255_12_lut (.I0(GND_net), .I1(n9956[9]), .I2(n837), .I3(n29064), 
            .O(n9942[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5255_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5255_12 (.CI(n29064), .I0(n9956[9]), .I1(n837), .CO(n29065));
    SB_LUT4 add_5255_11_lut (.I0(GND_net), .I1(n9956[8]), .I2(n764), .I3(n29063), 
            .O(n9942[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5255_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5255_11 (.CI(n29063), .I0(n9956[8]), .I1(n764), .CO(n29064));
    SB_LUT4 add_5255_10_lut (.I0(GND_net), .I1(n9956[7]), .I2(n691), .I3(n29062), 
            .O(n9942[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5255_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5255_10 (.CI(n29062), .I0(n9956[7]), .I1(n691), .CO(n29063));
    SB_LUT4 add_5255_9_lut (.I0(GND_net), .I1(n9956[6]), .I2(n618), .I3(n29061), 
            .O(n9942[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5255_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5255_9 (.CI(n29061), .I0(n9956[6]), .I1(n618), .CO(n29062));
    SB_LUT4 add_5255_8_lut (.I0(GND_net), .I1(n9956[5]), .I2(n545), .I3(n29060), 
            .O(n9942[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5255_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5255_8 (.CI(n29060), .I0(n9956[5]), .I1(n545), .CO(n29061));
    SB_LUT4 add_5255_7_lut (.I0(GND_net), .I1(n9956[4]), .I2(n472), .I3(n29059), 
            .O(n9942[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5255_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5255_7 (.CI(n29059), .I0(n9956[4]), .I1(n472), .CO(n29060));
    SB_LUT4 add_5255_6_lut (.I0(GND_net), .I1(n9956[3]), .I2(n399), .I3(n29058), 
            .O(n9942[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5255_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5255_6 (.CI(n29058), .I0(n9956[3]), .I1(n399), .CO(n29059));
    SB_LUT4 add_5255_5_lut (.I0(GND_net), .I1(n9956[2]), .I2(n326), .I3(n29057), 
            .O(n9942[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5255_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5255_5 (.CI(n29057), .I0(n9956[2]), .I1(n326), .CO(n29058));
    SB_LUT4 add_5255_4_lut (.I0(GND_net), .I1(n9956[1]), .I2(n253), .I3(n29056), 
            .O(n9942[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5255_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5255_4 (.CI(n29056), .I0(n9956[1]), .I1(n253), .CO(n29057));
    SB_LUT4 add_5255_3_lut (.I0(GND_net), .I1(n9956[0]), .I2(n180), .I3(n29055), 
            .O(n9942[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5255_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5255_3 (.CI(n29055), .I0(n9956[0]), .I1(n180), .CO(n29056));
    SB_LUT4 add_5255_2_lut (.I0(GND_net), .I1(n38), .I2(n107), .I3(GND_net), 
            .O(n9942[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5255_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5255_2 (.CI(GND_net), .I0(n38), .I1(n107), .CO(n29055));
    SB_LUT4 add_5254_14_lut (.I0(GND_net), .I1(n9942[11]), .I2(n980), 
            .I3(n29054), .O(n9927[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5254_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5254_13_lut (.I0(GND_net), .I1(n9942[10]), .I2(n907), 
            .I3(n29053), .O(n9927[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5254_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5254_13 (.CI(n29053), .I0(n9942[10]), .I1(n907), .CO(n29054));
    SB_LUT4 add_5254_12_lut (.I0(GND_net), .I1(n9942[9]), .I2(n834), .I3(n29052), 
            .O(n9927[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5254_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5254_12 (.CI(n29052), .I0(n9942[9]), .I1(n834), .CO(n29053));
    SB_LUT4 add_5254_11_lut (.I0(GND_net), .I1(n9942[8]), .I2(n761), .I3(n29051), 
            .O(n9927[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5254_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5254_11 (.CI(n29051), .I0(n9942[8]), .I1(n761), .CO(n29052));
    SB_LUT4 add_5254_10_lut (.I0(GND_net), .I1(n9942[7]), .I2(n688), .I3(n29050), 
            .O(n9927[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5254_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5254_10 (.CI(n29050), .I0(n9942[7]), .I1(n688), .CO(n29051));
    SB_LUT4 add_5254_9_lut (.I0(GND_net), .I1(n9942[6]), .I2(n615), .I3(n29049), 
            .O(n9927[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5254_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5254_9 (.CI(n29049), .I0(n9942[6]), .I1(n615), .CO(n29050));
    SB_LUT4 add_5254_8_lut (.I0(GND_net), .I1(n9942[5]), .I2(n542), .I3(n29048), 
            .O(n9927[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5254_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5254_8 (.CI(n29048), .I0(n9942[5]), .I1(n542), .CO(n29049));
    SB_LUT4 add_5254_7_lut (.I0(GND_net), .I1(n9942[4]), .I2(n469), .I3(n29047), 
            .O(n9927[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5254_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5254_7 (.CI(n29047), .I0(n9942[4]), .I1(n469), .CO(n29048));
    SB_LUT4 add_5254_6_lut (.I0(GND_net), .I1(n9942[3]), .I2(n396), .I3(n29046), 
            .O(n9927[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5254_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5254_6 (.CI(n29046), .I0(n9942[3]), .I1(n396), .CO(n29047));
    SB_LUT4 add_5254_5_lut (.I0(GND_net), .I1(n9942[2]), .I2(n323), .I3(n29045), 
            .O(n9927[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5254_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5254_5 (.CI(n29045), .I0(n9942[2]), .I1(n323), .CO(n29046));
    SB_LUT4 add_5254_4_lut (.I0(GND_net), .I1(n9942[1]), .I2(n250), .I3(n29044), 
            .O(n9927[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5254_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5254_4 (.CI(n29044), .I0(n9942[1]), .I1(n250), .CO(n29045));
    SB_LUT4 add_5254_3_lut (.I0(GND_net), .I1(n9942[0]), .I2(n177), .I3(n29043), 
            .O(n9927[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5254_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5254_3 (.CI(n29043), .I0(n9942[0]), .I1(n177), .CO(n29044));
    SB_LUT4 add_5254_2_lut (.I0(GND_net), .I1(n35), .I2(n104), .I3(GND_net), 
            .O(n9927[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5254_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5254_2 (.CI(GND_net), .I0(n35), .I1(n104), .CO(n29043));
    SB_LUT4 add_5253_15_lut (.I0(GND_net), .I1(n9927[12]), .I2(n1050), 
            .I3(n29042), .O(n9911[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5253_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5253_14_lut (.I0(GND_net), .I1(n9927[11]), .I2(n977), 
            .I3(n29041), .O(n9911[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5253_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5253_14 (.CI(n29041), .I0(n9927[11]), .I1(n977), .CO(n29042));
    SB_LUT4 add_5253_13_lut (.I0(GND_net), .I1(n9927[10]), .I2(n904), 
            .I3(n29040), .O(n9911[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5253_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5253_13 (.CI(n29040), .I0(n9927[10]), .I1(n904), .CO(n29041));
    SB_LUT4 add_5253_12_lut (.I0(GND_net), .I1(n9927[9]), .I2(n831), .I3(n29039), 
            .O(n9911[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5253_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5253_12 (.CI(n29039), .I0(n9927[9]), .I1(n831), .CO(n29040));
    SB_LUT4 add_5253_11_lut (.I0(GND_net), .I1(n9927[8]), .I2(n758), .I3(n29038), 
            .O(n9911[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5253_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5253_11 (.CI(n29038), .I0(n9927[8]), .I1(n758), .CO(n29039));
    SB_LUT4 add_5253_10_lut (.I0(GND_net), .I1(n9927[7]), .I2(n685), .I3(n29037), 
            .O(n9911[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5253_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5253_10 (.CI(n29037), .I0(n9927[7]), .I1(n685), .CO(n29038));
    SB_LUT4 add_5253_9_lut (.I0(GND_net), .I1(n9927[6]), .I2(n612), .I3(n29036), 
            .O(n9911[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5253_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5253_9 (.CI(n29036), .I0(n9927[6]), .I1(n612), .CO(n29037));
    SB_LUT4 add_5253_8_lut (.I0(GND_net), .I1(n9927[5]), .I2(n539), .I3(n29035), 
            .O(n9911[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5253_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5253_8 (.CI(n29035), .I0(n9927[5]), .I1(n539), .CO(n29036));
    SB_LUT4 add_5253_7_lut (.I0(GND_net), .I1(n9927[4]), .I2(n466), .I3(n29034), 
            .O(n9911[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5253_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5253_7 (.CI(n29034), .I0(n9927[4]), .I1(n466), .CO(n29035));
    SB_LUT4 add_5253_6_lut (.I0(GND_net), .I1(n9927[3]), .I2(n393), .I3(n29033), 
            .O(n9911[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5253_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5253_6 (.CI(n29033), .I0(n9927[3]), .I1(n393), .CO(n29034));
    SB_LUT4 add_5253_5_lut (.I0(GND_net), .I1(n9927[2]), .I2(n320), .I3(n29032), 
            .O(n9911[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5253_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5253_5 (.CI(n29032), .I0(n9927[2]), .I1(n320), .CO(n29033));
    SB_LUT4 add_5253_4_lut (.I0(GND_net), .I1(n9927[1]), .I2(n247), .I3(n29031), 
            .O(n9911[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5253_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5253_4 (.CI(n29031), .I0(n9927[1]), .I1(n247), .CO(n29032));
    SB_LUT4 add_5253_3_lut (.I0(GND_net), .I1(n9927[0]), .I2(n174), .I3(n29030), 
            .O(n9911[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5253_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5253_3 (.CI(n29030), .I0(n9927[0]), .I1(n174), .CO(n29031));
    SB_LUT4 add_5253_2_lut (.I0(GND_net), .I1(n32), .I2(n101), .I3(GND_net), 
            .O(n9911[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5253_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5253_2 (.CI(GND_net), .I0(n32), .I1(n101), .CO(n29030));
    SB_LUT4 add_5252_16_lut (.I0(GND_net), .I1(n9911[13]), .I2(n1120), 
            .I3(n29029), .O(n9894[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5252_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5252_15_lut (.I0(GND_net), .I1(n9911[12]), .I2(n1047), 
            .I3(n29028), .O(n9894[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5252_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5252_15 (.CI(n29028), .I0(n9911[12]), .I1(n1047), .CO(n29029));
    SB_LUT4 add_5252_14_lut (.I0(GND_net), .I1(n9911[11]), .I2(n974), 
            .I3(n29027), .O(n9894[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5252_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5252_14 (.CI(n29027), .I0(n9911[11]), .I1(n974), .CO(n29028));
    SB_LUT4 add_5252_13_lut (.I0(GND_net), .I1(n9911[10]), .I2(n901), 
            .I3(n29026), .O(n9894[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5252_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5252_13 (.CI(n29026), .I0(n9911[10]), .I1(n901), .CO(n29027));
    SB_LUT4 add_5252_12_lut (.I0(GND_net), .I1(n9911[9]), .I2(n828), .I3(n29025), 
            .O(n9894[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5252_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5252_12 (.CI(n29025), .I0(n9911[9]), .I1(n828), .CO(n29026));
    SB_LUT4 add_5252_11_lut (.I0(GND_net), .I1(n9911[8]), .I2(n755), .I3(n29024), 
            .O(n9894[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5252_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5252_11 (.CI(n29024), .I0(n9911[8]), .I1(n755), .CO(n29025));
    SB_LUT4 add_5252_10_lut (.I0(GND_net), .I1(n9911[7]), .I2(n682), .I3(n29023), 
            .O(n9894[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5252_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5252_10 (.CI(n29023), .I0(n9911[7]), .I1(n682), .CO(n29024));
    SB_LUT4 add_5252_9_lut (.I0(GND_net), .I1(n9911[6]), .I2(n609), .I3(n29022), 
            .O(n9894[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5252_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5252_9 (.CI(n29022), .I0(n9911[6]), .I1(n609), .CO(n29023));
    SB_LUT4 add_5252_8_lut (.I0(GND_net), .I1(n9911[5]), .I2(n536), .I3(n29021), 
            .O(n9894[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5252_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5252_8 (.CI(n29021), .I0(n9911[5]), .I1(n536), .CO(n29022));
    SB_DFF result_i2 (.Q(duty[2]), .C(clk32MHz), .D(duty_23__N_3522[2]));   // verilog/motorControl.v(29[14] 48[8])
    SB_LUT4 add_5252_7_lut (.I0(GND_net), .I1(n9911[4]), .I2(n463), .I3(n29020), 
            .O(n9894[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5252_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5252_7 (.CI(n29020), .I0(n9911[4]), .I1(n463), .CO(n29021));
    SB_LUT4 add_5252_6_lut (.I0(GND_net), .I1(n9911[3]), .I2(n390), .I3(n29019), 
            .O(n9894[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5252_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5252_6 (.CI(n29019), .I0(n9911[3]), .I1(n390), .CO(n29020));
    SB_LUT4 add_5252_5_lut (.I0(GND_net), .I1(n9911[2]), .I2(n317), .I3(n29018), 
            .O(n9894[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5252_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i302_2_lut (.I0(\Kp[6] ), .I1(n28[3]), .I2(GND_net), 
            .I3(GND_net), .O(n448_adj_4688));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i302_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5252_5 (.CI(n29018), .I0(n9911[2]), .I1(n317), .CO(n29019));
    SB_LUT4 add_5252_4_lut (.I0(GND_net), .I1(n9911[1]), .I2(n244), .I3(n29017), 
            .O(n9894[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5252_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5252_4 (.CI(n29017), .I0(n9911[1]), .I1(n244), .CO(n29018));
    SB_LUT4 add_5252_3_lut (.I0(GND_net), .I1(n9911[0]), .I2(n171), .I3(n29016), 
            .O(n9894[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5252_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5252_3 (.CI(n29016), .I0(n9911[0]), .I1(n171), .CO(n29017));
    SB_LUT4 mult_10_i351_2_lut (.I0(\Kp[7] ), .I1(n28[3]), .I2(GND_net), 
            .I3(GND_net), .O(n521_adj_4689));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i351_2_lut.LUT_INIT = 16'h8888;
    SB_DFF result_i3 (.Q(duty[3]), .C(clk32MHz), .D(duty_23__N_3522[3]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i4 (.Q(duty[4]), .C(clk32MHz), .D(duty_23__N_3522[4]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i5 (.Q(duty[5]), .C(clk32MHz), .D(duty_23__N_3522[5]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i6 (.Q(duty[6]), .C(clk32MHz), .D(duty_23__N_3522[6]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i7 (.Q(duty[7]), .C(clk32MHz), .D(duty_23__N_3522[7]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i8 (.Q(duty[8]), .C(clk32MHz), .D(duty_23__N_3522[8]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i9 (.Q(duty[9]), .C(clk32MHz), .D(duty_23__N_3522[9]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i10 (.Q(duty[10]), .C(clk32MHz), .D(duty_23__N_3522[10]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i11 (.Q(duty[11]), .C(clk32MHz), .D(duty_23__N_3522[11]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i12 (.Q(duty[12]), .C(clk32MHz), .D(duty_23__N_3522[12]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i13 (.Q(duty[13]), .C(clk32MHz), .D(duty_23__N_3522[13]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i14 (.Q(duty[14]), .C(clk32MHz), .D(duty_23__N_3522[14]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i15 (.Q(duty[15]), .C(clk32MHz), .D(duty_23__N_3522[15]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i16 (.Q(duty[16]), .C(clk32MHz), .D(duty_23__N_3522[16]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i17 (.Q(duty[17]), .C(clk32MHz), .D(duty_23__N_3522[17]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i18 (.Q(duty[18]), .C(clk32MHz), .D(duty_23__N_3522[18]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i19 (.Q(duty[19]), .C(clk32MHz), .D(duty_23__N_3522[19]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i20 (.Q(duty[20]), .C(clk32MHz), .D(duty_23__N_3522[20]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i21 (.Q(duty[21]), .C(clk32MHz), .D(duty_23__N_3522[21]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i22 (.Q(duty[22]), .C(clk32MHz), .D(duty_23__N_3522[22]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i23 (.Q(duty[23]), .C(clk32MHz), .D(duty_23__N_3522[23]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.integral_i1  (.Q(\PID_CONTROLLER.integral [1]), 
           .C(clk32MHz), .D(\PID_CONTROLLER.integral_23__N_3546 [1]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.integral_i2  (.Q(\PID_CONTROLLER.integral [2]), 
           .C(clk32MHz), .D(\PID_CONTROLLER.integral_23__N_3546 [2]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.integral_i3  (.Q(\PID_CONTROLLER.integral [3]), 
           .C(clk32MHz), .D(\PID_CONTROLLER.integral_23__N_3546 [3]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.integral_i4  (.Q(\PID_CONTROLLER.integral [4]), 
           .C(clk32MHz), .D(\PID_CONTROLLER.integral_23__N_3546 [4]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.integral_i5  (.Q(\PID_CONTROLLER.integral [5]), 
           .C(clk32MHz), .D(\PID_CONTROLLER.integral_23__N_3546 [5]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.integral_i6  (.Q(\PID_CONTROLLER.integral [6]), 
           .C(clk32MHz), .D(\PID_CONTROLLER.integral_23__N_3546 [6]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.integral_i7  (.Q(\PID_CONTROLLER.integral [7]), 
           .C(clk32MHz), .D(\PID_CONTROLLER.integral_23__N_3546 [7]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.integral_i8  (.Q(\PID_CONTROLLER.integral [8]), 
           .C(clk32MHz), .D(\PID_CONTROLLER.integral_23__N_3546 [8]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.integral_i9  (.Q(\PID_CONTROLLER.integral [9]), 
           .C(clk32MHz), .D(\PID_CONTROLLER.integral_23__N_3546 [9]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.integral_i10  (.Q(\PID_CONTROLLER.integral [10]), 
           .C(clk32MHz), .D(\PID_CONTROLLER.integral_23__N_3546 [10]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.integral_i11  (.Q(\PID_CONTROLLER.integral [11]), 
           .C(clk32MHz), .D(\PID_CONTROLLER.integral_23__N_3546 [11]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.integral_i12  (.Q(\PID_CONTROLLER.integral [12]), 
           .C(clk32MHz), .D(\PID_CONTROLLER.integral_23__N_3546 [12]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.integral_i13  (.Q(\PID_CONTROLLER.integral [13]), 
           .C(clk32MHz), .D(\PID_CONTROLLER.integral_23__N_3546 [13]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.integral_i14  (.Q(\PID_CONTROLLER.integral [14]), 
           .C(clk32MHz), .D(\PID_CONTROLLER.integral_23__N_3546 [14]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.integral_i15  (.Q(\PID_CONTROLLER.integral [15]), 
           .C(clk32MHz), .D(\PID_CONTROLLER.integral_23__N_3546 [15]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.integral_i16  (.Q(\PID_CONTROLLER.integral [16]), 
           .C(clk32MHz), .D(\PID_CONTROLLER.integral_23__N_3546 [16]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.integral_i17  (.Q(\PID_CONTROLLER.integral [17]), 
           .C(clk32MHz), .D(\PID_CONTROLLER.integral_23__N_3546 [17]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.integral_i18  (.Q(\PID_CONTROLLER.integral [18]), 
           .C(clk32MHz), .D(\PID_CONTROLLER.integral_23__N_3546 [18]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.integral_i19  (.Q(\PID_CONTROLLER.integral [19]), 
           .C(clk32MHz), .D(\PID_CONTROLLER.integral_23__N_3546 [19]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.integral_i20  (.Q(\PID_CONTROLLER.integral [20]), 
           .C(clk32MHz), .D(\PID_CONTROLLER.integral_23__N_3546 [20]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.integral_i21  (.Q(\PID_CONTROLLER.integral [21]), 
           .C(clk32MHz), .D(\PID_CONTROLLER.integral_23__N_3546 [21]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.integral_i22  (.Q(\PID_CONTROLLER.integral [22]), 
           .C(clk32MHz), .D(\PID_CONTROLLER.integral_23__N_3546 [22]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.integral_i23  (.Q(\PID_CONTROLLER.integral [23]), 
           .C(clk32MHz), .D(\PID_CONTROLLER.integral_23__N_3546 [23]));   // verilog/motorControl.v(29[14] 48[8])
    SB_LUT4 add_5252_2_lut (.I0(GND_net), .I1(n29), .I2(n98), .I3(GND_net), 
            .O(n9894[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5252_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5252_2 (.CI(GND_net), .I0(n29), .I1(n98), .CO(n29016));
    SB_LUT4 add_5251_17_lut (.I0(GND_net), .I1(n9894[14]), .I2(GND_net), 
            .I3(n29015), .O(n9876[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5251_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5251_16_lut (.I0(GND_net), .I1(n9894[13]), .I2(n1117), 
            .I3(n29014), .O(n9876[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5251_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5251_16 (.CI(n29014), .I0(n9894[13]), .I1(n1117), .CO(n29015));
    SB_LUT4 add_5251_15_lut (.I0(GND_net), .I1(n9894[12]), .I2(n1044), 
            .I3(n29013), .O(n9876[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5251_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5251_15 (.CI(n29013), .I0(n9894[12]), .I1(n1044), .CO(n29014));
    SB_LUT4 add_5251_14_lut (.I0(GND_net), .I1(n9894[11]), .I2(n971), 
            .I3(n29012), .O(n9876[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5251_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5251_14 (.CI(n29012), .I0(n9894[11]), .I1(n971), .CO(n29013));
    SB_LUT4 add_5251_13_lut (.I0(GND_net), .I1(n9894[10]), .I2(n898), 
            .I3(n29011), .O(n9876[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5251_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5251_13 (.CI(n29011), .I0(n9894[10]), .I1(n898), .CO(n29012));
    SB_LUT4 add_5251_12_lut (.I0(GND_net), .I1(n9894[9]), .I2(n825), .I3(n29010), 
            .O(n9876[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5251_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i400_2_lut (.I0(\Kp[8] ), .I1(n28[3]), .I2(GND_net), 
            .I3(GND_net), .O(n594_adj_4690));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i400_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5251_12 (.CI(n29010), .I0(n9894[9]), .I1(n825), .CO(n29011));
    SB_LUT4 add_5251_11_lut (.I0(GND_net), .I1(n9894[8]), .I2(n752), .I3(n29009), 
            .O(n9876[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5251_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5251_11 (.CI(n29009), .I0(n9894[8]), .I1(n752), .CO(n29010));
    SB_LUT4 add_5251_10_lut (.I0(GND_net), .I1(n9894[7]), .I2(n679), .I3(n29008), 
            .O(n9876[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5251_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5251_10 (.CI(n29008), .I0(n9894[7]), .I1(n679), .CO(n29009));
    SB_LUT4 add_5251_9_lut (.I0(GND_net), .I1(n9894[6]), .I2(n606), .I3(n29007), 
            .O(n9876[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5251_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5251_9 (.CI(n29007), .I0(n9894[6]), .I1(n606), .CO(n29008));
    SB_LUT4 mult_10_i449_2_lut (.I0(\Kp[9] ), .I1(n28[3]), .I2(GND_net), 
            .I3(GND_net), .O(n667_adj_4691));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i449_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5251_8_lut (.I0(GND_net), .I1(n9894[5]), .I2(n533), .I3(n29006), 
            .O(n9876[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5251_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5251_8 (.CI(n29006), .I0(n9894[5]), .I1(n533), .CO(n29007));
    SB_LUT4 add_5251_7_lut (.I0(GND_net), .I1(n9894[4]), .I2(n460), .I3(n29005), 
            .O(n9876[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5251_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5251_7 (.CI(n29005), .I0(n9894[4]), .I1(n460), .CO(n29006));
    SB_LUT4 add_5251_6_lut (.I0(GND_net), .I1(n9894[3]), .I2(n387), .I3(n29004), 
            .O(n9876[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5251_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5251_6 (.CI(n29004), .I0(n9894[3]), .I1(n387), .CO(n29005));
    SB_LUT4 add_5251_5_lut (.I0(GND_net), .I1(n9894[2]), .I2(n314), .I3(n29003), 
            .O(n9876[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5251_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5251_5 (.CI(n29003), .I0(n9894[2]), .I1(n314), .CO(n29004));
    SB_LUT4 add_5251_4_lut (.I0(GND_net), .I1(n9894[1]), .I2(n241), .I3(n29002), 
            .O(n9876[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5251_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5251_4 (.CI(n29002), .I0(n9894[1]), .I1(n241), .CO(n29003));
    SB_LUT4 add_5251_3_lut (.I0(GND_net), .I1(n9894[0]), .I2(n168), .I3(n29001), 
            .O(n9876[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5251_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5251_3 (.CI(n29001), .I0(n9894[0]), .I1(n168), .CO(n29002));
    SB_LUT4 add_5251_2_lut (.I0(GND_net), .I1(n26_adj_4313), .I2(n95), 
            .I3(GND_net), .O(n9876[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5251_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5251_2 (.CI(GND_net), .I0(n26_adj_4313), .I1(n95), .CO(n29001));
    SB_LUT4 add_5250_18_lut (.I0(GND_net), .I1(n9876[15]), .I2(GND_net), 
            .I3(n29000), .O(n9857[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5250_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5250_17_lut (.I0(GND_net), .I1(n9876[14]), .I2(GND_net), 
            .I3(n28999), .O(n9857[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5250_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5250_17 (.CI(n28999), .I0(n9876[14]), .I1(GND_net), .CO(n29000));
    SB_LUT4 add_5250_16_lut (.I0(GND_net), .I1(n9876[13]), .I2(n1114), 
            .I3(n28998), .O(n9857[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5250_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5250_16 (.CI(n28998), .I0(n9876[13]), .I1(n1114), .CO(n28999));
    SB_LUT4 add_5250_15_lut (.I0(GND_net), .I1(n9876[12]), .I2(n1041), 
            .I3(n28997), .O(n9857[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5250_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5250_15 (.CI(n28997), .I0(n9876[12]), .I1(n1041), .CO(n28998));
    SB_LUT4 add_5250_14_lut (.I0(GND_net), .I1(n9876[11]), .I2(n968), 
            .I3(n28996), .O(n9857[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5250_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5250_14 (.CI(n28996), .I0(n9876[11]), .I1(n968), .CO(n28997));
    SB_LUT4 add_5250_13_lut (.I0(GND_net), .I1(n9876[10]), .I2(n895), 
            .I3(n28995), .O(n9857[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5250_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5250_13 (.CI(n28995), .I0(n9876[10]), .I1(n895), .CO(n28996));
    SB_LUT4 add_5250_12_lut (.I0(GND_net), .I1(n9876[9]), .I2(n822), .I3(n28994), 
            .O(n9857[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5250_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5250_12 (.CI(n28994), .I0(n9876[9]), .I1(n822), .CO(n28995));
    SB_LUT4 add_5250_11_lut (.I0(GND_net), .I1(n9876[8]), .I2(n749), .I3(n28993), 
            .O(n9857[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5250_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5250_11 (.CI(n28993), .I0(n9876[8]), .I1(n749), .CO(n28994));
    SB_LUT4 add_5250_10_lut (.I0(GND_net), .I1(n9876[7]), .I2(n676), .I3(n28992), 
            .O(n9857[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5250_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5250_10 (.CI(n28992), .I0(n9876[7]), .I1(n676), .CO(n28993));
    SB_LUT4 add_5250_9_lut (.I0(GND_net), .I1(n9876[6]), .I2(n603), .I3(n28991), 
            .O(n9857[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5250_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5250_9 (.CI(n28991), .I0(n9876[6]), .I1(n603), .CO(n28992));
    SB_LUT4 add_5250_8_lut (.I0(GND_net), .I1(n9876[5]), .I2(n530), .I3(n28990), 
            .O(n9857[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5250_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5250_8 (.CI(n28990), .I0(n9876[5]), .I1(n530), .CO(n28991));
    SB_LUT4 add_5250_7_lut (.I0(GND_net), .I1(n9876[4]), .I2(n457), .I3(n28989), 
            .O(n9857[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5250_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5250_7 (.CI(n28989), .I0(n9876[4]), .I1(n457), .CO(n28990));
    SB_LUT4 add_5250_6_lut (.I0(GND_net), .I1(n9876[3]), .I2(n384), .I3(n28988), 
            .O(n9857[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5250_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5250_6 (.CI(n28988), .I0(n9876[3]), .I1(n384), .CO(n28989));
    SB_LUT4 add_5250_5_lut (.I0(GND_net), .I1(n9876[2]), .I2(n311), .I3(n28987), 
            .O(n9857[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5250_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5250_5 (.CI(n28987), .I0(n9876[2]), .I1(n311), .CO(n28988));
    SB_LUT4 add_5250_4_lut (.I0(GND_net), .I1(n9876[1]), .I2(n238), .I3(n28986), 
            .O(n9857[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5250_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5250_4 (.CI(n28986), .I0(n9876[1]), .I1(n238), .CO(n28987));
    SB_LUT4 add_5250_3_lut (.I0(GND_net), .I1(n9876[0]), .I2(n165), .I3(n28985), 
            .O(n9857[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5250_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5250_3 (.CI(n28985), .I0(n9876[0]), .I1(n165), .CO(n28986));
    SB_LUT4 add_5250_2_lut (.I0(GND_net), .I1(n23), .I2(n92), .I3(GND_net), 
            .O(n9857[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5250_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5250_2 (.CI(GND_net), .I0(n23), .I1(n92), .CO(n28985));
    SB_LUT4 add_5249_19_lut (.I0(GND_net), .I1(n9857[16]), .I2(GND_net), 
            .I3(n28984), .O(n9837[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5249_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5249_18_lut (.I0(GND_net), .I1(n9857[15]), .I2(GND_net), 
            .I3(n28983), .O(n9837[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5249_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5249_18 (.CI(n28983), .I0(n9857[15]), .I1(GND_net), .CO(n28984));
    SB_LUT4 add_5249_17_lut (.I0(GND_net), .I1(n9857[14]), .I2(GND_net), 
            .I3(n28982), .O(n9837[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5249_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5249_17 (.CI(n28982), .I0(n9857[14]), .I1(GND_net), .CO(n28983));
    SB_LUT4 add_5249_16_lut (.I0(GND_net), .I1(n9857[13]), .I2(n1111), 
            .I3(n28981), .O(n9837[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5249_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5249_16 (.CI(n28981), .I0(n9857[13]), .I1(n1111), .CO(n28982));
    SB_LUT4 add_5249_15_lut (.I0(GND_net), .I1(n9857[12]), .I2(n1038), 
            .I3(n28980), .O(n9837[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5249_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5249_15 (.CI(n28980), .I0(n9857[12]), .I1(n1038), .CO(n28981));
    SB_LUT4 add_5249_14_lut (.I0(GND_net), .I1(n9857[11]), .I2(n965), 
            .I3(n28979), .O(n9837[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5249_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5249_14 (.CI(n28979), .I0(n9857[11]), .I1(n965), .CO(n28980));
    SB_LUT4 add_5249_13_lut (.I0(GND_net), .I1(n9857[10]), .I2(n892), 
            .I3(n28978), .O(n9837[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5249_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5249_13 (.CI(n28978), .I0(n9857[10]), .I1(n892), .CO(n28979));
    SB_LUT4 add_5249_12_lut (.I0(GND_net), .I1(n9857[9]), .I2(n819), .I3(n28977), 
            .O(n9837[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5249_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5249_12 (.CI(n28977), .I0(n9857[9]), .I1(n819), .CO(n28978));
    SB_LUT4 add_5249_11_lut (.I0(GND_net), .I1(n9857[8]), .I2(n746), .I3(n28976), 
            .O(n9837[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5249_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5249_11 (.CI(n28976), .I0(n9857[8]), .I1(n746), .CO(n28977));
    SB_LUT4 add_5249_10_lut (.I0(GND_net), .I1(n9857[7]), .I2(n673), .I3(n28975), 
            .O(n9837[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5249_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5249_10 (.CI(n28975), .I0(n9857[7]), .I1(n673), .CO(n28976));
    SB_LUT4 add_5249_9_lut (.I0(GND_net), .I1(n9857[6]), .I2(n600), .I3(n28974), 
            .O(n9837[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5249_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5249_9 (.CI(n28974), .I0(n9857[6]), .I1(n600), .CO(n28975));
    SB_LUT4 add_5249_8_lut (.I0(GND_net), .I1(n9857[5]), .I2(n527), .I3(n28973), 
            .O(n9837[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5249_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5249_8 (.CI(n28973), .I0(n9857[5]), .I1(n527), .CO(n28974));
    SB_LUT4 add_5249_7_lut (.I0(GND_net), .I1(n9857[4]), .I2(n454), .I3(n28972), 
            .O(n9837[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5249_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5249_7 (.CI(n28972), .I0(n9857[4]), .I1(n454), .CO(n28973));
    SB_LUT4 add_5249_6_lut (.I0(GND_net), .I1(n9857[3]), .I2(n381), .I3(n28971), 
            .O(n9837[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5249_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5249_6 (.CI(n28971), .I0(n9857[3]), .I1(n381), .CO(n28972));
    SB_LUT4 add_5249_5_lut (.I0(GND_net), .I1(n9857[2]), .I2(n308), .I3(n28970), 
            .O(n9837[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5249_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i498_2_lut (.I0(\Kp[10] ), .I1(n28[3]), .I2(GND_net), 
            .I3(GND_net), .O(n740_adj_4692));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i498_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i547_2_lut (.I0(\Kp[11] ), .I1(n28[3]), .I2(GND_net), 
            .I3(GND_net), .O(n813_adj_4693));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i547_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_16_inv_0_i16_1_lut (.I0(PWMLimit[15]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4735[15]));   // verilog/motorControl.v(39[18:27])
    defparam unary_minus_16_inv_0_i16_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i596_2_lut (.I0(\Kp[12] ), .I1(n28[3]), .I2(GND_net), 
            .I3(GND_net), .O(n886_adj_4695));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i596_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i645_2_lut (.I0(\Kp[13] ), .I1(n28[3]), .I2(GND_net), 
            .I3(GND_net), .O(n959_adj_4696));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i645_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_16_inv_0_i17_1_lut (.I0(PWMLimit[16]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4735[16]));   // verilog/motorControl.v(39[18:27])
    defparam unary_minus_16_inv_0_i17_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i694_2_lut (.I0(\Kp[14] ), .I1(n28[3]), .I2(GND_net), 
            .I3(GND_net), .O(n1032_adj_4698));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i694_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i743_2_lut (.I0(\Kp[15] ), .I1(n28[3]), .I2(GND_net), 
            .I3(GND_net), .O(n1105_adj_4699));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i743_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i59_2_lut (.I0(\Kp[1] ), .I1(n28[4]), .I2(GND_net), 
            .I3(GND_net), .O(n86_adj_4700));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i59_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i12_2_lut (.I0(\Kp[0] ), .I1(n28[5]), .I2(GND_net), 
            .I3(GND_net), .O(n17_adj_4701));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i12_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_16_inv_0_i18_1_lut (.I0(PWMLimit[17]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4735[17]));   // verilog/motorControl.v(39[18:27])
    defparam unary_minus_16_inv_0_i18_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i108_2_lut (.I0(\Kp[2] ), .I1(n28[4]), .I2(GND_net), 
            .I3(GND_net), .O(n159_adj_4703));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i108_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_16_inv_0_i19_1_lut (.I0(PWMLimit[18]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4735[18]));   // verilog/motorControl.v(39[18:27])
    defparam unary_minus_16_inv_0_i19_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_16_inv_0_i20_1_lut (.I0(PWMLimit[19]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4735[19]));   // verilog/motorControl.v(39[18:27])
    defparam unary_minus_16_inv_0_i20_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_16_inv_0_i21_1_lut (.I0(PWMLimit[20]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4735[20]));   // verilog/motorControl.v(39[18:27])
    defparam unary_minus_16_inv_0_i21_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_5249_5 (.CI(n28970), .I0(n9857[2]), .I1(n308), .CO(n28971));
    SB_LUT4 add_5249_4_lut (.I0(GND_net), .I1(n9857[1]), .I2(n235), .I3(n28969), 
            .O(n9837[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5249_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5249_4 (.CI(n28969), .I0(n9857[1]), .I1(n235), .CO(n28970));
    SB_LUT4 add_5249_3_lut (.I0(GND_net), .I1(n9857[0]), .I2(n162), .I3(n28968), 
            .O(n9837[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5249_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5249_3 (.CI(n28968), .I0(n9857[0]), .I1(n162), .CO(n28969));
    SB_LUT4 add_5249_2_lut (.I0(GND_net), .I1(n20_adj_4707), .I2(n89_adj_4708), 
            .I3(GND_net), .O(n9837[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5249_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5249_2 (.CI(GND_net), .I0(n20_adj_4707), .I1(n89_adj_4708), 
            .CO(n28968));
    SB_LUT4 add_5248_20_lut (.I0(GND_net), .I1(n9837[17]), .I2(GND_net), 
            .I3(n28967), .O(n9816[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5248_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5248_19_lut (.I0(GND_net), .I1(n9837[16]), .I2(GND_net), 
            .I3(n28966), .O(n9816[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5248_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5248_19 (.CI(n28966), .I0(n9837[16]), .I1(GND_net), .CO(n28967));
    SB_LUT4 add_5248_18_lut (.I0(GND_net), .I1(n9837[15]), .I2(GND_net), 
            .I3(n28965), .O(n9816[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5248_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5248_18 (.CI(n28965), .I0(n9837[15]), .I1(GND_net), .CO(n28966));
    SB_LUT4 add_5248_17_lut (.I0(GND_net), .I1(n9837[14]), .I2(GND_net), 
            .I3(n28964), .O(n9816[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5248_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5248_17 (.CI(n28964), .I0(n9837[14]), .I1(GND_net), .CO(n28965));
    SB_LUT4 add_5248_16_lut (.I0(GND_net), .I1(n9837[13]), .I2(n1108_adj_4709), 
            .I3(n28963), .O(n9816[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5248_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5248_16 (.CI(n28963), .I0(n9837[13]), .I1(n1108_adj_4709), 
            .CO(n28964));
    SB_LUT4 add_5248_15_lut (.I0(GND_net), .I1(n9837[12]), .I2(n1035_adj_4710), 
            .I3(n28962), .O(n9816[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5248_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5248_15 (.CI(n28962), .I0(n9837[12]), .I1(n1035_adj_4710), 
            .CO(n28963));
    SB_LUT4 add_5248_14_lut (.I0(GND_net), .I1(n9837[11]), .I2(n962_adj_4711), 
            .I3(n28961), .O(n9816[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5248_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5248_14 (.CI(n28961), .I0(n9837[11]), .I1(n962_adj_4711), 
            .CO(n28962));
    SB_LUT4 add_5248_13_lut (.I0(GND_net), .I1(n9837[10]), .I2(n889_adj_4712), 
            .I3(n28960), .O(n9816[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5248_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5248_13 (.CI(n28960), .I0(n9837[10]), .I1(n889_adj_4712), 
            .CO(n28961));
    SB_LUT4 add_5248_12_lut (.I0(GND_net), .I1(n9837[9]), .I2(n816_adj_4713), 
            .I3(n28959), .O(n9816[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5248_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5248_12 (.CI(n28959), .I0(n9837[9]), .I1(n816_adj_4713), 
            .CO(n28960));
    SB_LUT4 add_5248_11_lut (.I0(GND_net), .I1(n9837[8]), .I2(n743_adj_4714), 
            .I3(n28958), .O(n9816[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5248_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5248_11 (.CI(n28958), .I0(n9837[8]), .I1(n743_adj_4714), 
            .CO(n28959));
    SB_LUT4 add_5248_10_lut (.I0(GND_net), .I1(n9837[7]), .I2(n670_adj_4715), 
            .I3(n28957), .O(n9816[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5248_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5248_10 (.CI(n28957), .I0(n9837[7]), .I1(n670_adj_4715), 
            .CO(n28958));
    SB_LUT4 add_5248_9_lut (.I0(GND_net), .I1(n9837[6]), .I2(n597_adj_4716), 
            .I3(n28956), .O(n9816[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5248_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5248_9 (.CI(n28956), .I0(n9837[6]), .I1(n597_adj_4716), 
            .CO(n28957));
    SB_LUT4 mult_10_i157_2_lut (.I0(\Kp[3] ), .I1(n28[4]), .I2(GND_net), 
            .I3(GND_net), .O(n232_adj_4717));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i157_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_16_inv_0_i22_1_lut (.I0(PWMLimit[21]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4735[21]));   // verilog/motorControl.v(39[18:27])
    defparam unary_minus_16_inv_0_i22_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_16_inv_0_i23_1_lut (.I0(PWMLimit[22]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4735[22]));   // verilog/motorControl.v(39[18:27])
    defparam unary_minus_16_inv_0_i23_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_16_inv_0_i24_1_lut (.I0(PWMLimit[23]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4735[23]));   // verilog/motorControl.v(39[18:27])
    defparam unary_minus_16_inv_0_i24_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i206_2_lut (.I0(\Kp[4] ), .I1(n28[4]), .I2(GND_net), 
            .I3(GND_net), .O(n305_adj_4721));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i206_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i19131_2_lut (.I0(n28[3]), .I1(\PID_CONTROLLER.integral_23__N_3594 ), 
            .I2(GND_net), .I3(GND_net), .O(n3302[3]));   // verilog/motorControl.v(31[7] 33[10])
    defparam i19131_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i610_2_lut (.I0(\Ki[12] ), .I1(\PID_CONTROLLER.integral_23__N_3546 [10]), 
            .I2(GND_net), .I3(GND_net), .O(n907_adj_4622));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i610_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i659_2_lut (.I0(\Ki[13] ), .I1(\PID_CONTROLLER.integral_23__N_3546 [10]), 
            .I2(GND_net), .I3(GND_net), .O(n980_adj_4621));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i659_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i73_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3546 [11]), 
            .I2(GND_net), .I3(GND_net), .O(n107_adj_4620));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i73_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i26_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3546 [12]), 
            .I2(GND_net), .I3(GND_net), .O(n38_adj_4619));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i26_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i122_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3546 [11]), 
            .I2(GND_net), .I3(GND_net), .O(n180_adj_4618));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i122_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i19132_2_lut (.I0(n28[4]), .I1(\PID_CONTROLLER.integral_23__N_3594 ), 
            .I2(GND_net), .I3(GND_net), .O(n3302[4]));   // verilog/motorControl.v(31[7] 33[10])
    defparam i19132_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i171_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3546 [11]), 
            .I2(GND_net), .I3(GND_net), .O(n253_adj_4617));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i171_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i19133_2_lut (.I0(n28[5]), .I1(\PID_CONTROLLER.integral_23__N_3594 ), 
            .I2(GND_net), .I3(GND_net), .O(n3302[5]));   // verilog/motorControl.v(31[7] 33[10])
    defparam i19133_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i30880_1_lut (.I0(duty[23]), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n37633));   // verilog/motorControl.v(29[14] 48[8])
    defparam i30880_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i22575_3_lut_4_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3546 [20]), 
            .I2(n27680), .I3(n10334[0]), .O(n4_adj_4722));   // verilog/motorControl.v(34[25:36])
    defparam i22575_3_lut_4_lut.LUT_INIT = 16'hf880;
    SB_LUT4 i2_3_lut_4_lut_adj_1490 (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3546 [20]), 
            .I2(n10334[0]), .I3(n27680), .O(n10329[1]));   // verilog/motorControl.v(34[25:36])
    defparam i2_3_lut_4_lut_adj_1490.LUT_INIT = 16'h8778;
    SB_LUT4 mult_11_i220_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3546 [11]), 
            .I2(GND_net), .I3(GND_net), .O(n326_adj_4615));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i220_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i22564_2_lut_3_lut_4_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3546 [21]), 
            .I2(\PID_CONTROLLER.integral_23__N_3546 [20]), .I3(\Ki[1] ), 
            .O(n27680));   // verilog/motorControl.v(34[25:36])
    defparam i22564_2_lut_3_lut_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 mult_11_i269_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3546 [11]), 
            .I2(GND_net), .I3(GND_net), .O(n399_adj_4614));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i269_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i22562_2_lut_3_lut_4_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3546 [21]), 
            .I2(\PID_CONTROLLER.integral_23__N_3546 [20]), .I3(\Ki[1] ), 
            .O(n10329[0]));   // verilog/motorControl.v(34[25:36])
    defparam i22562_2_lut_3_lut_4_lut.LUT_INIT = 16'h7888;
    SB_LUT4 i19134_2_lut (.I0(n28[6]), .I1(\PID_CONTROLLER.integral_23__N_3594 ), 
            .I2(GND_net), .I3(GND_net), .O(n3302[6]));   // verilog/motorControl.v(31[7] 33[10])
    defparam i19134_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i318_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3546 [11]), 
            .I2(GND_net), .I3(GND_net), .O(n472_adj_4612));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i318_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i367_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3546 [11]), 
            .I2(GND_net), .I3(GND_net), .O(n545_adj_4611));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i367_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5248_8_lut (.I0(GND_net), .I1(n9837[5]), .I2(n524_adj_4723), 
            .I3(n28955), .O(n9816[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5248_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5248_8 (.CI(n28955), .I0(n9837[5]), .I1(n524_adj_4723), 
            .CO(n28956));
    SB_LUT4 add_5248_7_lut (.I0(GND_net), .I1(n9837[4]), .I2(n451_adj_4724), 
            .I3(n28954), .O(n9816[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5248_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i416_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3546 [11]), 
            .I2(GND_net), .I3(GND_net), .O(n618_adj_4609));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i416_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i22544_3_lut_4_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3546 [19]), 
            .I2(n27646), .I3(n10329[0]), .O(n4_adj_4725));   // verilog/motorControl.v(34[25:36])
    defparam i22544_3_lut_4_lut.LUT_INIT = 16'hf880;
    SB_LUT4 mult_11_i465_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral_23__N_3546 [11]), 
            .I2(GND_net), .I3(GND_net), .O(n691_adj_4608));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i465_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i514_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral_23__N_3546 [11]), 
            .I2(GND_net), .I3(GND_net), .O(n764_adj_4607));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i514_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i563_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral_23__N_3546 [11]), 
            .I2(GND_net), .I3(GND_net), .O(n837_adj_4606));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i563_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i2_3_lut_4_lut_adj_1491 (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3546 [19]), 
            .I2(n10329[0]), .I3(n27646), .O(n10323[1]));   // verilog/motorControl.v(34[25:36])
    defparam i2_3_lut_4_lut_adj_1491.LUT_INIT = 16'h8778;
    SB_CARRY add_5248_7 (.CI(n28954), .I0(n9837[4]), .I1(n451_adj_4724), 
            .CO(n28955));
    SB_LUT4 mult_11_i612_2_lut (.I0(\Ki[12] ), .I1(\PID_CONTROLLER.integral_23__N_3546 [11]), 
            .I2(GND_net), .I3(GND_net), .O(n910_adj_4605));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i612_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i75_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3546 [12]), 
            .I2(GND_net), .I3(GND_net), .O(n110_adj_4604));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i75_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5248_6_lut (.I0(GND_net), .I1(n9837[3]), .I2(n378_adj_4726), 
            .I3(n28953), .O(n9816[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5248_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i28_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3546 [13]), 
            .I2(GND_net), .I3(GND_net), .O(n41_adj_4603));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i28_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i22531_2_lut_3_lut_4_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3546 [20]), 
            .I2(\PID_CONTROLLER.integral_23__N_3546 [19]), .I3(\Ki[1] ), 
            .O(n10323[0]));   // verilog/motorControl.v(34[25:36])
    defparam i22531_2_lut_3_lut_4_lut.LUT_INIT = 16'h7888;
    SB_LUT4 i22533_2_lut_3_lut_4_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3546 [20]), 
            .I2(\PID_CONTROLLER.integral_23__N_3546 [19]), .I3(\Ki[1] ), 
            .O(n27646));   // verilog/motorControl.v(34[25:36])
    defparam i22533_2_lut_3_lut_4_lut.LUT_INIT = 16'h8000;
    SB_CARRY add_5248_6 (.CI(n28953), .I0(n9837[3]), .I1(n378_adj_4726), 
            .CO(n28954));
    SB_LUT4 i22513_3_lut_4_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3546 [18]), 
            .I2(n4_adj_4727), .I3(n10323[1]), .O(n6_adj_4728));   // verilog/motorControl.v(34[25:36])
    defparam i22513_3_lut_4_lut.LUT_INIT = 16'hf880;
    SB_LUT4 mult_11_i124_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3546 [12]), 
            .I2(GND_net), .I3(GND_net), .O(n183_adj_4602));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i124_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i173_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3546 [12]), 
            .I2(GND_net), .I3(GND_net), .O(n256_adj_4601));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i173_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i222_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3546 [12]), 
            .I2(GND_net), .I3(GND_net), .O(n329_adj_4600));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i222_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5248_5_lut (.I0(GND_net), .I1(n9837[2]), .I2(n305_adj_4721), 
            .I3(n28952), .O(n9816[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5248_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i271_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3546 [12]), 
            .I2(GND_net), .I3(GND_net), .O(n402_adj_4599));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i271_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i2_3_lut_4_lut_adj_1492 (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3546 [18]), 
            .I2(n10323[1]), .I3(n4_adj_4727), .O(n10316[2]));   // verilog/motorControl.v(34[25:36])
    defparam i2_3_lut_4_lut_adj_1492.LUT_INIT = 16'h8778;
    SB_LUT4 mult_11_i320_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3546 [12]), 
            .I2(GND_net), .I3(GND_net), .O(n475_adj_4598));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i320_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i2_3_lut_4_lut_adj_1493 (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3546 [18]), 
            .I2(n10323[0]), .I3(n27603), .O(n10316[1]));   // verilog/motorControl.v(34[25:36])
    defparam i2_3_lut_4_lut_adj_1493.LUT_INIT = 16'h8778;
    SB_LUT4 unary_minus_5_inv_0_i23_1_lut (.I0(IntegralLimit[22]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[22]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i23_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_11_i369_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3546 [12]), 
            .I2(GND_net), .I3(GND_net), .O(n548_adj_4597));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i369_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i418_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3546 [12]), 
            .I2(GND_net), .I3(GND_net), .O(n621_adj_4596));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i418_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i467_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral_23__N_3546 [12]), 
            .I2(GND_net), .I3(GND_net), .O(n694_adj_4595));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i467_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i516_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral_23__N_3546 [12]), 
            .I2(GND_net), .I3(GND_net), .O(n767_adj_4594));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i516_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i565_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral_23__N_3546 [12]), 
            .I2(GND_net), .I3(GND_net), .O(n840_adj_4593));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i565_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i22505_3_lut_4_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3546 [18]), 
            .I2(n27603), .I3(n10323[0]), .O(n4_adj_4727));   // verilog/motorControl.v(34[25:36])
    defparam i22505_3_lut_4_lut.LUT_INIT = 16'hf880;
    SB_LUT4 i22494_2_lut_3_lut_4_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3546 [19]), 
            .I2(\PID_CONTROLLER.integral_23__N_3546 [18]), .I3(\Ki[1] ), 
            .O(n27603));   // verilog/motorControl.v(34[25:36])
    defparam i22494_2_lut_3_lut_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 unary_minus_16_add_3_25_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4735[23]), 
            .I3(n28049), .O(n257[23])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i77_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3546 [13]), 
            .I2(GND_net), .I3(GND_net), .O(n113_adj_4592));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i77_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i30_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3546 [14]), 
            .I2(GND_net), .I3(GND_net), .O(n44_adj_4591));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i30_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i126_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3546 [13]), 
            .I2(GND_net), .I3(GND_net), .O(n186_adj_4589));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i126_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_16_add_3_24_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4735[22]), 
            .I3(n28048), .O(n257[22])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5248_5 (.CI(n28952), .I0(n9837[2]), .I1(n305_adj_4721), 
            .CO(n28953));
    SB_CARRY unary_minus_16_add_3_24 (.CI(n28048), .I0(GND_net), .I1(n1_adj_4735[22]), 
            .CO(n28049));
    SB_LUT4 mult_11_i175_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3546 [13]), 
            .I2(GND_net), .I3(GND_net), .O(n259_adj_4588));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i175_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i22492_2_lut_3_lut_4_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3546 [19]), 
            .I2(\PID_CONTROLLER.integral_23__N_3546 [18]), .I3(\Ki[1] ), 
            .O(n10316[0]));   // verilog/motorControl.v(34[25:36])
    defparam i22492_2_lut_3_lut_4_lut.LUT_INIT = 16'h7888;
    SB_LUT4 mult_11_i224_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3546 [13]), 
            .I2(GND_net), .I3(GND_net), .O(n332_adj_4587));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i224_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_16_add_3_23_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4735[21]), 
            .I3(n28047), .O(n257[21])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i273_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3546 [13]), 
            .I2(GND_net), .I3(GND_net), .O(n405_adj_4586));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i273_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5248_4_lut (.I0(GND_net), .I1(n9837[1]), .I2(n232_adj_4717), 
            .I3(n28951), .O(n9816[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5248_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i322_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3546 [13]), 
            .I2(GND_net), .I3(GND_net), .O(n478_adj_4585));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i322_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i371_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3546 [13]), 
            .I2(GND_net), .I3(GND_net), .O(n551_adj_4584));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i371_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i420_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3546 [13]), 
            .I2(GND_net), .I3(GND_net), .O(n624_adj_4582));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i420_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i469_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral_23__N_3546 [13]), 
            .I2(GND_net), .I3(GND_net), .O(n697_adj_4581));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i469_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY unary_minus_16_add_3_23 (.CI(n28047), .I0(GND_net), .I1(n1_adj_4735[21]), 
            .CO(n28048));
    SB_CARRY add_5248_4 (.CI(n28951), .I0(n9837[1]), .I1(n232_adj_4717), 
            .CO(n28952));
    SB_LUT4 unary_minus_16_add_3_22_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4735[20]), 
            .I3(n28046), .O(n257[20])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_22 (.CI(n28046), .I0(GND_net), .I1(n1_adj_4735[20]), 
            .CO(n28047));
    SB_LUT4 unary_minus_16_add_3_21_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4735[19]), 
            .I3(n28045), .O(n257[19])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i255_2_lut (.I0(\Kp[5] ), .I1(n28[4]), .I2(GND_net), 
            .I3(GND_net), .O(n378_adj_4726));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i255_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i29618_2_lut_4_lut (.I0(duty_23__N_3646[21]), .I1(n257[21]), 
            .I2(duty_23__N_3646[9]), .I3(n257[9]), .O(n36373));
    defparam i29618_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 i29630_2_lut_4_lut (.I0(duty_23__N_3646[16]), .I1(n257[16]), 
            .I2(duty_23__N_3646[7]), .I3(n257[7]), .O(n36385));
    defparam i29630_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_CARRY unary_minus_16_add_3_21 (.CI(n28045), .I0(GND_net), .I1(n1_adj_4735[19]), 
            .CO(n28046));
    SB_LUT4 i29655_2_lut_4_lut (.I0(PWMLimit[21]), .I1(duty_23__N_3646[21]), 
            .I2(PWMLimit[9]), .I3(duty_23__N_3646[9]), .O(n36410));
    defparam i29655_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 unary_minus_16_add_3_20_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4735[18]), 
            .I3(n28044), .O(n257[18])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_20 (.CI(n28044), .I0(GND_net), .I1(n1_adj_4735[18]), 
            .CO(n28045));
    SB_LUT4 i29665_2_lut_4_lut (.I0(PWMLimit[16]), .I1(duty_23__N_3646[16]), 
            .I2(PWMLimit[7]), .I3(duty_23__N_3646[7]), .O(n36420));
    defparam i29665_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 mult_11_i518_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral_23__N_3546 [13]), 
            .I2(GND_net), .I3(GND_net), .O(n770_adj_4580));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i518_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5248_3_lut (.I0(GND_net), .I1(n9837[0]), .I2(n159_adj_4703), 
            .I3(n28950), .O(n9816[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5248_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i19135_2_lut (.I0(n28[7]), .I1(\PID_CONTROLLER.integral_23__N_3594 ), 
            .I2(GND_net), .I3(GND_net), .O(n3302[7]));   // verilog/motorControl.v(31[7] 33[10])
    defparam i19135_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i79_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3546 [14]), 
            .I2(GND_net), .I3(GND_net), .O(n116_adj_4577));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i79_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i32_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3546 [15]), 
            .I2(GND_net), .I3(GND_net), .O(n47_adj_4576));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i32_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5248_3 (.CI(n28950), .I0(n9837[0]), .I1(n159_adj_4703), 
            .CO(n28951));
    SB_LUT4 unary_minus_16_add_3_19_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4735[17]), 
            .I3(n28043), .O(n257[17])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5248_2_lut (.I0(GND_net), .I1(n17_adj_4701), .I2(n86_adj_4700), 
            .I3(GND_net), .O(n9816[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5248_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5248_2 (.CI(GND_net), .I0(n17_adj_4701), .I1(n86_adj_4700), 
            .CO(n28950));
    SB_LUT4 add_5247_21_lut (.I0(GND_net), .I1(n9816[18]), .I2(GND_net), 
            .I3(n28949), .O(n9794[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5247_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5247_20_lut (.I0(GND_net), .I1(n9816[17]), .I2(GND_net), 
            .I3(n28948), .O(n9794[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5247_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_19 (.CI(n28043), .I0(GND_net), .I1(n1_adj_4735[17]), 
            .CO(n28044));
    SB_CARRY add_5247_20 (.CI(n28948), .I0(n9816[17]), .I1(GND_net), .CO(n28949));
    SB_LUT4 add_5247_19_lut (.I0(GND_net), .I1(n9816[16]), .I2(GND_net), 
            .I3(n28947), .O(n9794[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5247_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5247_19 (.CI(n28947), .I0(n9816[16]), .I1(GND_net), .CO(n28948));
    SB_LUT4 add_5247_18_lut (.I0(GND_net), .I1(n9816[15]), .I2(GND_net), 
            .I3(n28946), .O(n9794[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5247_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5247_18 (.CI(n28946), .I0(n9816[15]), .I1(GND_net), .CO(n28947));
    SB_LUT4 add_5247_17_lut (.I0(GND_net), .I1(n9816[14]), .I2(GND_net), 
            .I3(n28945), .O(n9794[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5247_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5247_17 (.CI(n28945), .I0(n9816[14]), .I1(GND_net), .CO(n28946));
    SB_LUT4 add_5247_16_lut (.I0(GND_net), .I1(n9816[13]), .I2(n1105_adj_4699), 
            .I3(n28944), .O(n9794[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5247_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5247_16 (.CI(n28944), .I0(n9816[13]), .I1(n1105_adj_4699), 
            .CO(n28945));
    SB_LUT4 add_5247_15_lut (.I0(GND_net), .I1(n9816[12]), .I2(n1032_adj_4698), 
            .I3(n28943), .O(n9794[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5247_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5247_15 (.CI(n28943), .I0(n9816[12]), .I1(n1032_adj_4698), 
            .CO(n28944));
    SB_LUT4 unary_minus_16_add_3_18_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4735[16]), 
            .I3(n28042), .O(n257[16])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5247_14_lut (.I0(GND_net), .I1(n9816[11]), .I2(n959_adj_4696), 
            .I3(n28942), .O(n9794[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5247_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5247_14 (.CI(n28942), .I0(n9816[11]), .I1(n959_adj_4696), 
            .CO(n28943));
    SB_LUT4 add_5247_13_lut (.I0(GND_net), .I1(n9816[10]), .I2(n886_adj_4695), 
            .I3(n28941), .O(n9794[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5247_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_18 (.CI(n28042), .I0(GND_net), .I1(n1_adj_4735[16]), 
            .CO(n28043));
    SB_LUT4 unary_minus_16_add_3_17_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4735[15]), 
            .I3(n28041), .O(n257[15])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5247_13 (.CI(n28941), .I0(n9816[10]), .I1(n886_adj_4695), 
            .CO(n28942));
    SB_LUT4 add_5247_12_lut (.I0(GND_net), .I1(n9816[9]), .I2(n813_adj_4693), 
            .I3(n28940), .O(n9794[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5247_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5247_12 (.CI(n28940), .I0(n9816[9]), .I1(n813_adj_4693), 
            .CO(n28941));
    SB_LUT4 add_5247_11_lut (.I0(GND_net), .I1(n9816[8]), .I2(n740_adj_4692), 
            .I3(n28939), .O(n9794[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5247_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5247_11 (.CI(n28939), .I0(n9816[8]), .I1(n740_adj_4692), 
            .CO(n28940));
    SB_LUT4 add_5247_10_lut (.I0(GND_net), .I1(n9816[7]), .I2(n667_adj_4691), 
            .I3(n28938), .O(n9794[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5247_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5247_10 (.CI(n28938), .I0(n9816[7]), .I1(n667_adj_4691), 
            .CO(n28939));
    SB_LUT4 add_5247_9_lut (.I0(GND_net), .I1(n9816[6]), .I2(n594_adj_4690), 
            .I3(n28937), .O(n9794[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5247_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5247_9 (.CI(n28937), .I0(n9816[6]), .I1(n594_adj_4690), 
            .CO(n28938));
    SB_LUT4 add_5247_8_lut (.I0(GND_net), .I1(n9816[5]), .I2(n521_adj_4689), 
            .I3(n28936), .O(n9794[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5247_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5247_8 (.CI(n28936), .I0(n9816[5]), .I1(n521_adj_4689), 
            .CO(n28937));
    SB_LUT4 add_5247_7_lut (.I0(GND_net), .I1(n9816[4]), .I2(n448_adj_4688), 
            .I3(n28935), .O(n9794[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5247_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5247_7 (.CI(n28935), .I0(n9816[4]), .I1(n448_adj_4688), 
            .CO(n28936));
    SB_LUT4 add_5247_6_lut (.I0(GND_net), .I1(n9816[3]), .I2(n375_adj_4685), 
            .I3(n28934), .O(n9794[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5247_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5247_6 (.CI(n28934), .I0(n9816[3]), .I1(n375_adj_4685), 
            .CO(n28935));
    SB_CARRY unary_minus_16_add_3_17 (.CI(n28041), .I0(GND_net), .I1(n1_adj_4735[15]), 
            .CO(n28042));
    SB_LUT4 add_5247_5_lut (.I0(GND_net), .I1(n9816[2]), .I2(n302_adj_4684), 
            .I3(n28933), .O(n9794[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5247_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5247_5 (.CI(n28933), .I0(n9816[2]), .I1(n302_adj_4684), 
            .CO(n28934));
    SB_LUT4 unary_minus_16_add_3_16_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4735[14]), 
            .I3(n28040), .O(n257[14])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5247_4_lut (.I0(GND_net), .I1(n9816[1]), .I2(n229_adj_4682), 
            .I3(n28932), .O(n9794[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5247_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5247_4 (.CI(n28932), .I0(n9816[1]), .I1(n229_adj_4682), 
            .CO(n28933));
    SB_LUT4 add_5247_3_lut (.I0(GND_net), .I1(n9816[0]), .I2(n156_adj_4681), 
            .I3(n28931), .O(n9794[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5247_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5247_3 (.CI(n28931), .I0(n9816[0]), .I1(n156_adj_4681), 
            .CO(n28932));
    SB_LUT4 add_5247_2_lut (.I0(GND_net), .I1(n14_adj_4680), .I2(n83_adj_4679), 
            .I3(GND_net), .O(n9794[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5247_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5247_2 (.CI(GND_net), .I0(n14_adj_4680), .I1(n83_adj_4679), 
            .CO(n28931));
    SB_LUT4 add_5246_22_lut (.I0(GND_net), .I1(n9794[19]), .I2(GND_net), 
            .I3(n28930), .O(n9771[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5246_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5246_21_lut (.I0(GND_net), .I1(n9794[18]), .I2(GND_net), 
            .I3(n28929), .O(n9771[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5246_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5246_21 (.CI(n28929), .I0(n9794[18]), .I1(GND_net), .CO(n28930));
    SB_LUT4 add_5246_20_lut (.I0(GND_net), .I1(n9794[17]), .I2(GND_net), 
            .I3(n28928), .O(n9771[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5246_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5246_20 (.CI(n28928), .I0(n9794[17]), .I1(GND_net), .CO(n28929));
    SB_LUT4 add_5246_19_lut (.I0(GND_net), .I1(n9794[16]), .I2(GND_net), 
            .I3(n28927), .O(n9771[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5246_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5246_19 (.CI(n28927), .I0(n9794[16]), .I1(GND_net), .CO(n28928));
    SB_LUT4 add_5246_18_lut (.I0(GND_net), .I1(n9794[15]), .I2(GND_net), 
            .I3(n28926), .O(n9771[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5246_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5246_18 (.CI(n28926), .I0(n9794[15]), .I1(GND_net), .CO(n28927));
    SB_LUT4 add_5246_17_lut (.I0(GND_net), .I1(n9794[14]), .I2(GND_net), 
            .I3(n28925), .O(n9771[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5246_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5246_17 (.CI(n28925), .I0(n9794[14]), .I1(GND_net), .CO(n28926));
    SB_LUT4 add_5246_16_lut (.I0(GND_net), .I1(n9794[13]), .I2(n1102_adj_4613), 
            .I3(n28924), .O(n9771[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5246_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5246_16 (.CI(n28924), .I0(n9794[13]), .I1(n1102_adj_4613), 
            .CO(n28925));
    SB_LUT4 add_5246_15_lut (.I0(GND_net), .I1(n9794[12]), .I2(n1029_adj_4610), 
            .I3(n28923), .O(n9771[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5246_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5246_15 (.CI(n28923), .I0(n9794[12]), .I1(n1029_adj_4610), 
            .CO(n28924));
    SB_LUT4 add_5246_14_lut (.I0(GND_net), .I1(n9794[11]), .I2(n956_adj_4590), 
            .I3(n28922), .O(n9771[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5246_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5246_14 (.CI(n28922), .I0(n9794[11]), .I1(n956_adj_4590), 
            .CO(n28923));
    SB_LUT4 add_5246_13_lut (.I0(GND_net), .I1(n9794[10]), .I2(n883_adj_4583), 
            .I3(n28921), .O(n9771[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5246_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5246_13 (.CI(n28921), .I0(n9794[10]), .I1(n883_adj_4583), 
            .CO(n28922));
    SB_LUT4 add_5246_12_lut (.I0(GND_net), .I1(n9794[9]), .I2(n810_adj_4579), 
            .I3(n28920), .O(n9771[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5246_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5246_12 (.CI(n28920), .I0(n9794[9]), .I1(n810_adj_4579), 
            .CO(n28921));
    SB_LUT4 add_5246_11_lut (.I0(GND_net), .I1(n9794[8]), .I2(n737_adj_4578), 
            .I3(n28919), .O(n9771[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5246_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5246_11 (.CI(n28919), .I0(n9794[8]), .I1(n737_adj_4578), 
            .CO(n28920));
    SB_LUT4 add_5246_10_lut (.I0(GND_net), .I1(n9794[7]), .I2(n664_adj_4575), 
            .I3(n28918), .O(n9771[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5246_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5246_10 (.CI(n28918), .I0(n9794[7]), .I1(n664_adj_4575), 
            .CO(n28919));
    SB_LUT4 add_5246_9_lut (.I0(GND_net), .I1(n9794[6]), .I2(n591_adj_4574), 
            .I3(n28917), .O(n9771[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5246_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5246_9 (.CI(n28917), .I0(n9794[6]), .I1(n591_adj_4574), 
            .CO(n28918));
    SB_LUT4 add_5246_8_lut (.I0(GND_net), .I1(n9794[5]), .I2(n518_adj_4573), 
            .I3(n28916), .O(n9771[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5246_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5246_8 (.CI(n28916), .I0(n9794[5]), .I1(n518_adj_4573), 
            .CO(n28917));
    SB_LUT4 add_5246_7_lut (.I0(GND_net), .I1(n9794[4]), .I2(n445_adj_4571), 
            .I3(n28915), .O(n9771[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5246_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5246_7 (.CI(n28915), .I0(n9794[4]), .I1(n445_adj_4571), 
            .CO(n28916));
    SB_LUT4 add_5246_6_lut (.I0(GND_net), .I1(n9794[3]), .I2(n372_adj_4570), 
            .I3(n28914), .O(n9771[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5246_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5246_6 (.CI(n28914), .I0(n9794[3]), .I1(n372_adj_4570), 
            .CO(n28915));
    SB_LUT4 add_5246_5_lut (.I0(GND_net), .I1(n9794[2]), .I2(n299_adj_4567), 
            .I3(n28913), .O(n9771[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5246_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5246_5 (.CI(n28913), .I0(n9794[2]), .I1(n299_adj_4567), 
            .CO(n28914));
    SB_CARRY unary_minus_16_add_3_16 (.CI(n28040), .I0(GND_net), .I1(n1_adj_4735[14]), 
            .CO(n28041));
    SB_LUT4 add_5246_4_lut (.I0(GND_net), .I1(n9794[1]), .I2(n226_adj_4565), 
            .I3(n28912), .O(n9771[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5246_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5246_4 (.CI(n28912), .I0(n9794[1]), .I1(n226_adj_4565), 
            .CO(n28913));
    SB_LUT4 add_5246_3_lut (.I0(GND_net), .I1(n9794[0]), .I2(n153_adj_4555), 
            .I3(n28911), .O(n9771[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5246_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5246_3 (.CI(n28911), .I0(n9794[0]), .I1(n153_adj_4555), 
            .CO(n28912));
    SB_LUT4 add_5246_2_lut (.I0(GND_net), .I1(n11_adj_4535), .I2(n80_adj_4533), 
            .I3(GND_net), .O(n9771[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5246_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5246_2 (.CI(GND_net), .I0(n11_adj_4535), .I1(n80_adj_4533), 
            .CO(n28911));
    SB_LUT4 mult_10_add_1225_24_lut (.I0(n28[23]), .I1(n9747[21]), .I2(GND_net), 
            .I3(n28910), .O(n8175[0])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_24_lut.LUT_INIT = 16'h6996;
    SB_LUT4 mult_10_add_1225_23_lut (.I0(GND_net), .I1(n9747[20]), .I2(GND_net), 
            .I3(n28909), .O(n106[22])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_1225_23 (.CI(n28909), .I0(n9747[20]), .I1(GND_net), 
            .CO(n28910));
    SB_LUT4 mult_10_add_1225_22_lut (.I0(GND_net), .I1(n9747[19]), .I2(GND_net), 
            .I3(n28908), .O(n106[21])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_1225_22 (.CI(n28908), .I0(n9747[19]), .I1(GND_net), 
            .CO(n28909));
    SB_LUT4 mult_10_add_1225_21_lut (.I0(GND_net), .I1(n9747[18]), .I2(GND_net), 
            .I3(n28907), .O(n106[20])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_1225_21 (.CI(n28907), .I0(n9747[18]), .I1(GND_net), 
            .CO(n28908));
    SB_LUT4 mult_10_add_1225_20_lut (.I0(GND_net), .I1(n9747[17]), .I2(GND_net), 
            .I3(n28906), .O(n106[19])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_1225_20 (.CI(n28906), .I0(n9747[17]), .I1(GND_net), 
            .CO(n28907));
    SB_LUT4 mult_10_add_1225_19_lut (.I0(GND_net), .I1(n9747[16]), .I2(GND_net), 
            .I3(n28905), .O(n106[18])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_1225_19 (.CI(n28905), .I0(n9747[16]), .I1(GND_net), 
            .CO(n28906));
    SB_LUT4 mult_10_add_1225_18_lut (.I0(GND_net), .I1(n9747[15]), .I2(GND_net), 
            .I3(n28904), .O(n106[17])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_1225_18 (.CI(n28904), .I0(n9747[15]), .I1(GND_net), 
            .CO(n28905));
    SB_LUT4 unary_minus_16_add_3_15_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4735[13]), 
            .I3(n28039), .O(n257[13])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_add_1225_17_lut (.I0(GND_net), .I1(n9747[14]), .I2(GND_net), 
            .I3(n28903), .O(n106[16])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_1225_17 (.CI(n28903), .I0(n9747[14]), .I1(GND_net), 
            .CO(n28904));
    SB_LUT4 mult_10_add_1225_16_lut (.I0(GND_net), .I1(n9747[13]), .I2(n1096_adj_4518), 
            .I3(n28902), .O(n106[15])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_1225_16 (.CI(n28902), .I0(n9747[13]), .I1(n1096_adj_4518), 
            .CO(n28903));
    SB_LUT4 mult_10_add_1225_15_lut (.I0(GND_net), .I1(n9747[12]), .I2(n1023_adj_4513), 
            .I3(n28901), .O(n106[14])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_1225_15 (.CI(n28901), .I0(n9747[12]), .I1(n1023_adj_4513), 
            .CO(n28902));
    SB_LUT4 mult_10_add_1225_14_lut (.I0(GND_net), .I1(n9747[11]), .I2(n950_adj_4503), 
            .I3(n28900), .O(n106[13])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_1225_14 (.CI(n28900), .I0(n9747[11]), .I1(n950_adj_4503), 
            .CO(n28901));
    SB_LUT4 mult_10_add_1225_13_lut (.I0(GND_net), .I1(n9747[10]), .I2(n877_adj_4500), 
            .I3(n28899), .O(n106[12])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_1225_13 (.CI(n28899), .I0(n9747[10]), .I1(n877_adj_4500), 
            .CO(n28900));
    SB_LUT4 mult_10_add_1225_12_lut (.I0(GND_net), .I1(n9747[9]), .I2(n804_adj_4499), 
            .I3(n28898), .O(n106[11])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_1225_12 (.CI(n28898), .I0(n9747[9]), .I1(n804_adj_4499), 
            .CO(n28899));
    SB_LUT4 mult_10_add_1225_11_lut (.I0(GND_net), .I1(n9747[8]), .I2(n731_adj_4493), 
            .I3(n28897), .O(n106[10])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_1225_11 (.CI(n28897), .I0(n9747[8]), .I1(n731_adj_4493), 
            .CO(n28898));
    SB_LUT4 mult_10_add_1225_10_lut (.I0(GND_net), .I1(n9747[7]), .I2(n658_adj_4491), 
            .I3(n28896), .O(n106[9])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_1225_10 (.CI(n28896), .I0(n9747[7]), .I1(n658_adj_4491), 
            .CO(n28897));
    SB_LUT4 mult_10_add_1225_9_lut (.I0(GND_net), .I1(n9747[6]), .I2(n585_adj_4490), 
            .I3(n28895), .O(n106[8])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_1225_9 (.CI(n28895), .I0(n9747[6]), .I1(n585_adj_4490), 
            .CO(n28896));
    SB_LUT4 mult_10_add_1225_8_lut (.I0(GND_net), .I1(n9747[5]), .I2(n512_adj_4489), 
            .I3(n28894), .O(n106[7])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_1225_8 (.CI(n28894), .I0(n9747[5]), .I1(n512_adj_4489), 
            .CO(n28895));
    SB_LUT4 mult_10_add_1225_7_lut (.I0(GND_net), .I1(n9747[4]), .I2(n439_adj_4483), 
            .I3(n28893), .O(n106[6])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_1225_7 (.CI(n28893), .I0(n9747[4]), .I1(n439_adj_4483), 
            .CO(n28894));
    SB_LUT4 mult_10_add_1225_6_lut (.I0(GND_net), .I1(n9747[3]), .I2(n366_adj_4478), 
            .I3(n28892), .O(n106[5])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_1225_6 (.CI(n28892), .I0(n9747[3]), .I1(n366_adj_4478), 
            .CO(n28893));
    SB_LUT4 mult_10_add_1225_5_lut (.I0(GND_net), .I1(n9747[2]), .I2(n293_adj_4475), 
            .I3(n28891), .O(n106[4])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_1225_5 (.CI(n28891), .I0(n9747[2]), .I1(n293_adj_4475), 
            .CO(n28892));
    SB_LUT4 mult_10_add_1225_4_lut (.I0(GND_net), .I1(n9747[1]), .I2(n220_adj_4472), 
            .I3(n28890), .O(n106[3])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_1225_4 (.CI(n28890), .I0(n9747[1]), .I1(n220_adj_4472), 
            .CO(n28891));
    SB_LUT4 mult_10_add_1225_3_lut (.I0(GND_net), .I1(n9747[0]), .I2(n147_adj_4469), 
            .I3(n28889), .O(n106[2])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_1225_3 (.CI(n28889), .I0(n9747[0]), .I1(n147_adj_4469), 
            .CO(n28890));
    SB_LUT4 mult_10_add_1225_2_lut (.I0(GND_net), .I1(n5_adj_4460), .I2(n74_adj_4458), 
            .I3(GND_net), .O(n106[1])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_1225_2 (.CI(GND_net), .I0(n5_adj_4460), .I1(n74_adj_4458), 
            .CO(n28889));
    SB_LUT4 add_5245_23_lut (.I0(GND_net), .I1(n9771[20]), .I2(GND_net), 
            .I3(n28888), .O(n9747[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5245_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5245_22_lut (.I0(GND_net), .I1(n9771[19]), .I2(GND_net), 
            .I3(n28887), .O(n9747[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5245_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5245_22 (.CI(n28887), .I0(n9771[19]), .I1(GND_net), .CO(n28888));
    SB_LUT4 add_5245_21_lut (.I0(GND_net), .I1(n9771[18]), .I2(GND_net), 
            .I3(n28886), .O(n9747[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5245_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5245_21 (.CI(n28886), .I0(n9771[18]), .I1(GND_net), .CO(n28887));
    SB_LUT4 add_5245_20_lut (.I0(GND_net), .I1(n9771[17]), .I2(GND_net), 
            .I3(n28885), .O(n9747[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5245_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5245_20 (.CI(n28885), .I0(n9771[17]), .I1(GND_net), .CO(n28886));
    SB_LUT4 add_5245_19_lut (.I0(GND_net), .I1(n9771[16]), .I2(GND_net), 
            .I3(n28884), .O(n9747[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5245_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5245_19 (.CI(n28884), .I0(n9771[16]), .I1(GND_net), .CO(n28885));
    SB_LUT4 add_5245_18_lut (.I0(GND_net), .I1(n9771[15]), .I2(GND_net), 
            .I3(n28883), .O(n9747[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5245_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5245_18 (.CI(n28883), .I0(n9771[15]), .I1(GND_net), .CO(n28884));
    SB_LUT4 add_5245_17_lut (.I0(GND_net), .I1(n9771[14]), .I2(GND_net), 
            .I3(n28882), .O(n9747[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5245_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5245_17 (.CI(n28882), .I0(n9771[14]), .I1(GND_net), .CO(n28883));
    SB_LUT4 add_5245_16_lut (.I0(GND_net), .I1(n9771[13]), .I2(n1099_adj_4438), 
            .I3(n28881), .O(n9747[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5245_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5245_16 (.CI(n28881), .I0(n9771[13]), .I1(n1099_adj_4438), 
            .CO(n28882));
    SB_LUT4 add_5245_15_lut (.I0(GND_net), .I1(n9771[12]), .I2(n1026_adj_4433), 
            .I3(n28880), .O(n9747[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5245_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5245_15 (.CI(n28880), .I0(n9771[12]), .I1(n1026_adj_4433), 
            .CO(n28881));
    SB_LUT4 add_5245_14_lut (.I0(GND_net), .I1(n9771[11]), .I2(n953_adj_4426), 
            .I3(n28879), .O(n9747[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5245_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5245_14 (.CI(n28879), .I0(n9771[11]), .I1(n953_adj_4426), 
            .CO(n28880));
    SB_LUT4 add_5245_13_lut (.I0(GND_net), .I1(n9771[10]), .I2(n880_adj_4423), 
            .I3(n28878), .O(n9747[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5245_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5245_13 (.CI(n28878), .I0(n9771[10]), .I1(n880_adj_4423), 
            .CO(n28879));
    SB_LUT4 add_5245_12_lut (.I0(GND_net), .I1(n9771[9]), .I2(n807_adj_4417), 
            .I3(n28877), .O(n9747[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5245_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5245_12 (.CI(n28877), .I0(n9771[9]), .I1(n807_adj_4417), 
            .CO(n28878));
    SB_LUT4 add_5245_11_lut (.I0(GND_net), .I1(n9771[8]), .I2(n734_adj_4414), 
            .I3(n28876), .O(n9747[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5245_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5245_11 (.CI(n28876), .I0(n9771[8]), .I1(n734_adj_4414), 
            .CO(n28877));
    SB_LUT4 add_5245_10_lut (.I0(GND_net), .I1(n9771[7]), .I2(n661_adj_4413), 
            .I3(n28875), .O(n9747[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5245_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5245_10 (.CI(n28875), .I0(n9771[7]), .I1(n661_adj_4413), 
            .CO(n28876));
    SB_LUT4 add_5245_9_lut (.I0(GND_net), .I1(n9771[6]), .I2(n588_adj_4412), 
            .I3(n28874), .O(n9747[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5245_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5245_9 (.CI(n28874), .I0(n9771[6]), .I1(n588_adj_4412), 
            .CO(n28875));
    SB_LUT4 add_5245_8_lut (.I0(GND_net), .I1(n9771[5]), .I2(n515_adj_4411), 
            .I3(n28873), .O(n9747[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5245_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5245_8 (.CI(n28873), .I0(n9771[5]), .I1(n515_adj_4411), 
            .CO(n28874));
    SB_LUT4 add_5245_7_lut (.I0(GND_net), .I1(n9771[4]), .I2(n442_adj_4410), 
            .I3(n28872), .O(n9747[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5245_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5245_7 (.CI(n28872), .I0(n9771[4]), .I1(n442_adj_4410), 
            .CO(n28873));
    SB_LUT4 add_5245_6_lut (.I0(GND_net), .I1(n9771[3]), .I2(n369_adj_4409), 
            .I3(n28871), .O(n9747[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5245_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5245_6 (.CI(n28871), .I0(n9771[3]), .I1(n369_adj_4409), 
            .CO(n28872));
    SB_LUT4 add_5245_5_lut (.I0(GND_net), .I1(n9771[2]), .I2(n296_adj_4408), 
            .I3(n28870), .O(n9747[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5245_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_12_25_lut (.I0(GND_net), .I1(n8175[0]), .I2(n8179[0]), 
            .I3(n27877), .O(duty_23__N_3646[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5245_5 (.CI(n28870), .I0(n9771[2]), .I1(n296_adj_4408), 
            .CO(n28871));
    SB_LUT4 add_5245_4_lut (.I0(GND_net), .I1(n9771[1]), .I2(n223_adj_4407), 
            .I3(n28869), .O(n9747[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5245_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i304_2_lut (.I0(\Kp[6] ), .I1(n28[4]), .I2(GND_net), 
            .I3(GND_net), .O(n451_adj_4724));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i304_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY unary_minus_16_add_3_15 (.CI(n28039), .I0(GND_net), .I1(n1_adj_4735[13]), 
            .CO(n28040));
    SB_CARRY add_5245_4 (.CI(n28869), .I0(n9771[1]), .I1(n223_adj_4407), 
            .CO(n28870));
    SB_LUT4 unary_minus_16_add_3_14_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4735[12]), 
            .I3(n28038), .O(n257[12])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i19136_2_lut (.I0(n28[8]), .I1(\PID_CONTROLLER.integral_23__N_3594 ), 
            .I2(GND_net), .I3(GND_net), .O(n3302[8]));   // verilog/motorControl.v(31[7] 33[10])
    defparam i19136_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5245_3_lut (.I0(GND_net), .I1(n9771[0]), .I2(n150_adj_4405), 
            .I3(n28868), .O(n9747[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5245_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5245_3 (.CI(n28868), .I0(n9771[0]), .I1(n150_adj_4405), 
            .CO(n28869));
    SB_LUT4 add_5245_2_lut (.I0(GND_net), .I1(n8_adj_4404), .I2(n77_adj_4402), 
            .I3(GND_net), .O(n9747[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5245_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5245_2 (.CI(GND_net), .I0(n8_adj_4404), .I1(n77_adj_4402), 
            .CO(n28868));
    SB_CARRY unary_minus_16_add_3_14 (.CI(n28038), .I0(GND_net), .I1(n1_adj_4735[12]), 
            .CO(n28039));
    SB_LUT4 unary_minus_16_add_3_13_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4735[11]), 
            .I3(n28037), .O(n257[11])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_12_24_lut (.I0(GND_net), .I1(n106[22]), .I2(n155[22]), 
            .I3(n27876), .O(duty_23__N_3646[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_13 (.CI(n28037), .I0(GND_net), .I1(n1_adj_4735[11]), 
            .CO(n28038));
    SB_LUT4 unary_minus_16_add_3_12_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4735[10]), 
            .I3(n28036), .O(n257[10])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_12 (.CI(n28036), .I0(GND_net), .I1(n1_adj_4735[10]), 
            .CO(n28037));
    SB_LUT4 unary_minus_16_add_3_11_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4735[9]), 
            .I3(n28035), .O(n257[9])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_11 (.CI(n28035), .I0(GND_net), .I1(n1_adj_4735[9]), 
            .CO(n28036));
    SB_LUT4 unary_minus_16_add_3_10_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4735[8]), 
            .I3(n28034), .O(n257[8])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_12_24 (.CI(n27876), .I0(n106[22]), .I1(n155[22]), .CO(n27877));
    SB_LUT4 mult_10_i353_2_lut (.I0(\Kp[7] ), .I1(n28[4]), .I2(GND_net), 
            .I3(GND_net), .O(n524_adj_4723));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i353_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY unary_minus_16_add_3_10 (.CI(n28034), .I0(GND_net), .I1(n1_adj_4735[8]), 
            .CO(n28035));
    SB_LUT4 add_12_23_lut (.I0(GND_net), .I1(n106[21]), .I2(n155[21]), 
            .I3(n27875), .O(duty_23__N_3646[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_16_add_3_9_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4735[7]), 
            .I3(n28033), .O(n257[7])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_9 (.CI(n28033), .I0(GND_net), .I1(n1_adj_4735[7]), 
            .CO(n28034));
    SB_LUT4 unary_minus_16_add_3_8_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4735[6]), 
            .I3(n28032), .O(n257[6])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i128_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3546 [14]), 
            .I2(GND_net), .I3(GND_net), .O(n189_adj_4572));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i128_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i177_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3546 [14]), 
            .I2(GND_net), .I3(GND_net), .O(n262_adj_4569));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i177_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_12_23 (.CI(n27875), .I0(n106[21]), .I1(n155[21]), .CO(n27876));
    SB_CARRY unary_minus_16_add_3_8 (.CI(n28032), .I0(GND_net), .I1(n1_adj_4735[6]), 
            .CO(n28033));
    SB_LUT4 add_12_22_lut (.I0(GND_net), .I1(n106[20]), .I2(n155[20]), 
            .I3(n27874), .O(duty_23__N_3646[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_16_add_3_7_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4735[5]), 
            .I3(n28031), .O(n257[5])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_12_22 (.CI(n27874), .I0(n106[20]), .I1(n155[20]), .CO(n27875));
    SB_LUT4 mult_11_i226_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3546 [14]), 
            .I2(GND_net), .I3(GND_net), .O(n335_adj_4568));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i226_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i275_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3546 [14]), 
            .I2(GND_net), .I3(GND_net), .O(n408_adj_4566));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i275_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY unary_minus_16_add_3_7 (.CI(n28031), .I0(GND_net), .I1(n1_adj_4735[5]), 
            .CO(n28032));
    SB_LUT4 unary_minus_16_add_3_6_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4735[4]), 
            .I3(n28030), .O(n257[4])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_12_21_lut (.I0(GND_net), .I1(n106[19]), .I2(n155[19]), 
            .I3(n27873), .O(duty_23__N_3646[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_12_21 (.CI(n27873), .I0(n106[19]), .I1(n155[19]), .CO(n27874));
    SB_LUT4 add_12_20_lut (.I0(GND_net), .I1(n106[18]), .I2(n155[18]), 
            .I3(n27872), .O(duty_23__N_3646[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_12_20 (.CI(n27872), .I0(n106[18]), .I1(n155[18]), .CO(n27873));
    SB_LUT4 add_12_19_lut (.I0(GND_net), .I1(n106[17]), .I2(n155[17]), 
            .I3(n27871), .O(duty_23__N_3646[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_12_19 (.CI(n27871), .I0(n106[17]), .I1(n155[17]), .CO(n27872));
    SB_CARRY unary_minus_16_add_3_6 (.CI(n28030), .I0(GND_net), .I1(n1_adj_4735[4]), 
            .CO(n28031));
    SB_LUT4 unary_minus_16_add_3_5_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4735[3]), 
            .I3(n28029), .O(n257[3])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_5 (.CI(n28029), .I0(GND_net), .I1(n1_adj_4735[3]), 
            .CO(n28030));
    SB_LUT4 mult_11_i324_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3546 [14]), 
            .I2(GND_net), .I3(GND_net), .O(n481_adj_4564));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i324_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_16_add_3_4_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4735[2]), 
            .I3(n28028), .O(n257[2])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_12_18_lut (.I0(GND_net), .I1(n106[16]), .I2(n155[16]), 
            .I3(n27870), .O(duty_23__N_3646[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_4 (.CI(n28028), .I0(GND_net), .I1(n1_adj_4735[2]), 
            .CO(n28029));
    SB_CARRY add_12_18 (.CI(n27870), .I0(n106[16]), .I1(n155[16]), .CO(n27871));
    SB_LUT4 mult_11_i373_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3546 [14]), 
            .I2(GND_net), .I3(GND_net), .O(n554_adj_4563));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i373_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i422_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3546 [14]), 
            .I2(GND_net), .I3(GND_net), .O(n627_adj_4562));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i422_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_12_17_lut (.I0(GND_net), .I1(n106[15]), .I2(n155[15]), 
            .I3(n27869), .O(duty_23__N_3646[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i19137_2_lut (.I0(n28[9]), .I1(\PID_CONTROLLER.integral_23__N_3594 ), 
            .I2(GND_net), .I3(GND_net), .O(n3302[9]));   // verilog/motorControl.v(31[7] 33[10])
    defparam i19137_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i471_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral_23__N_3546 [14]), 
            .I2(GND_net), .I3(GND_net), .O(n700_adj_4561));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i471_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_12_17 (.CI(n27869), .I0(n106[15]), .I1(n155[15]), .CO(n27870));
    SB_LUT4 mult_11_i81_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3546 [15]), 
            .I2(GND_net), .I3(GND_net), .O(n119_adj_4560));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i81_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i34_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3546 [16]), 
            .I2(GND_net), .I3(GND_net), .O(n50_adj_4559));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i34_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_16_add_3_3_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4735[1]), 
            .I3(n28027), .O(n257[1])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_3 (.CI(n28027), .I0(GND_net), .I1(n1_adj_4735[1]), 
            .CO(n28028));
    SB_LUT4 unary_minus_16_add_3_2_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4735[0]), 
            .I3(VCC_net), .O(n257[0])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_2 (.CI(VCC_net), .I0(GND_net), .I1(n1_adj_4735[0]), 
            .CO(n28027));
    SB_LUT4 unary_minus_5_add_3_25_lut (.I0(GND_net), .I1(GND_net), .I2(n1[23]), 
            .I3(n28026), .O(\PID_CONTROLLER.integral_23__N_3597 [23])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i130_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3546 [15]), 
            .I2(GND_net), .I3(GND_net), .O(n192_adj_4558));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i130_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i179_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3546 [15]), 
            .I2(GND_net), .I3(GND_net), .O(n265_adj_4557));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i179_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i19138_2_lut (.I0(n28[10]), .I1(\PID_CONTROLLER.integral_23__N_3594 ), 
            .I2(GND_net), .I3(GND_net), .O(n3302[10]));   // verilog/motorControl.v(31[7] 33[10])
    defparam i19138_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i228_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3546 [15]), 
            .I2(GND_net), .I3(GND_net), .O(n338_adj_4556));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i228_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i277_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3546 [15]), 
            .I2(GND_net), .I3(GND_net), .O(n411_adj_4554));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i277_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i326_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3546 [15]), 
            .I2(GND_net), .I3(GND_net), .O(n484_adj_4553));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i326_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i375_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3546 [15]), 
            .I2(GND_net), .I3(GND_net), .O(n557_adj_4552));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i375_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i424_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3546 [15]), 
            .I2(GND_net), .I3(GND_net), .O(n630_adj_4551));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i424_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i83_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3546 [16]), 
            .I2(GND_net), .I3(GND_net), .O(n122_adj_4550));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i83_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i36_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3546 [17]), 
            .I2(GND_net), .I3(GND_net), .O(n53_adj_4549));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i36_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i132_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3546 [16]), 
            .I2(GND_net), .I3(GND_net), .O(n195_adj_4548));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i132_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i181_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3546 [16]), 
            .I2(GND_net), .I3(GND_net), .O(n268_adj_4547));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i181_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i230_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3546 [16]), 
            .I2(GND_net), .I3(GND_net), .O(n341_adj_4546));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i230_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i279_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3546 [16]), 
            .I2(GND_net), .I3(GND_net), .O(n414_adj_4545));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i279_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i328_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3546 [16]), 
            .I2(GND_net), .I3(GND_net), .O(n487_adj_4544));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i328_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i377_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3546 [16]), 
            .I2(GND_net), .I3(GND_net), .O(n560_adj_4543));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i377_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i85_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3546 [17]), 
            .I2(GND_net), .I3(GND_net), .O(n125_adj_4542));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i85_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i38_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3546 [18]), 
            .I2(GND_net), .I3(GND_net), .O(n56_adj_4541));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i38_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i134_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3546 [17]), 
            .I2(GND_net), .I3(GND_net), .O(n198_adj_4540));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i134_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i183_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3546 [17]), 
            .I2(GND_net), .I3(GND_net), .O(n271_adj_4539));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i183_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i232_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3546 [17]), 
            .I2(GND_net), .I3(GND_net), .O(n344_adj_4538));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i232_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i281_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3546 [17]), 
            .I2(GND_net), .I3(GND_net), .O(n417_adj_4537));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i281_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i2_4_lut_adj_1494 (.I0(n6_adj_4728), .I1(\Ki[4] ), .I2(n10323[2]), 
            .I3(\PID_CONTROLLER.integral_23__N_3546 [18]), .O(n10316[3]));   // verilog/motorControl.v(34[25:36])
    defparam i2_4_lut_adj_1494.LUT_INIT = 16'h965a;
    SB_LUT4 IntegralLimit_23__I_0_i8_3_lut_3_lut (.I0(IntegralLimit[4]), .I1(IntegralLimit[8]), 
            .I2(\PID_CONTROLLER.integral [8]), .I3(GND_net), .O(n8_adj_4335));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i8_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i22585_4_lut (.I0(\Ki[0] ), .I1(\Ki[1] ), .I2(\PID_CONTROLLER.integral_23__N_3546 [22]), 
            .I3(\PID_CONTROLLER.integral_23__N_3546 [21]), .O(n10334[0]));   // verilog/motorControl.v(34[25:36])
    defparam i22585_4_lut.LUT_INIT = 16'h6ca0;
    SB_LUT4 i2_4_lut_adj_1495 (.I0(n4_adj_4725), .I1(\Ki[3] ), .I2(n10329[1]), 
            .I3(\PID_CONTROLLER.integral_23__N_3546 [19]), .O(n10323[2]));   // verilog/motorControl.v(34[25:36])
    defparam i2_4_lut_adj_1495.LUT_INIT = 16'h965a;
    SB_LUT4 mult_11_i330_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3546 [17]), 
            .I2(GND_net), .I3(GND_net), .O(n490_adj_4536));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i330_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i2_4_lut_adj_1496 (.I0(\Ki[0] ), .I1(\Ki[3] ), .I2(\PID_CONTROLLER.integral_23__N_3546 [23]), 
            .I3(\PID_CONTROLLER.integral_23__N_3546 [20]), .O(n12_adj_4729));   // verilog/motorControl.v(34[25:36])
    defparam i2_4_lut_adj_1496.LUT_INIT = 16'h9c50;
    SB_LUT4 i22521_4_lut (.I0(n10323[2]), .I1(\Ki[4] ), .I2(n6_adj_4728), 
            .I3(\PID_CONTROLLER.integral_23__N_3546 [18]), .O(n8_adj_4730));   // verilog/motorControl.v(34[25:36])
    defparam i22521_4_lut.LUT_INIT = 16'he8a0;
    SB_LUT4 i1_4_lut_adj_1497 (.I0(\Ki[4] ), .I1(\Ki[2] ), .I2(\PID_CONTROLLER.integral_23__N_3546 [19]), 
            .I3(\PID_CONTROLLER.integral_23__N_3546 [21]), .O(n11_adj_4731));   // verilog/motorControl.v(34[25:36])
    defparam i1_4_lut_adj_1497.LUT_INIT = 16'h6ca0;
    SB_LUT4 i22552_4_lut (.I0(n10329[1]), .I1(\Ki[3] ), .I2(n4_adj_4725), 
            .I3(\PID_CONTROLLER.integral_23__N_3546 [19]), .O(n6_adj_4732));   // verilog/motorControl.v(34[25:36])
    defparam i22552_4_lut.LUT_INIT = 16'he8a0;
    SB_LUT4 i22587_4_lut (.I0(\Ki[0] ), .I1(\Ki[1] ), .I2(\PID_CONTROLLER.integral_23__N_3546 [22]), 
            .I3(\PID_CONTROLLER.integral_23__N_3546 [21]), .O(n27705));   // verilog/motorControl.v(34[25:36])
    defparam i22587_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i8_4_lut_adj_1498 (.I0(n6_adj_4732), .I1(n11_adj_4731), .I2(n8_adj_4730), 
            .I3(n12_adj_4729), .O(n18_adj_4733));   // verilog/motorControl.v(34[25:36])
    defparam i8_4_lut_adj_1498.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1499 (.I0(\Ki[5] ), .I1(\Ki[1] ), .I2(\PID_CONTROLLER.integral_23__N_3546 [18]), 
            .I3(\PID_CONTROLLER.integral_23__N_3546 [22]), .O(n13_adj_4734));   // verilog/motorControl.v(34[25:36])
    defparam i3_4_lut_adj_1499.LUT_INIT = 16'h6ca0;
    SB_LUT4 i9_4_lut_adj_1500 (.I0(n13_adj_4734), .I1(n18_adj_4733), .I2(n27705), 
            .I3(n4_adj_4722), .O(n34185));   // verilog/motorControl.v(34[25:36])
    defparam i9_4_lut_adj_1500.LUT_INIT = 16'h6996;
    SB_LUT4 i29653_3_lut_4_lut (.I0(duty_23__N_3646[3]), .I1(n257[3]), .I2(n257[2]), 
            .I3(duty_23__N_3646[2]), .O(n36408));   // verilog/motorControl.v(38[19:35])
    defparam i29653_3_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 LessThan_15_i6_3_lut_3_lut (.I0(duty_23__N_3646[3]), .I1(n257[3]), 
            .I2(n257[2]), .I3(GND_net), .O(n6_adj_4674));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i6_3_lut_3_lut.LUT_INIT = 16'hd4d4;
    SB_LUT4 i29687_3_lut_4_lut (.I0(PWMLimit[3]), .I1(duty_23__N_3646[3]), 
            .I2(duty_23__N_3646[2]), .I3(PWMLimit[2]), .O(n36442));   // verilog/motorControl.v(36[10:25])
    defparam i29687_3_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 duty_23__I_831_i6_3_lut_3_lut (.I0(PWMLimit[3]), .I1(duty_23__N_3646[3]), 
            .I2(duty_23__N_3646[2]), .I3(GND_net), .O(n6_adj_4646));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_831_i6_3_lut_3_lut.LUT_INIT = 16'hd4d4;
    SB_LUT4 i19139_2_lut (.I0(n28[11]), .I1(\PID_CONTROLLER.integral_23__N_3594 ), 
            .I2(GND_net), .I3(GND_net), .O(n3302[11]));   // verilog/motorControl.v(31[7] 33[10])
    defparam i19139_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i19140_2_lut (.I0(n28[12]), .I1(\PID_CONTROLLER.integral_23__N_3594 ), 
            .I2(GND_net), .I3(GND_net), .O(n3302[12]));   // verilog/motorControl.v(31[7] 33[10])
    defparam i19140_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i19141_2_lut (.I0(n28[13]), .I1(\PID_CONTROLLER.integral_23__N_3594 ), 
            .I2(GND_net), .I3(GND_net), .O(n3302[13]));   // verilog/motorControl.v(31[7] 33[10])
    defparam i19141_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i19142_2_lut (.I0(n28[14]), .I1(\PID_CONTROLLER.integral_23__N_3594 ), 
            .I2(GND_net), .I3(GND_net), .O(n3302[14]));   // verilog/motorControl.v(31[7] 33[10])
    defparam i19142_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i19143_2_lut (.I0(n28[15]), .I1(\PID_CONTROLLER.integral_23__N_3594 ), 
            .I2(GND_net), .I3(GND_net), .O(n3302[15]));   // verilog/motorControl.v(31[7] 33[10])
    defparam i19143_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i19144_2_lut (.I0(n28[16]), .I1(\PID_CONTROLLER.integral_23__N_3594 ), 
            .I2(GND_net), .I3(GND_net), .O(n3302[16]));   // verilog/motorControl.v(31[7] 33[10])
    defparam i19144_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i19145_2_lut (.I0(n28[17]), .I1(\PID_CONTROLLER.integral_23__N_3594 ), 
            .I2(GND_net), .I3(GND_net), .O(n3302[17]));   // verilog/motorControl.v(31[7] 33[10])
    defparam i19145_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i19146_2_lut (.I0(n28[18]), .I1(\PID_CONTROLLER.integral_23__N_3594 ), 
            .I2(GND_net), .I3(GND_net), .O(n3302[18]));   // verilog/motorControl.v(31[7] 33[10])
    defparam i19146_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i402_2_lut (.I0(\Kp[8] ), .I1(n28[4]), .I2(GND_net), 
            .I3(GND_net), .O(n597_adj_4716));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i402_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i451_2_lut (.I0(\Kp[9] ), .I1(n28[4]), .I2(GND_net), 
            .I3(GND_net), .O(n670_adj_4715));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i451_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i500_2_lut (.I0(\Kp[10] ), .I1(n28[4]), .I2(GND_net), 
            .I3(GND_net), .O(n743_adj_4714));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i500_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i549_2_lut (.I0(\Kp[11] ), .I1(n28[4]), .I2(GND_net), 
            .I3(GND_net), .O(n816_adj_4713));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i549_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i598_2_lut (.I0(\Kp[12] ), .I1(n28[4]), .I2(GND_net), 
            .I3(GND_net), .O(n889_adj_4712));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i598_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i647_2_lut (.I0(\Kp[13] ), .I1(n28[4]), .I2(GND_net), 
            .I3(GND_net), .O(n962_adj_4711));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i647_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i696_2_lut (.I0(\Kp[14] ), .I1(n28[4]), .I2(GND_net), 
            .I3(GND_net), .O(n1035_adj_4710));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i696_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i745_2_lut (.I0(\Kp[15] ), .I1(n28[4]), .I2(GND_net), 
            .I3(GND_net), .O(n1108_adj_4709));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i745_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i61_2_lut (.I0(\Kp[1] ), .I1(n28[5]), .I2(GND_net), 
            .I3(GND_net), .O(n89_adj_4708));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i61_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i14_2_lut (.I0(\Kp[0] ), .I1(n28[6]), .I2(GND_net), 
            .I3(GND_net), .O(n20_adj_4707));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i14_2_lut.LUT_INIT = 16'h8888;
    
endmodule
//
// Verilog Description of module coms
//

module coms (n63, n771, n10417, GND_net, \data_out_frame[19] , \data_out_frame[23] , 
            \data_out_frame[24] , \data_out_frame[17] , n3303, n123, 
            \FRAME_MATCHER.state_31__N_2662[1] , clk32MHz, \data_out_frame[15] , 
            \data_out_frame[20] , \data_out_frame[13] , \data_in_frame[4] , 
            \data_in_frame[1] , \data_out_frame[18] , \data_out_frame[25] , 
            \data_out_frame[16] , \data_in_frame[3] , \data_out_frame[10] , 
            \data_out_frame[8] , \data_out_frame[6] , \data_out_frame[12] , 
            n33567, \data_out_frame[11] , \data_out_frame[5] , \data_out_frame[14] , 
            \data_out_frame[7] , \data_in_frame[13] , \data_in_frame[9] , 
            \data_out_frame[9] , \data_out_frame[4] , \data_in_frame[6] , 
            \data_in_frame[5] , \data_in_frame[8] , rx_data, \data_in_frame[12] , 
            \FRAME_MATCHER.state , \data_in_frame[2] , \FRAME_MATCHER.state[0] , 
            n63_adj_8, n2970, n14711, n39, \data_in[1] , \data_in[0] , 
            \data_in[3] , \data_in[2] , n4452, \data_in_frame[10] , 
            \data_in_frame[11] , rx_data_ready, setpoint, \state[2] , 
            \state[3] , n10, \data_in_frame[21] , n3, n7, ID, n17474, 
            n17552, n17476, n5592, tx_active, n19101, n19100, n19099, 
            n19098, n19097, n19096, n19095, n19094, n19093, control_mode, 
            n19092, n19091, n19090, n19089, n19088, n19087, n19086, 
            PWMLimit, n19085, n19084, n19083, n19082, n19081, n19080, 
            n19079, n19078, n19077, n19076, n19075, n19074, n19073, 
            n19072, n19071, n19070, n19069, n19068, n19067, n19066, 
            n19065, n19064, n38205, n38206, n32009, n19047, n19046, 
            n19044, neopxl_color, LED_c, n19043, \Ki[0] , n19042, 
            \Kp[0] , n19041, n32173, DE_c, n19581, IntegralLimit, 
            n19580, n19579, n19578, n19577, n19576, n19575, n19574, 
            n19573, n19572, n19571, n19570, n19569, n19568, n19567, 
            n19566, n19565, n19564, n19563, n19562, n19561, n19560, 
            n19559, n19520, n19519, n19518, n19517, n19516, n19515, 
            n19514, n19513, n19512, n19511, n19510, n19509, n19508, 
            n19507, n19506, n19505, n19504, n19503, n19502, n19501, 
            n19500, n19499, n19498, n19497, n19496, n19495, n19494, 
            n19493, n19492, n19491, n19490, n19489, \Kp[1] , n19488, 
            \Kp[2] , n19487, \Kp[3] , n19486, \Kp[4] , n19485, \Kp[5] , 
            n19484, \Kp[6] , n19483, \Kp[7] , n19482, \Kp[8] , n19481, 
            \Kp[9] , n19480, \Kp[10] , n19479, \Kp[11] , n19478, 
            \Kp[12] , n19477, \Kp[13] , n19476, \Kp[14] , n19475, 
            \Kp[15] , n19474, \Ki[1] , n19473, \Ki[2] , n19472, 
            \Ki[3] , n19471, \Ki[4] , n19470, \Ki[5] , n19469, \Ki[6] , 
            n19468, \Ki[7] , n19467, \Ki[8] , n19466, \Ki[9] , n19465, 
            \Ki[10] , n19464, \Ki[11] , n19463, \Ki[12] , n19462, 
            \Ki[13] , n19461, \Ki[14] , n19452, \Ki[15] , n19451, 
            n19450, n19449, n19448, n19447, n19446, n19445, n19444, 
            n19443, n19442, n19441, n19440, n19439, n19438, n19437, 
            n19436, n19435, n19434, n19433, n19432, n19431, n19430, 
            n19429, n19428, n19427, n19426, n19425, n19424, n19423, 
            n19422, n19421, n19420, n19419, n19418, n19417, n19416, 
            n19415, n19414, n19413, n19412, n19411, n19410, n19409, 
            n19408, n19407, n19406, n19405, n19404, n19403, n19402, 
            n19401, n19400, n19399, n19398, n19397, n19396, n19395, 
            n19394, n19393, n19392, n19391, n19390, n19389, n19388, 
            n19387, n19386, n19385, n19384, n19383, \state[0] , 
            n5690, n19382, n19381, n32, n19380, n19379, n19378, 
            n19377, n19376, n19375, n19374, n19373, n19372, n19371, 
            n19370, n19369, n19368, n19367, n19366, n19365, n19364, 
            n19363, n19362, n19361, n19360, n19359, n19358, n19357, 
            n19356, n19355, n19354, n19353, n19352, n19351, n19350, 
            n19349, n19348, n19347, n19346, n19345, n19344, n19343, 
            n19342, n19341, n19340, n19339, n19338, n19337, n19336, 
            n19335, n19334, n19333, n19332, n19331, n19330, n19329, 
            n19328, n19327, n19326, n19325, n19324, n19323, n19322, 
            n19321, n19320, n19319, n19318, n19317, n19316, n19315, 
            n19314, n19313, n19312, n19023, n19311, n19310, n19309, 
            n19308, n19307, n19306, n19305, n19304, n19303, n19302, 
            n19301, n19300, n19299, n19298, n19297, n19296, n19295, 
            n19294, n19293, n19292, n19291, n19290, n19289, n19288, 
            n19287, n19286, n19285, n19284, n19283, n19282, n19281, 
            n19280, n19279, n19278, n19277, n19276, n19275, n19274, 
            n14867, n19273, n19272, n19271, n19270, n19269, n19229, 
            n19228, n19227, n19226, n19225, n19224, n19223, n19222, 
            n19165, n19164, n19163, n19162, n19161, n19160, n19159, 
            n19158, n32667, n32679, n32660, n17504, n20830, n5, 
            n38579, n18738, n18956, tx_o, r_SM_Main, VCC_net, \r_SM_Main_2__N_3487[1] , 
            n4, \r_Bit_Index[0] , n19052, n19460, n38214, tx_enable, 
            n10524, n18732, n18954, r_Rx_Data, RX_N_10, \r_Bit_Index[0]_adj_9 , 
            n23879, n4_adj_10, n4_adj_11, n17539, n19524, n19583, 
            n19035, n19034, n19033, n19032, n19031, n19030, n19029, 
            n17534, n4_adj_12) /* synthesis syn_module_defined=1 */ ;
    output n63;
    output n771;
    output n10417;
    input GND_net;
    output [7:0]\data_out_frame[19] ;
    output [7:0]\data_out_frame[23] ;
    output [7:0]\data_out_frame[24] ;
    output [7:0]\data_out_frame[17] ;
    output n3303;
    output n123;
    output \FRAME_MATCHER.state_31__N_2662[1] ;
    input clk32MHz;
    output [7:0]\data_out_frame[15] ;
    output [7:0]\data_out_frame[20] ;
    output [7:0]\data_out_frame[13] ;
    output [7:0]\data_in_frame[4] ;
    output [7:0]\data_in_frame[1] ;
    output [7:0]\data_out_frame[18] ;
    output [7:0]\data_out_frame[25] ;
    output [7:0]\data_out_frame[16] ;
    output [7:0]\data_in_frame[3] ;
    output [7:0]\data_out_frame[10] ;
    output [7:0]\data_out_frame[8] ;
    output [7:0]\data_out_frame[6] ;
    output [7:0]\data_out_frame[12] ;
    output n33567;
    output [7:0]\data_out_frame[11] ;
    output [7:0]\data_out_frame[5] ;
    output [7:0]\data_out_frame[14] ;
    output [7:0]\data_out_frame[7] ;
    output [7:0]\data_in_frame[13] ;
    output [7:0]\data_in_frame[9] ;
    output [7:0]\data_out_frame[9] ;
    output [7:0]\data_out_frame[4] ;
    output [7:0]\data_in_frame[6] ;
    output [7:0]\data_in_frame[5] ;
    output [7:0]\data_in_frame[8] ;
    output [7:0]rx_data;
    output [7:0]\data_in_frame[12] ;
    output [31:0]\FRAME_MATCHER.state ;
    output [7:0]\data_in_frame[2] ;
    output \FRAME_MATCHER.state[0] ;
    output n63_adj_8;
    output n2970;
    output n14711;
    output n39;
    output [7:0]\data_in[1] ;
    output [7:0]\data_in[0] ;
    output [7:0]\data_in[3] ;
    output [7:0]\data_in[2] ;
    output n4452;
    output [7:0]\data_in_frame[10] ;
    output [7:0]\data_in_frame[11] ;
    output rx_data_ready;
    output [23:0]setpoint;
    input \state[2] ;
    input \state[3] ;
    output n10;
    output [7:0]\data_in_frame[21] ;
    output n3;
    output n7;
    input [7:0]ID;
    output n17474;
    output n17552;
    output n17476;
    output n5592;
    output tx_active;
    input n19101;
    input n19100;
    input n19099;
    input n19098;
    input n19097;
    input n19096;
    input n19095;
    input n19094;
    input n19093;
    output [7:0]control_mode;
    input n19092;
    input n19091;
    input n19090;
    input n19089;
    input n19088;
    input n19087;
    input n19086;
    output [23:0]PWMLimit;
    input n19085;
    input n19084;
    input n19083;
    input n19082;
    input n19081;
    input n19080;
    input n19079;
    input n19078;
    input n19077;
    input n19076;
    input n19075;
    input n19074;
    input n19073;
    input n19072;
    input n19071;
    input n19070;
    input n19069;
    input n19068;
    input n19067;
    input n19066;
    input n19065;
    input n19064;
    input n38205;
    input n38206;
    input n32009;
    input n19047;
    input n19046;
    input n19044;
    output [23:0]neopxl_color;
    output LED_c;
    input n19043;
    output \Ki[0] ;
    input n19042;
    output \Kp[0] ;
    input n19041;
    input n32173;
    output DE_c;
    input n19581;
    output [23:0]IntegralLimit;
    input n19580;
    input n19579;
    input n19578;
    input n19577;
    input n19576;
    input n19575;
    input n19574;
    input n19573;
    input n19572;
    input n19571;
    input n19570;
    input n19569;
    input n19568;
    input n19567;
    input n19566;
    input n19565;
    input n19564;
    input n19563;
    input n19562;
    input n19561;
    input n19560;
    input n19559;
    input n19520;
    input n19519;
    input n19518;
    input n19517;
    input n19516;
    input n19515;
    input n19514;
    input n19513;
    input n19512;
    input n19511;
    input n19510;
    input n19509;
    input n19508;
    input n19507;
    input n19506;
    input n19505;
    input n19504;
    input n19503;
    input n19502;
    input n19501;
    input n19500;
    input n19499;
    input n19498;
    input n19497;
    input n19496;
    input n19495;
    input n19494;
    input n19493;
    input n19492;
    input n19491;
    input n19490;
    input n19489;
    output \Kp[1] ;
    input n19488;
    output \Kp[2] ;
    input n19487;
    output \Kp[3] ;
    input n19486;
    output \Kp[4] ;
    input n19485;
    output \Kp[5] ;
    input n19484;
    output \Kp[6] ;
    input n19483;
    output \Kp[7] ;
    input n19482;
    output \Kp[8] ;
    input n19481;
    output \Kp[9] ;
    input n19480;
    output \Kp[10] ;
    input n19479;
    output \Kp[11] ;
    input n19478;
    output \Kp[12] ;
    input n19477;
    output \Kp[13] ;
    input n19476;
    output \Kp[14] ;
    input n19475;
    output \Kp[15] ;
    input n19474;
    output \Ki[1] ;
    input n19473;
    output \Ki[2] ;
    input n19472;
    output \Ki[3] ;
    input n19471;
    output \Ki[4] ;
    input n19470;
    output \Ki[5] ;
    input n19469;
    output \Ki[6] ;
    input n19468;
    output \Ki[7] ;
    input n19467;
    output \Ki[8] ;
    input n19466;
    output \Ki[9] ;
    input n19465;
    output \Ki[10] ;
    input n19464;
    output \Ki[11] ;
    input n19463;
    output \Ki[12] ;
    input n19462;
    output \Ki[13] ;
    input n19461;
    output \Ki[14] ;
    input n19452;
    output \Ki[15] ;
    input n19451;
    input n19450;
    input n19449;
    input n19448;
    input n19447;
    input n19446;
    input n19445;
    input n19444;
    input n19443;
    input n19442;
    input n19441;
    input n19440;
    input n19439;
    input n19438;
    input n19437;
    input n19436;
    input n19435;
    input n19434;
    input n19433;
    input n19432;
    input n19431;
    input n19430;
    input n19429;
    input n19428;
    input n19427;
    input n19426;
    input n19425;
    input n19424;
    input n19423;
    input n19422;
    input n19421;
    input n19420;
    input n19419;
    input n19418;
    input n19417;
    input n19416;
    input n19415;
    input n19414;
    input n19413;
    input n19412;
    input n19411;
    input n19410;
    input n19409;
    input n19408;
    input n19407;
    input n19406;
    input n19405;
    input n19404;
    input n19403;
    input n19402;
    input n19401;
    input n19400;
    input n19399;
    input n19398;
    input n19397;
    input n19396;
    input n19395;
    input n19394;
    input n19393;
    input n19392;
    input n19391;
    input n19390;
    input n19389;
    input n19388;
    input n19387;
    input n19386;
    input n19385;
    input n19384;
    input n19383;
    input \state[0] ;
    output n5690;
    input n19382;
    input n19381;
    output n32;
    input n19380;
    input n19379;
    input n19378;
    input n19377;
    input n19376;
    input n19375;
    input n19374;
    input n19373;
    input n19372;
    input n19371;
    input n19370;
    input n19369;
    input n19368;
    input n19367;
    input n19366;
    input n19365;
    input n19364;
    input n19363;
    input n19362;
    input n19361;
    input n19360;
    input n19359;
    input n19358;
    input n19357;
    input n19356;
    input n19355;
    input n19354;
    input n19353;
    input n19352;
    input n19351;
    input n19350;
    input n19349;
    input n19348;
    input n19347;
    input n19346;
    input n19345;
    input n19344;
    input n19343;
    input n19342;
    input n19341;
    input n19340;
    input n19339;
    input n19338;
    input n19337;
    input n19336;
    input n19335;
    input n19334;
    input n19333;
    input n19332;
    input n19331;
    input n19330;
    input n19329;
    input n19328;
    input n19327;
    input n19326;
    input n19325;
    input n19324;
    input n19323;
    input n19322;
    input n19321;
    input n19320;
    input n19319;
    input n19318;
    input n19317;
    input n19316;
    input n19315;
    input n19314;
    input n19313;
    input n19312;
    input n19023;
    input n19311;
    input n19310;
    input n19309;
    input n19308;
    input n19307;
    input n19306;
    input n19305;
    input n19304;
    input n19303;
    input n19302;
    input n19301;
    input n19300;
    input n19299;
    input n19298;
    input n19297;
    input n19296;
    input n19295;
    input n19294;
    input n19293;
    input n19292;
    input n19291;
    input n19290;
    input n19289;
    input n19288;
    input n19287;
    input n19286;
    input n19285;
    input n19284;
    input n19283;
    input n19282;
    input n19281;
    input n19280;
    input n19279;
    input n19278;
    input n19277;
    input n19276;
    input n19275;
    input n19274;
    output n14867;
    input n19273;
    input n19272;
    input n19271;
    input n19270;
    input n19269;
    input n19229;
    input n19228;
    input n19227;
    input n19226;
    input n19225;
    input n19224;
    input n19223;
    input n19222;
    input n19165;
    input n19164;
    input n19163;
    input n19162;
    input n19161;
    input n19160;
    input n19159;
    input n19158;
    output n32667;
    output n32679;
    output n32660;
    output n17504;
    output n20830;
    output n5;
    output n38579;
    output n18738;
    output n18956;
    output tx_o;
    output [2:0]r_SM_Main;
    input VCC_net;
    output \r_SM_Main_2__N_3487[1] ;
    output n4;
    output \r_Bit_Index[0] ;
    input n19052;
    input n19460;
    input n38214;
    output tx_enable;
    output n10524;
    output n18732;
    output n18954;
    output r_Rx_Data;
    input RX_N_10;
    output \r_Bit_Index[0]_adj_9 ;
    output n23879;
    output n4_adj_10;
    output n4_adj_11;
    output n17539;
    input n19524;
    input n19583;
    input n19035;
    input n19034;
    input n19033;
    input n19032;
    input n19031;
    input n19030;
    input n19029;
    output n17534;
    output n4_adj_12;
    
    wire clk32MHz /* synthesis SET_AS_NETWORK=clk32MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(33[6:14])
    
    wire n7_c, n30170, n34061, n33296, n34391, n17126, n30116, 
        n32975, n30174, n14, n10_c, n30895, n33752, n30219, n34362, 
        n30870, n32870, n17098, n19154;
    wire [7:0]\data_in_frame[14] ;   // verilog/coms.v(96[12:25])
    
    wire n33230, n32884, n33064, n33007, n33034, n10_adj_4021, n32991, 
        n32926, n17084, n17604, n17885, Kp_23__N_1175, n8, n32759, 
        n30624, n18086, n2;
    wire [31:0]\FRAME_MATCHER.i ;   // verilog/coms.v(115[11:12])
    
    wire n27820, n2312, n32756, n6, Kp_23__N_1063, n2_adj_4022, 
        n3_c, n19153, n30866, n10_adj_4023, n19152, n32787, n30139, 
        n30073, n33133, n10_adj_4024, n30948, n34865, n30823, n33020, 
        n30058, n31000, n33890, n33156, n18019, n33259, n19151, 
        n18241, n32943, n17086, n32981, n33239, n30108, n51, n56, 
        n32997, n54, n32861, n18437, n18363, n55, n53, n32713, 
        n32994, n18330, n50, n33086, n40, n58, n62, n33088, 
        n33251, n49, n33326, n33218, n10_adj_4025, n33245, n32816, 
        n30049, n33085, n30874, n33130, n34449, n33224, n17070, 
        n33281, n10_adj_4026, n32902, n30145, n30986, n6_adj_4027, 
        n32984, n30858, n17161, n34371, n32887, n10_adj_4028;
    wire [7:0]\data_in_frame[19] ;   // verilog/coms.v(96[12:25])
    
    wire n5454, n5456, n30141, n32753, n17112, n32987, n32988, 
        n33193, n4_c, n30957, n33031, n30885, n30995, n33003, 
        n32881, n17232, n33043, n32939, n7_adj_4029, n30902, n33865, 
        n30908, n33248, n33249, n6_adj_4030, n18450, n32963, n17820, 
        n17615, n33172, n6_adj_4031, n33227, n33228, n32735, n32738, 
        n1668, n12, n33148, n1835, n33175, n17566, n32841, n18, 
        n4_adj_4032, n14993, n31, n17548, n33105, n32743, n20, 
        n16, n32908, n33278, n16_adj_4033, n1247, n17, n17622, 
        n32949, Kp_23__N_1195;
    wire [7:0]\data_in_frame[16] ;   // verilog/coms.v(96[12:25])
    
    wire n33317, n33181, n32912, n12_adj_4034, n18075, n33178, n18397, 
        n33290, n17569, n14_adj_4035, n10_adj_4036, n32829, n32864, 
        n12_adj_4037, n18424, n33187, n18503, n18496, n32844, n10_adj_4038, 
        n1168, n17243, n33028, n30018, n10_adj_4039, n32718, n10_adj_4040, 
        n33074, n17768, n33311;
    wire [7:0]n8825;
    
    wire n18619;
    wire [7:0]byte_transmit_counter;   // verilog/coms.v(102[12:33])
    
    wire n18939, n18434, n33069, n6_adj_4041, Kp_23__N_804, n8_adj_4042, 
        n32732, n8_adj_4043, n18431, n32729, n17676, n12_adj_4044, 
        n32894, n17858, n33350;
    wire [7:0]\data_in_frame[7] ;   // verilog/coms.v(96[12:25])
    
    wire n32794, n6_adj_4045, n17846, n33082, n33197, n18105, n12_adj_4046, 
        n33314, n34545, n33320, n33102, n32852, n32807, n1191, 
        n32920, n17563, n18119, n33215, n33265, n30, n33093, n33332, 
        n34, n32_c, n33, n31_adj_4047, n33120, n18275, n6_adj_4048, 
        n35042, n14_adj_4049, n33287, n33206, n15, n33308, n43, 
        n19150, n33356, n18_adj_4050, n19, n30860, n33046, n42, 
        n17_adj_4051, n31_adj_4052, n40_adj_4053, n46, n39_c, n38, 
        n47, n35183, n40_adj_4054, n38_adj_4055, n39_adj_4056, n37, 
        n42_adj_4057, n5_c, n46_adj_4058, n41, n32849, n15_adj_4059, 
        n14_adj_4060, n31008, n8_adj_4061, n33096, n10_adj_4062, n12_adj_4063, 
        n33323, n12_adj_4064, n32878, n32960, n6_adj_4065, n8_adj_4066, 
        n32666, n19166, n17582, n16_adj_4067, n17_adj_4068, n14_adj_4069, 
        n10_adj_4070, n36285, n33889, n6_adj_4071, n36284, n33256, 
        n33453, n32564, n16_adj_4072, n10_adj_4073, n17_adj_4074, 
        n36274, n36273, n16_adj_4075, n17_adj_4076, n36271, n36270, 
        n18_adj_4077;
    wire [7:0]\data_in_frame[0] ;   // verilog/coms.v(96[12:25])
    
    wire n22, n32776, n28, n18264, n17794, n30_adj_4078, Kp_23__N_843, 
        n33066, n23, n19_adj_4079, n31_adj_4080, n35326;
    wire [31:0]\FRAME_MATCHER.state_31__N_2598 ;
    
    wire n17553, n32677, n32231;
    wire [31:0]\FRAME_MATCHER.state_c ;   // verilog/coms.v(112[11:16])
    
    wire n6_adj_4081, n32021, n17551, n2_adj_4082, n4_adj_4083, n32177, 
        n32139, n32135, n32131, n32127, n32123, n32041, n32119, 
        n32115, n32111, n32107, n32103, n3_adj_4084, n1, n2_adj_4085, 
        n32027, n32099, n32095, n32091, n32087, n32005, n32083, 
        n32079, n32075, n32071, n32067, n5_adj_4086, n5534, n27821, 
        n19149;
    wire [7:0]\data_in_frame[15] ;   // verilog/coms.v(96[12:25])
    
    wire n17559, n63_adj_4087, n10_adj_4089, n24499, n17471, n17373, 
        n8_adj_4090, n24763, n11316, tx_transmit_N_3387, n44, n42_adj_4092, 
        n43_adj_4093, n41_adj_4094, n40_adj_4095, n39_adj_4096, n50_adj_4097, 
        n45, n16_adj_4098, n17_adj_4099, n17468, n17465, n18_adj_4100, 
        n20_adj_4101, n15_adj_4102, n63_adj_4103, n17384, n16_adj_4104, 
        n17_adj_4105, n63_adj_4106, n10_adj_4107, n17528, n14_adj_4108, 
        n15_adj_4109, n10_adj_4110, n14_adj_4111, n20_adj_4112, n19_adj_4113, 
        n35352, n8_adj_4114, n32063, n19148, n19147, n19146, n19145, 
        n2_adj_4115, n27819, n19167, n4_adj_4116, n33117, n33111, 
        n10_adj_4117, n19168, n19169, n18293, n33013, n33090, n12_adj_4118, 
        n30037, n33236, n30850, n33879, n16400, n30596, n28_adj_4119, 
        n30653, n32773, n33305, n18268, n26, n30008, n33293, n33338, 
        n32858, n27, n30545, n33353, n32966, n25, n33284, n6_adj_4120, 
        n32978, n33329, n33040, n14_adj_4121;
    wire [7:0]\data_in_frame[17] ;   // verilog/coms.v(96[12:25])
    
    wire n10_adj_4122, n32766, n18312, n6_adj_4123;
    wire [7:0]\data_in_frame[18] ;   // verilog/coms.v(96[12:25])
    
    wire n17901, n32873, n17863, n16_adj_4124, n33123, n17_adj_4125, 
        n30920, n35067, n33203, n17595, n18440, n10_adj_4126, n33253, 
        n6_adj_4127, n33169, n12_adj_4128, n33302, n34447, n30132, 
        n30106, n10_adj_4129, n29976, n18168, n17894, n28_adj_4130, 
        n32940, n26_adj_4131, n33344, n33166, n27_adj_4132, n30872, 
        n25_adj_4133, n35078, n54_adj_4134, n33145, n33099, n32969, 
        n52, n17704, n53_adj_4135, n33341, n30114, n33184, n51_adj_4136, 
        n33242, n32954, n30095, n48, n33010, n50_adj_4137, n49_adj_4138, 
        n60, Kp_23__N_1372, n33347, n55_adj_4139, n19144, n30666, 
        n33200, n12_adj_4140, n15914, n34344, n30093, n12_adj_4141, 
        n33262, n16_adj_4142, n17719, n33051, n12_adj_4143, n19143, 
        n30089, n17652, n29957, n17_adj_4144, n36303, n19170, n36302, 
        n16_adj_4145, n33212, n17983, n12_adj_4146, n31003, n33271, 
        n7_adj_4147, n12_adj_4148, n17_adj_4149, n19171;
    wire [0:0]n3598;
    wire [2:0]r_SM_Main_2__N_3490;
    
    wire n33511, n36306, n36305, n16_adj_4150, n6_adj_4151, n19172, 
        n19173, n17_adj_4152, n36300, n36299, \FRAME_MATCHER.rx_data_ready_prev , 
        n30900, Kp_23__N_1630, n8_adj_4153, Kp_23__N_735, n6_adj_4154, 
        n33054, n17811, n18506, n6_adj_4155, n30880, n33023, n33079, 
        n10_adj_4156, n35280, n19142, n2_adj_4157, n27818, n19141, 
        n5455, n18646, n19140, n32923, n14_adj_4158, n33162, n32824, 
        n30946, n6_adj_4159, n19139, n35440, n35438, n37877, n37751, 
        n14_adj_4160, n33108, n20_adj_4161, n37901, n36248, n17714, 
        n17827, n32749, n19_adj_4162, n29786, n17738, n21, n35434, 
        n35432, n37859, n37841, n14_adj_4164, n30876, n30939, n12_adj_4165, 
        n37907, n36272, n32899, n35427, n35428, n35426, Kp_23__N_1204, 
        n12_adj_4166, n8_adj_4167, n18460, n33114, n32746, n16_adj_4168, 
        n10_adj_4169, n37853, n37889, n14_adj_4170, n37913, n36279, 
        n34364, n30950, n33136, n2_adj_4171, n27817, n32797, n33299, 
        n33268, n12_adj_4172, n35421, n35422, n35420, n37847, n37727, 
        n14_adj_4173, n37919, n36290, n33159, n35127, n35415, n35416, 
        n35414, n18285, n17_adj_4174, n37835, n37925, n14_adj_4175, 
        n33335, n37655, n36293, n35409, n35410, n35408, n37817, 
        n37931, n14_adj_4176, n37649, n36298, n31_adj_4177, n35400, 
        n35401, n30848, n35399, n37871, n37865, n14_adj_4178, n37721, 
        n36304, n4_adj_4179, n17101, n15_adj_4180, n14_adj_4181, n10_adj_4182, 
        n34498, Kp_23__N_1069, n17730, n14_adj_4183, n10_adj_4184, 
        n12_adj_4185, n32905, n32791, n33127, n10_adj_4186, n14_adj_4187, 
        n30853, n33057, n10_adj_4188;
    wire [7:0]\data_in_frame[20] ;   // verilog/coms.v(96[12:25])
    
    wire n33708, n12_adj_4189, n18058, n6_adj_4190, n17843, n32784, 
        n33142, n27_adj_4191, n10_adj_4192, n2_adj_4193, n27816, n10_adj_4194, 
        n2_adj_4195, n27815, n19138, n19137, n5_adj_4196, n2_adj_4197, 
        n27814, n35404, n35402, n15965, n7_adj_4198, n34273, n37805, 
        n37799, n14_adj_4199, n33707, n6_adj_4200, n35054, n32702, 
        n34290, n34316, n34619, n37661, n36301, n2_adj_4201, n27813, 
        n33768, n6_adj_4202, n38349, n2_adj_4203, n27812, n10_adj_4204, 
        n32227, n32225, n32223, n32221, n32219, n32217, n32215, 
        n32213, n32211, n32209, n32207, n32205, n32203, n32201, 
        n32199, n32197, n32195, n23755, n24510, n23753, n24508, 
        n7_adj_4205, n31999, n32233, n32193, n32191, n32145, n24506, 
        n32189, n32185, n32181, n32017, n18682;
    wire [7:0]\data_out_frame[27] ;   // verilog/coms.v(97[12:26])
    
    wire n2_adj_4206, n27811, n30031, n35169, n34941, n24, n22_adj_4207, 
        n23_adj_4208, n21_adj_4209, n8_adj_4210, n33979;
    wire [7:0]\data_out_frame[26] ;   // verilog/coms.v(97[12:26])
    
    wire n32982, n33700, n33784, n32947, n34053, n18_adj_4211, n2_adj_4212, 
        n3_adj_4213, Kp_23__N_894, n27854, n26_adj_4215, n27853, n2_adj_4216, 
        n3_adj_4217, n2_adj_4218, n3_adj_4219, n2_adj_4220, n3_adj_4221, 
        n2_adj_4222, n3_adj_4223, n3_adj_4224, n3_adj_4225, n6_adj_4226, 
        Kp_23__N_862, n14_adj_4227, n10_adj_4228, n17784, n32781, 
        n32813, n17749, n18235, n32934, n32710, n6_adj_4229, n30_adj_4230, 
        n3_adj_4231, n2_adj_4232, n27810, n3_adj_4233, n3_adj_4234, 
        n3_adj_4235, n17_adj_4236, n3_adj_4237, n3_adj_4238, n3_adj_4239, 
        n3_adj_4240, n3_adj_4241, n2_adj_4242, n3_adj_4243, n2_adj_4244, 
        n3_adj_4245, n2_adj_4246, n3_adj_4247, n2_adj_4248, n3_adj_4249, 
        n2_adj_4250, n3_adj_4251, n2_adj_4252, n3_adj_4253, n2_adj_4254, 
        n3_adj_4255, n27852, n2_adj_4256, n3_adj_4257, n2_adj_4258, 
        n3_adj_4259, n2_adj_4260, n3_adj_4261, n2_adj_4262, n3_adj_4263, 
        n2_adj_4264, n3_adj_4265, n2_adj_4266, n3_adj_4267, n2_adj_4268, 
        n3_adj_4269, n2_adj_4270, n3_adj_4271, n27851, n27809, n27808, 
        n27807, n27850, n27806, n27849, n2_adj_4272, n27848, n32931, 
        n32655, n14574, n12_adj_4274, n10_adj_4275, n11, n9, n8_adj_4276, 
        n19136, n23788, n32678, n19135, n19134, n19133, n19132, 
        n19131, n19130, n19129, n19128, n19127, n19126, n19125, 
        n19124, n19123, n19122, n19121, n19120, n19119, n19118, 
        n19117, n19116, n19115, n19114, n28_adj_4277, n26_adj_4278, 
        n27_adj_4279, n25_adj_4280, n32685, n24511, n32549, n24587, 
        n27805, n32653, n161, n19113, n27804, n19112, n2994, n18858, 
        n1_adj_4281, n5_adj_4282, n24295, n19111, n17503, n23740, 
        n24226, n34406, n27803, n6_adj_4283, n37673, n37934, n7_adj_4284;
    wire [7:0]tx_data;   // verilog/coms.v(105[13:20])
    
    wire n37928, n37922, n37916, n37910, n37904, n37898, n27802, 
        n37886, n37874, n37868, n37862, n37856, n37850, n37844, 
        n37838, n37832, n27801, n37814, n37802, n37796, n33000, 
        n37679, n37790, n7_adj_4285, n37685, n37784, n7_adj_4286, 
        n37691, n37778, n7_adj_4287, n37697, n37772, n7_adj_4288, 
        n37703, n37766, n7_adj_4289, n37709, n37760, n7_adj_4290, 
        n37715, n37754, n7_adj_4291, n37748, n37724, n32769, n37718, 
        n27800, n27799, n27798, n19110, n37712, n37706, n37700, 
        n19109, n33139, n19108, n27797, n19107, n27796, n19106, 
        n19105, n19104, n19103, n19102, n5457, n27795, n36291, 
        n36292, n37694, n5458, n5459, n5460, n5461, n5462, n5463, 
        n5464, n5465, n5466, n5467, n5468, n5469, n5470, n5471, 
        n5472, n5473, n5474, n5475, n5476, n5477, n5478, n23_adj_4292, 
        n31_adj_4293, n19045, n36, n32657, n19262, n32597, n33587, 
        n19263, n19264, n19265, n19266, n19267, n19268, n35, n32916, 
        n33_adj_4294, n34_adj_4295, n17_adj_4296, n16_adj_4297, n36296, 
        n36297, n37688, n17_adj_4298, n16_adj_4299, n8_adj_4300, n8_adj_4302, 
        n8_adj_4303, n35330, n14557, n19261, n19260, n19259, n19258, 
        n19257, n15920, n19256, n19255, n19254, n19253, n19252, 
        n19251, n19250, n19249, n19248, n19247, n19246, n19245, 
        n19244, n19243, n19242, n19241, n19240, n19239, n19238, 
        n19237, n19236, n19235, n19234, n19233, n19232, n19231, 
        n19230, n19221, n19220, n19219, n19218, n19217, n19216, 
        n19215, n19214, n19213, n19212, n19211, n19210, n19209, 
        n19208, n19207, n19206, n19205, n19204, n19203, n19202, 
        n19201, n19200, n19199, n19198, n19197, n19196, n19195, 
        n19194, n19193, n19192, n19191, n19190, n19189, n19188, 
        n19187, n19186, n19185, n19184, n19183, n19182, n19181, 
        n19180, n19179, n19178, n19177, n19176, n19175, n19174, 
        n8_adj_4304, n19155, n27825, n27824, n27823, n19156, n19157, 
        n27822, n24559, n37682, n18333, n4_adj_4305, n37676, n37670, 
        n6_adj_4306, n37658, n37652, n37646;
    
    SB_LUT4 i4_4_lut (.I0(n7_c), .I1(n30170), .I2(n34061), .I3(n33296), 
            .O(n34391));
    defparam i4_4_lut.LUT_INIT = 16'h9669;
    SB_LUT4 i5366_2_lut (.I0(n63), .I1(n771), .I2(GND_net), .I3(GND_net), 
            .O(n10417));   // verilog/coms.v(157[6] 159[9])
    defparam i5366_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i2_3_lut (.I0(\data_out_frame[19] [2]), .I1(n17126), .I2(\data_out_frame[23] [6]), 
            .I3(GND_net), .O(n30116));
    defparam i2_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 i6_4_lut (.I0(n32975), .I1(n30174), .I2(n30116), .I3(\data_out_frame[19] [5]), 
            .O(n14));
    defparam i6_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut (.I0(\data_out_frame[24] [1]), .I1(n14), .I2(n10_c), 
            .I3(n30895), .O(n33752));
    defparam i7_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_846 (.I0(\data_out_frame[17] [5]), .I1(\data_out_frame[19] [7]), 
            .I2(n30219), .I3(GND_net), .O(n34362));
    defparam i2_3_lut_adj_846.LUT_INIT = 16'h9696;
    SB_LUT4 i3_4_lut (.I0(n30870), .I1(n34362), .I2(n32870), .I3(n17098), 
            .O(n30174));
    defparam i3_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_847 (.I0(n63), .I1(n3303), .I2(n123), .I3(GND_net), 
            .O(\FRAME_MATCHER.state_31__N_2662[1] ));
    defparam i2_3_lut_adj_847.LUT_INIT = 16'hfdfd;
    SB_DFF data_in_frame_0__i116 (.Q(\data_in_frame[14] [3]), .C(clk32MHz), 
           .D(n19154));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i3_4_lut_adj_848 (.I0(\data_out_frame[17] [3]), .I1(n33230), 
            .I2(n32884), .I3(\data_out_frame[15] [2]), .O(n30895));
    defparam i3_4_lut_adj_848.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_849 (.I0(n30895), .I1(n33064), .I2(\data_out_frame[19] [5]), 
            .I3(GND_net), .O(n30870));
    defparam i2_3_lut_adj_849.LUT_INIT = 16'h6969;
    SB_LUT4 i4_4_lut_adj_850 (.I0(n33007), .I1(\data_out_frame[20] [1]), 
            .I2(n30219), .I3(n33034), .O(n10_adj_4021));
    defparam i4_4_lut_adj_850.LUT_INIT = 16'h6996;
    SB_LUT4 i5_3_lut (.I0(n32991), .I1(n10_adj_4021), .I2(n30870), .I3(GND_net), 
            .O(n34061));
    defparam i5_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_adj_851 (.I0(\data_out_frame[15] [5]), .I1(n32926), 
            .I2(\data_out_frame[15] [4]), .I3(GND_net), .O(n17098));
    defparam i2_3_lut_adj_851.LUT_INIT = 16'h9696;
    SB_LUT4 i3_4_lut_adj_852 (.I0(\data_out_frame[13] [0]), .I1(\data_out_frame[15] [2]), 
            .I2(n17084), .I3(n17604), .O(n32991));
    defparam i3_4_lut_adj_852.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_853 (.I0(n32991), .I1(\data_out_frame[17] [4]), 
            .I2(\data_out_frame[15] [3]), .I3(GND_net), .O(n33064));
    defparam i2_3_lut_adj_853.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_4_lut (.I0(n17885), .I1(Kp_23__N_1175), .I2(n8), 
            .I3(n32759), .O(n30624));
    defparam i2_3_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_854 (.I0(n32975), .I1(n33064), .I2(n32870), .I3(GND_net), 
            .O(n18086));   // verilog/coms.v(71[16:27])
    defparam i2_3_lut_adj_854.LUT_INIT = 16'h9696;
    SB_LUT4 add_43_28_lut (.I0(n2312), .I1(\FRAME_MATCHER.i [26]), .I2(GND_net), 
            .I3(n27820), .O(n2)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_28_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i4_4_lut_adj_855 (.I0(\data_in_frame[4] [0]), .I1(\data_in_frame[1] [4]), 
            .I2(n32756), .I3(n6), .O(Kp_23__N_1063));   // verilog/coms.v(78[16:27])
    defparam i4_4_lut_adj_855.LUT_INIT = 16'h6996;
    SB_DFFSS \FRAME_MATCHER.i_i0  (.Q(\FRAME_MATCHER.i [0]), .C(clk32MHz), 
            .D(n2_adj_4022), .S(n3_c));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i117 (.Q(\data_in_frame[14] [4]), .C(clk32MHz), 
           .D(n19153));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i4_4_lut_adj_856 (.I0(\data_out_frame[20] [1]), .I1(\data_out_frame[19] [7]), 
            .I2(n30866), .I3(n33034), .O(n10_adj_4023));
    defparam i4_4_lut_adj_856.LUT_INIT = 16'h6996;
    SB_DFF data_in_frame_0__i118 (.Q(\data_in_frame[14] [5]), .C(clk32MHz), 
           .D(n19152));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i4_4_lut_adj_857 (.I0(n32787), .I1(n30139), .I2(n30073), .I3(n33133), 
            .O(n10_adj_4024));
    defparam i4_4_lut_adj_857.LUT_INIT = 16'h6996;
    SB_LUT4 i5_3_lut_adj_858 (.I0(n30948), .I1(n10_adj_4024), .I2(\data_out_frame[24] [5]), 
            .I3(GND_net), .O(n34865));
    defparam i5_3_lut_adj_858.LUT_INIT = 16'h6969;
    SB_LUT4 i3_4_lut_adj_859 (.I0(n30823), .I1(n33020), .I2(n30058), .I3(n31000), 
            .O(n33890));
    defparam i3_4_lut_adj_859.LUT_INIT = 16'h9669;
    SB_LUT4 i3_4_lut_adj_860 (.I0(\data_out_frame[23] [5]), .I1(n33156), 
            .I2(n18019), .I3(\data_out_frame[24] [0]), .O(n33296));
    defparam i3_4_lut_adj_860.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut (.I0(\data_out_frame[18] [0]), .I1(\data_out_frame[15] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n33259));
    defparam i1_2_lut.LUT_INIT = 16'h6666;
    SB_DFF data_in_frame_0__i119 (.Q(\data_in_frame[14] [6]), .C(clk32MHz), 
           .D(n19151));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i3_4_lut_adj_861 (.I0(n18241), .I1(n32943), .I2(\data_out_frame[13] [1]), 
            .I3(n17086), .O(n30219));
    defparam i3_4_lut_adj_861.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_862 (.I0(\data_out_frame[24] [5]), .I1(\data_out_frame[24] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n32981));
    defparam i1_2_lut_adj_862.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_863 (.I0(\data_out_frame[17] [6]), .I1(\data_out_frame[20] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n32870));   // verilog/coms.v(71[16:27])
    defparam i1_2_lut_adj_863.LUT_INIT = 16'h6666;
    SB_LUT4 i19_4_lut (.I0(\data_out_frame[24] [7]), .I1(n33239), .I2(n30108), 
            .I3(n32870), .O(n51));
    defparam i19_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i24_4_lut (.I0(\data_out_frame[24] [3]), .I1(\data_out_frame[23] [6]), 
            .I2(\data_out_frame[23] [3]), .I3(\data_out_frame[23] [7]), 
            .O(n56));
    defparam i24_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i22_4_lut (.I0(\data_out_frame[20] [1]), .I1(n32981), .I2(n32997), 
            .I3(n32926), .O(n54));
    defparam i22_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i23_4_lut (.I0(n32861), .I1(\data_out_frame[20] [7]), .I2(n18437), 
            .I3(n18363), .O(n55));
    defparam i23_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i21_4_lut (.I0(n30866), .I1(n30073), .I2(n30219), .I3(n33259), 
            .O(n53));
    defparam i21_4_lut.LUT_INIT = 16'h9669;
    SB_LUT4 i18_4_lut (.I0(n32713), .I1(n32994), .I2(\data_out_frame[25] [1]), 
            .I3(n18330), .O(n50));
    defparam i18_4_lut.LUT_INIT = 16'h9669;
    SB_LUT4 i26_4_lut (.I0(n51), .I1(n33086), .I2(n40), .I3(\data_out_frame[24] [6]), 
            .O(n58));
    defparam i26_4_lut.LUT_INIT = 16'h9669;
    SB_LUT4 i30_4_lut (.I0(n53), .I1(n55), .I2(n54), .I3(n56), .O(n62));
    defparam i30_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i17_4_lut (.I0(n33088), .I1(\data_out_frame[25] [7]), .I2(n33296), 
            .I3(n33251), .O(n49));
    defparam i17_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i31_4_lut (.I0(n49), .I1(n62), .I2(n58), .I3(n50), .O(n30948));
    defparam i31_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_864 (.I0(\data_out_frame[17] [7]), .I1(\data_out_frame[15] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n32994));   // verilog/coms.v(74[16:43])
    defparam i1_2_lut_adj_864.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_865 (.I0(\data_out_frame[20] [2]), .I1(n33326), 
            .I2(n33218), .I3(\data_out_frame[18] [0]), .O(n10_adj_4025));
    defparam i4_4_lut_adj_865.LUT_INIT = 16'h6996;
    SB_LUT4 i5_3_lut_adj_866 (.I0(n33245), .I1(n10_adj_4025), .I2(\data_out_frame[17] [6]), 
            .I3(GND_net), .O(n32816));
    defparam i5_3_lut_adj_866.LUT_INIT = 16'h9696;
    SB_LUT4 i1_4_lut (.I0(\data_out_frame[25] [0]), .I1(n30049), .I2(n33085), 
            .I3(n30874), .O(n33133));
    defparam i1_4_lut.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_adj_867 (.I0(n30866), .I1(n32816), .I2(GND_net), 
            .I3(GND_net), .O(n33156));
    defparam i1_2_lut_adj_867.LUT_INIT = 16'h9999;
    SB_LUT4 i3_4_lut_adj_868 (.I0(\data_out_frame[25] [1]), .I1(n33130), 
            .I2(n33020), .I3(n30073), .O(n34449));
    defparam i3_4_lut_adj_868.LUT_INIT = 16'h9669;
    SB_LUT4 i4_4_lut_adj_869 (.I0(n33224), .I1(n18241), .I2(n17070), .I3(n33281), 
            .O(n10_adj_4026));
    defparam i4_4_lut_adj_869.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_870 (.I0(\data_out_frame[18] [1]), .I1(n32902), 
            .I2(n10_adj_4026), .I3(n30145), .O(n33245));
    defparam i1_4_lut_adj_870.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_adj_871 (.I0(\data_out_frame[23] [0]), .I1(n30986), 
            .I2(GND_net), .I3(GND_net), .O(n32787));
    defparam i1_2_lut_adj_871.LUT_INIT = 16'h9999;
    SB_LUT4 i1_4_lut_adj_872 (.I0(\data_out_frame[20] [3]), .I1(\data_out_frame[16] [1]), 
            .I2(n6_adj_4027), .I3(n32984), .O(n30866));
    defparam i1_4_lut_adj_872.LUT_INIT = 16'h9669;
    SB_LUT4 i2_3_lut_adj_873 (.I0(n30858), .I1(n33130), .I2(n30058), .I3(GND_net), 
            .O(n17161));
    defparam i2_3_lut_adj_873.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_adj_874 (.I0(n33088), .I1(n17161), .I2(\data_out_frame[25] [1]), 
            .I3(GND_net), .O(n34371));
    defparam i2_3_lut_adj_874.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_adj_875 (.I0(\data_out_frame[16] [0]), .I1(\data_out_frame[13] [6]), 
            .I2(\data_out_frame[13] [4]), .I3(GND_net), .O(n32902));   // verilog/coms.v(75[16:43])
    defparam i2_3_lut_adj_875.LUT_INIT = 16'h9696;
    SB_LUT4 i4_4_lut_adj_876 (.I0(\data_out_frame[18] [2]), .I1(n32902), 
            .I2(n17070), .I3(n32887), .O(n10_adj_4028));
    defparam i4_4_lut_adj_876.LUT_INIT = 16'h6996;
    SB_LUT4 mux_1387_i2_3_lut (.I0(\data_in_frame[19] [1]), .I1(\data_in_frame[3] [1]), 
            .I2(n5454), .I3(GND_net), .O(n5456));
    defparam mux_1387_i2_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3_4_lut_adj_877 (.I0(\data_out_frame[20] [4]), .I1(n30141), 
            .I2(n32984), .I3(\data_out_frame[18] [3]), .O(n30049));
    defparam i3_4_lut_adj_877.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_878 (.I0(n30874), .I1(n30049), .I2(\data_out_frame[23] [1]), 
            .I3(\data_out_frame[23] [0]), .O(n33239));
    defparam i1_4_lut_adj_878.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_879 (.I0(\data_in_frame[3] [6]), .I1(\data_in_frame[3] [5]), 
            .I2(\data_in_frame[3] [7]), .I3(\data_in_frame[4] [0]), .O(n32753));   // verilog/coms.v(76[16:43])
    defparam i3_4_lut_adj_879.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_880 (.I0(\data_out_frame[25] [2]), .I1(n17112), 
            .I2(n33239), .I3(\data_out_frame[20] [6]), .O(n33088));
    defparam i3_4_lut_adj_880.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_881 (.I0(n33088), .I1(n32987), .I2(GND_net), 
            .I3(GND_net), .O(n32988));
    defparam i1_2_lut_adj_881.LUT_INIT = 16'h6666;
    SB_LUT4 i2_4_lut (.I0(\data_out_frame[15] [7]), .I1(\data_out_frame[13] [7]), 
            .I2(n33193), .I3(n4_c), .O(n30145));
    defparam i2_4_lut.LUT_INIT = 16'h9669;
    SB_LUT4 i2_3_lut_adj_882 (.I0(n30957), .I1(n33031), .I2(n30145), .I3(GND_net), 
            .O(n30885));
    defparam i2_3_lut_adj_882.LUT_INIT = 16'h6969;
    SB_LUT4 i1_2_lut_adj_883 (.I0(n30874), .I1(n33086), .I2(GND_net), 
            .I3(GND_net), .O(n30995));
    defparam i1_2_lut_adj_883.LUT_INIT = 16'h9999;
    SB_LUT4 i1_2_lut_adj_884 (.I0(\data_out_frame[23] [2]), .I1(n30885), 
            .I2(GND_net), .I3(GND_net), .O(n32997));
    defparam i1_2_lut_adj_884.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_885 (.I0(\data_out_frame[25] [3]), .I1(\data_out_frame[23] [1]), 
            .I2(n32997), .I3(n30995), .O(n32987));
    defparam i3_4_lut_adj_885.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_adj_886 (.I0(n32987), .I1(n33003), .I2(GND_net), 
            .I3(GND_net), .O(n33251));
    defparam i1_2_lut_adj_886.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_887 (.I0(n32881), .I1(\data_out_frame[16] [2]), 
            .I2(n17232), .I3(GND_net), .O(n30141));   // verilog/coms.v(71[16:27])
    defparam i2_3_lut_adj_887.LUT_INIT = 16'h9696;
    SB_LUT4 i3_4_lut_adj_888 (.I0(n30141), .I1(n33043), .I2(n32939), .I3(\data_out_frame[18] [4]), 
            .O(n30874));
    defparam i3_4_lut_adj_888.LUT_INIT = 16'h9669;
    SB_LUT4 i4_4_lut_adj_889 (.I0(n7_adj_4029), .I1(\data_out_frame[20] [6]), 
            .I2(\data_out_frame[20] [7]), .I3(n30874), .O(n30858));   // verilog/coms.v(78[16:27])
    defparam i4_4_lut_adj_889.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_adj_890 (.I0(n30073), .I1(n30858), .I2(GND_net), 
            .I3(GND_net), .O(n31000));
    defparam i1_2_lut_adj_890.LUT_INIT = 16'h6666;
    SB_LUT4 i1_4_lut_adj_891 (.I0(\data_out_frame[25] [4]), .I1(\data_out_frame[23] [2]), 
            .I2(n31000), .I3(n30902), .O(n33003));
    defparam i1_4_lut_adj_891.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut (.I0(n17126), .I1(n33865), .I2(n30908), .I3(\data_out_frame[20] [7]), 
            .O(n30073));
    defparam i1_2_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_892 (.I0(n33003), .I1(n33248), .I2(GND_net), 
            .I3(GND_net), .O(n33249));
    defparam i1_2_lut_adj_892.LUT_INIT = 16'h9999;
    SB_LUT4 i1_2_lut_adj_893 (.I0(n17084), .I1(\data_out_frame[15] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n32884));
    defparam i1_2_lut_adj_893.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_894 (.I0(\data_out_frame[17] [2]), .I1(\data_out_frame[13] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_4030));
    defparam i1_2_lut_adj_894.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_895 (.I0(\data_out_frame[15] [0]), .I1(n18450), 
            .I2(n32884), .I3(n6_adj_4030), .O(n32963));
    defparam i4_4_lut_adj_895.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_896 (.I0(n17820), .I1(n17615), .I2(n33172), .I3(n6_adj_4031), 
            .O(n17126));   // verilog/coms.v(75[16:43])
    defparam i4_4_lut_adj_896.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_897 (.I0(\data_out_frame[16] [7]), .I1(n33227), 
            .I2(GND_net), .I3(GND_net), .O(n33228));
    defparam i1_2_lut_adj_897.LUT_INIT = 16'h6666;
    SB_LUT4 i5_4_lut (.I0(n32735), .I1(n32738), .I2(n1668), .I3(\data_out_frame[10] [4]), 
            .O(n12));   // verilog/coms.v(76[16:43])
    defparam i5_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_898 (.I0(\data_out_frame[8] [3]), .I1(n12), .I2(n33148), 
            .I3(\data_out_frame[6] [0]), .O(n17084));   // verilog/coms.v(76[16:43])
    defparam i6_4_lut_adj_898.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_899 (.I0(\data_out_frame[16] [3]), .I1(\data_out_frame[16] [1]), 
            .I2(\data_out_frame[18] [4]), .I3(\data_out_frame[18] [3]), 
            .O(n33031));
    defparam i3_4_lut_adj_899.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_900 (.I0(\data_out_frame[18] [5]), .I1(\data_out_frame[16] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n33043));
    defparam i1_2_lut_adj_900.LUT_INIT = 16'h6666;
    SB_LUT4 i1047_2_lut (.I0(\data_out_frame[15] [7]), .I1(\data_out_frame[15] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n1835));   // verilog/coms.v(71[16:27])
    defparam i1047_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_901 (.I0(\data_out_frame[17] [7]), .I1(\data_out_frame[15] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n33224));
    defparam i1_2_lut_adj_901.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_902 (.I0(\data_out_frame[15] [3]), .I1(\data_out_frame[15] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n32943));
    defparam i1_2_lut_adj_902.LUT_INIT = 16'h6666;
    SB_LUT4 i7_4_lut_adj_903 (.I0(n33175), .I1(\data_out_frame[12] [7]), 
            .I2(n17566), .I3(n32841), .O(n18));   // verilog/coms.v(74[16:43])
    defparam i7_4_lut_adj_903.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_904 (.I0(n4_adj_4032), .I1(n14993), .I2(n31), 
            .I3(n17548), .O(n33567));
    defparam i3_4_lut_adj_904.LUT_INIT = 16'hfffe;
    SB_LUT4 i9_4_lut (.I0(n33105), .I1(n18), .I2(n32743), .I3(\data_out_frame[11] [0]), 
            .O(n20));   // verilog/coms.v(74[16:43])
    defparam i9_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i10_4_lut (.I0(\data_out_frame[8] [4]), .I1(n20), .I2(n16), 
            .I3(\data_out_frame[5] [7]), .O(n17086));   // verilog/coms.v(74[16:43])
    defparam i10_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_905 (.I0(\data_out_frame[14] [7]), .I1(n32908), 
            .I2(\data_out_frame[7] [7]), .I3(n33278), .O(n16_adj_4033));   // verilog/coms.v(85[17:70])
    defparam i6_4_lut_adj_905.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut_adj_906 (.I0(\data_out_frame[5] [5]), .I1(n1247), .I2(\data_out_frame[12] [7]), 
            .I3(n32738), .O(n17));   // verilog/coms.v(85[17:70])
    defparam i7_4_lut_adj_906.LUT_INIT = 16'h6996;
    SB_LUT4 i9_4_lut_adj_907 (.I0(n17), .I1(n17622), .I2(n16_adj_4033), 
            .I3(\data_out_frame[12] [5]), .O(n32949));   // verilog/coms.v(85[17:70])
    defparam i9_4_lut_adj_907.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_908 (.I0(\data_out_frame[13] [1]), .I1(n17086), 
            .I2(GND_net), .I3(GND_net), .O(n18437));
    defparam i1_2_lut_adj_908.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_4_lut_adj_909 (.I0(\data_in_frame[13] [5]), .I1(Kp_23__N_1195), 
            .I2(\data_in_frame[9] [1]), .I3(\data_in_frame[16] [0]), .O(n33317));   // verilog/coms.v(74[16:43])
    defparam i1_2_lut_4_lut_adj_909.LUT_INIT = 16'h6996;
    SB_LUT4 i5_4_lut_adj_910 (.I0(\data_out_frame[11] [4]), .I1(n33181), 
            .I2(\data_out_frame[11] [3]), .I3(n32912), .O(n12_adj_4034));
    defparam i5_4_lut_adj_910.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_911 (.I0(n18075), .I1(n12_adj_4034), .I2(\data_out_frame[13] [5]), 
            .I3(n33178), .O(n30108));
    defparam i6_4_lut_adj_911.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_912 (.I0(\data_out_frame[10] [5]), .I1(\data_out_frame[8] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n33175));   // verilog/coms.v(76[16:43])
    defparam i1_2_lut_adj_912.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_913 (.I0(\data_out_frame[9] [0]), .I1(\data_out_frame[4] [4]), 
            .I2(\data_out_frame[4] [5]), .I3(GND_net), .O(n18397));   // verilog/coms.v(76[16:27])
    defparam i2_3_lut_adj_913.LUT_INIT = 16'h9696;
    SB_LUT4 i6_4_lut_adj_914 (.I0(n33290), .I1(n17569), .I2(n32738), .I3(n18397), 
            .O(n14_adj_4035));   // verilog/coms.v(85[17:28])
    defparam i6_4_lut_adj_914.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut_adj_915 (.I0(\data_out_frame[13] [2]), .I1(n14_adj_4035), 
            .I2(n10_adj_4036), .I3(\data_out_frame[8] [4]), .O(n17604));   // verilog/coms.v(85[17:28])
    defparam i7_4_lut_adj_915.LUT_INIT = 16'h6996;
    SB_LUT4 i5_4_lut_adj_916 (.I0(n32829), .I1(n32864), .I2(\data_out_frame[8] [7]), 
            .I3(n18397), .O(n12_adj_4037));
    defparam i5_4_lut_adj_916.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_917 (.I0(n18424), .I1(n12_adj_4037), .I2(n33187), 
            .I3(n18503), .O(n17070));
    defparam i6_4_lut_adj_917.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_918 (.I0(\data_out_frame[8] [5]), .I1(\data_out_frame[10] [7]), 
            .I2(n18503), .I3(n1247), .O(n32841));
    defparam i3_4_lut_adj_918.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_919 (.I0(\data_out_frame[9] [1]), .I1(n18496), 
            .I2(\data_out_frame[8] [7]), .I3(GND_net), .O(n33178));
    defparam i2_3_lut_adj_919.LUT_INIT = 16'h9696;
    SB_LUT4 i4_4_lut_adj_920 (.I0(n32844), .I1(\data_out_frame[11] [1]), 
            .I2(\data_out_frame[13] [3]), .I3(n33178), .O(n10_adj_4038));
    defparam i4_4_lut_adj_920.LUT_INIT = 16'h6996;
    SB_LUT4 i5_3_lut_adj_921 (.I0(n32841), .I1(n10_adj_4038), .I2(\data_out_frame[11] [2]), 
            .I3(GND_net), .O(n18241));
    defparam i5_3_lut_adj_921.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_adj_922 (.I0(n17070), .I1(n17604), .I2(\data_out_frame[13] [4]), 
            .I3(GND_net), .O(n32926));
    defparam i2_3_lut_adj_922.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_923 (.I0(n32926), .I1(n18241), .I2(GND_net), 
            .I3(GND_net), .O(n33326));
    defparam i1_2_lut_adj_923.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_924 (.I0(\data_out_frame[4] [7]), .I1(\data_out_frame[7] [1]), 
            .I2(n1168), .I3(GND_net), .O(n32829));   // verilog/coms.v(71[16:69])
    defparam i2_3_lut_adj_924.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_925 (.I0(\data_out_frame[9] [3]), .I1(n32829), 
            .I2(GND_net), .I3(GND_net), .O(n33181));
    defparam i1_2_lut_adj_925.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_926 (.I0(\data_out_frame[11] [5]), .I1(n17243), 
            .I2(GND_net), .I3(GND_net), .O(n33193));
    defparam i1_2_lut_adj_926.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_4_lut_adj_927 (.I0(\data_out_frame[19] [4]), .I1(n30895), 
            .I2(n32963), .I3(n18086), .O(n33028));
    defparam i1_2_lut_4_lut_adj_927.LUT_INIT = 16'h9669;
    SB_LUT4 i880_2_lut (.I0(\data_out_frame[12] [7]), .I1(\data_out_frame[12] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n1668));   // verilog/coms.v(85[17:28])
    defparam i880_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_928 (.I0(\data_out_frame[11] [3]), .I1(\data_out_frame[11] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n33187));
    defparam i1_2_lut_adj_928.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_929 (.I0(n1668), .I1(n30018), .I2(\data_out_frame[12] [0]), 
            .I3(\data_out_frame[12] [1]), .O(n10_adj_4039));
    defparam i4_4_lut_adj_929.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_930 (.I0(\data_out_frame[11] [1]), .I1(\data_out_frame[11] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n33290));   // verilog/coms.v(85[17:28])
    defparam i1_2_lut_adj_930.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_931 (.I0(\data_out_frame[5] [7]), .I1(\data_out_frame[8] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n33278));   // verilog/coms.v(75[16:27])
    defparam i1_2_lut_adj_931.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_932 (.I0(n18496), .I1(n32718), .I2(\data_out_frame[6] [7]), 
            .I3(\data_out_frame[6] [6]), .O(n10_adj_4040));   // verilog/coms.v(85[17:70])
    defparam i4_4_lut_adj_932.LUT_INIT = 16'h6996;
    SB_LUT4 i5_3_lut_adj_933 (.I0(\data_out_frame[4] [4]), .I1(n10_adj_4040), 
            .I2(\data_out_frame[9] [2]), .I3(GND_net), .O(n32864));   // verilog/coms.v(85[17:70])
    defparam i5_3_lut_adj_933.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_adj_934 (.I0(\data_out_frame[14] [0]), .I1(n33074), 
            .I2(n17768), .I3(GND_net), .O(n33311));
    defparam i2_3_lut_adj_934.LUT_INIT = 16'h9696;
    SB_LUT4 i3_4_lut_adj_935 (.I0(\data_out_frame[11] [4]), .I1(\data_out_frame[9] [3]), 
            .I2(n32912), .I3(n32864), .O(n32887));
    defparam i3_4_lut_adj_935.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_936 (.I0(n32887), .I1(n33311), .I2(\data_out_frame[13] [7]), 
            .I3(GND_net), .O(n33281));   // verilog/coms.v(71[16:27])
    defparam i2_3_lut_adj_936.LUT_INIT = 16'h9696;
    SB_DFFESR byte_transmit_counter_i0_i7 (.Q(byte_transmit_counter[7]), .C(clk32MHz), 
            .E(n18619), .D(n8825[7]), .R(n18939));   // verilog/coms.v(127[12] 300[6])
    SB_DFFESR byte_transmit_counter_i0_i6 (.Q(byte_transmit_counter[6]), .C(clk32MHz), 
            .E(n18619), .D(n8825[6]), .R(n18939));   // verilog/coms.v(127[12] 300[6])
    SB_DFFESR byte_transmit_counter_i0_i5 (.Q(byte_transmit_counter[5]), .C(clk32MHz), 
            .E(n18619), .D(n8825[5]), .R(n18939));   // verilog/coms.v(127[12] 300[6])
    SB_DFFESR byte_transmit_counter_i0_i4 (.Q(byte_transmit_counter[4]), .C(clk32MHz), 
            .E(n18619), .D(n8825[4]), .R(n18939));   // verilog/coms.v(127[12] 300[6])
    SB_DFFESR byte_transmit_counter_i0_i3 (.Q(byte_transmit_counter[3]), .C(clk32MHz), 
            .E(n18619), .D(n8825[3]), .R(n18939));   // verilog/coms.v(127[12] 300[6])
    SB_DFFESR byte_transmit_counter_i0_i2 (.Q(byte_transmit_counter[2]), .C(clk32MHz), 
            .E(n18619), .D(n8825[2]), .R(n18939));   // verilog/coms.v(127[12] 300[6])
    SB_DFFESR byte_transmit_counter_i0_i1 (.Q(byte_transmit_counter[1]), .C(clk32MHz), 
            .E(n18619), .D(n8825[1]), .R(n18939));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i4_4_lut_adj_937 (.I0(n18434), .I1(\data_out_frame[7] [5]), 
            .I2(n33069), .I3(n6_adj_4041), .O(n17615));   // verilog/coms.v(75[16:27])
    defparam i4_4_lut_adj_937.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_938 (.I0(n17885), .I1(Kp_23__N_804), .I2(n8_adj_4042), 
            .I3(n32732), .O(n8_adj_4043));
    defparam i1_4_lut_adj_938.LUT_INIT = 16'hd77d;
    SB_LUT4 i2_3_lut_adj_939 (.I0(n18431), .I1(n32729), .I2(n17615), .I3(GND_net), 
            .O(n17676));   // verilog/coms.v(85[17:70])
    defparam i2_3_lut_adj_939.LUT_INIT = 16'h9696;
    SB_LUT4 i5_4_lut_adj_940 (.I0(\data_in_frame[6] [0]), .I1(n32753), .I2(\data_in_frame[6] [1]), 
            .I3(\data_in_frame[5] [6]), .O(n12_adj_4044));   // verilog/coms.v(76[16:43])
    defparam i5_4_lut_adj_940.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_941 (.I0(\data_in_frame[8] [2]), .I1(n12_adj_4044), 
            .I2(n32894), .I3(\data_in_frame[1] [6]), .O(n17858));   // verilog/coms.v(76[16:43])
    defparam i6_4_lut_adj_941.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_942 (.I0(\data_out_frame[13] [6]), .I1(n33281), 
            .I2(\data_out_frame[14] [1]), .I3(GND_net), .O(n32881));   // verilog/coms.v(71[16:27])
    defparam i2_3_lut_adj_942.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_943 (.I0(\data_out_frame[10] [7]), .I1(\data_out_frame[10] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n33350));
    defparam i1_2_lut_adj_943.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_944 (.I0(\data_out_frame[10] [4]), .I1(\data_out_frame[10] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n32908));   // verilog/coms.v(85[17:63])
    defparam i1_2_lut_adj_944.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_945 (.I0(\data_in_frame[7] [1]), .I1(\data_in_frame[6] [7]), 
            .I2(n32794), .I3(n6_adj_4045), .O(n17846));   // verilog/coms.v(70[16:27])
    defparam i4_4_lut_adj_945.LUT_INIT = 16'h6996;
    SB_LUT4 i5_4_lut_adj_946 (.I0(n33082), .I1(n33197), .I2(\data_out_frame[9] [3]), 
            .I3(n18105), .O(n12_adj_4046));
    defparam i5_4_lut_adj_946.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_947 (.I0(\data_out_frame[9] [4]), .I1(n12_adj_4046), 
            .I2(n33314), .I3(n1247), .O(n34545));
    defparam i6_4_lut_adj_947.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_948 (.I0(n1247), .I1(\data_out_frame[10] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n33320));   // verilog/coms.v(85[17:63])
    defparam i1_2_lut_adj_948.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_949 (.I0(\data_out_frame[8] [5]), .I1(\data_out_frame[10] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n32738));   // verilog/coms.v(85[17:70])
    defparam i1_2_lut_adj_949.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_950 (.I0(\data_out_frame[8] [7]), .I1(\data_out_frame[8] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n33102));   // verilog/coms.v(85[17:28])
    defparam i1_2_lut_adj_950.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_951 (.I0(\data_out_frame[4] [4]), .I1(\data_out_frame[6] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n32852));
    defparam i1_2_lut_adj_951.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_952 (.I0(\data_out_frame[4] [2]), .I1(\data_out_frame[6] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n33105));   // verilog/coms.v(74[16:43])
    defparam i1_2_lut_adj_952.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_953 (.I0(\data_out_frame[6] [6]), .I1(n32844), 
            .I2(GND_net), .I3(GND_net), .O(n18424));
    defparam i1_2_lut_adj_953.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_954 (.I0(\data_out_frame[4] [3]), .I1(\data_out_frame[6] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n32807));   // verilog/coms.v(75[16:43])
    defparam i1_2_lut_adj_954.LUT_INIT = 16'h6666;
    SB_LUT4 i375_2_lut (.I0(\data_out_frame[5] [7]), .I1(\data_out_frame[5] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n1191));   // verilog/coms.v(71[16:27])
    defparam i375_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_955 (.I0(\data_out_frame[5] [3]), .I1(n32920), 
            .I2(n17563), .I3(n1191), .O(n1168));   // verilog/coms.v(71[16:62])
    defparam i3_4_lut_adj_955.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_956 (.I0(\data_out_frame[5] [0]), .I1(n1168), .I2(GND_net), 
            .I3(GND_net), .O(n32718));   // verilog/coms.v(85[17:70])
    defparam i1_2_lut_adj_956.LUT_INIT = 16'h6666;
    SB_LUT4 i11_4_lut (.I0(n18119), .I1(\data_out_frame[8] [0]), .I2(n33215), 
            .I3(n33265), .O(n30));   // verilog/coms.v(75[16:27])
    defparam i11_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i15_4_lut (.I0(n18496), .I1(n30), .I2(n33093), .I3(n33332), 
            .O(n34));   // verilog/coms.v(75[16:27])
    defparam i15_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i13_4_lut (.I0(n32807), .I1(n18424), .I2(n33105), .I3(n17566), 
            .O(n32_c));   // verilog/coms.v(75[16:27])
    defparam i13_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i14_4_lut (.I0(n32852), .I1(\data_out_frame[4] [7]), .I2(\data_out_frame[4] [6]), 
            .I3(\data_out_frame[5] [5]), .O(n33));   // verilog/coms.v(75[16:27])
    defparam i14_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i12_4_lut (.I0(n33102), .I1(\data_out_frame[6] [0]), .I2(\data_out_frame[7] [1]), 
            .I3(n32735), .O(n31_adj_4047));   // verilog/coms.v(75[16:27])
    defparam i12_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_adj_957 (.I0(\data_in_frame[13] [5]), .I1(Kp_23__N_1195), 
            .I2(\data_in_frame[9] [1]), .I3(n33120), .O(n18275));   // verilog/coms.v(74[16:43])
    defparam i1_2_lut_4_lut_adj_957.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_958 (.I0(\data_out_frame[9] [0]), .I1(\data_out_frame[9] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_4048));
    defparam i1_2_lut_adj_958.LUT_INIT = 16'h6666;
    SB_LUT4 i18_4_lut_adj_959 (.I0(n31_adj_4047), .I1(n33), .I2(n32_c), 
            .I3(n34), .O(n35042));   // verilog/coms.v(75[16:27])
    defparam i18_4_lut_adj_959.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_960 (.I0(\data_out_frame[9] [1]), .I1(\data_out_frame[9] [2]), 
            .I2(n35042), .I3(n6_adj_4048), .O(n33082));
    defparam i4_4_lut_adj_960.LUT_INIT = 16'h6996;
    SB_LUT4 i5_3_lut_adj_961 (.I0(\data_out_frame[11] [5]), .I1(n30018), 
            .I2(n33082), .I3(GND_net), .O(n14_adj_4049));
    defparam i5_3_lut_adj_961.LUT_INIT = 16'h9696;
    SB_LUT4 i6_4_lut_adj_962 (.I0(n33287), .I1(\data_out_frame[13] [7]), 
            .I2(n32829), .I3(n33206), .O(n15));
    defparam i6_4_lut_adj_962.LUT_INIT = 16'h6996;
    SB_LUT4 i8_4_lut (.I0(n15), .I1(n32844), .I2(n14_adj_4049), .I3(n32738), 
            .O(n17232));
    defparam i8_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_963 (.I0(\data_out_frame[16] [7]), .I1(\data_out_frame[16] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n17820));   // verilog/coms.v(85[17:28])
    defparam i1_2_lut_adj_963.LUT_INIT = 16'h6666;
    SB_LUT4 i18_4_lut_adj_964 (.I0(n33290), .I1(n33308), .I2(\data_out_frame[12] [3]), 
            .I3(n33187), .O(n43));
    defparam i18_4_lut_adj_964.LUT_INIT = 16'h6996;
    SB_DFF data_in_frame_0__i120 (.Q(\data_in_frame[14] [7]), .C(clk32MHz), 
           .D(n19150));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i7_4_lut_adj_965 (.I0(n33069), .I1(n33356), .I2(n33320), .I3(n33193), 
            .O(n18_adj_4050));
    defparam i7_4_lut_adj_965.LUT_INIT = 16'h6996;
    SB_LUT4 i8_4_lut_adj_966 (.I0(n34545), .I1(n33308), .I2(n33350), .I3(n33175), 
            .O(n19));
    defparam i8_4_lut_adj_966.LUT_INIT = 16'h9669;
    SB_LUT4 i17_4_lut_adj_967 (.I0(n1668), .I1(\data_out_frame[11] [4]), 
            .I2(n30860), .I3(n33046), .O(n42));
    defparam i17_4_lut_adj_967.LUT_INIT = 16'h9669;
    SB_LUT4 i6_4_lut_adj_968 (.I0(n19), .I1(\data_out_frame[14] [6]), .I2(n17_adj_4051), 
            .I3(n18_adj_4050), .O(n31_adj_4052));
    defparam i6_4_lut_adj_968.LUT_INIT = 16'h6996;
    SB_LUT4 i15_4_lut_adj_969 (.I0(n30108), .I1(\data_out_frame[14] [2]), 
            .I2(\data_out_frame[15] [1]), .I3(\data_out_frame[13] [0]), 
            .O(n40_adj_4053));
    defparam i15_4_lut_adj_969.LUT_INIT = 16'h6996;
    SB_LUT4 i21_4_lut_adj_970 (.I0(n31_adj_4052), .I1(n42), .I2(n33230), 
            .I3(\data_out_frame[14] [3]), .O(n46));
    defparam i21_4_lut_adj_970.LUT_INIT = 16'h6996;
    SB_LUT4 i14_4_lut_adj_971 (.I0(n32943), .I1(n33224), .I2(n1835), .I3(\data_out_frame[15] [2]), 
            .O(n39_c));
    defparam i14_4_lut_adj_971.LUT_INIT = 16'h6996;
    SB_LUT4 i22_4_lut_adj_972 (.I0(n43), .I1(\data_out_frame[11] [6]), .I2(n38), 
            .I3(n17243), .O(n47));
    defparam i22_4_lut_adj_972.LUT_INIT = 16'h6996;
    SB_LUT4 i24_4_lut_adj_973 (.I0(n47), .I1(n39_c), .I2(n46), .I3(n40_adj_4053), 
            .O(n35183));
    defparam i24_4_lut_adj_973.LUT_INIT = 16'h6996;
    SB_LUT4 i16_4_lut (.I0(n33043), .I1(\data_out_frame[16] [5]), .I2(n33007), 
            .I3(\data_out_frame[18] [6]), .O(n40_adj_4054));
    defparam i16_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i14_4_lut_adj_974 (.I0(n35183), .I1(n33031), .I2(\data_out_frame[19] [5]), 
            .I3(\data_out_frame[18] [1]), .O(n38_adj_4055));
    defparam i14_4_lut_adj_974.LUT_INIT = 16'h9669;
    SB_LUT4 i15_4_lut_adj_975 (.I0(\data_out_frame[16] [0]), .I1(\data_out_frame[17] [5]), 
            .I2(\data_out_frame[19] [2]), .I3(\data_out_frame[17] [2]), 
            .O(n39_adj_4056));
    defparam i15_4_lut_adj_975.LUT_INIT = 16'h6996;
    SB_LUT4 i13_4_lut_adj_976 (.I0(\data_out_frame[16] [2]), .I1(\data_out_frame[19] [1]), 
            .I2(n33228), .I3(\data_out_frame[18] [7]), .O(n37));
    defparam i13_4_lut_adj_976.LUT_INIT = 16'h9669;
    SB_LUT4 i18_4_lut_adj_977 (.I0(n17676), .I1(n17820), .I2(\data_out_frame[19] [4]), 
            .I3(\data_out_frame[19] [3]), .O(n42_adj_4057));
    defparam i18_4_lut_adj_977.LUT_INIT = 16'h6996;
    SB_LUT4 equal_1577_i5_2_lut (.I0(Kp_23__N_1063), .I1(\data_in_frame[8] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n5_c));   // verilog/coms.v(236[9:81])
    defparam equal_1577_i5_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i22_4_lut_adj_978 (.I0(n37), .I1(n39_adj_4056), .I2(n38_adj_4055), 
            .I3(n40_adj_4054), .O(n46_adj_4058));
    defparam i22_4_lut_adj_978.LUT_INIT = 16'h6996;
    SB_LUT4 i17_4_lut_adj_979 (.I0(\data_out_frame[17] [0]), .I1(\data_out_frame[18] [2]), 
            .I2(\data_out_frame[17] [6]), .I3(\data_out_frame[17] [3]), 
            .O(n41));
    defparam i17_4_lut_adj_979.LUT_INIT = 16'h6996;
    SB_LUT4 i23_3_lut (.I0(n41), .I1(n46_adj_4058), .I2(n42_adj_4057), 
            .I3(GND_net), .O(n30908));
    defparam i23_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 i6_4_lut_adj_980 (.I0(n33227), .I1(n18363), .I2(\data_out_frame[18] [5]), 
            .I3(n32849), .O(n15_adj_4059));
    defparam i6_4_lut_adj_980.LUT_INIT = 16'h6996;
    SB_LUT4 i8_4_lut_adj_981 (.I0(n15_adj_4059), .I1(\data_out_frame[16] [3]), 
            .I2(n14_adj_4060), .I3(\data_out_frame[17] [1]), .O(n30986));
    defparam i8_4_lut_adj_981.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_982 (.I0(n30073), .I1(n30986), .I2(GND_net), 
            .I3(GND_net), .O(n31008));
    defparam i1_2_lut_adj_982.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_983 (.I0(\data_out_frame[23] [3]), .I1(n18363), 
            .I2(n18019), .I3(n31008), .O(n30902));
    defparam i3_4_lut_adj_983.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_adj_984 (.I0(\data_out_frame[7] [5]), .I1(\data_out_frame[8] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n18105));
    defparam i1_2_lut_adj_984.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_985 (.I0(\data_out_frame[5] [3]), .I1(\data_out_frame[9] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n33197));
    defparam i1_2_lut_adj_985.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_986 (.I0(\data_out_frame[8] [5]), .I1(\data_out_frame[11] [7]), 
            .I2(\data_out_frame[10] [0]), .I3(GND_net), .O(n33046));   // verilog/coms.v(76[16:43])
    defparam i2_3_lut_adj_986.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_987 (.I0(\data_out_frame[5] [3]), .I1(\data_out_frame[9] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n18434));   // verilog/coms.v(75[16:27])
    defparam i1_2_lut_adj_987.LUT_INIT = 16'h6666;
    SB_LUT4 i3_3_lut (.I0(\data_out_frame[5] [5]), .I1(n17768), .I2(n33265), 
            .I3(GND_net), .O(n8_adj_4061));
    defparam i3_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 i1_4_lut_adj_988 (.I0(\data_out_frame[12] [1]), .I1(n18434), 
            .I2(n8_adj_4061), .I3(n33046), .O(n33096));
    defparam i1_4_lut_adj_988.LUT_INIT = 16'h9669;
    SB_LUT4 i2_3_lut_adj_989 (.I0(\data_out_frame[5] [0]), .I1(\data_out_frame[7] [2]), 
            .I2(\data_out_frame[4] [6]), .I3(GND_net), .O(n33332));   // verilog/coms.v(85[17:28])
    defparam i2_3_lut_adj_989.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_990 (.I0(\data_out_frame[5] [2]), .I1(\data_out_frame[5] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n17563));   // verilog/coms.v(73[16:34])
    defparam i1_2_lut_adj_990.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_991 (.I0(\data_out_frame[5] [4]), .I1(\data_out_frame[9] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n33314));
    defparam i1_2_lut_adj_991.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_992 (.I0(\data_out_frame[12] [0]), .I1(\data_out_frame[11] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n33287));
    defparam i1_2_lut_adj_992.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_993 (.I0(n33287), .I1(n33074), .I2(\data_out_frame[7] [5]), 
            .I3(n33314), .O(n10_adj_4062));
    defparam i4_4_lut_adj_993.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_994 (.I0(\data_out_frame[7] [5]), .I1(\data_out_frame[7] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n18119));   // verilog/coms.v(74[16:27])
    defparam i1_2_lut_adj_994.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_995 (.I0(\data_out_frame[6] [0]), .I1(\data_out_frame[10] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n17622));   // verilog/coms.v(72[16:27])
    defparam i1_2_lut_adj_995.LUT_INIT = 16'h6666;
    SB_LUT4 i5_4_lut_adj_996 (.I0(n17622), .I1(\data_out_frame[6] [1]), 
            .I2(\data_out_frame[4] [0]), .I3(\data_out_frame[12] [4]), .O(n12_adj_4063));   // verilog/coms.v(74[16:27])
    defparam i5_4_lut_adj_996.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_997 (.I0(\data_out_frame[14] [5]), .I1(n12_adj_4063), 
            .I2(n33323), .I3(\data_out_frame[5] [4]), .O(n32729));   // verilog/coms.v(74[16:27])
    defparam i6_4_lut_adj_997.LUT_INIT = 16'h6996;
    SB_LUT4 i5_4_lut_adj_998 (.I0(\data_out_frame[5] [6]), .I1(\data_out_frame[10] [0]), 
            .I2(\data_out_frame[5] [2]), .I3(\data_out_frame[9] [6]), .O(n12_adj_4064));   // verilog/coms.v(74[16:27])
    defparam i5_4_lut_adj_998.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_999 (.I0(n18119), .I1(n12_adj_4064), .I2(\data_out_frame[10] [1]), 
            .I3(\data_out_frame[12] [2]), .O(n32878));   // verilog/coms.v(74[16:27])
    defparam i6_4_lut_adj_999.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1000 (.I0(\data_out_frame[18] [7]), .I1(\data_out_frame[14] [4]), 
            .I2(n32878), .I3(n32729), .O(n32960));   // verilog/coms.v(74[16:27])
    defparam i3_4_lut_adj_1000.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1001 (.I0(\data_out_frame[18] [6]), .I1(n32960), 
            .I2(GND_net), .I3(GND_net), .O(n32849));
    defparam i1_2_lut_adj_1001.LUT_INIT = 16'h6666;
    SB_LUT4 i1_4_lut_adj_1002 (.I0(\data_out_frame[19] [0]), .I1(\data_out_frame[16] [6]), 
            .I2(n6_adj_4065), .I3(n32939), .O(n18363));
    defparam i1_4_lut_adj_1002.LUT_INIT = 16'h9669;
    SB_LUT4 i14024_3_lut_4_lut (.I0(n8_adj_4066), .I1(n32666), .I2(rx_data[7]), 
            .I3(\data_in_frame[12] [7]), .O(n19166));
    defparam i14024_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_1003 (.I0(\data_out_frame[4] [0]), .I1(\data_out_frame[6] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n32743));   // verilog/coms.v(74[16:43])
    defparam i1_2_lut_adj_1003.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1004 (.I0(\data_out_frame[12] [5]), .I1(\data_out_frame[12] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n17582));   // verilog/coms.v(85[17:63])
    defparam i1_2_lut_adj_1004.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1005 (.I0(\data_out_frame[5] [5]), .I1(\data_out_frame[5] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n32920));   // verilog/coms.v(71[16:62])
    defparam i1_2_lut_adj_1005.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1006 (.I0(\data_out_frame[8] [2]), .I1(\data_out_frame[10] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n33323));   // verilog/coms.v(85[17:70])
    defparam i1_2_lut_adj_1006.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_1007 (.I0(\data_out_frame[8] [1]), .I1(\data_out_frame[7] [7]), 
            .I2(\data_out_frame[8] [3]), .I3(GND_net), .O(n33215));   // verilog/coms.v(72[16:27])
    defparam i2_3_lut_adj_1007.LUT_INIT = 16'h9696;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_5_i16_3_lut (.I0(\data_out_frame[16] [5]), 
            .I1(\data_out_frame[17] [5]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n16_adj_4067));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_5_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_5_i17_3_lut (.I0(\data_out_frame[18] [5]), 
            .I1(\data_out_frame[19] [5]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n17_adj_4068));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_5_i17_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i6_4_lut_adj_1008 (.I0(n33323), .I1(\data_out_frame[10] [4]), 
            .I2(n32920), .I3(n17582), .O(n14_adj_4069));   // verilog/coms.v(85[17:70])
    defparam i6_4_lut_adj_1008.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut_adj_1009 (.I0(\data_out_frame[14] [6]), .I1(n14_adj_4069), 
            .I2(n10_adj_4070), .I3(n17569), .O(n18450));   // verilog/coms.v(85[17:70])
    defparam i7_4_lut_adj_1009.LUT_INIT = 16'h6996;
    SB_LUT4 i29824_2_lut (.I0(\data_out_frame[23] [5]), .I1(byte_transmit_counter[0]), 
            .I2(GND_net), .I3(GND_net), .O(n36285));
    defparam i29824_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i4_4_lut_adj_1010 (.I0(n33889), .I1(\data_out_frame[16] [7]), 
            .I2(n32960), .I3(n6_adj_4071), .O(n33865));
    defparam i4_4_lut_adj_1010.LUT_INIT = 16'h9669;
    SB_LUT4 i29804_2_lut (.I0(\data_out_frame[20] [5]), .I1(byte_transmit_counter[0]), 
            .I2(GND_net), .I3(GND_net), .O(n36284));
    defparam i29804_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i1_2_lut_adj_1011 (.I0(\data_out_frame[19] [1]), .I1(n33865), 
            .I2(GND_net), .I3(GND_net), .O(n18019));
    defparam i1_2_lut_adj_1011.LUT_INIT = 16'h9999;
    SB_LUT4 i2_3_lut_adj_1012 (.I0(n33256), .I1(\data_out_frame[25] [5]), 
            .I2(n30902), .I3(GND_net), .O(n33248));
    defparam i2_3_lut_adj_1012.LUT_INIT = 16'h6969;
    SB_LUT4 i1_2_lut_adj_1013 (.I0(\FRAME_MATCHER.state [3]), .I1(n33453), 
            .I2(GND_net), .I3(GND_net), .O(n32564));
    defparam i1_2_lut_adj_1013.LUT_INIT = 16'h2222;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_6_i16_3_lut (.I0(\data_out_frame[16] [6]), 
            .I1(\data_out_frame[17] [6]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n16_adj_4072));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_6_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4_4_lut_adj_1014 (.I0(n33248), .I1(n32861), .I2(\data_out_frame[25] [6]), 
            .I3(n18019), .O(n10_adj_4073));
    defparam i4_4_lut_adj_1014.LUT_INIT = 16'h6996;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_6_i17_3_lut (.I0(\data_out_frame[18] [6]), 
            .I1(\data_out_frame[19] [6]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n17_adj_4074));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_6_i17_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i29827_2_lut (.I0(\data_out_frame[23] [6]), .I1(byte_transmit_counter[0]), 
            .I2(GND_net), .I3(GND_net), .O(n36274));
    defparam i29827_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i29829_2_lut (.I0(\data_out_frame[20] [6]), .I1(byte_transmit_counter[0]), 
            .I2(GND_net), .I3(GND_net), .O(n36273));
    defparam i29829_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_7_i16_3_lut (.I0(\data_out_frame[16] [7]), 
            .I1(\data_out_frame[17] [7]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n16_adj_4075));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_7_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_7_i17_3_lut (.I0(\data_out_frame[18] [7]), 
            .I1(\data_out_frame[19] [7]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n17_adj_4076));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_7_i17_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i29830_2_lut (.I0(\data_out_frame[23] [7]), .I1(byte_transmit_counter[0]), 
            .I2(GND_net), .I3(GND_net), .O(n36271));
    defparam i29830_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i29803_2_lut (.I0(\data_out_frame[20] [7]), .I1(byte_transmit_counter[0]), 
            .I2(GND_net), .I3(GND_net), .O(n36270));
    defparam i29803_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i1_2_lut_adj_1015 (.I0(\data_in_frame[1] [5]), .I1(\data_in_frame[1] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n18_adj_4077));
    defparam i1_2_lut_adj_1015.LUT_INIT = 16'h8888;
    SB_LUT4 i11_4_lut_adj_1016 (.I0(\data_in_frame[0] [7]), .I1(n22), .I2(\data_in_frame[1] [1]), 
            .I3(n32776), .O(n28));
    defparam i11_4_lut_adj_1016.LUT_INIT = 16'h0480;
    SB_LUT4 i13_4_lut_adj_1017 (.I0(n18264), .I1(n17794), .I2(n14993), 
            .I3(n18_adj_4077), .O(n30_adj_4078));
    defparam i13_4_lut_adj_1017.LUT_INIT = 16'h0100;
    SB_LUT4 i6_4_lut_adj_1018 (.I0(\data_in_frame[2] [7]), .I1(Kp_23__N_843), 
            .I2(n33066), .I3(\data_in_frame[2] [1]), .O(n23));
    defparam i6_4_lut_adj_1018.LUT_INIT = 16'h2184;
    SB_LUT4 i14_4_lut_adj_1019 (.I0(n19_adj_4079), .I1(n28), .I2(\data_in_frame[1] [2]), 
            .I3(\data_in_frame[1] [3]), .O(n31_adj_4080));
    defparam i14_4_lut_adj_1019.LUT_INIT = 16'h8000;
    SB_LUT4 i16_4_lut_adj_1020 (.I0(n31_adj_4080), .I1(n23), .I2(n30_adj_4078), 
            .I3(n35326), .O(\FRAME_MATCHER.state_31__N_2598 [3]));
    defparam i16_4_lut_adj_1020.LUT_INIT = 16'h0080;
    SB_LUT4 i1_4_lut_adj_1021 (.I0(\FRAME_MATCHER.state_31__N_2598 [3]), .I1(\FRAME_MATCHER.state [3]), 
            .I2(n17553), .I3(n32677), .O(n32231));
    defparam i1_4_lut_adj_1021.LUT_INIT = 16'hce0a;
    SB_LUT4 i1_2_lut_adj_1022 (.I0(\FRAME_MATCHER.state_c [4]), .I1(n6_adj_4081), 
            .I2(GND_net), .I3(GND_net), .O(n32021));
    defparam i1_2_lut_adj_1022.LUT_INIT = 16'h8888;
    SB_LUT4 i1_4_lut_adj_1023 (.I0(\FRAME_MATCHER.state_c [4]), .I1(n17551), 
            .I2(n2_adj_4082), .I3(n4_adj_4083), .O(n32177));
    defparam i1_4_lut_adj_1023.LUT_INIT = 16'ha2a0;
    SB_LUT4 i1_2_lut_adj_1024 (.I0(\FRAME_MATCHER.state_c [5]), .I1(n6_adj_4081), 
            .I2(GND_net), .I3(GND_net), .O(n32139));
    defparam i1_2_lut_adj_1024.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_1025 (.I0(\FRAME_MATCHER.state_c [6]), .I1(n6_adj_4081), 
            .I2(GND_net), .I3(GND_net), .O(n32135));
    defparam i1_2_lut_adj_1025.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_1026 (.I0(\FRAME_MATCHER.state_c [7]), .I1(n6_adj_4081), 
            .I2(GND_net), .I3(GND_net), .O(n32131));
    defparam i1_2_lut_adj_1026.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_1027 (.I0(\FRAME_MATCHER.state_c [9]), .I1(n6_adj_4081), 
            .I2(GND_net), .I3(GND_net), .O(n32127));
    defparam i1_2_lut_adj_1027.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_1028 (.I0(\FRAME_MATCHER.state_c [10]), .I1(n6_adj_4081), 
            .I2(GND_net), .I3(GND_net), .O(n32123));
    defparam i1_2_lut_adj_1028.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_1029 (.I0(\FRAME_MATCHER.state_c [11]), .I1(n6_adj_4081), 
            .I2(GND_net), .I3(GND_net), .O(n32041));
    defparam i1_2_lut_adj_1029.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_1030 (.I0(\FRAME_MATCHER.state_c [15]), .I1(n6_adj_4081), 
            .I2(GND_net), .I3(GND_net), .O(n32119));
    defparam i1_2_lut_adj_1030.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_1031 (.I0(\FRAME_MATCHER.state_c [16]), .I1(n6_adj_4081), 
            .I2(GND_net), .I3(GND_net), .O(n32115));
    defparam i1_2_lut_adj_1031.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_1032 (.I0(\FRAME_MATCHER.state_c [17]), .I1(n6_adj_4081), 
            .I2(GND_net), .I3(GND_net), .O(n32111));
    defparam i1_2_lut_adj_1032.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_1033 (.I0(\FRAME_MATCHER.state_c [18]), .I1(n6_adj_4081), 
            .I2(GND_net), .I3(GND_net), .O(n32107));
    defparam i1_2_lut_adj_1033.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_1034 (.I0(\FRAME_MATCHER.state_c [19]), .I1(n6_adj_4081), 
            .I2(GND_net), .I3(GND_net), .O(n32103));
    defparam i1_2_lut_adj_1034.LUT_INIT = 16'h8888;
    SB_LUT4 i1_4_lut_adj_1035 (.I0(\FRAME_MATCHER.state_c [20]), .I1(n3_adj_4084), 
            .I2(n1), .I3(n2_adj_4085), .O(n32027));
    defparam i1_4_lut_adj_1035.LUT_INIT = 16'haaa8;
    SB_LUT4 i1_2_lut_adj_1036 (.I0(\FRAME_MATCHER.state_c [21]), .I1(n6_adj_4081), 
            .I2(GND_net), .I3(GND_net), .O(n32099));
    defparam i1_2_lut_adj_1036.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_1037 (.I0(\FRAME_MATCHER.state_c [22]), .I1(n6_adj_4081), 
            .I2(GND_net), .I3(GND_net), .O(n32095));
    defparam i1_2_lut_adj_1037.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_1038 (.I0(\FRAME_MATCHER.state_c [23]), .I1(n6_adj_4081), 
            .I2(GND_net), .I3(GND_net), .O(n32091));
    defparam i1_2_lut_adj_1038.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_1039 (.I0(\FRAME_MATCHER.state_c [24]), .I1(n6_adj_4081), 
            .I2(GND_net), .I3(GND_net), .O(n32087));
    defparam i1_2_lut_adj_1039.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_1040 (.I0(\FRAME_MATCHER.state_c [25]), .I1(n6_adj_4081), 
            .I2(GND_net), .I3(GND_net), .O(n32005));
    defparam i1_2_lut_adj_1040.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_1041 (.I0(\FRAME_MATCHER.state_c [26]), .I1(n6_adj_4081), 
            .I2(GND_net), .I3(GND_net), .O(n32083));
    defparam i1_2_lut_adj_1041.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_1042 (.I0(\FRAME_MATCHER.state_c [27]), .I1(n6_adj_4081), 
            .I2(GND_net), .I3(GND_net), .O(n32079));
    defparam i1_2_lut_adj_1042.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_1043 (.I0(\FRAME_MATCHER.state_c [28]), .I1(n6_adj_4081), 
            .I2(GND_net), .I3(GND_net), .O(n32075));
    defparam i1_2_lut_adj_1043.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_1044 (.I0(\FRAME_MATCHER.state_c [29]), .I1(n6_adj_4081), 
            .I2(GND_net), .I3(GND_net), .O(n32071));
    defparam i1_2_lut_adj_1044.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_1045 (.I0(\FRAME_MATCHER.state_c [30]), .I1(n6_adj_4081), 
            .I2(GND_net), .I3(GND_net), .O(n32067));
    defparam i1_2_lut_adj_1045.LUT_INIT = 16'h8888;
    SB_LUT4 i18790_4_lut (.I0(n5_adj_4086), .I1(\FRAME_MATCHER.i [31]), 
            .I2(\FRAME_MATCHER.i [2]), .I3(\FRAME_MATCHER.i [3]), .O(n771));   // verilog/coms.v(157[9:60])
    defparam i18790_4_lut.LUT_INIT = 16'h3332;
    SB_LUT4 i1435_2_lut (.I0(\FRAME_MATCHER.state[0] ), .I1(\FRAME_MATCHER.state_c [1]), 
            .I2(GND_net), .I3(GND_net), .O(n5534));   // verilog/coms.v(145[4] 299[11])
    defparam i1435_2_lut.LUT_INIT = 16'hbbbb;
    SB_CARRY add_43_28 (.CI(n27820), .I0(\FRAME_MATCHER.i [26]), .I1(GND_net), 
            .CO(n27821));
    SB_DFF data_in_frame_0__i121 (.Q(\data_in_frame[15] [0]), .C(clk32MHz), 
           .D(n19149));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i1_2_lut_adj_1046 (.I0(\FRAME_MATCHER.state[0] ), .I1(n17551), 
            .I2(GND_net), .I3(GND_net), .O(n17553));   // verilog/coms.v(161[5:29])
    defparam i1_2_lut_adj_1046.LUT_INIT = 16'heeee;
    SB_LUT4 i1_2_lut_adj_1047 (.I0(\FRAME_MATCHER.state[0] ), .I1(\FRAME_MATCHER.state_c [2]), 
            .I2(GND_net), .I3(GND_net), .O(n4_adj_4032));   // verilog/coms.v(263[5:27])
    defparam i1_2_lut_adj_1047.LUT_INIT = 16'hbbbb;
    SB_LUT4 i4_4_lut_adj_1048 (.I0(n17559), .I1(n17553), .I2(n63_adj_4087), 
            .I3(n63_adj_8), .O(n10_adj_4089));
    defparam i4_4_lut_adj_1048.LUT_INIT = 16'h8000;
    SB_LUT4 i5_4_lut_adj_1049 (.I0(n17548), .I1(n10_adj_4089), .I2(n24499), 
            .I3(n4_adj_4032), .O(n2970));
    defparam i5_4_lut_adj_1049.LUT_INIT = 16'hc080;
    SB_LUT4 i1_2_lut_adj_1050 (.I0(\FRAME_MATCHER.i [4]), .I1(n17471), .I2(GND_net), 
            .I3(GND_net), .O(n17373));   // verilog/coms.v(154[7:23])
    defparam i1_2_lut_adj_1050.LUT_INIT = 16'heeee;
    SB_LUT4 i18791_4_lut (.I0(n8_adj_4090), .I1(\FRAME_MATCHER.i [31]), 
            .I2(n17373), .I3(\FRAME_MATCHER.i [3]), .O(n3303));   // verilog/coms.v(227[9:54])
    defparam i18791_4_lut.LUT_INIT = 16'h3230;
    SB_LUT4 i1_3_lut (.I0(n14711), .I1(n39), .I2(n3303), .I3(GND_net), 
            .O(n3_adj_4084));
    defparam i1_3_lut.LUT_INIT = 16'h0202;
    SB_LUT4 i1_2_lut_adj_1051 (.I0(n2970), .I1(n14711), .I2(GND_net), 
            .I3(GND_net), .O(n1));
    defparam i1_2_lut_adj_1051.LUT_INIT = 16'h8888;
    SB_LUT4 i30542_2_lut (.I0(n24763), .I1(n11316), .I2(GND_net), .I3(GND_net), 
            .O(tx_transmit_N_3387));
    defparam i30542_2_lut.LUT_INIT = 16'h1111;
    SB_LUT4 i18_4_lut_adj_1052 (.I0(\FRAME_MATCHER.i [30]), .I1(\FRAME_MATCHER.i [21]), 
            .I2(\FRAME_MATCHER.i [24]), .I3(\FRAME_MATCHER.i [17]), .O(n44));   // verilog/coms.v(154[7:23])
    defparam i18_4_lut_adj_1052.LUT_INIT = 16'hfffe;
    SB_LUT4 i16_4_lut_adj_1053 (.I0(\FRAME_MATCHER.i [29]), .I1(\FRAME_MATCHER.i [6]), 
            .I2(\FRAME_MATCHER.i [18]), .I3(\FRAME_MATCHER.i [23]), .O(n42_adj_4092));   // verilog/coms.v(154[7:23])
    defparam i16_4_lut_adj_1053.LUT_INIT = 16'hfffe;
    SB_LUT4 i17_4_lut_adj_1054 (.I0(\FRAME_MATCHER.i [7]), .I1(\FRAME_MATCHER.i [20]), 
            .I2(\FRAME_MATCHER.i [12]), .I3(\FRAME_MATCHER.i [14]), .O(n43_adj_4093));   // verilog/coms.v(154[7:23])
    defparam i17_4_lut_adj_1054.LUT_INIT = 16'hfffe;
    SB_LUT4 i15_4_lut_adj_1055 (.I0(\FRAME_MATCHER.i [22]), .I1(\FRAME_MATCHER.i [11]), 
            .I2(\FRAME_MATCHER.i [26]), .I3(\FRAME_MATCHER.i [16]), .O(n41_adj_4094));   // verilog/coms.v(154[7:23])
    defparam i15_4_lut_adj_1055.LUT_INIT = 16'hfffe;
    SB_LUT4 i14_4_lut_adj_1056 (.I0(\FRAME_MATCHER.i [13]), .I1(\FRAME_MATCHER.i [15]), 
            .I2(\FRAME_MATCHER.i [10]), .I3(\FRAME_MATCHER.i [28]), .O(n40_adj_4095));   // verilog/coms.v(154[7:23])
    defparam i14_4_lut_adj_1056.LUT_INIT = 16'hfffe;
    SB_LUT4 i13_2_lut (.I0(\FRAME_MATCHER.i [9]), .I1(\FRAME_MATCHER.i [27]), 
            .I2(GND_net), .I3(GND_net), .O(n39_adj_4096));   // verilog/coms.v(154[7:23])
    defparam i13_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i24_4_lut_adj_1057 (.I0(n41_adj_4094), .I1(n43_adj_4093), .I2(n42_adj_4092), 
            .I3(n44), .O(n50_adj_4097));   // verilog/coms.v(154[7:23])
    defparam i24_4_lut_adj_1057.LUT_INIT = 16'hfffe;
    SB_LUT4 i19_4_lut_adj_1058 (.I0(\FRAME_MATCHER.i [8]), .I1(\FRAME_MATCHER.i [25]), 
            .I2(\FRAME_MATCHER.i [5]), .I3(\FRAME_MATCHER.i [19]), .O(n45));   // verilog/coms.v(154[7:23])
    defparam i19_4_lut_adj_1058.LUT_INIT = 16'hfffe;
    SB_LUT4 i25_4_lut (.I0(n45), .I1(n50_adj_4097), .I2(n39_adj_4096), 
            .I3(n40_adj_4095), .O(n17471));   // verilog/coms.v(154[7:23])
    defparam i25_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i6_4_lut_adj_1059 (.I0(\data_in[1] [3]), .I1(\data_in[0] [1]), 
            .I2(\data_in[3] [2]), .I3(\data_in[0] [5]), .O(n16_adj_4098));
    defparam i6_4_lut_adj_1059.LUT_INIT = 16'hfffe;
    SB_LUT4 i7_4_lut_adj_1060 (.I0(\data_in[2] [6]), .I1(\data_in[2] [5]), 
            .I2(\data_in[2] [0]), .I3(\data_in[1] [2]), .O(n17_adj_4099));
    defparam i7_4_lut_adj_1060.LUT_INIT = 16'hfffd;
    SB_LUT4 i9_4_lut_adj_1061 (.I0(n17_adj_4099), .I1(\data_in[1] [6]), 
            .I2(n16_adj_4098), .I3(\data_in[3] [7]), .O(n17468));
    defparam i9_4_lut_adj_1061.LUT_INIT = 16'hfbff;
    SB_LUT4 i7_4_lut_adj_1062 (.I0(\data_in[2] [4]), .I1(\data_in[2] [2]), 
            .I2(n17465), .I3(\data_in[1] [0]), .O(n18_adj_4100));
    defparam i7_4_lut_adj_1062.LUT_INIT = 16'hfffd;
    SB_LUT4 i9_4_lut_adj_1063 (.I0(\data_in[1] [4]), .I1(n18_adj_4100), 
            .I2(\data_in[1] [5]), .I3(\data_in[0] [3]), .O(n20_adj_4101));
    defparam i9_4_lut_adj_1063.LUT_INIT = 16'hfffd;
    SB_LUT4 i10_4_lut_adj_1064 (.I0(n15_adj_4102), .I1(n20_adj_4101), .I2(n17468), 
            .I3(\data_in[0] [6]), .O(n63_adj_4103));
    defparam i10_4_lut_adj_1064.LUT_INIT = 16'hfeff;
    SB_LUT4 i6_4_lut_adj_1065 (.I0(n17384), .I1(\data_in[0] [7]), .I2(\data_in[2] [1]), 
            .I3(\data_in[2] [3]), .O(n16_adj_4104));
    defparam i6_4_lut_adj_1065.LUT_INIT = 16'hefff;
    SB_LUT4 i7_4_lut_adj_1066 (.I0(\data_in[0] [2]), .I1(\data_in[3] [6]), 
            .I2(\data_in[3] [1]), .I3(n17468), .O(n17_adj_4105));
    defparam i7_4_lut_adj_1066.LUT_INIT = 16'hffdf;
    SB_LUT4 i9_4_lut_adj_1067 (.I0(n17_adj_4105), .I1(\data_in[3] [3]), 
            .I2(n16_adj_4104), .I3(\data_in[3] [5]), .O(n63_adj_4106));
    defparam i9_4_lut_adj_1067.LUT_INIT = 16'hfbff;
    SB_LUT4 i4_4_lut_adj_1068 (.I0(\data_in[1] [7]), .I1(\data_in[0] [0]), 
            .I2(\data_in[1] [1]), .I3(\data_in[0] [4]), .O(n10_adj_4107));
    defparam i4_4_lut_adj_1068.LUT_INIT = 16'hfdff;
    SB_LUT4 i5_3_lut_adj_1069 (.I0(\data_in[3] [4]), .I1(n10_adj_4107), 
            .I2(\data_in[2] [7]), .I3(GND_net), .O(n17528));
    defparam i5_3_lut_adj_1069.LUT_INIT = 16'hdfdf;
    SB_LUT4 i5_3_lut_adj_1070 (.I0(\data_in[0] [3]), .I1(\data_in[1] [4]), 
            .I2(\data_in[1] [5]), .I3(GND_net), .O(n14_adj_4108));
    defparam i5_3_lut_adj_1070.LUT_INIT = 16'hdfdf;
    SB_LUT4 i6_4_lut_adj_1071 (.I0(\data_in[0] [6]), .I1(n17528), .I2(\data_in[2] [4]), 
            .I3(\data_in[1] [0]), .O(n15_adj_4109));
    defparam i6_4_lut_adj_1071.LUT_INIT = 16'hfeff;
    SB_LUT4 i8_4_lut_adj_1072 (.I0(n15_adj_4109), .I1(\data_in[2] [2]), 
            .I2(n14_adj_4108), .I3(\data_in[3] [0]), .O(n17384));
    defparam i8_4_lut_adj_1072.LUT_INIT = 16'hfbff;
    SB_LUT4 i2_2_lut (.I0(\data_in[2] [3]), .I1(\data_in[3] [5]), .I2(GND_net), 
            .I3(GND_net), .O(n10_adj_4110));
    defparam i2_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i6_4_lut_adj_1073 (.I0(\data_in[0] [2]), .I1(\data_in[3] [3]), 
            .I2(\data_in[3] [1]), .I3(\data_in[0] [7]), .O(n14_adj_4111));
    defparam i6_4_lut_adj_1073.LUT_INIT = 16'hfeff;
    SB_LUT4 i7_4_lut_adj_1074 (.I0(\data_in[3] [6]), .I1(n14_adj_4111), 
            .I2(n10_adj_4110), .I3(\data_in[2] [1]), .O(n17465));
    defparam i7_4_lut_adj_1074.LUT_INIT = 16'hfffd;
    SB_LUT4 i8_4_lut_adj_1075 (.I0(n17465), .I1(\data_in[1] [3]), .I2(n17384), 
            .I3(\data_in[2] [0]), .O(n20_adj_4112));
    defparam i8_4_lut_adj_1075.LUT_INIT = 16'hfbff;
    SB_LUT4 i7_4_lut_adj_1076 (.I0(\data_in[2] [6]), .I1(\data_in[1] [6]), 
            .I2(\data_in[3] [7]), .I3(\data_in[0] [1]), .O(n19_adj_4113));
    defparam i7_4_lut_adj_1076.LUT_INIT = 16'hfeff;
    SB_LUT4 i28598_4_lut (.I0(\data_in[1] [2]), .I1(\data_in[3] [2]), .I2(\data_in[2] [5]), 
            .I3(\data_in[0] [5]), .O(n35352));
    defparam i28598_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i11_3_lut (.I0(n35352), .I1(n19_adj_4113), .I2(n20_adj_4112), 
            .I3(GND_net), .O(n63));
    defparam i11_3_lut.LUT_INIT = 16'hfdfd;
    SB_LUT4 i18792_4_lut (.I0(n8_adj_4114), .I1(\FRAME_MATCHER.i [31]), 
            .I2(n17471), .I3(\FRAME_MATCHER.i [4]), .O(n4452));   // verilog/coms.v(259[9:58])
    defparam i18792_4_lut.LUT_INIT = 16'h3230;
    SB_LUT4 i1_2_lut_adj_1077 (.I0(\FRAME_MATCHER.state_c [31]), .I1(n6_adj_4081), 
            .I2(GND_net), .I3(GND_net), .O(n32063));
    defparam i1_2_lut_adj_1077.LUT_INIT = 16'h8888;
    SB_DFF data_in_frame_0__i122 (.Q(\data_in_frame[15] [1]), .C(clk32MHz), 
           .D(n19148));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i123 (.Q(\data_in_frame[15] [2]), .C(clk32MHz), 
           .D(n19147));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i124 (.Q(\data_in_frame[15] [3]), .C(clk32MHz), 
           .D(n19146));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i125 (.Q(\data_in_frame[15] [4]), .C(clk32MHz), 
           .D(n19145));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 add_43_27_lut (.I0(n2312), .I1(\FRAME_MATCHER.i [25]), .I2(GND_net), 
            .I3(n27819), .O(n2_adj_4115)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_27_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i14025_3_lut_4_lut (.I0(n8_adj_4066), .I1(n32666), .I2(rx_data[6]), 
            .I3(\data_in_frame[12] [6]), .O(n19167));
    defparam i14025_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i4_4_lut_adj_1078 (.I0(n4_adj_4116), .I1(\data_in_frame[8] [5]), 
            .I2(n33117), .I3(n33111), .O(n10_adj_4117));   // verilog/coms.v(78[16:27])
    defparam i4_4_lut_adj_1078.LUT_INIT = 16'h6996;
    SB_LUT4 i14026_3_lut_4_lut (.I0(n8_adj_4066), .I1(n32666), .I2(rx_data[5]), 
            .I3(\data_in_frame[12] [5]), .O(n19168));
    defparam i14026_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i14027_3_lut_4_lut (.I0(n8_adj_4066), .I1(n32666), .I2(rx_data[4]), 
            .I3(\data_in_frame[12] [4]), .O(n19169));
    defparam i14027_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i5_3_lut_adj_1079 (.I0(\data_in_frame[1] [5]), .I1(n10_adj_4117), 
            .I2(\data_in_frame[4] [1]), .I3(GND_net), .O(n18293));   // verilog/coms.v(78[16:27])
    defparam i5_3_lut_adj_1079.LUT_INIT = 16'h9696;
    SB_LUT4 i5_4_lut_adj_1080 (.I0(n33013), .I1(n33090), .I2(\data_in_frame[19] [0]), 
            .I3(\data_in_frame[16] [4]), .O(n12_adj_4118));
    defparam i5_4_lut_adj_1080.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_1081 (.I0(n30037), .I1(n12_adj_4118), .I2(n33236), 
            .I3(n30850), .O(n33879));
    defparam i6_4_lut_adj_1081.LUT_INIT = 16'h6996;
    SB_LUT4 i12_4_lut_adj_1082 (.I0(n16400), .I1(\data_in_frame[7] [1]), 
            .I2(\data_in_frame[9] [5]), .I3(n30596), .O(n28_adj_4119));
    defparam i12_4_lut_adj_1082.LUT_INIT = 16'h6996;
    SB_LUT4 i10_4_lut_adj_1083 (.I0(n30653), .I1(n32773), .I2(n33305), 
            .I3(n18268), .O(n26));
    defparam i10_4_lut_adj_1083.LUT_INIT = 16'h6996;
    SB_LUT4 i11_4_lut_adj_1084 (.I0(n30008), .I1(n33293), .I2(n33338), 
            .I3(n32858), .O(n27));
    defparam i11_4_lut_adj_1084.LUT_INIT = 16'h6996;
    SB_LUT4 i9_4_lut_adj_1085 (.I0(\data_in_frame[14] [2]), .I1(n30545), 
            .I2(n33353), .I3(n32966), .O(n25));
    defparam i9_4_lut_adj_1085.LUT_INIT = 16'h6996;
    SB_LUT4 i15_4_lut_adj_1086 (.I0(n25), .I1(n27), .I2(n26), .I3(n28_adj_4119), 
            .O(n30037));
    defparam i15_4_lut_adj_1086.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_1087 (.I0(n33284), .I1(\data_in_frame[16] [2]), 
            .I2(n30037), .I3(n6_adj_4120), .O(n32978));
    defparam i4_4_lut_adj_1087.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_1088 (.I0(n33329), .I1(\data_in_frame[15] [2]), 
            .I2(n33040), .I3(\data_in_frame[15] [1]), .O(n14_adj_4121));
    defparam i6_4_lut_adj_1088.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut_adj_1089 (.I0(\data_in_frame[17] [3]), .I1(n14_adj_4121), 
            .I2(n10_adj_4122), .I3(n32766), .O(n18312));
    defparam i7_4_lut_adj_1089.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1090 (.I0(\data_in_frame[16] [0]), .I1(\data_in_frame[15] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_4123));   // verilog/coms.v(70[16:27])
    defparam i1_2_lut_adj_1090.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1091 (.I0(\data_in_frame[18] [0]), .I1(\data_in_frame[15] [6]), 
            .I2(n17901), .I3(n6_adj_4123), .O(n32873));   // verilog/coms.v(70[16:27])
    defparam i4_4_lut_adj_1091.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1092 (.I0(\data_in_frame[12] [6]), .I1(\data_in_frame[14] [7]), 
            .I2(\data_in_frame[12] [5]), .I3(GND_net), .O(n32766));
    defparam i2_3_lut_adj_1092.LUT_INIT = 16'h9696;
    SB_LUT4 i6_4_lut_adj_1093 (.I0(n17863), .I1(\data_in_frame[17] [1]), 
            .I2(n32766), .I3(n5_c), .O(n16_adj_4124));
    defparam i6_4_lut_adj_1093.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut_adj_1094 (.I0(\data_in_frame[16] [7]), .I1(\data_in_frame[15] [0]), 
            .I2(n33123), .I3(\data_in_frame[12] [3]), .O(n17_adj_4125));
    defparam i7_4_lut_adj_1094.LUT_INIT = 16'h6996;
    SB_LUT4 i9_4_lut_adj_1095 (.I0(n17_adj_4125), .I1(\data_in_frame[14] [5]), 
            .I2(n16_adj_4124), .I3(n30920), .O(n35067));
    defparam i9_4_lut_adj_1095.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_1096 (.I0(\data_in_frame[18] [4]), .I1(n33203), 
            .I2(n17595), .I3(n18440), .O(n10_adj_4126));   // verilog/coms.v(74[16:43])
    defparam i4_4_lut_adj_1096.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1097 (.I0(\data_in_frame[12] [6]), .I1(\data_in_frame[13] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n33253));
    defparam i1_2_lut_adj_1097.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1098 (.I0(\data_in_frame[15] [0]), .I1(n18293), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_4127));
    defparam i1_2_lut_adj_1098.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1099 (.I0(\data_in_frame[12] [5]), .I1(\data_in_frame[10] [6]), 
            .I2(\data_in_frame[14] [6]), .I3(n6_adj_4127), .O(n33169));
    defparam i4_4_lut_adj_1099.LUT_INIT = 16'h6996;
    SB_LUT4 i5_4_lut_adj_1100 (.I0(n33169), .I1(n33253), .I2(\data_in_frame[17] [2]), 
            .I3(n5_c), .O(n12_adj_4128));
    defparam i5_4_lut_adj_1100.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_1101 (.I0(\data_in_frame[15] [1]), .I1(n12_adj_4128), 
            .I2(n33302), .I3(\data_in_frame[12] [7]), .O(n34447));
    defparam i6_4_lut_adj_1101.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1102 (.I0(n30132), .I1(\data_in_frame[18] [6]), 
            .I2(n30106), .I3(GND_net), .O(n33013));
    defparam i2_3_lut_adj_1102.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_adj_1103 (.I0(\data_in_frame[10] [5]), .I1(\data_in_frame[12] [4]), 
            .I2(\data_in_frame[10] [1]), .I3(GND_net), .O(n33123));
    defparam i2_3_lut_adj_1103.LUT_INIT = 16'h9696;
    SB_LUT4 i4_4_lut_adj_1104 (.I0(\data_in_frame[11] [6]), .I1(\data_in_frame[12] [1]), 
            .I2(\data_in_frame[9] [6]), .I3(\data_in_frame[9] [5]), .O(n10_adj_4129));
    defparam i4_4_lut_adj_1104.LUT_INIT = 16'h6996;
    SB_LUT4 i5_3_lut_adj_1105 (.I0(\data_in_frame[12] [0]), .I1(n10_adj_4129), 
            .I2(n29976), .I3(GND_net), .O(n33305));
    defparam i5_3_lut_adj_1105.LUT_INIT = 16'h9696;
    SB_LUT4 i12_4_lut_adj_1106 (.I0(n18168), .I1(\data_in_frame[11] [7]), 
            .I2(n17894), .I3(\data_in_frame[12] [7]), .O(n28_adj_4130));
    defparam i12_4_lut_adj_1106.LUT_INIT = 16'h6996;
    SB_LUT4 i10_4_lut_adj_1107 (.I0(n33305), .I1(\data_in_frame[10] [6]), 
            .I2(n32940), .I3(\data_in_frame[12] [6]), .O(n26_adj_4131));
    defparam i10_4_lut_adj_1107.LUT_INIT = 16'h6996;
    SB_LUT4 i11_4_lut_adj_1108 (.I0(n33344), .I1(n33120), .I2(n33166), 
            .I3(n32759), .O(n27_adj_4132));
    defparam i11_4_lut_adj_1108.LUT_INIT = 16'h6996;
    SB_LUT4 i9_4_lut_adj_1109 (.I0(n30872), .I1(n33123), .I2(\data_in_frame[11] [0]), 
            .I3(\data_in_frame[10] [3]), .O(n25_adj_4133));
    defparam i9_4_lut_adj_1109.LUT_INIT = 16'h9669;
    SB_LUT4 i15_4_lut_adj_1110 (.I0(n25_adj_4133), .I1(n27_adj_4132), .I2(n26_adj_4131), 
            .I3(n28_adj_4130), .O(n35078));
    defparam i15_4_lut_adj_1110.LUT_INIT = 16'h6996;
    SB_LUT4 i23_4_lut_adj_1111 (.I0(\data_in_frame[17] [3]), .I1(n34447), 
            .I2(\data_in_frame[14] [2]), .I3(\data_in_frame[17] [5]), .O(n54_adj_4134));
    defparam i23_4_lut_adj_1111.LUT_INIT = 16'h9669;
    SB_LUT4 i21_4_lut_adj_1112 (.I0(n33145), .I1(n33013), .I2(n33099), 
            .I3(n32969), .O(n52));
    defparam i21_4_lut_adj_1112.LUT_INIT = 16'h6996;
    SB_LUT4 i22_4_lut_adj_1113 (.I0(n30920), .I1(\data_in_frame[15] [7]), 
            .I2(n17704), .I3(n35078), .O(n53_adj_4135));
    defparam i22_4_lut_adj_1113.LUT_INIT = 16'h6996;
    SB_LUT4 i20_4_lut (.I0(\data_in_frame[18] [1]), .I1(n33341), .I2(n30114), 
            .I3(n33184), .O(n51_adj_4136));
    defparam i20_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1114 (.I0(\data_in_frame[18] [2]), .I1(n33242), 
            .I2(GND_net), .I3(GND_net), .O(n32954));
    defparam i1_2_lut_adj_1114.LUT_INIT = 16'h6666;
    SB_LUT4 i17_4_lut_adj_1115 (.I0(n30095), .I1(n33169), .I2(Kp_23__N_1195), 
            .I3(n32954), .O(n48));
    defparam i17_4_lut_adj_1115.LUT_INIT = 16'h6996;
    SB_LUT4 i19_4_lut_adj_1116 (.I0(n33010), .I1(\data_in_frame[14] [3]), 
            .I2(\data_in_frame[13] [3]), .I3(\data_in_frame[15] [4]), .O(n50_adj_4137));
    defparam i19_4_lut_adj_1116.LUT_INIT = 16'h6996;
    SB_LUT4 i18_4_lut_adj_1117 (.I0(\data_in_frame[13] [1]), .I1(n33284), 
            .I2(\data_in_frame[18] [7]), .I3(n33123), .O(n49_adj_4138));
    defparam i18_4_lut_adj_1117.LUT_INIT = 16'h6996;
    SB_LUT4 i29_4_lut (.I0(n51_adj_4136), .I1(n53_adj_4135), .I2(n52), 
            .I3(n54_adj_4134), .O(n60));
    defparam i29_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i24_4_lut_adj_1118 (.I0(Kp_23__N_1372), .I1(n48), .I2(n33347), 
            .I3(n35067), .O(n55_adj_4139));
    defparam i24_4_lut_adj_1118.LUT_INIT = 16'h9669;
    SB_DFF data_in_frame_0__i126 (.Q(\data_in_frame[15] [5]), .C(clk32MHz), 
           .D(n19144));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i30_4_lut_adj_1119 (.I0(n55_adj_4139), .I1(n60), .I2(n49_adj_4138), 
            .I3(n50_adj_4137), .O(n30666));
    defparam i30_4_lut_adj_1119.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1120 (.I0(\data_in_frame[9] [7]), .I1(n33200), 
            .I2(n30596), .I3(GND_net), .O(n30920));
    defparam i2_3_lut_adj_1120.LUT_INIT = 16'h9696;
    SB_LUT4 i5_4_lut_adj_1121 (.I0(n30920), .I1(\data_in_frame[10] [1]), 
            .I2(\data_in_frame[12] [4]), .I3(\data_in_frame[10] [3]), .O(n12_adj_4140));
    defparam i5_4_lut_adj_1121.LUT_INIT = 16'h9669;
    SB_LUT4 i6_4_lut_adj_1122 (.I0(n15914), .I1(n12_adj_4140), .I2(\data_in_frame[14] [5]), 
            .I3(\data_in_frame[12] [3]), .O(n30132));
    defparam i6_4_lut_adj_1122.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1123 (.I0(\data_in_frame[16] [6]), .I1(n34344), 
            .I2(GND_net), .I3(GND_net), .O(n33090));
    defparam i1_2_lut_adj_1123.LUT_INIT = 16'h9999;
    SB_LUT4 i3_4_lut_adj_1124 (.I0(\data_in_frame[16] [5]), .I1(n33090), 
            .I2(n30132), .I3(n30093), .O(n30106));
    defparam i3_4_lut_adj_1124.LUT_INIT = 16'h6996;
    SB_LUT4 i5_4_lut_adj_1125 (.I0(\data_in_frame[15] [3]), .I1(\data_in_frame[10] [4]), 
            .I2(\data_in_frame[12] [7]), .I3(\data_in_frame[17] [4]), .O(n12_adj_4141));
    defparam i5_4_lut_adj_1125.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_1126 (.I0(n17858), .I1(n12_adj_4141), .I2(\data_in_frame[15] [2]), 
            .I3(\data_in_frame[13] [2]), .O(n33010));
    defparam i6_4_lut_adj_1126.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1127 (.I0(\data_in_frame[12] [7]), .I1(\data_in_frame[13] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n33262));
    defparam i1_2_lut_adj_1127.LUT_INIT = 16'h6666;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_1_i16_3_lut (.I0(\data_out_frame[16] [1]), 
            .I1(\data_out_frame[17] [1]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n16_adj_4142));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_1_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_adj_1128 (.I0(n17863), .I1(n18293), .I2(GND_net), 
            .I3(GND_net), .O(n17719));   // verilog/coms.v(75[16:43])
    defparam i1_2_lut_adj_1128.LUT_INIT = 16'h6666;
    SB_LUT4 i5_4_lut_adj_1129 (.I0(n17719), .I1(n33051), .I2(\data_in_frame[17] [5]), 
            .I3(\data_in_frame[10] [5]), .O(n12_adj_4143));
    defparam i5_4_lut_adj_1129.LUT_INIT = 16'h6996;
    SB_DFF data_in_frame_0__i127 (.Q(\data_in_frame[15] [6]), .C(clk32MHz), 
           .D(n19143));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i6_4_lut_adj_1130 (.I0(n30089), .I1(n12_adj_4143), .I2(n33262), 
            .I3(\data_in_frame[15] [3]), .O(n17652));
    defparam i6_4_lut_adj_1130.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1131 (.I0(\data_in_frame[10] [2]), .I1(n29957), 
            .I2(GND_net), .I3(GND_net), .O(n33099));
    defparam i1_2_lut_adj_1131.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1132 (.I0(\data_in_frame[12] [5]), .I1(\data_in_frame[10] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n33166));
    defparam i1_2_lut_adj_1132.LUT_INIT = 16'h6666;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_1_i17_3_lut (.I0(\data_out_frame[18] [1]), 
            .I1(\data_out_frame[19] [1]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n17_adj_4144));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_1_i17_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i29810_2_lut (.I0(\data_out_frame[23] [1]), .I1(byte_transmit_counter[0]), 
            .I2(GND_net), .I3(GND_net), .O(n36303));
    defparam i29810_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i14028_3_lut_4_lut (.I0(n8_adj_4066), .I1(n32666), .I2(rx_data[3]), 
            .I3(\data_in_frame[12] [3]), .O(n19170));
    defparam i14028_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i29812_2_lut (.I0(\data_out_frame[20] [1]), .I1(byte_transmit_counter[0]), 
            .I2(GND_net), .I3(GND_net), .O(n36302));
    defparam i29812_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_0_i16_3_lut (.I0(\data_out_frame[16] [0]), 
            .I1(\data_out_frame[17] [0]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n16_adj_4145));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_0_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i5_4_lut_adj_1133 (.I0(n32732), .I1(n33212), .I2(n17983), 
            .I3(\data_in_frame[6] [0]), .O(n12_adj_4146));
    defparam i5_4_lut_adj_1133.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_1134 (.I0(n31003), .I1(n12_adj_4146), .I2(n33271), 
            .I3(\data_in_frame[7] [6]), .O(n29957));
    defparam i6_4_lut_adj_1134.LUT_INIT = 16'h9669;
    SB_LUT4 i5_4_lut_adj_1135 (.I0(n17983), .I1(n7_adj_4147), .I2(n17894), 
            .I3(n30545), .O(n12_adj_4148));
    defparam i5_4_lut_adj_1135.LUT_INIT = 16'hdfff;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_0_i17_3_lut (.I0(\data_out_frame[18] [0]), 
            .I1(\data_out_frame[19] [0]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n17_adj_4149));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_0_i17_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14029_3_lut_4_lut (.I0(n8_adj_4066), .I1(n32666), .I2(rx_data[2]), 
            .I3(\data_in_frame[12] [2]), .O(n19171));
    defparam i14029_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFFSR tx_transmit_3871 (.Q(r_SM_Main_2__N_3490[0]), .C(clk32MHz), 
            .D(n3598[0]), .R(n33511));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i2_3_lut_adj_1136 (.I0(\data_in_frame[12] [3]), .I1(n33341), 
            .I2(\data_in_frame[10] [2]), .I3(GND_net), .O(n32940));
    defparam i2_3_lut_adj_1136.LUT_INIT = 16'h9696;
    SB_LUT4 i29774_2_lut (.I0(\data_out_frame[23] [0]), .I1(byte_transmit_counter[0]), 
            .I2(GND_net), .I3(GND_net), .O(n36306));
    defparam i29774_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i29761_2_lut (.I0(\data_out_frame[20] [0]), .I1(byte_transmit_counter[0]), 
            .I2(GND_net), .I3(GND_net), .O(n36305));
    defparam i29761_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_2_i16_3_lut (.I0(\data_out_frame[16] [2]), 
            .I1(\data_out_frame[17] [2]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n16_adj_4150));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_2_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4_4_lut_adj_1137 (.I0(\data_in_frame[14] [6]), .I1(n17858), 
            .I2(n33166), .I3(n6_adj_4151), .O(n30850));
    defparam i4_4_lut_adj_1137.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1138 (.I0(n30850), .I1(\data_in_frame[14] [4]), 
            .I2(n32940), .I3(n29957), .O(n33236));
    defparam i3_4_lut_adj_1138.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_adj_1139 (.I0(\data_in_frame[16] [7]), .I1(\data_in_frame[16] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n32969));
    defparam i1_2_lut_adj_1139.LUT_INIT = 16'h6666;
    SB_LUT4 i14030_3_lut_4_lut (.I0(n8_adj_4066), .I1(n32666), .I2(rx_data[1]), 
            .I3(\data_in_frame[12] [1]), .O(n19172));
    defparam i14030_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i14031_3_lut_4_lut (.I0(n8_adj_4066), .I1(n32666), .I2(rx_data[0]), 
            .I3(\data_in_frame[12] [0]), .O(n19173));
    defparam i14031_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_2_i17_3_lut (.I0(\data_out_frame[18] [2]), 
            .I1(\data_out_frame[19] [2]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n17_adj_4152));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_2_i17_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i29813_2_lut (.I0(\data_out_frame[23] [2]), .I1(byte_transmit_counter[0]), 
            .I2(GND_net), .I3(GND_net), .O(n36300));
    defparam i29813_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i29815_2_lut (.I0(\data_out_frame[20] [2]), .I1(byte_transmit_counter[0]), 
            .I2(GND_net), .I3(GND_net), .O(n36299));
    defparam i29815_2_lut.LUT_INIT = 16'h2222;
    SB_DFF \FRAME_MATCHER.rx_data_ready_prev_3872  (.Q(\FRAME_MATCHER.rx_data_ready_prev ), 
           .C(clk32MHz), .D(rx_data_ready));   // verilog/coms.v(127[12] 300[6])
    SB_CARRY add_43_27 (.CI(n27819), .I0(\FRAME_MATCHER.i [25]), .I1(GND_net), 
            .CO(n27820));
    SB_LUT4 i1_2_lut_adj_1140 (.I0(n17652), .I1(n30900), .I2(GND_net), 
            .I3(GND_net), .O(Kp_23__N_1630));
    defparam i1_2_lut_adj_1140.LUT_INIT = 16'h9999;
    SB_LUT4 i28573_3_lut_4_lut (.I0(\data_in_frame[0] [5]), .I1(\data_in_frame[0] [4]), 
            .I2(\data_in_frame[2] [6]), .I3(n18268), .O(n35326));   // verilog/coms.v(76[16:27])
    defparam i28573_3_lut_4_lut.LUT_INIT = 16'hff96;
    SB_LUT4 i3_4_lut_adj_1141 (.I0(\data_in_frame[19] [6]), .I1(\data_in_frame[19] [1]), 
            .I2(\data_in_frame[19] [2]), .I3(\data_in_frame[19] [3]), .O(n8_adj_4153));   // verilog/coms.v(268[9:85])
    defparam i3_4_lut_adj_1141.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_1142 (.I0(\data_in_frame[19] [7]), .I1(n8_adj_4153), 
            .I2(\data_in_frame[19] [4]), .I3(\data_in_frame[19] [5]), .O(Kp_23__N_735));   // verilog/coms.v(268[9:85])
    defparam i4_4_lut_adj_1142.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1143 (.I0(n33010), .I1(n33329), .I2(GND_net), 
            .I3(GND_net), .O(n6_adj_4154));
    defparam i1_2_lut_adj_1143.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1144 (.I0(n30624), .I1(n17719), .I2(n33253), 
            .I3(n6_adj_4154), .O(n30900));
    defparam i4_4_lut_adj_1144.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1145 (.I0(\data_in_frame[18] [7]), .I1(n30106), 
            .I2(GND_net), .I3(GND_net), .O(n33054));
    defparam i1_2_lut_adj_1145.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1146 (.I0(n17811), .I1(\data_in_frame[8] [0]), 
            .I2(n18506), .I3(n6_adj_4155), .O(n33200));
    defparam i4_4_lut_adj_1146.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1147 (.I0(n30880), .I1(n33023), .I2(\data_in_frame[9] [2]), 
            .I3(GND_net), .O(n30114));
    defparam i2_3_lut_adj_1147.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1148 (.I0(n30114), .I1(\data_in_frame[14] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n33079));
    defparam i1_2_lut_adj_1148.LUT_INIT = 16'h6666;
    SB_LUT4 i2_2_lut_adj_1149 (.I0(\data_in_frame[12] [2]), .I1(n30545), 
            .I2(GND_net), .I3(GND_net), .O(n10_adj_4156));
    defparam i2_2_lut_adj_1149.LUT_INIT = 16'h6666;
    SB_LUT4 i6_4_lut_adj_1150 (.I0(n31003), .I1(n12_adj_4148), .I2(n8_adj_4043), 
            .I3(\data_in_frame[7] [7]), .O(n35280));
    defparam i6_4_lut_adj_1150.LUT_INIT = 16'hfefd;
    SB_DFF data_in_frame_0__i128 (.Q(\data_in_frame[15] [7]), .C(clk32MHz), 
           .D(n19142));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 add_43_26_lut (.I0(n2312), .I1(\FRAME_MATCHER.i [24]), .I2(GND_net), 
            .I3(n27818), .O(n2_adj_4157)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_26_lut.LUT_INIT = 16'h8228;
    SB_DFF data_in_frame_0__i129 (.Q(\data_in_frame[16] [0]), .C(clk32MHz), 
           .D(n19141));   // verilog/coms.v(127[12] 300[6])
    SB_CARRY add_43_26 (.CI(n27818), .I0(\FRAME_MATCHER.i [24]), .I1(GND_net), 
            .CO(n27819));
    SB_DFFE setpoint__i0 (.Q(setpoint[0]), .C(clk32MHz), .E(n18646), .D(n5455));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i130 (.Q(\data_in_frame[16] [1]), .C(clk32MHz), 
           .D(n19140));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i6_4_lut_adj_1151 (.I0(\data_in_frame[11] [7]), .I1(\data_in_frame[12] [1]), 
            .I2(n32923), .I3(\data_in_frame[10] [1]), .O(n14_adj_4158));
    defparam i6_4_lut_adj_1151.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut_adj_1152 (.I0(\data_in_frame[14] [3]), .I1(n14_adj_4158), 
            .I2(n10_adj_4156), .I3(n33200), .O(n34344));
    defparam i7_4_lut_adj_1152.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1153 (.I0(\data_in_frame[11] [4]), .I1(n33162), 
            .I2(n32824), .I3(n30880), .O(n30946));
    defparam i3_4_lut_adj_1153.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1154 (.I0(\data_in_frame[18] [5]), .I1(\data_in_frame[16] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_4159));
    defparam i1_2_lut_adj_1154.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1155 (.I0(\data_in_frame[16] [4]), .I1(n34344), 
            .I2(n33079), .I3(n6_adj_4159), .O(n30095));
    defparam i4_4_lut_adj_1155.LUT_INIT = 16'h9669;
    SB_DFF data_in_frame_0__i131 (.Q(\data_in_frame[16] [2]), .C(clk32MHz), 
           .D(n19139));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i28685_4_lut (.I0(\data_out_frame[6] [7]), .I1(byte_transmit_counter[0]), 
            .I2(byte_transmit_counter[2]), .I3(\data_out_frame[7] [7]), 
            .O(n35440));
    defparam i28685_4_lut.LUT_INIT = 16'hec2c;
    SB_LUT4 i28683_3_lut (.I0(\data_out_frame[4] [7]), .I1(\data_out_frame[5] [7]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n35438));
    defparam i28683_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1982151_i1_3_lut (.I0(n37877), .I1(n37751), .I2(byte_transmit_counter[2]), 
            .I3(GND_net), .O(n14_adj_4160));
    defparam i1982151_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8_4_lut_adj_1156 (.I0(\data_in_frame[9] [0]), .I1(n33108), 
            .I2(\data_in_frame[8] [2]), .I3(\data_in_frame[9] [1]), .O(n20_adj_4161));   // verilog/coms.v(72[16:41])
    defparam i8_4_lut_adj_1156.LUT_INIT = 16'h6996;
    SB_LUT4 i29792_2_lut (.I0(n37901), .I1(byte_transmit_counter[2]), .I2(GND_net), 
            .I3(GND_net), .O(n36248));
    defparam i29792_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i7_4_lut_adj_1157 (.I0(n17714), .I1(\data_in_frame[8] [3]), 
            .I2(n17827), .I3(n32749), .O(n19_adj_4162));   // verilog/coms.v(72[16:41])
    defparam i7_4_lut_adj_1157.LUT_INIT = 16'h6996;
    SB_LUT4 i9_4_lut_adj_1158 (.I0(\data_in_frame[0] [0]), .I1(\data_in_frame[8] [1]), 
            .I2(n29786), .I3(n17738), .O(n21));   // verilog/coms.v(72[16:41])
    defparam i9_4_lut_adj_1158.LUT_INIT = 16'h6996;
    SB_LUT4 i11_3_lut_adj_1159 (.I0(n21), .I1(n19_adj_4162), .I2(n20_adj_4161), 
            .I3(GND_net), .O(n30653));   // verilog/coms.v(72[16:41])
    defparam i11_3_lut_adj_1159.LUT_INIT = 16'h9696;
    SB_LUT4 i28679_4_lut (.I0(\data_out_frame[6] [6]), .I1(byte_transmit_counter[0]), 
            .I2(byte_transmit_counter[2]), .I3(\data_out_frame[7] [6]), 
            .O(n35434));
    defparam i28679_4_lut.LUT_INIT = 16'hec2c;
    SB_LUT4 i28677_3_lut (.I0(\data_out_frame[4] [6]), .I1(\data_out_frame[5] [6]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n35432));
    defparam i28677_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i18689_2_lut (.I0(\state[2] ), .I1(\state[3] ), .I2(GND_net), 
            .I3(GND_net), .O(n10));
    defparam i18689_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i1982754_i1_3_lut (.I0(n37859), .I1(n37841), .I2(byte_transmit_counter[2]), 
            .I3(GND_net), .O(n14_adj_4164));
    defparam i1982754_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3_4_lut_adj_1160 (.I0(n30596), .I1(n30876), .I2(\data_in_frame[9] [6]), 
            .I3(Kp_23__N_1175), .O(n29976));
    defparam i3_4_lut_adj_1160.LUT_INIT = 16'h6996;
    SB_LUT4 i5_4_lut_adj_1161 (.I0(n29976), .I1(n30939), .I2(\data_in_frame[4] [1]), 
            .I3(\data_in_frame[12] [0]), .O(n12_adj_4165));
    defparam i5_4_lut_adj_1161.LUT_INIT = 16'h9669;
    SB_LUT4 i6_4_lut_adj_1162 (.I0(\data_in_frame[11] [7]), .I1(n12_adj_4165), 
            .I2(n30653), .I3(\data_in_frame[13] [7]), .O(n33023));
    defparam i6_4_lut_adj_1162.LUT_INIT = 16'h6996;
    SB_LUT4 i29831_2_lut (.I0(n37907), .I1(byte_transmit_counter[2]), .I2(GND_net), 
            .I3(GND_net), .O(n36272));
    defparam i29831_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i1_2_lut_adj_1163 (.I0(\data_in_frame[11] [4]), .I1(\data_in_frame[14] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n32899));   // verilog/coms.v(74[16:43])
    defparam i1_2_lut_adj_1163.LUT_INIT = 16'h6666;
    SB_LUT4 i28672_3_lut (.I0(\data_out_frame[6] [5]), .I1(\data_out_frame[7] [5]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n35427));
    defparam i28672_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i28673_4_lut (.I0(n35427), .I1(byte_transmit_counter[1]), .I2(byte_transmit_counter[2]), 
            .I3(byte_transmit_counter[0]), .O(n35428));
    defparam i28673_4_lut.LUT_INIT = 16'ha3a0;
    SB_LUT4 i28671_3_lut (.I0(\data_out_frame[4] [5]), .I1(\data_out_frame[5] [5]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n35426));
    defparam i28671_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i5_4_lut_adj_1164 (.I0(n32899), .I1(n33023), .I2(\data_in_frame[16] [2]), 
            .I3(Kp_23__N_1204), .O(n12_adj_4166));
    defparam i5_4_lut_adj_1164.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1165 (.I0(\data_in_frame[18] [3]), .I1(n18275), 
            .I2(n12_adj_4166), .I3(n8_adj_4167), .O(n33242));
    defparam i1_4_lut_adj_1165.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_adj_1166 (.I0(\data_in_frame[3] [5]), .I1(\data_in_frame[5] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n17811));   // verilog/coms.v(78[16:27])
    defparam i1_2_lut_adj_1166.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1167 (.I0(n18440), .I1(n18460), .I2(GND_net), 
            .I3(GND_net), .O(n33145));   // verilog/coms.v(72[16:41])
    defparam i1_2_lut_adj_1167.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_1168 (.I0(\data_in_frame[3] [6]), .I1(n33114), 
            .I2(\data_in_frame[8] [1]), .I3(GND_net), .O(n32746));   // verilog/coms.v(76[16:43])
    defparam i2_3_lut_adj_1168.LUT_INIT = 16'h9696;
    SB_LUT4 i6_4_lut_adj_1169 (.I0(n18293), .I1(n5_c), .I2(n17846), .I3(n17858), 
            .O(n16_adj_4168));
    defparam i6_4_lut_adj_1169.LUT_INIT = 16'hfffe;
    SB_LUT4 i2_3_lut_adj_1170 (.I0(\data_in_frame[13] [6]), .I1(\data_in_frame[14] [0]), 
            .I2(\data_in_frame[13] [7]), .I3(GND_net), .O(n33203));   // verilog/coms.v(70[16:27])
    defparam i2_3_lut_adj_1170.LUT_INIT = 16'h9696;
    SB_LUT4 i4_4_lut_adj_1171 (.I0(n33203), .I1(\data_in_frame[13] [4]), 
            .I2(\data_in_frame[16] [1]), .I3(n33317), .O(n10_adj_4169));   // verilog/coms.v(72[16:41])
    defparam i4_4_lut_adj_1171.LUT_INIT = 16'h6996;
    SB_LUT4 i1983357_i1_3_lut (.I0(n37853), .I1(n37889), .I2(byte_transmit_counter[2]), 
            .I3(GND_net), .O(n14_adj_4170));
    defparam i1983357_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i29809_2_lut (.I0(n37913), .I1(byte_transmit_counter[2]), .I2(GND_net), 
            .I3(GND_net), .O(n36279));
    defparam i29809_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i3_4_lut_adj_1172 (.I0(n34364), .I1(\data_in_frame[11] [1]), 
            .I2(\data_in_frame[10] [7]), .I3(n30950), .O(n32759));
    defparam i3_4_lut_adj_1172.LUT_INIT = 16'h9669;
    SB_LUT4 i2_3_lut_adj_1173 (.I0(\data_in_frame[13] [2]), .I1(n30624), 
            .I2(\data_in_frame[10] [6]), .I3(GND_net), .O(n33051));
    defparam i2_3_lut_adj_1173.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_4_lut_adj_1174 (.I0(\data_in_frame[0] [5]), .I1(\data_in_frame[0] [4]), 
            .I2(\data_in_frame[3] [0]), .I3(n16400), .O(n33136));   // verilog/coms.v(76[16:27])
    defparam i2_3_lut_4_lut_adj_1174.LUT_INIT = 16'h6996;
    SB_LUT4 add_43_25_lut (.I0(n2312), .I1(\FRAME_MATCHER.i [23]), .I2(GND_net), 
            .I3(n27817), .O(n2_adj_4171)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_25_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i2_3_lut_adj_1175 (.I0(\data_in_frame[11] [3]), .I1(n17704), 
            .I2(\data_in_frame[11] [4]), .I3(GND_net), .O(n33120));   // verilog/coms.v(74[16:43])
    defparam i2_3_lut_adj_1175.LUT_INIT = 16'h9696;
    SB_LUT4 i2_2_lut_adj_1176 (.I0(n17827), .I1(n8), .I2(GND_net), .I3(GND_net), 
            .O(Kp_23__N_1195));   // verilog/coms.v(85[17:70])
    defparam i2_2_lut_adj_1176.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_1177 (.I0(n33136), .I1(n33338), .I2(n32797), 
            .I3(GND_net), .O(n17885));
    defparam i2_3_lut_adj_1177.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1178 (.I0(\data_in_frame[9] [4]), .I1(\data_in_frame[13] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n33162));
    defparam i1_2_lut_adj_1178.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1179 (.I0(\data_in_frame[15] [5]), .I1(n30880), 
            .I2(GND_net), .I3(GND_net), .O(n33347));
    defparam i1_2_lut_adj_1179.LUT_INIT = 16'h9999;
    SB_LUT4 i5_4_lut_adj_1180 (.I0(n33299), .I1(n33317), .I2(\data_in_frame[17] [7]), 
            .I3(n33268), .O(n12_adj_4172));
    defparam i5_4_lut_adj_1180.LUT_INIT = 16'h6996;
    SB_LUT4 i28666_3_lut (.I0(\data_out_frame[6] [4]), .I1(\data_out_frame[7] [4]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n35421));
    defparam i28666_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i28667_4_lut (.I0(n35421), .I1(byte_transmit_counter[1]), .I2(byte_transmit_counter[2]), 
            .I3(byte_transmit_counter[0]), .O(n35422));
    defparam i28667_4_lut.LUT_INIT = 16'haca3;
    SB_LUT4 i28665_3_lut (.I0(\data_out_frame[4] [4]), .I1(\data_out_frame[5] [4]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n35420));
    defparam i28665_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1983960_i1_3_lut (.I0(n37847), .I1(n37727), .I2(byte_transmit_counter[2]), 
            .I3(GND_net), .O(n14_adj_4173));
    defparam i1983960_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i29847_2_lut (.I0(n37919), .I1(byte_transmit_counter[2]), .I2(GND_net), 
            .I3(GND_net), .O(n36290));
    defparam i29847_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i6_4_lut_adj_1181 (.I0(\data_in_frame[10] [7]), .I1(n12_adj_4172), 
            .I2(n33347), .I3(n33159), .O(n35127));
    defparam i6_4_lut_adj_1181.LUT_INIT = 16'h6996;
    SB_LUT4 i28660_3_lut (.I0(\data_out_frame[6] [3]), .I1(\data_out_frame[7] [3]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n35415));
    defparam i28660_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i28661_4_lut (.I0(n35415), .I1(byte_transmit_counter[1]), .I2(byte_transmit_counter[2]), 
            .I3(byte_transmit_counter[0]), .O(n35416));
    defparam i28661_4_lut.LUT_INIT = 16'hafa3;
    SB_LUT4 i28659_3_lut (.I0(\data_out_frame[4] [3]), .I1(\data_out_frame[5] [3]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n35414));
    defparam i28659_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_adj_1182 (.I0(\data_in_frame[9] [0]), .I1(\data_in_frame[11] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n33344));
    defparam i1_2_lut_adj_1182.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1183 (.I0(n29786), .I1(\data_in_frame[10] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n30008));
    defparam i1_2_lut_adj_1183.LUT_INIT = 16'h6666;
    SB_LUT4 i7_4_lut_adj_1184 (.I0(n30596), .I1(n8), .I2(n35280), .I3(n18285), 
            .O(n17_adj_4174));
    defparam i7_4_lut_adj_1184.LUT_INIT = 16'hfffe;
    SB_LUT4 i1984563_i1_3_lut (.I0(n37835), .I1(n37925), .I2(byte_transmit_counter[2]), 
            .I3(GND_net), .O(n14_adj_4175));
    defparam i1984563_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_adj_1185 (.I0(\data_in_frame[11] [0]), .I1(\data_in_frame[8] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n33335));
    defparam i1_2_lut_adj_1185.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1186 (.I0(\data_in_frame[9] [4]), .I1(\data_in_frame[9] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n33184));   // verilog/coms.v(75[16:43])
    defparam i1_2_lut_adj_1186.LUT_INIT = 16'h6666;
    SB_LUT4 i29821_2_lut (.I0(n37655), .I1(byte_transmit_counter[2]), .I2(GND_net), 
            .I3(GND_net), .O(n36293));
    defparam i29821_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i1_2_lut_adj_1187 (.I0(\data_in_frame[9] [2]), .I1(\data_in_frame[9] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n32858));   // verilog/coms.v(75[16:43])
    defparam i1_2_lut_adj_1187.LUT_INIT = 16'h6666;
    SB_LUT4 i28654_3_lut (.I0(\data_out_frame[6] [2]), .I1(\data_out_frame[7] [2]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n35409));
    defparam i28654_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i28655_4_lut (.I0(n35409), .I1(byte_transmit_counter[0]), .I2(byte_transmit_counter[2]), 
            .I3(byte_transmit_counter[1]), .O(n35410));
    defparam i28655_4_lut.LUT_INIT = 16'ha0a3;
    SB_LUT4 i28653_3_lut (.I0(\data_out_frame[4] [2]), .I1(\data_out_frame[5] [2]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n35408));
    defparam i28653_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_adj_1188 (.I0(n18168), .I1(n32923), .I2(GND_net), 
            .I3(GND_net), .O(Kp_23__N_1175));   // verilog/coms.v(85[17:63])
    defparam i1_2_lut_adj_1188.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_1189 (.I0(\data_in_frame[9] [0]), .I1(n34364), 
            .I2(n18293), .I3(GND_net), .O(n30876));
    defparam i2_3_lut_adj_1189.LUT_INIT = 16'h6969;
    SB_LUT4 i2_3_lut_adj_1190 (.I0(\data_in_frame[5] [2]), .I1(\data_in_frame[3] [0]), 
            .I2(\data_in_frame[4] [1]), .I3(GND_net), .O(n33293));
    defparam i2_3_lut_adj_1190.LUT_INIT = 16'h9696;
    SB_LUT4 i1985166_i1_3_lut (.I0(n37817), .I1(n37931), .I2(byte_transmit_counter[2]), 
            .I3(GND_net), .O(n14_adj_4176));
    defparam i1985166_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i29818_2_lut (.I0(n37649), .I1(byte_transmit_counter[2]), .I2(GND_net), 
            .I3(GND_net), .O(n36298));
    defparam i29818_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i9_4_lut_adj_1191 (.I0(n17_adj_4174), .I1(n17863), .I2(n16_adj_4168), 
            .I3(n17827), .O(n31_adj_4177));
    defparam i9_4_lut_adj_1191.LUT_INIT = 16'hfffe;
    SB_LUT4 i2_3_lut_adj_1192 (.I0(n17846), .I1(n18285), .I2(\data_in_frame[9] [3]), 
            .I3(GND_net), .O(n17704));   // verilog/coms.v(74[16:43])
    defparam i2_3_lut_adj_1192.LUT_INIT = 16'h9696;
    SB_LUT4 i28645_3_lut (.I0(\data_out_frame[6] [0]), .I1(\data_out_frame[7] [0]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n35400));
    defparam i28645_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i28646_4_lut (.I0(n35400), .I1(byte_transmit_counter[1]), .I2(byte_transmit_counter[2]), 
            .I3(byte_transmit_counter[0]), .O(n35401));
    defparam i28646_4_lut.LUT_INIT = 16'ha3a0;
    SB_LUT4 i1_2_lut_adj_1193 (.I0(n30545), .I1(n17885), .I2(GND_net), 
            .I3(GND_net), .O(n30848));
    defparam i1_2_lut_adj_1193.LUT_INIT = 16'h6666;
    SB_LUT4 i28644_3_lut (.I0(\data_out_frame[4] [0]), .I1(\data_out_frame[5] [0]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n35399));
    defparam i28644_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1987578_i1_3_lut (.I0(n37871), .I1(n37865), .I2(byte_transmit_counter[2]), 
            .I3(GND_net), .O(n14_adj_4178));
    defparam i1987578_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3_4_lut_adj_1194 (.I0(n17858), .I1(n32746), .I2(\data_in_frame[6] [0]), 
            .I3(n17738), .O(n15914));   // verilog/coms.v(76[16:43])
    defparam i3_4_lut_adj_1194.LUT_INIT = 16'h6996;
    SB_LUT4 i29811_2_lut (.I0(n37721), .I1(byte_transmit_counter[2]), .I2(GND_net), 
            .I3(GND_net), .O(n36304));
    defparam i29811_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i1_2_lut_adj_1195 (.I0(n18293), .I1(n15914), .I2(GND_net), 
            .I3(GND_net), .O(n33040));
    defparam i1_2_lut_adj_1195.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1196 (.I0(n17827), .I1(n17846), .I2(GND_net), 
            .I3(GND_net), .O(Kp_23__N_1204));   // verilog/coms.v(72[16:41])
    defparam i1_2_lut_adj_1196.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_4_lut_adj_1197 (.I0(n33212), .I1(n4_adj_4179), .I2(\data_in_frame[1] [5]), 
            .I3(\data_in_frame[7] [7]), .O(n17738));
    defparam i2_3_lut_4_lut_adj_1197.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_1198 (.I0(n33108), .I1(n17101), .I2(Kp_23__N_1204), 
            .I3(n33040), .O(n15_adj_4180));
    defparam i6_4_lut_adj_1198.LUT_INIT = 16'h6996;
    SB_LUT4 i8_4_lut_adj_1199 (.I0(n15_adj_4180), .I1(n30848), .I2(n14_adj_4181), 
            .I3(n17863), .O(n34364));
    defparam i8_4_lut_adj_1199.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_1200 (.I0(n34364), .I1(\data_in_frame[11] [1]), 
            .I2(\data_in_frame[13] [3]), .I3(n30950), .O(n10_adj_4182));
    defparam i4_4_lut_adj_1200.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut (.I0(n33212), .I1(n4_adj_4179), .I2(n30939), 
            .I3(GND_net), .O(n31003));
    defparam i1_2_lut_3_lut.LUT_INIT = 16'h9696;
    SB_CARRY add_43_25 (.CI(n27817), .I0(\FRAME_MATCHER.i [23]), .I1(GND_net), 
            .CO(n27818));
    SB_LUT4 i2_3_lut_4_lut_adj_1201 (.I0(n17652), .I1(n32873), .I2(\data_in_frame[19] [7]), 
            .I3(n30946), .O(n34498));
    defparam i2_3_lut_4_lut_adj_1201.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1202 (.I0(Kp_23__N_1069), .I1(\data_in_frame[8] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n17730));   // verilog/coms.v(71[16:27])
    defparam i1_2_lut_adj_1202.LUT_INIT = 16'h6666;
    SB_LUT4 i6_4_lut_adj_1203 (.I0(n17730), .I1(Kp_23__N_1063), .I2(n33268), 
            .I3(n17595), .O(n14_adj_4183));
    defparam i6_4_lut_adj_1203.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut_adj_1204 (.I0(\data_in_frame[15] [4]), .I1(n14_adj_4183), 
            .I2(n10_adj_4184), .I3(n33335), .O(n30089));
    defparam i7_4_lut_adj_1204.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1205 (.I0(\data_in_frame[11] [3]), .I1(n33159), 
            .I2(n18460), .I3(GND_net), .O(n17901));   // verilog/coms.v(73[16:42])
    defparam i2_3_lut_adj_1205.LUT_INIT = 16'h9696;
    SB_LUT4 data_in_frame_17__7__I_0_3899_2_lut (.I0(\data_in_frame[17] [7]), 
            .I1(\data_in_frame[17] [6]), .I2(GND_net), .I3(GND_net), .O(Kp_23__N_1372));   // verilog/coms.v(70[16:27])
    defparam data_in_frame_17__7__I_0_3899_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i5_4_lut_adj_1206 (.I0(Kp_23__N_1372), .I1(n17901), .I2(\data_in_frame[18] [0]), 
            .I3(n30089), .O(n12_adj_4185));
    defparam i5_4_lut_adj_1206.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_1207 (.I0(\data_in_frame[15] [6]), .I1(n12_adj_4185), 
            .I2(n18275), .I3(n35127), .O(n32905));
    defparam i6_4_lut_adj_1207.LUT_INIT = 16'h9669;
    SB_LUT4 i4_4_lut_adj_1208 (.I0(n32791), .I1(n18264), .I2(\data_in_frame[7] [0]), 
            .I3(n33127), .O(n10_adj_4186));   // verilog/coms.v(74[16:43])
    defparam i4_4_lut_adj_1208.LUT_INIT = 16'h6996;
    SB_LUT4 i5_3_lut_adj_1209 (.I0(\data_in_frame[6] [6]), .I1(n10_adj_4186), 
            .I2(\data_in_frame[6] [7]), .I3(GND_net), .O(n17827));   // verilog/coms.v(74[16:43])
    defparam i5_3_lut_adj_1209.LUT_INIT = 16'h9696;
    SB_LUT4 i6_4_lut_adj_1210 (.I0(n33114), .I1(\data_in_frame[4] [1]), 
            .I2(\data_in_frame[1] [7]), .I3(\data_in_frame[8] [3]), .O(n14_adj_4187));   // verilog/coms.v(75[16:27])
    defparam i6_4_lut_adj_1210.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_1211 (.I0(n17652), .I1(n32873), .I2(n30666), 
            .I3(n30946), .O(n30853));
    defparam i2_3_lut_4_lut_adj_1211.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_adj_1212 (.I0(\data_in_frame[5] [4]), .I1(n33057), 
            .I2(GND_net), .I3(GND_net), .O(n33271));
    defparam i1_2_lut_adj_1212.LUT_INIT = 16'h6666;
    SB_LUT4 i7_4_lut_adj_1213 (.I0(\data_in_frame[6] [1]), .I1(n14_adj_4187), 
            .I2(n10_adj_4188), .I3(\data_in_frame[3] [7]), .O(n17863));   // verilog/coms.v(75[16:27])
    defparam i7_4_lut_adj_1213.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1214 (.I0(\data_in_frame[20] [2]), .I1(n32905), 
            .I2(\data_in_frame[18] [1]), .I3(GND_net), .O(n33708));
    defparam i2_3_lut_adj_1214.LUT_INIT = 16'h9696;
    SB_LUT4 i5_4_lut_adj_1215 (.I0(n32791), .I1(n33136), .I2(\data_in_frame[7] [2]), 
            .I3(\data_in_frame[2] [6]), .O(n12_adj_4189));
    defparam i5_4_lut_adj_1215.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_1216 (.I0(\data_in_frame[5] [1]), .I1(n12_adj_4189), 
            .I2(n18058), .I3(\data_in_frame[5] [0]), .O(n18285));
    defparam i6_4_lut_adj_1216.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1217 (.I0(\data_in_frame[6] [6]), .I1(\data_in_frame[8] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_4190));   // verilog/coms.v(75[16:43])
    defparam i1_2_lut_adj_1217.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1218 (.I0(n17843), .I1(n33127), .I2(n32784), 
            .I3(n6_adj_4190), .O(n8));   // verilog/coms.v(75[16:43])
    defparam i4_4_lut_adj_1218.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_1219 (.I0(n33142), .I1(\data_in_frame[3] [3]), 
            .I2(\data_in_frame[7] [5]), .I3(n27_adj_4191), .O(n10_adj_4192));
    defparam i4_4_lut_adj_1219.LUT_INIT = 16'h6996;
    SB_LUT4 i5_3_lut_adj_1220 (.I0(\data_in_frame[3] [1]), .I1(n10_adj_4192), 
            .I2(\data_in_frame[5] [4]), .I3(GND_net), .O(n30596));
    defparam i5_3_lut_adj_1220.LUT_INIT = 16'h9696;
    SB_LUT4 add_43_24_lut (.I0(n2312), .I1(\FRAME_MATCHER.i [22]), .I2(GND_net), 
            .I3(n27816), .O(n2_adj_4193)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_24_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i2_3_lut_adj_1221 (.I0(\data_in_frame[6] [3]), .I1(\data_in_frame[2] [1]), 
            .I2(\data_in_frame[3] [7]), .I3(GND_net), .O(n32749));   // verilog/coms.v(72[16:41])
    defparam i2_3_lut_adj_1221.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1222 (.I0(\data_in_frame[3] [6]), .I1(\data_in_frame[6] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n32756));   // verilog/coms.v(75[16:27])
    defparam i1_2_lut_adj_1222.LUT_INIT = 16'h6666;
    SB_CARRY add_43_24 (.CI(n27816), .I0(\FRAME_MATCHER.i [22]), .I1(GND_net), 
            .CO(n27817));
    SB_LUT4 i4_4_lut_adj_1223 (.I0(\data_in_frame[6] [6]), .I1(\data_in_frame[6] [1]), 
            .I2(\data_in_frame[6] [3]), .I3(\data_in_frame[6] [4]), .O(n10_adj_4194));   // verilog/coms.v(85[17:28])
    defparam i4_4_lut_adj_1223.LUT_INIT = 16'h6996;
    SB_LUT4 add_43_23_lut (.I0(n2312), .I1(\FRAME_MATCHER.i [21]), .I2(GND_net), 
            .I3(n27815), .O(n2_adj_4195)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_23_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_43_23 (.CI(n27815), .I0(\FRAME_MATCHER.i [21]), .I1(GND_net), 
            .CO(n27816));
    SB_DFF data_in_frame_0__i132 (.Q(\data_in_frame[16] [3]), .C(clk32MHz), 
           .D(n19138));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i133 (.Q(\data_in_frame[16] [4]), .C(clk32MHz), 
           .D(n19137));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i1_3_lut_adj_1224 (.I0(\data_in_frame[19] [4]), .I1(\data_in_frame[21] [6]), 
            .I2(\data_in_frame[19] [5]), .I3(GND_net), .O(n5_adj_4196));
    defparam i1_3_lut_adj_1224.LUT_INIT = 16'h9696;
    SB_LUT4 add_43_22_lut (.I0(n2312), .I1(\FRAME_MATCHER.i [20]), .I2(GND_net), 
            .I3(n27814), .O(n2_adj_4197)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_22_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i28649_4_lut (.I0(\data_out_frame[6] [1]), .I1(byte_transmit_counter[0]), 
            .I2(byte_transmit_counter[2]), .I3(\data_out_frame[7] [1]), 
            .O(n35404));
    defparam i28649_4_lut.LUT_INIT = 16'hec2c;
    SB_LUT4 i28647_3_lut (.I0(\data_out_frame[4] [1]), .I1(\data_out_frame[5] [1]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n35402));
    defparam i28647_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2_2_lut_adj_1225 (.I0(\data_in_frame[20] [3]), .I1(n15965), 
            .I2(GND_net), .I3(GND_net), .O(n7_adj_4198));
    defparam i2_2_lut_adj_1225.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1226 (.I0(n7_adj_4198), .I1(\data_in_frame[18] [1]), 
            .I2(n35127), .I3(\data_in_frame[18] [2]), .O(n34273));
    defparam i4_4_lut_adj_1226.LUT_INIT = 16'h9669;
    SB_LUT4 i1985769_i1_3_lut (.I0(n37805), .I1(n37799), .I2(byte_transmit_counter[2]), 
            .I3(GND_net), .O(n14_adj_4199));
    defparam i1985769_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2_4_lut_adj_1227 (.I0(n15965), .I1(\data_in_frame[18] [2]), 
            .I2(\data_in_frame[20] [4]), .I3(n33242), .O(n33707));
    defparam i2_4_lut_adj_1227.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1228 (.I0(\data_in_frame[19] [3]), .I1(\data_in_frame[19] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_4200));
    defparam i1_2_lut_adj_1228.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_1229 (.I0(n30095), .I1(\data_in_frame[20] [7]), 
            .I2(\data_in_frame[19] [0]), .I3(n30946), .O(n35054));
    defparam i3_4_lut_adj_1229.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1230 (.I0(n30853), .I1(n33054), .I2(n32702), 
            .I3(\data_in_frame[21] [1]), .O(n34290));
    defparam i3_4_lut_adj_1230.LUT_INIT = 16'h9669;
    SB_LUT4 i3_4_lut_adj_1231 (.I0(n32873), .I1(n30666), .I2(n35054), 
            .I3(Kp_23__N_735), .O(n34316));
    defparam i3_4_lut_adj_1231.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_1232 (.I0(\data_in_frame[21] [5]), .I1(n35067), 
            .I2(n18312), .I3(n6_adj_4200), .O(n34619));
    defparam i4_4_lut_adj_1232.LUT_INIT = 16'h9669;
    SB_LUT4 i29814_2_lut (.I0(n37661), .I1(byte_transmit_counter[2]), .I2(GND_net), 
            .I3(GND_net), .O(n36301));
    defparam i29814_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i2_3_lut_4_lut_adj_1233 (.I0(\data_out_frame[17] [1]), .I1(n33228), 
            .I2(\data_out_frame[19] [3]), .I3(n32963), .O(n18330));
    defparam i2_3_lut_4_lut_adj_1233.LUT_INIT = 16'h9669;
    SB_CARRY add_43_22 (.CI(n27814), .I0(\FRAME_MATCHER.i [20]), .I1(GND_net), 
            .CO(n27815));
    SB_LUT4 add_43_21_lut (.I0(n2312), .I1(\FRAME_MATCHER.i [19]), .I2(GND_net), 
            .I3(n27813), .O(n2_adj_4201)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_21_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i2_3_lut_adj_1234 (.I0(n30095), .I1(n32978), .I2(\data_in_frame[20] [6]), 
            .I3(GND_net), .O(n33768));
    defparam i2_3_lut_adj_1234.LUT_INIT = 16'h9696;
    SB_LUT4 i5_3_lut_adj_1235 (.I0(\data_in_frame[6] [2]), .I1(n10_adj_4194), 
            .I2(\data_in_frame[6] [5]), .I3(GND_net), .O(n32773));   // verilog/coms.v(85[17:28])
    defparam i5_3_lut_adj_1235.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1236 (.I0(\data_in_frame[20] [0]), .I1(n32905), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_4202));
    defparam i1_2_lut_adj_1236.LUT_INIT = 16'h6666;
    SB_LUT4 i1_rep_67_2_lut (.I0(\data_in_frame[19] [2]), .I1(\data_in_frame[19] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n38349));   // verilog/coms.v(268[9:85])
    defparam i1_rep_67_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_43_21 (.CI(n27813), .I0(\FRAME_MATCHER.i [19]), .I1(GND_net), 
            .CO(n27814));
    SB_LUT4 add_43_20_lut (.I0(n2312), .I1(\FRAME_MATCHER.i [18]), .I2(GND_net), 
            .I3(n27812), .O(n2_adj_4203)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_20_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i4_4_lut_adj_1237 (.I0(\data_in_frame[19] [1]), .I1(\data_in_frame[19] [2]), 
            .I2(\data_in_frame[21] [3]), .I3(n33054), .O(n10_adj_4204));
    defparam i4_4_lut_adj_1237.LUT_INIT = 16'h6996;
    SB_DFFSS \FRAME_MATCHER.state_i31  (.Q(\FRAME_MATCHER.state_c [31]), .C(clk32MHz), 
            .D(n32227), .S(n32063));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i30  (.Q(\FRAME_MATCHER.state_c [30]), .C(clk32MHz), 
            .D(n32225), .S(n32067));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i29  (.Q(\FRAME_MATCHER.state_c [29]), .C(clk32MHz), 
            .D(n32223), .S(n32071));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i28  (.Q(\FRAME_MATCHER.state_c [28]), .C(clk32MHz), 
            .D(n32221), .S(n32075));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i27  (.Q(\FRAME_MATCHER.state_c [27]), .C(clk32MHz), 
            .D(n32219), .S(n32079));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i26  (.Q(\FRAME_MATCHER.state_c [26]), .C(clk32MHz), 
            .D(n32217), .S(n32083));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i25  (.Q(\FRAME_MATCHER.state_c [25]), .C(clk32MHz), 
            .D(n32215), .S(n32005));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i24  (.Q(\FRAME_MATCHER.state_c [24]), .C(clk32MHz), 
            .D(n32213), .S(n32087));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i23  (.Q(\FRAME_MATCHER.state_c [23]), .C(clk32MHz), 
            .D(n32211), .S(n32091));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i22  (.Q(\FRAME_MATCHER.state_c [22]), .C(clk32MHz), 
            .D(n32209), .S(n32095));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i21  (.Q(\FRAME_MATCHER.state_c [21]), .C(clk32MHz), 
            .D(n32207), .S(n32099));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i20  (.Q(\FRAME_MATCHER.state_c [20]), .C(clk32MHz), 
            .D(n32205), .S(n32027));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i19  (.Q(\FRAME_MATCHER.state_c [19]), .C(clk32MHz), 
            .D(n32203), .S(n32103));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i18  (.Q(\FRAME_MATCHER.state_c [18]), .C(clk32MHz), 
            .D(n32201), .S(n32107));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i17  (.Q(\FRAME_MATCHER.state_c [17]), .C(clk32MHz), 
            .D(n32199), .S(n32111));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i16  (.Q(\FRAME_MATCHER.state_c [16]), .C(clk32MHz), 
            .D(n32197), .S(n32115));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i15  (.Q(\FRAME_MATCHER.state_c [15]), .C(clk32MHz), 
            .D(n32195), .S(n32119));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i14  (.Q(\FRAME_MATCHER.state_c [14]), .C(clk32MHz), 
            .D(n23755), .S(n24510));   // verilog/coms.v(127[12] 300[6])
    SB_CARRY add_43_20 (.CI(n27812), .I0(\FRAME_MATCHER.i [18]), .I1(GND_net), 
            .CO(n27813));
    SB_DFFSS \FRAME_MATCHER.state_i13  (.Q(\FRAME_MATCHER.state_c [13]), .C(clk32MHz), 
            .D(n23753), .S(n24508));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i12  (.Q(\FRAME_MATCHER.state_c [12]), .C(clk32MHz), 
            .D(n7_adj_4205), .S(n31999));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i11  (.Q(\FRAME_MATCHER.state_c [11]), .C(clk32MHz), 
            .D(n32233), .S(n32041));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i10  (.Q(\FRAME_MATCHER.state_c [10]), .C(clk32MHz), 
            .D(n32193), .S(n32123));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i9  (.Q(\FRAME_MATCHER.state_c [9]), .C(clk32MHz), 
            .D(n32191), .S(n32127));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i8  (.Q(\FRAME_MATCHER.state_c [8]), .C(clk32MHz), 
            .D(n32145), .S(n24506));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i7  (.Q(\FRAME_MATCHER.state_c [7]), .C(clk32MHz), 
            .D(n32189), .S(n32131));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i6  (.Q(\FRAME_MATCHER.state_c [6]), .C(clk32MHz), 
            .D(n32185), .S(n32135));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i5  (.Q(\FRAME_MATCHER.state_c [5]), .C(clk32MHz), 
            .D(n32181), .S(n32139));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i4  (.Q(\FRAME_MATCHER.state_c [4]), .C(clk32MHz), 
            .D(n32177), .S(n32021));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i3  (.Q(\FRAME_MATCHER.state [3]), .C(clk32MHz), 
            .D(n32017), .S(n32231));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE data_out_frame_0___i224 (.Q(\data_out_frame[27] [7]), .C(clk32MHz), 
            .E(n18682), .D(n32713));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 add_43_19_lut (.I0(n2312), .I1(\FRAME_MATCHER.i [17]), .I2(GND_net), 
            .I3(n27811), .O(n2_adj_4206)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_19_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i1_2_lut_adj_1238 (.I0(\data_in_frame[6] [0]), .I1(n30031), 
            .I2(GND_net), .I3(GND_net), .O(n32966));
    defparam i1_2_lut_adj_1238.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_1239 (.I0(n38349), .I1(n34447), .I2(\data_in_frame[21] [4]), 
            .I3(n30093), .O(n35169));
    defparam i3_4_lut_adj_1239.LUT_INIT = 16'h9669;
    SB_LUT4 i4_4_lut_adj_1240 (.I0(\data_in_frame[19] [6]), .I1(n34498), 
            .I2(Kp_23__N_1630), .I3(n6_adj_4202), .O(n34941));
    defparam i4_4_lut_adj_1240.LUT_INIT = 16'h9669;
    SB_LUT4 i8_4_lut_adj_1241 (.I0(n5_adj_4196), .I1(n33708), .I2(n30900), 
            .I3(n34447), .O(n24));
    defparam i8_4_lut_adj_1241.LUT_INIT = 16'h7bb7;
    SB_LUT4 i6_4_lut_adj_1242 (.I0(n34273), .I1(\data_in_frame[19] [1]), 
            .I2(\data_in_frame[21] [2]), .I3(n33879), .O(n22_adj_4207));
    defparam i6_4_lut_adj_1242.LUT_INIT = 16'h7dd7;
    SB_LUT4 i7_4_lut_adj_1243 (.I0(n35067), .I1(n35169), .I2(n10_adj_4204), 
            .I3(n30093), .O(n23_adj_4208));
    defparam i7_4_lut_adj_1243.LUT_INIT = 16'hdeed;
    SB_LUT4 i5_4_lut_adj_1244 (.I0(n34941), .I1(\data_in_frame[20] [1]), 
            .I2(n35127), .I3(n34498), .O(n21_adj_4209));
    defparam i5_4_lut_adj_1244.LUT_INIT = 16'hbeeb;
    SB_LUT4 i3_3_lut_adj_1245 (.I0(n17652), .I1(\data_in_frame[19] [6]), 
            .I2(\data_in_frame[19] [5]), .I3(GND_net), .O(n8_adj_4210));
    defparam i3_3_lut_adj_1245.LUT_INIT = 16'h9696;
    SB_LUT4 i3_4_lut_adj_1246 (.I0(n30853), .I1(n32702), .I2(n33879), 
            .I3(\data_in_frame[21] [0]), .O(n33979));
    defparam i3_4_lut_adj_1246.LUT_INIT = 16'h9669;
    SB_DFFE data_out_frame_0___i223 (.Q(\data_out_frame[27] [6]), .C(clk32MHz), 
            .E(n18682), .D(n33249));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE data_out_frame_0___i222 (.Q(\data_out_frame[27] [5]), .C(clk32MHz), 
            .E(n18682), .D(n33251));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE data_out_frame_0___i221 (.Q(\data_out_frame[27] [4]), .C(clk32MHz), 
            .E(n18682), .D(n32988));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE data_out_frame_0___i220 (.Q(\data_out_frame[27] [3]), .C(clk32MHz), 
            .E(n18682), .D(n34371));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE data_out_frame_0___i219 (.Q(\data_out_frame[27] [2]), .C(clk32MHz), 
            .E(n18682), .D(n34449));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE data_out_frame_0___i218 (.Q(\data_out_frame[27] [1]), .C(clk32MHz), 
            .E(n18682), .D(n30823));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE data_out_frame_0___i217 (.Q(\data_out_frame[27] [0]), .C(clk32MHz), 
            .E(n18682), .D(n33890));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE data_out_frame_0___i216 (.Q(\data_out_frame[26] [7]), .C(clk32MHz), 
            .E(n18682), .D(n34865));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE data_out_frame_0___i215 (.Q(\data_out_frame[26] [6]), .C(clk32MHz), 
            .E(n18682), .D(n32982));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE data_out_frame_0___i214 (.Q(\data_out_frame[26] [5]), .C(clk32MHz), 
            .E(n18682), .D(n33700));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE data_out_frame_0___i213 (.Q(\data_out_frame[26] [4]), .C(clk32MHz), 
            .E(n18682), .D(n33784));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE data_out_frame_0___i212 (.Q(\data_out_frame[26] [3]), .C(clk32MHz), 
            .E(n18682), .D(n32947));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE data_out_frame_0___i211 (.Q(\data_out_frame[26] [2]), .C(clk32MHz), 
            .E(n18682), .D(n33752));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE data_out_frame_0___i210 (.Q(\data_out_frame[26] [1]), .C(clk32MHz), 
            .E(n18682), .D(n34391));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE data_out_frame_0___i209 (.Q(\data_out_frame[26] [0]), .C(clk32MHz), 
            .E(n18682), .D(n34053));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i2_4_lut_adj_1247 (.I0(n33707), .I1(n32978), .I2(n33242), 
            .I3(\data_in_frame[20] [5]), .O(n18_adj_4211));
    defparam i2_4_lut_adj_1247.LUT_INIT = 16'hbeeb;
    SB_LUT4 i1387_2_lut_3_lut (.I0(n31_adj_4177), .I1(n14993), .I2(\FRAME_MATCHER.state_c [1]), 
            .I3(GND_net), .O(n5454));
    defparam i1387_2_lut_3_lut.LUT_INIT = 16'h1010;
    SB_DFFSS \FRAME_MATCHER.i_i31  (.Q(\FRAME_MATCHER.i [31]), .C(clk32MHz), 
            .D(n2_adj_4212), .S(n3_adj_4213));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 equal_442_i3_2_lut_3_lut (.I0(n31_adj_4177), .I1(n14993), .I2(n63_adj_4087), 
            .I3(GND_net), .O(n3));
    defparam equal_442_i3_2_lut_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i1_2_lut_adj_1248 (.I0(\data_in_frame[1] [2]), .I1(\data_in_frame[3] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n32894));
    defparam i1_2_lut_adj_1248.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_1249 (.I0(Kp_23__N_894), .I1(n32966), .I2(\data_in_frame[4] [5]), 
            .I3(Kp_23__N_804), .O(n30939));
    defparam i3_4_lut_adj_1249.LUT_INIT = 16'h6996;
    SB_LUT4 add_3971_9_lut (.I0(GND_net), .I1(byte_transmit_counter[7]), 
            .I2(GND_net), .I3(n27854), .O(n8825[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3971_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i10_4_lut_adj_1250 (.I0(n33768), .I1(n34619), .I2(n34316), 
            .I3(n34290), .O(n26_adj_4215));
    defparam i10_4_lut_adj_1250.LUT_INIT = 16'hffbf;
    SB_CARRY add_43_19 (.CI(n27811), .I0(\FRAME_MATCHER.i [17]), .I1(GND_net), 
            .CO(n27812));
    SB_LUT4 add_3971_8_lut (.I0(GND_net), .I1(byte_transmit_counter[6]), 
            .I2(GND_net), .I3(n27853), .O(n8825[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3971_8_lut.LUT_INIT = 16'hC33C;
    SB_DFFSS \FRAME_MATCHER.i_i30  (.Q(\FRAME_MATCHER.i [30]), .C(clk32MHz), 
            .D(n2_adj_4216), .S(n3_adj_4217));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i29  (.Q(\FRAME_MATCHER.i [29]), .C(clk32MHz), 
            .D(n2_adj_4218), .S(n3_adj_4219));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i28  (.Q(\FRAME_MATCHER.i [28]), .C(clk32MHz), 
            .D(n2_adj_4220), .S(n3_adj_4221));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i27  (.Q(\FRAME_MATCHER.i [27]), .C(clk32MHz), 
            .D(n2_adj_4222), .S(n3_adj_4223));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i26  (.Q(\FRAME_MATCHER.i [26]), .C(clk32MHz), 
            .D(n2), .S(n3_adj_4224));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i25  (.Q(\FRAME_MATCHER.i [25]), .C(clk32MHz), 
            .D(n2_adj_4115), .S(n3_adj_4225));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i4_4_lut_adj_1251 (.I0(\data_in_frame[5] [6]), .I1(n30939), 
            .I2(\data_in_frame[3] [5]), .I3(n6_adj_4226), .O(n17101));
    defparam i4_4_lut_adj_1251.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_adj_1252 (.I0(\data_in_frame[5] [2]), .I1(\data_in_frame[2] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n32797));   // verilog/coms.v(85[17:70])
    defparam i1_2_lut_adj_1252.LUT_INIT = 16'h6666;
    SB_LUT4 i6_4_lut_adj_1253 (.I0(\data_in_frame[7] [3]), .I1(Kp_23__N_862), 
            .I2(\data_in_frame[0] [7]), .I3(n18058), .O(n14_adj_4227));   // verilog/coms.v(71[16:69])
    defparam i6_4_lut_adj_1253.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut_adj_1254 (.I0(n32797), .I1(n14_adj_4227), .I2(n10_adj_4228), 
            .I3(n17784), .O(n30545));   // verilog/coms.v(71[16:69])
    defparam i7_4_lut_adj_1254.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1255 (.I0(\data_in_frame[7] [6]), .I1(n32781), 
            .I2(GND_net), .I3(GND_net), .O(n17894));
    defparam i1_2_lut_adj_1255.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1256 (.I0(\data_in_frame[8] [0]), .I1(n17101), 
            .I2(GND_net), .I3(GND_net), .O(n17983));
    defparam i1_2_lut_adj_1256.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1257 (.I0(\data_in_frame[1] [7]), .I1(\data_in_frame[0] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n32813));   // verilog/coms.v(70[16:69])
    defparam i1_2_lut_adj_1257.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1258 (.I0(\data_in_frame[6] [4]), .I1(\data_in_frame[4] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n33111));   // verilog/coms.v(73[16:42])
    defparam i1_2_lut_adj_1258.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_1259 (.I0(\data_in_frame[6] [5]), .I1(n32813), 
            .I2(n17749), .I3(n18235), .O(n17843));   // verilog/coms.v(74[16:43])
    defparam i3_4_lut_adj_1259.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1260 (.I0(n17843), .I1(n33111), .I2(n32934), 
            .I3(n17714), .O(Kp_23__N_1069));   // verilog/coms.v(73[16:42])
    defparam i3_4_lut_adj_1260.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1261 (.I0(\data_in_frame[0] [2]), .I1(\data_in_frame[0] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n32710));   // verilog/coms.v(166[9:87])
    defparam i1_2_lut_adj_1261.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1262 (.I0(\data_in_frame[0] [6]), .I1(\data_in_frame[0] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n33066));   // verilog/coms.v(77[16:27])
    defparam i1_2_lut_adj_1262.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1263 (.I0(\data_in_frame[0] [4]), .I1(\data_in_frame[0] [7]), 
            .I2(n32710), .I3(n6_adj_4229), .O(Kp_23__N_843));   // verilog/coms.v(70[16:27])
    defparam i4_4_lut_adj_1263.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1264 (.I0(\data_in_frame[2] [0]), .I1(n4_adj_4116), 
            .I2(GND_net), .I3(GND_net), .O(n32934));   // verilog/coms.v(73[16:42])
    defparam i1_2_lut_adj_1264.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1265 (.I0(\data_in_frame[2] [1]), .I1(n18264), 
            .I2(GND_net), .I3(GND_net), .O(n17749));   // verilog/coms.v(74[16:43])
    defparam i1_2_lut_adj_1265.LUT_INIT = 16'h6666;
    SB_LUT4 i14_4_lut_adj_1266 (.I0(n21_adj_4209), .I1(n23_adj_4208), .I2(n22_adj_4207), 
            .I3(n24), .O(n30_adj_4230));
    defparam i14_4_lut_adj_1266.LUT_INIT = 16'hfffe;
    SB_DFFSS \FRAME_MATCHER.i_i24  (.Q(\FRAME_MATCHER.i [24]), .C(clk32MHz), 
            .D(n2_adj_4157), .S(n3_adj_4231));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 add_43_18_lut (.I0(n2312), .I1(\FRAME_MATCHER.i [16]), .I2(GND_net), 
            .I3(n27810), .O(n2_adj_4232)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_18_lut.LUT_INIT = 16'h8228;
    SB_DFFSS \FRAME_MATCHER.i_i23  (.Q(\FRAME_MATCHER.i [23]), .C(clk32MHz), 
            .D(n2_adj_4171), .S(n3_adj_4233));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i22  (.Q(\FRAME_MATCHER.i [22]), .C(clk32MHz), 
            .D(n2_adj_4193), .S(n3_adj_4234));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i21  (.Q(\FRAME_MATCHER.i [21]), .C(clk32MHz), 
            .D(n2_adj_4195), .S(n3_adj_4235));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i1_4_lut_adj_1267 (.I0(n33979), .I1(\data_in_frame[21] [7]), 
            .I2(n8_adj_4210), .I3(n18312), .O(n17_adj_4236));
    defparam i1_4_lut_adj_1267.LUT_INIT = 16'hd77d;
    SB_DFFSS \FRAME_MATCHER.i_i20  (.Q(\FRAME_MATCHER.i [20]), .C(clk32MHz), 
            .D(n2_adj_4197), .S(n3_adj_4237));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i19  (.Q(\FRAME_MATCHER.i [19]), .C(clk32MHz), 
            .D(n2_adj_4201), .S(n3_adj_4238));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i18  (.Q(\FRAME_MATCHER.i [18]), .C(clk32MHz), 
            .D(n2_adj_4203), .S(n3_adj_4239));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i17  (.Q(\FRAME_MATCHER.i [17]), .C(clk32MHz), 
            .D(n2_adj_4206), .S(n3_adj_4240));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i15_4_lut_adj_1268 (.I0(n17_adj_4236), .I1(n30_adj_4230), .I2(n26_adj_4215), 
            .I3(n18_adj_4211), .O(n31));
    defparam i15_4_lut_adj_1268.LUT_INIT = 16'hfffe;
    SB_DFFSS \FRAME_MATCHER.i_i16  (.Q(\FRAME_MATCHER.i [16]), .C(clk32MHz), 
            .D(n2_adj_4232), .S(n3_adj_4241));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i15  (.Q(\FRAME_MATCHER.i [15]), .C(clk32MHz), 
            .D(n2_adj_4242), .S(n3_adj_4243));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i14  (.Q(\FRAME_MATCHER.i [14]), .C(clk32MHz), 
            .D(n2_adj_4244), .S(n3_adj_4245));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i13  (.Q(\FRAME_MATCHER.i [13]), .C(clk32MHz), 
            .D(n2_adj_4246), .S(n3_adj_4247));   // verilog/coms.v(127[12] 300[6])
    SB_CARRY add_3971_8 (.CI(n27853), .I0(byte_transmit_counter[6]), .I1(GND_net), 
            .CO(n27854));
    SB_DFFSS \FRAME_MATCHER.i_i12  (.Q(\FRAME_MATCHER.i [12]), .C(clk32MHz), 
            .D(n2_adj_4248), .S(n3_adj_4249));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i11  (.Q(\FRAME_MATCHER.i [11]), .C(clk32MHz), 
            .D(n2_adj_4250), .S(n3_adj_4251));   // verilog/coms.v(127[12] 300[6])
    SB_CARRY add_43_18 (.CI(n27810), .I0(\FRAME_MATCHER.i [16]), .I1(GND_net), 
            .CO(n27811));
    SB_DFFSS \FRAME_MATCHER.i_i10  (.Q(\FRAME_MATCHER.i [10]), .C(clk32MHz), 
            .D(n2_adj_4252), .S(n3_adj_4253));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i9  (.Q(\FRAME_MATCHER.i [9]), .C(clk32MHz), 
            .D(n2_adj_4254), .S(n3_adj_4255));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 add_3971_7_lut (.I0(GND_net), .I1(byte_transmit_counter[5]), 
            .I2(GND_net), .I3(n27852), .O(n8825[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3971_7_lut.LUT_INIT = 16'hC33C;
    SB_DFFSS \FRAME_MATCHER.i_i8  (.Q(\FRAME_MATCHER.i [8]), .C(clk32MHz), 
            .D(n2_adj_4256), .S(n3_adj_4257));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i7  (.Q(\FRAME_MATCHER.i [7]), .C(clk32MHz), 
            .D(n2_adj_4258), .S(n3_adj_4259));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i6  (.Q(\FRAME_MATCHER.i [6]), .C(clk32MHz), 
            .D(n2_adj_4260), .S(n3_adj_4261));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i5  (.Q(\FRAME_MATCHER.i [5]), .C(clk32MHz), 
            .D(n2_adj_4262), .S(n3_adj_4263));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i4  (.Q(\FRAME_MATCHER.i [4]), .C(clk32MHz), 
            .D(n2_adj_4264), .S(n3_adj_4265));   // verilog/coms.v(127[12] 300[6])
    SB_CARRY add_3971_7 (.CI(n27852), .I0(byte_transmit_counter[5]), .I1(GND_net), 
            .CO(n27853));
    SB_DFFSS \FRAME_MATCHER.i_i3  (.Q(\FRAME_MATCHER.i [3]), .C(clk32MHz), 
            .D(n2_adj_4266), .S(n3_adj_4267));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i2  (.Q(\FRAME_MATCHER.i [2]), .C(clk32MHz), 
            .D(n2_adj_4268), .S(n3_adj_4269));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i1  (.Q(\FRAME_MATCHER.i [1]), .C(clk32MHz), 
            .D(n2_adj_4270), .S(n3_adj_4271));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 add_3971_6_lut (.I0(GND_net), .I1(byte_transmit_counter[4]), 
            .I2(GND_net), .I3(n27851), .O(n8825[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3971_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_43_17_lut (.I0(n2312), .I1(\FRAME_MATCHER.i [15]), .I2(GND_net), 
            .I3(n27809), .O(n2_adj_4242)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_17_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_43_17 (.CI(n27809), .I0(\FRAME_MATCHER.i [15]), .I1(GND_net), 
            .CO(n27810));
    SB_LUT4 add_43_16_lut (.I0(n2312), .I1(\FRAME_MATCHER.i [14]), .I2(GND_net), 
            .I3(n27808), .O(n2_adj_4244)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_16_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_3971_6 (.CI(n27851), .I0(byte_transmit_counter[4]), .I1(GND_net), 
            .CO(n27852));
    SB_CARRY add_43_16 (.CI(n27808), .I0(\FRAME_MATCHER.i [14]), .I1(GND_net), 
            .CO(n27809));
    SB_LUT4 add_43_15_lut (.I0(n2312), .I1(\FRAME_MATCHER.i [13]), .I2(GND_net), 
            .I3(n27807), .O(n2_adj_4246)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_15_lut.LUT_INIT = 16'h8228;
    SB_LUT4 add_3971_5_lut (.I0(GND_net), .I1(byte_transmit_counter[3]), 
            .I2(GND_net), .I3(n27850), .O(n8825[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3971_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_43_15 (.CI(n27807), .I0(\FRAME_MATCHER.i [13]), .I1(GND_net), 
            .CO(n27808));
    SB_CARRY add_3971_5 (.CI(n27850), .I0(byte_transmit_counter[3]), .I1(GND_net), 
            .CO(n27851));
    SB_LUT4 add_43_14_lut (.I0(n2312), .I1(\FRAME_MATCHER.i [12]), .I2(GND_net), 
            .I3(n27806), .O(n2_adj_4248)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_14_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_43_14 (.CI(n27806), .I0(\FRAME_MATCHER.i [12]), .I1(GND_net), 
            .CO(n27807));
    SB_LUT4 add_3971_4_lut (.I0(GND_net), .I1(byte_transmit_counter[2]), 
            .I2(GND_net), .I3(n27849), .O(n8825[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3971_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_2_lut_3_lut_adj_1269 (.I0(n2_adj_4082), .I1(n2_adj_4272), 
            .I2(\FRAME_MATCHER.state_c [5]), .I3(GND_net), .O(n32181));
    defparam i1_2_lut_3_lut_adj_1269.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_2_lut_3_lut_adj_1270 (.I0(n2_adj_4082), .I1(n2_adj_4272), 
            .I2(\FRAME_MATCHER.state_c [6]), .I3(GND_net), .O(n32185));
    defparam i1_2_lut_3_lut_adj_1270.LUT_INIT = 16'he0e0;
    SB_CARRY add_3971_4 (.CI(n27849), .I0(byte_transmit_counter[2]), .I1(GND_net), 
            .CO(n27850));
    SB_LUT4 i1_2_lut_3_lut_adj_1271 (.I0(n2_adj_4082), .I1(n2_adj_4272), 
            .I2(\FRAME_MATCHER.state_c [7]), .I3(GND_net), .O(n32189));
    defparam i1_2_lut_3_lut_adj_1271.LUT_INIT = 16'he0e0;
    SB_LUT4 add_3971_3_lut (.I0(GND_net), .I1(byte_transmit_counter[1]), 
            .I2(GND_net), .I3(n27848), .O(n8825[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3971_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_2_lut_3_lut_adj_1272 (.I0(n2_adj_4082), .I1(n2_adj_4272), 
            .I2(\FRAME_MATCHER.state_c [8]), .I3(GND_net), .O(n32145));
    defparam i1_2_lut_3_lut_adj_1272.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_2_lut_3_lut_adj_1273 (.I0(n2_adj_4082), .I1(n2_adj_4272), 
            .I2(\FRAME_MATCHER.state_c [9]), .I3(GND_net), .O(n32191));
    defparam i1_2_lut_3_lut_adj_1273.LUT_INIT = 16'he0e0;
    SB_CARRY add_3971_3 (.CI(n27848), .I0(byte_transmit_counter[1]), .I1(GND_net), 
            .CO(n27849));
    SB_LUT4 i1_2_lut_3_lut_adj_1274 (.I0(n2_adj_4082), .I1(n2_adj_4272), 
            .I2(\FRAME_MATCHER.state_c [10]), .I3(GND_net), .O(n32193));
    defparam i1_2_lut_3_lut_adj_1274.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_3_lut_4_lut (.I0(\data_out_frame[24] [2]), .I1(\data_out_frame[24] [1]), 
            .I2(n32931), .I3(n18330), .O(n32947));   // verilog/coms.v(78[16:27])
    defparam i1_3_lut_4_lut.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_3_lut_adj_1275 (.I0(n2_adj_4082), .I1(n2_adj_4272), 
            .I2(\FRAME_MATCHER.state_c [11]), .I3(GND_net), .O(n32233));
    defparam i1_2_lut_3_lut_adj_1275.LUT_INIT = 16'he0e0;
    SB_LUT4 i8_2_lut_3_lut (.I0(\data_out_frame[24] [2]), .I1(\data_out_frame[24] [1]), 
            .I2(n30866), .I3(GND_net), .O(n40));   // verilog/coms.v(78[16:27])
    defparam i8_2_lut_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1276 (.I0(n2_adj_4082), .I1(n2_adj_4272), 
            .I2(\FRAME_MATCHER.state_c [12]), .I3(GND_net), .O(n7_adj_4205));
    defparam i1_2_lut_3_lut_adj_1276.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_2_lut_adj_1277 (.I0(\FRAME_MATCHER.state[0] ), .I1(n32655), 
            .I2(GND_net), .I3(GND_net), .O(n7));
    defparam i1_2_lut_adj_1277.LUT_INIT = 16'heeee;
    SB_LUT4 i9331_3_lut (.I0(n31), .I1(n31_adj_4177), .I2(\FRAME_MATCHER.state_c [1]), 
            .I3(GND_net), .O(n14574));   // verilog/coms.v(145[4] 299[11])
    defparam i9331_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4_4_lut_adj_1278 (.I0(\data_in_frame[0] [4]), .I1(\data_in_frame[0] [6]), 
            .I2(ID[4]), .I3(ID[6]), .O(n12_adj_4274));   // verilog/coms.v(238[12:32])
    defparam i4_4_lut_adj_1278.LUT_INIT = 16'h7bde;
    SB_LUT4 i2_4_lut_adj_1279 (.I0(\data_in_frame[0] [1]), .I1(\data_in_frame[0] [2]), 
            .I2(ID[1]), .I3(ID[2]), .O(n10_adj_4275));   // verilog/coms.v(238[12:32])
    defparam i2_4_lut_adj_1279.LUT_INIT = 16'h7bde;
    SB_LUT4 i3_4_lut_adj_1280 (.I0(\data_in_frame[0] [7]), .I1(\data_in_frame[0] [5]), 
            .I2(ID[7]), .I3(ID[5]), .O(n11));   // verilog/coms.v(238[12:32])
    defparam i3_4_lut_adj_1280.LUT_INIT = 16'h7bde;
    SB_LUT4 i1_4_lut_adj_1281 (.I0(\data_in_frame[0] [0]), .I1(\data_in_frame[0] [3]), 
            .I2(ID[0]), .I3(ID[3]), .O(n9));   // verilog/coms.v(238[12:32])
    defparam i1_4_lut_adj_1281.LUT_INIT = 16'h7bde;
    SB_LUT4 i7_4_lut_adj_1282 (.I0(n9), .I1(n11), .I2(n10_adj_4275), .I3(n12_adj_4274), 
            .O(n14993));   // verilog/coms.v(238[12:32])
    defparam i7_4_lut_adj_1282.LUT_INIT = 16'hfffe;
    SB_LUT4 i2_2_lut_adj_1283 (.I0(n14993), .I1(\FRAME_MATCHER.state [3]), 
            .I2(GND_net), .I3(GND_net), .O(n8_adj_4276));
    defparam i2_2_lut_adj_1283.LUT_INIT = 16'heeee;
    SB_LUT4 i30402_4_lut (.I0(n14574), .I1(n7), .I2(\FRAME_MATCHER.state_c [2]), 
            .I3(n8_adj_4276), .O(n18646));
    defparam i30402_4_lut.LUT_INIT = 16'h0010;
    SB_LUT4 i18627_2_lut_3_lut (.I0(n2_adj_4082), .I1(n2_adj_4272), .I2(\FRAME_MATCHER.state_c [13]), 
            .I3(GND_net), .O(n23753));
    defparam i18627_2_lut_3_lut.LUT_INIT = 16'he0e0;
    SB_LUT4 mux_1387_i1_3_lut (.I0(\data_in_frame[19] [0]), .I1(\data_in_frame[3] [0]), 
            .I2(n5454), .I3(GND_net), .O(n5455));
    defparam mux_1387_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i18628_2_lut_3_lut (.I0(n2_adj_4082), .I1(n2_adj_4272), .I2(\FRAME_MATCHER.state_c [14]), 
            .I3(GND_net), .O(n23755));
    defparam i18628_2_lut_3_lut.LUT_INIT = 16'he0e0;
    SB_LUT4 add_3971_2_lut (.I0(GND_net), .I1(byte_transmit_counter[0]), 
            .I2(tx_transmit_N_3387), .I3(GND_net), .O(n8825[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3971_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_2_lut_3_lut_adj_1284 (.I0(n2_adj_4082), .I1(n2_adj_4272), 
            .I2(\FRAME_MATCHER.state_c [15]), .I3(GND_net), .O(n32195));
    defparam i1_2_lut_3_lut_adj_1284.LUT_INIT = 16'he0e0;
    SB_DFF data_in_frame_0__i134 (.Q(\data_in_frame[16] [5]), .C(clk32MHz), 
           .D(n19136));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i3_4_lut_adj_1285 (.I0(n23788), .I1(\FRAME_MATCHER.i [5]), .I2(\FRAME_MATCHER.i [4]), 
            .I3(\FRAME_MATCHER.i [3]), .O(n32678));   // verilog/coms.v(154[7:23])
    defparam i3_4_lut_adj_1285.LUT_INIT = 16'hffdf;
    SB_DFF data_in_frame_0__i135 (.Q(\data_in_frame[16] [6]), .C(clk32MHz), 
           .D(n19135));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i136 (.Q(\data_in_frame[16] [7]), .C(clk32MHz), 
           .D(n19134));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i137 (.Q(\data_in_frame[17] [0]), .C(clk32MHz), 
           .D(n19133));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i138 (.Q(\data_in_frame[17] [1]), .C(clk32MHz), 
           .D(n19132));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i139 (.Q(\data_in_frame[17] [2]), .C(clk32MHz), 
           .D(n19131));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i140 (.Q(\data_in_frame[17] [3]), .C(clk32MHz), 
           .D(n19130));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i141 (.Q(\data_in_frame[17] [4]), .C(clk32MHz), 
           .D(n19129));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i142 (.Q(\data_in_frame[17] [5]), .C(clk32MHz), 
           .D(n19128));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i143 (.Q(\data_in_frame[17] [6]), .C(clk32MHz), 
           .D(n19127));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i144 (.Q(\data_in_frame[17] [7]), .C(clk32MHz), 
           .D(n19126));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i145 (.Q(\data_in_frame[18] [0]), .C(clk32MHz), 
           .D(n19125));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i146 (.Q(\data_in_frame[18] [1]), .C(clk32MHz), 
           .D(n19124));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i147 (.Q(\data_in_frame[18] [2]), .C(clk32MHz), 
           .D(n19123));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i148 (.Q(\data_in_frame[18] [3]), .C(clk32MHz), 
           .D(n19122));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i149 (.Q(\data_in_frame[18] [4]), .C(clk32MHz), 
           .D(n19121));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i150 (.Q(\data_in_frame[18] [5]), .C(clk32MHz), 
           .D(n19120));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i151 (.Q(\data_in_frame[18] [6]), .C(clk32MHz), 
           .D(n19119));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i152 (.Q(\data_in_frame[18] [7]), .C(clk32MHz), 
           .D(n19118));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i153 (.Q(\data_in_frame[19] [0]), .C(clk32MHz), 
           .D(n19117));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i154 (.Q(\data_in_frame[19] [1]), .C(clk32MHz), 
           .D(n19116));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i155 (.Q(\data_in_frame[19] [2]), .C(clk32MHz), 
           .D(n19115));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i156 (.Q(\data_in_frame[19] [3]), .C(clk32MHz), 
           .D(n19114));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i1_2_lut_adj_1286 (.I0(\FRAME_MATCHER.state_c [1]), .I1(\FRAME_MATCHER.state_c [2]), 
            .I2(GND_net), .I3(GND_net), .O(n17474));
    defparam i1_2_lut_adj_1286.LUT_INIT = 16'heeee;
    SB_LUT4 i12_4_lut_adj_1287 (.I0(\FRAME_MATCHER.state_c [19]), .I1(\FRAME_MATCHER.state_c [23]), 
            .I2(\FRAME_MATCHER.state_c [26]), .I3(\FRAME_MATCHER.state_c [27]), 
            .O(n28_adj_4277));
    defparam i12_4_lut_adj_1287.LUT_INIT = 16'hfffe;
    SB_LUT4 i10_4_lut_adj_1288 (.I0(\FRAME_MATCHER.state_c [17]), .I1(\FRAME_MATCHER.state_c [31]), 
            .I2(\FRAME_MATCHER.state_c [20]), .I3(\FRAME_MATCHER.state_c [16]), 
            .O(n26_adj_4278));
    defparam i10_4_lut_adj_1288.LUT_INIT = 16'hfffe;
    SB_LUT4 i11_4_lut_adj_1289 (.I0(\FRAME_MATCHER.state_c [29]), .I1(\FRAME_MATCHER.state_c [30]), 
            .I2(\FRAME_MATCHER.state_c [22]), .I3(\FRAME_MATCHER.state_c [18]), 
            .O(n27_adj_4279));
    defparam i11_4_lut_adj_1289.LUT_INIT = 16'hfffe;
    SB_LUT4 i9_4_lut_adj_1290 (.I0(\FRAME_MATCHER.state_c [25]), .I1(\FRAME_MATCHER.state_c [21]), 
            .I2(\FRAME_MATCHER.state_c [28]), .I3(\FRAME_MATCHER.state_c [24]), 
            .O(n25_adj_4280));
    defparam i9_4_lut_adj_1290.LUT_INIT = 16'hfffe;
    SB_LUT4 i3_4_lut_adj_1291 (.I0(\FRAME_MATCHER.state_c [12]), .I1(\FRAME_MATCHER.state_c [10]), 
            .I2(\FRAME_MATCHER.state_c [14]), .I3(\FRAME_MATCHER.state_c [13]), 
            .O(n32685));   // verilog/coms.v(127[12] 300[6])
    defparam i3_4_lut_adj_1291.LUT_INIT = 16'hfffe;
    SB_LUT4 i3_4_lut_adj_1292 (.I0(\FRAME_MATCHER.state_c [6]), .I1(\FRAME_MATCHER.state_c [7]), 
            .I2(\FRAME_MATCHER.state_c [4]), .I3(\FRAME_MATCHER.state_c [5]), 
            .O(n24511));
    defparam i3_4_lut_adj_1292.LUT_INIT = 16'hfffe;
    SB_LUT4 i3_4_lut_adj_1293 (.I0(\FRAME_MATCHER.state_c [15]), .I1(\FRAME_MATCHER.state_c [11]), 
            .I2(\FRAME_MATCHER.state_c [8]), .I3(\FRAME_MATCHER.state_c [9]), 
            .O(n32549));
    defparam i3_4_lut_adj_1293.LUT_INIT = 16'hfffe;
    SB_LUT4 i15_4_lut_adj_1294 (.I0(n25_adj_4280), .I1(n27_adj_4279), .I2(n26_adj_4278), 
            .I3(n28_adj_4277), .O(n24587));
    defparam i15_4_lut_adj_1294.LUT_INIT = 16'hfffe;
    SB_LUT4 i2_4_lut_adj_1295 (.I0(n24587), .I1(n32549), .I2(n24511), 
            .I3(n32685), .O(n32655));   // verilog/coms.v(201[5:24])
    defparam i2_4_lut_adj_1295.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_adj_1296 (.I0(\FRAME_MATCHER.state[0] ), .I1(n17551), 
            .I2(GND_net), .I3(GND_net), .O(n17552));   // verilog/coms.v(254[5:25])
    defparam i1_2_lut_adj_1296.LUT_INIT = 16'hdddd;
    SB_CARRY add_3971_2 (.CI(GND_net), .I0(byte_transmit_counter[0]), .I1(tx_transmit_N_3387), 
            .CO(n27848));
    SB_LUT4 add_43_13_lut (.I0(n2312), .I1(\FRAME_MATCHER.i [11]), .I2(GND_net), 
            .I3(n27805), .O(n2_adj_4250)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_13_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_43_13 (.CI(n27805), .I0(\FRAME_MATCHER.i [11]), .I1(GND_net), 
            .CO(n27806));
    SB_LUT4 i1_2_lut_adj_1297 (.I0(\FRAME_MATCHER.state[0] ), .I1(n32653), 
            .I2(GND_net), .I3(GND_net), .O(n17476));   // verilog/coms.v(151[5:27])
    defparam i1_2_lut_adj_1297.LUT_INIT = 16'hdddd;
    SB_LUT4 i14_2_lut (.I0(rx_data_ready), .I1(\FRAME_MATCHER.rx_data_ready_prev ), 
            .I2(GND_net), .I3(GND_net), .O(n161));   // verilog/coms.v(153[9:50])
    defparam i14_2_lut.LUT_INIT = 16'h2222;
    SB_DFF data_in_frame_0__i157 (.Q(\data_in_frame[19] [4]), .C(clk32MHz), 
           .D(n19113));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 add_43_12_lut (.I0(n2312), .I1(\FRAME_MATCHER.i [10]), .I2(GND_net), 
            .I3(n27804), .O(n2_adj_4252)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_12_lut.LUT_INIT = 16'h8228;
    SB_DFF data_in_frame_0__i158 (.Q(\data_in_frame[19] [5]), .C(clk32MHz), 
           .D(n19112));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 select_422_Select_0_i3_2_lut (.I0(\FRAME_MATCHER.i [0]), .I1(n2994), 
            .I2(GND_net), .I3(GND_net), .O(n3_c));
    defparam select_422_Select_0_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i30409_2_lut_3_lut (.I0(\FRAME_MATCHER.state_c [1]), .I1(\FRAME_MATCHER.state_c [2]), 
            .I2(\FRAME_MATCHER.state[0] ), .I3(GND_net), .O(n18858));
    defparam i30409_2_lut_3_lut.LUT_INIT = 16'h0e0e;
    SB_LUT4 i1_4_lut_4_lut (.I0(\FRAME_MATCHER.state[0] ), .I1(\FRAME_MATCHER.state_c [2]), 
            .I2(n1_adj_4281), .I3(\FRAME_MATCHER.state_c [1]), .O(n5_adj_4282));
    defparam i1_4_lut_4_lut.LUT_INIT = 16'h6273;
    SB_LUT4 i18822_2_lut_4_lut (.I0(n14993), .I1(n31), .I2(n31_adj_4177), 
            .I3(\FRAME_MATCHER.state_c [1]), .O(n1_adj_4281));
    defparam i18822_2_lut_4_lut.LUT_INIT = 16'hfaee;
    SB_LUT4 i2_3_lut_adj_1298 (.I0(byte_transmit_counter[5]), .I1(byte_transmit_counter[7]), 
            .I2(byte_transmit_counter[6]), .I3(GND_net), .O(n11316));   // verilog/coms.v(214[11:56])
    defparam i2_3_lut_adj_1298.LUT_INIT = 16'hfefe;
    SB_LUT4 i19162_2_lut (.I0(byte_transmit_counter[0]), .I1(byte_transmit_counter[1]), 
            .I2(GND_net), .I3(GND_net), .O(n24295));
    defparam i19162_2_lut.LUT_INIT = 16'h8888;
    SB_DFF data_in_frame_0__i159 (.Q(\data_in_frame[19] [6]), .C(clk32MHz), 
           .D(n19111));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i2_4_lut_adj_1299 (.I0(byte_transmit_counter[3]), .I1(byte_transmit_counter[4]), 
            .I2(n24295), .I3(byte_transmit_counter[2]), .O(n24763));
    defparam i2_4_lut_adj_1299.LUT_INIT = 16'h8880;
    SB_LUT4 i1_3_lut_4_lut_adj_1300 (.I0(\FRAME_MATCHER.state [3]), .I1(n32655), 
            .I2(n33453), .I3(n5592), .O(n17503));
    defparam i1_3_lut_4_lut_adj_1300.LUT_INIT = 16'hecee;
    SB_LUT4 i26762_3_lut (.I0(\FRAME_MATCHER.state [3]), .I1(n32655), .I2(n33453), 
            .I3(GND_net), .O(n33511));
    defparam i26762_3_lut.LUT_INIT = 16'hecec;
    SB_LUT4 i3_4_lut_adj_1301 (.I0(n24763), .I1(n23740), .I2(n24226), 
            .I3(n11316), .O(n34406));
    defparam i3_4_lut_adj_1301.LUT_INIT = 16'hffef;
    SB_LUT4 mux_911_i1_3_lut (.I0(n34406), .I1(\FRAME_MATCHER.state [3]), 
            .I2(n5592), .I3(GND_net), .O(n3598[0]));   // verilog/coms.v(145[4] 299[11])
    defparam mux_911_i1_3_lut.LUT_INIT = 16'h5c5c;
    SB_DFFESR byte_transmit_counter_i0_i0 (.Q(byte_transmit_counter[0]), .C(clk32MHz), 
            .E(n18619), .D(n8825[0]), .R(n18939));   // verilog/coms.v(127[12] 300[6])
    SB_CARRY add_43_12 (.CI(n27804), .I0(\FRAME_MATCHER.i [10]), .I1(GND_net), 
            .CO(n27805));
    SB_LUT4 i5_2_lut_3_lut_4_lut (.I0(\data_out_frame[4] [3]), .I1(\data_out_frame[4] [4]), 
            .I2(\data_out_frame[6] [5]), .I3(\data_out_frame[4] [0]), .O(n16));   // verilog/coms.v(74[16:43])
    defparam i5_2_lut_3_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i18615_2_lut (.I0(tx_active), .I1(r_SM_Main_2__N_3490[0]), .I2(GND_net), 
            .I3(GND_net), .O(n23740));
    defparam i18615_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 add_43_11_lut (.I0(n2312), .I1(\FRAME_MATCHER.i [9]), .I2(GND_net), 
            .I3(n27803), .O(n2_adj_4254)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_11_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i3_4_lut_adj_1302 (.I0(\FRAME_MATCHER.state[0] ), .I1(n17474), 
            .I2(\FRAME_MATCHER.state [3]), .I3(n32655), .O(n63_adj_8));   // verilog/coms.v(201[5:24])
    defparam i3_4_lut_adj_1302.LUT_INIT = 16'hffef;
    SB_LUT4 i1_2_lut_3_lut_4_lut (.I0(\data_out_frame[6] [1]), .I1(\data_out_frame[4] [1]), 
            .I2(\data_out_frame[4] [0]), .I3(\data_out_frame[6] [2]), .O(n17566));   // verilog/coms.v(73[16:42])
    defparam i1_2_lut_3_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i13802_2_lut (.I0(n18619), .I1(n17559), .I2(GND_net), .I3(GND_net), 
            .O(n18939));   // verilog/coms.v(127[12] 300[6])
    defparam i13802_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1303 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(n32655), .I2(\FRAME_MATCHER.state_c [1]), .I3(\FRAME_MATCHER.state_c [2]), 
            .O(n32653));   // verilog/coms.v(212[5:16])
    defparam i1_2_lut_3_lut_4_lut_adj_1303.LUT_INIT = 16'hfffe;
    SB_LUT4 i2_4_lut_4_lut_4_lut (.I0(\FRAME_MATCHER.state_c [2]), .I1(\FRAME_MATCHER.state[0] ), 
            .I2(\FRAME_MATCHER.state_31__N_2598 [3]), .I3(\FRAME_MATCHER.state_c [1]), 
            .O(n6_adj_4283));
    defparam i2_4_lut_4_lut_4_lut.LUT_INIT = 16'h8988;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1304 (.I0(\FRAME_MATCHER.state[0] ), 
            .I1(n17551), .I2(n39), .I3(n32653), .O(n24499));
    defparam i1_2_lut_3_lut_4_lut_adj_1304.LUT_INIT = 16'hd050;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1305 (.I0(\FRAME_MATCHER.state[0] ), 
            .I1(n17551), .I2(n39), .I3(n32653), .O(n2994));
    defparam i1_2_lut_3_lut_4_lut_adj_1305.LUT_INIT = 16'hd000;
    SB_LUT4 i1_2_lut_3_lut_adj_1306 (.I0(n2_adj_4082), .I1(n2_adj_4272), 
            .I2(\FRAME_MATCHER.state_c [16]), .I3(GND_net), .O(n32197));
    defparam i1_2_lut_3_lut_adj_1306.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_2_lut_3_lut_adj_1307 (.I0(n2_adj_4082), .I1(n2_adj_4272), 
            .I2(\FRAME_MATCHER.state_c [17]), .I3(GND_net), .O(n32199));
    defparam i1_2_lut_3_lut_adj_1307.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_2_lut_3_lut_adj_1308 (.I0(n2_adj_4082), .I1(n2_adj_4272), 
            .I2(\FRAME_MATCHER.state_c [18]), .I3(GND_net), .O(n32201));
    defparam i1_2_lut_3_lut_adj_1308.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_2_lut_3_lut_adj_1309 (.I0(n2_adj_4082), .I1(n2_adj_4272), 
            .I2(\FRAME_MATCHER.state_c [19]), .I3(GND_net), .O(n32203));
    defparam i1_2_lut_3_lut_adj_1309.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1310 (.I0(\data_out_frame[7] [7]), .I1(\data_out_frame[7] [6]), 
            .I2(\data_out_frame[5] [7]), .I3(\data_out_frame[8] [1]), .O(n6_adj_4041));   // verilog/coms.v(85[17:70])
    defparam i1_2_lut_3_lut_4_lut_adj_1310.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1311 (.I0(\data_in_frame[15] [7]), .I1(\data_in_frame[9] [4]), 
            .I2(\data_in_frame[13] [6]), .I3(\data_in_frame[16] [1]), .O(n8_adj_4167));
    defparam i1_2_lut_3_lut_4_lut_adj_1311.LUT_INIT = 16'h6996;
    SB_LUT4 byte_transmit_counter_3__bdd_4_lut (.I0(byte_transmit_counter[3]), 
            .I1(n37673), .I2(n36301), .I3(byte_transmit_counter[4]), .O(n37934));
    defparam byte_transmit_counter_3__bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_LUT4 n37934_bdd_4_lut (.I0(n37934), .I1(n14_adj_4199), .I2(n7_adj_4284), 
            .I3(byte_transmit_counter[4]), .O(tx_data[1]));
    defparam n37934_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[14] [2]), .I2(\data_out_frame[15] [2]), 
            .I3(byte_transmit_counter[1]), .O(n37928));
    defparam byte_transmit_counter_0__bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_LUT4 n37928_bdd_4_lut (.I0(n37928), .I1(\data_out_frame[13] [2]), 
            .I2(\data_out_frame[12] [2]), .I3(byte_transmit_counter[1]), 
            .O(n37931));
    defparam n37928_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_31125 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[14] [3]), .I2(\data_out_frame[15] [3]), 
            .I3(byte_transmit_counter[1]), .O(n37922));
    defparam byte_transmit_counter_0__bdd_4_lut_31125.LUT_INIT = 16'he4aa;
    SB_CARRY add_43_11 (.CI(n27803), .I0(\FRAME_MATCHER.i [9]), .I1(GND_net), 
            .CO(n27804));
    SB_LUT4 n37922_bdd_4_lut (.I0(n37922), .I1(\data_out_frame[13] [3]), 
            .I2(\data_out_frame[12] [3]), .I3(byte_transmit_counter[1]), 
            .O(n37925));
    defparam n37922_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_31120 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[26] [4]), .I2(\data_out_frame[27] [4]), 
            .I3(byte_transmit_counter[1]), .O(n37916));
    defparam byte_transmit_counter_0__bdd_4_lut_31120.LUT_INIT = 16'he4aa;
    SB_LUT4 n37916_bdd_4_lut (.I0(n37916), .I1(\data_out_frame[25] [4]), 
            .I2(\data_out_frame[24] [4]), .I3(byte_transmit_counter[1]), 
            .O(n37919));
    defparam n37916_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_31115 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[26] [5]), .I2(\data_out_frame[27] [5]), 
            .I3(byte_transmit_counter[1]), .O(n37910));
    defparam byte_transmit_counter_0__bdd_4_lut_31115.LUT_INIT = 16'he4aa;
    SB_LUT4 n37910_bdd_4_lut (.I0(n37910), .I1(\data_out_frame[25] [5]), 
            .I2(\data_out_frame[24] [5]), .I3(byte_transmit_counter[1]), 
            .O(n37913));
    defparam n37910_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_31110 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[26] [6]), .I2(\data_out_frame[27] [6]), 
            .I3(byte_transmit_counter[1]), .O(n37904));
    defparam byte_transmit_counter_0__bdd_4_lut_31110.LUT_INIT = 16'he4aa;
    SB_LUT4 n37904_bdd_4_lut (.I0(n37904), .I1(\data_out_frame[25] [6]), 
            .I2(\data_out_frame[24] [6]), .I3(byte_transmit_counter[1]), 
            .O(n37907));
    defparam n37904_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_31105 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[26] [7]), .I2(\data_out_frame[27] [7]), 
            .I3(byte_transmit_counter[1]), .O(n37898));
    defparam byte_transmit_counter_0__bdd_4_lut_31105.LUT_INIT = 16'he4aa;
    SB_LUT4 n37898_bdd_4_lut (.I0(n37898), .I1(\data_out_frame[25] [7]), 
            .I2(\data_out_frame[24] [7]), .I3(byte_transmit_counter[1]), 
            .O(n37901));
    defparam n37898_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 add_43_10_lut (.I0(n2312), .I1(\FRAME_MATCHER.i [8]), .I2(GND_net), 
            .I3(n27802), .O(n2_adj_4256)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_10_lut.LUT_INIT = 16'h8228;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_31100 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[14] [5]), .I2(\data_out_frame[15] [5]), 
            .I3(byte_transmit_counter[1]), .O(n37886));
    defparam byte_transmit_counter_0__bdd_4_lut_31100.LUT_INIT = 16'he4aa;
    SB_LUT4 n37886_bdd_4_lut (.I0(n37886), .I1(\data_out_frame[13] [5]), 
            .I2(\data_out_frame[12] [5]), .I3(byte_transmit_counter[1]), 
            .O(n37889));
    defparam n37886_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_31090 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[10] [7]), .I2(\data_out_frame[11] [7]), 
            .I3(byte_transmit_counter[1]), .O(n37874));
    defparam byte_transmit_counter_0__bdd_4_lut_31090.LUT_INIT = 16'he4aa;
    SB_LUT4 n37874_bdd_4_lut (.I0(n37874), .I1(\data_out_frame[9] [7]), 
            .I2(\data_out_frame[8] [7]), .I3(byte_transmit_counter[1]), 
            .O(n37877));
    defparam n37874_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_31080 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[10] [0]), .I2(\data_out_frame[11] [0]), 
            .I3(byte_transmit_counter[1]), .O(n37868));
    defparam byte_transmit_counter_0__bdd_4_lut_31080.LUT_INIT = 16'he4aa;
    SB_LUT4 n37868_bdd_4_lut (.I0(n37868), .I1(\data_out_frame[9] [0]), 
            .I2(\data_out_frame[8] [0]), .I3(byte_transmit_counter[1]), 
            .O(n37871));
    defparam n37868_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_31075 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[14] [0]), .I2(\data_out_frame[15] [0]), 
            .I3(byte_transmit_counter[1]), .O(n37862));
    defparam byte_transmit_counter_0__bdd_4_lut_31075.LUT_INIT = 16'he4aa;
    SB_LUT4 n37862_bdd_4_lut (.I0(n37862), .I1(\data_out_frame[13] [0]), 
            .I2(\data_out_frame[12] [0]), .I3(byte_transmit_counter[1]), 
            .O(n37865));
    defparam n37862_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_31070 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[10] [6]), .I2(\data_out_frame[11] [6]), 
            .I3(byte_transmit_counter[1]), .O(n37856));
    defparam byte_transmit_counter_0__bdd_4_lut_31070.LUT_INIT = 16'he4aa;
    SB_LUT4 n37856_bdd_4_lut (.I0(n37856), .I1(\data_out_frame[9] [6]), 
            .I2(\data_out_frame[8] [6]), .I3(byte_transmit_counter[1]), 
            .O(n37859));
    defparam n37856_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_CARRY add_43_10 (.CI(n27802), .I0(\FRAME_MATCHER.i [8]), .I1(GND_net), 
            .CO(n27803));
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_31065 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[10] [5]), .I2(\data_out_frame[11] [5]), 
            .I3(byte_transmit_counter[1]), .O(n37850));
    defparam byte_transmit_counter_0__bdd_4_lut_31065.LUT_INIT = 16'he4aa;
    SB_LUT4 n37850_bdd_4_lut (.I0(n37850), .I1(\data_out_frame[9] [5]), 
            .I2(\data_out_frame[8] [5]), .I3(byte_transmit_counter[1]), 
            .O(n37853));
    defparam n37850_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_2_lut_3_lut_adj_1312 (.I0(n2_adj_4082), .I1(n2_adj_4272), 
            .I2(\FRAME_MATCHER.state_c [20]), .I3(GND_net), .O(n32205));
    defparam i1_2_lut_3_lut_adj_1312.LUT_INIT = 16'he0e0;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_31060 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[10] [4]), .I2(\data_out_frame[11] [4]), 
            .I3(byte_transmit_counter[1]), .O(n37844));
    defparam byte_transmit_counter_0__bdd_4_lut_31060.LUT_INIT = 16'he4aa;
    SB_LUT4 n37844_bdd_4_lut (.I0(n37844), .I1(\data_out_frame[9] [4]), 
            .I2(\data_out_frame[8] [4]), .I3(byte_transmit_counter[1]), 
            .O(n37847));
    defparam n37844_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_31055 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[14] [6]), .I2(\data_out_frame[15] [6]), 
            .I3(byte_transmit_counter[1]), .O(n37838));
    defparam byte_transmit_counter_0__bdd_4_lut_31055.LUT_INIT = 16'he4aa;
    SB_LUT4 n37838_bdd_4_lut (.I0(n37838), .I1(\data_out_frame[13] [6]), 
            .I2(\data_out_frame[12] [6]), .I3(byte_transmit_counter[1]), 
            .O(n37841));
    defparam n37838_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i19364_1_lut (.I0(n24499), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n2312));
    defparam i19364_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_31050 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[10] [3]), .I2(\data_out_frame[11] [3]), 
            .I3(byte_transmit_counter[1]), .O(n37832));
    defparam byte_transmit_counter_0__bdd_4_lut_31050.LUT_INIT = 16'he4aa;
    SB_LUT4 n37832_bdd_4_lut (.I0(n37832), .I1(\data_out_frame[9] [3]), 
            .I2(\data_out_frame[8] [3]), .I3(byte_transmit_counter[1]), 
            .O(n37835));
    defparam n37832_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_2_lut_3_lut_adj_1313 (.I0(n2_adj_4082), .I1(n2_adj_4272), 
            .I2(\FRAME_MATCHER.state_c [21]), .I3(GND_net), .O(n32207));
    defparam i1_2_lut_3_lut_adj_1313.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_4_lut_adj_1314 (.I0(\data_in_frame[1] [0]), .I1(\data_in_frame[2] [7]), 
            .I2(Kp_23__N_862), .I3(\data_in_frame[0] [5]), .O(n18058));
    defparam i1_4_lut_adj_1314.LUT_INIT = 16'h6996;
    SB_LUT4 add_43_9_lut (.I0(n2312), .I1(\FRAME_MATCHER.i [7]), .I2(GND_net), 
            .I3(n27801), .O(n2_adj_4258)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_9_lut.LUT_INIT = 16'h8228;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_31045 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[10] [2]), .I2(\data_out_frame[11] [2]), 
            .I3(byte_transmit_counter[1]), .O(n37814));
    defparam byte_transmit_counter_0__bdd_4_lut_31045.LUT_INIT = 16'he4aa;
    SB_LUT4 n37814_bdd_4_lut (.I0(n37814), .I1(\data_out_frame[9] [2]), 
            .I2(\data_out_frame[8] [2]), .I3(byte_transmit_counter[1]), 
            .O(n37817));
    defparam n37814_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_2_lut_3_lut_adj_1315 (.I0(n2_adj_4082), .I1(n2_adj_4272), 
            .I2(\FRAME_MATCHER.state_c [22]), .I3(GND_net), .O(n32209));
    defparam i1_2_lut_3_lut_adj_1315.LUT_INIT = 16'he0e0;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_31030 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[10] [1]), .I2(\data_out_frame[11] [1]), 
            .I3(byte_transmit_counter[1]), .O(n37802));
    defparam byte_transmit_counter_0__bdd_4_lut_31030.LUT_INIT = 16'he4aa;
    SB_LUT4 n37802_bdd_4_lut (.I0(n37802), .I1(\data_out_frame[9] [1]), 
            .I2(\data_out_frame[8] [1]), .I3(byte_transmit_counter[1]), 
            .O(n37805));
    defparam n37802_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_31020 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[14] [1]), .I2(\data_out_frame[15] [1]), 
            .I3(byte_transmit_counter[1]), .O(n37796));
    defparam byte_transmit_counter_0__bdd_4_lut_31020.LUT_INIT = 16'he4aa;
    SB_LUT4 n37796_bdd_4_lut (.I0(n37796), .I1(\data_out_frame[13] [1]), 
            .I2(\data_out_frame[12] [1]), .I3(byte_transmit_counter[1]), 
            .O(n37799));
    defparam n37796_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i2_3_lut_4_lut_adj_1316 (.I0(n18086), .I1(n32816), .I2(\data_out_frame[24] [4]), 
            .I3(n33000), .O(n33700));
    defparam i2_3_lut_4_lut_adj_1316.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1317 (.I0(\data_in_frame[13] [4]), .I1(\data_in_frame[9] [2]), 
            .I2(n17827), .I3(n17846), .O(n33159));   // verilog/coms.v(73[16:42])
    defparam i1_2_lut_3_lut_4_lut_adj_1317.LUT_INIT = 16'h6996;
    SB_LUT4 byte_transmit_counter_3__bdd_4_lut_31130 (.I0(byte_transmit_counter[3]), 
            .I1(n37679), .I2(n36304), .I3(byte_transmit_counter[4]), .O(n37790));
    defparam byte_transmit_counter_3__bdd_4_lut_31130.LUT_INIT = 16'he4aa;
    SB_LUT4 n37790_bdd_4_lut (.I0(n37790), .I1(n14_adj_4178), .I2(n7_adj_4285), 
            .I3(byte_transmit_counter[4]), .O(tx_data[0]));
    defparam n37790_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_3__bdd_4_lut_31010 (.I0(byte_transmit_counter[3]), 
            .I1(n37685), .I2(n36298), .I3(byte_transmit_counter[4]), .O(n37784));
    defparam byte_transmit_counter_3__bdd_4_lut_31010.LUT_INIT = 16'he4aa;
    SB_LUT4 n37784_bdd_4_lut (.I0(n37784), .I1(n14_adj_4176), .I2(n7_adj_4286), 
            .I3(byte_transmit_counter[4]), .O(tx_data[2]));
    defparam n37784_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_3__bdd_4_lut_31005 (.I0(byte_transmit_counter[3]), 
            .I1(n37691), .I2(n36293), .I3(byte_transmit_counter[4]), .O(n37778));
    defparam byte_transmit_counter_3__bdd_4_lut_31005.LUT_INIT = 16'he4aa;
    SB_LUT4 n37778_bdd_4_lut (.I0(n37778), .I1(n14_adj_4175), .I2(n7_adj_4287), 
            .I3(byte_transmit_counter[4]), .O(tx_data[3]));
    defparam n37778_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_3__bdd_4_lut_31000 (.I0(byte_transmit_counter[3]), 
            .I1(n37697), .I2(n36290), .I3(byte_transmit_counter[4]), .O(n37772));
    defparam byte_transmit_counter_3__bdd_4_lut_31000.LUT_INIT = 16'he4aa;
    SB_LUT4 n37772_bdd_4_lut (.I0(n37772), .I1(n14_adj_4173), .I2(n7_adj_4288), 
            .I3(byte_transmit_counter[4]), .O(tx_data[4]));
    defparam n37772_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_2_lut_3_lut_adj_1318 (.I0(n2_adj_4082), .I1(n2_adj_4272), 
            .I2(\FRAME_MATCHER.state_c [23]), .I3(GND_net), .O(n32211));
    defparam i1_2_lut_3_lut_adj_1318.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_2_lut_3_lut_adj_1319 (.I0(n2_adj_4082), .I1(n2_adj_4272), 
            .I2(\FRAME_MATCHER.state_c [24]), .I3(GND_net), .O(n32213));
    defparam i1_2_lut_3_lut_adj_1319.LUT_INIT = 16'he0e0;
    SB_LUT4 byte_transmit_counter_3__bdd_4_lut_30995 (.I0(byte_transmit_counter[3]), 
            .I1(n37703), .I2(n36279), .I3(byte_transmit_counter[4]), .O(n37766));
    defparam byte_transmit_counter_3__bdd_4_lut_30995.LUT_INIT = 16'he4aa;
    SB_LUT4 n37766_bdd_4_lut (.I0(n37766), .I1(n14_adj_4170), .I2(n7_adj_4289), 
            .I3(byte_transmit_counter[4]), .O(tx_data[5]));
    defparam n37766_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_3__bdd_4_lut_30990 (.I0(byte_transmit_counter[3]), 
            .I1(n37709), .I2(n36272), .I3(byte_transmit_counter[4]), .O(n37760));
    defparam byte_transmit_counter_3__bdd_4_lut_30990.LUT_INIT = 16'he4aa;
    SB_LUT4 n37760_bdd_4_lut (.I0(n37760), .I1(n14_adj_4164), .I2(n7_adj_4290), 
            .I3(byte_transmit_counter[4]), .O(tx_data[6]));
    defparam n37760_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_3__bdd_4_lut_30985 (.I0(byte_transmit_counter[3]), 
            .I1(n37715), .I2(n36248), .I3(byte_transmit_counter[4]), .O(n37754));
    defparam byte_transmit_counter_3__bdd_4_lut_30985.LUT_INIT = 16'he4aa;
    SB_LUT4 n37754_bdd_4_lut (.I0(n37754), .I1(n14_adj_4160), .I2(n7_adj_4291), 
            .I3(byte_transmit_counter[4]), .O(tx_data[7]));
    defparam n37754_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_31015 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[14] [7]), .I2(\data_out_frame[15] [7]), 
            .I3(byte_transmit_counter[1]), .O(n37748));
    defparam byte_transmit_counter_0__bdd_4_lut_31015.LUT_INIT = 16'he4aa;
    SB_LUT4 n37748_bdd_4_lut (.I0(n37748), .I1(\data_out_frame[13] [7]), 
            .I2(\data_out_frame[12] [7]), .I3(byte_transmit_counter[1]), 
            .O(n37751));
    defparam n37748_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_CARRY add_43_9 (.CI(n27801), .I0(\FRAME_MATCHER.i [7]), .I1(GND_net), 
            .CO(n27802));
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_30976 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[14] [4]), .I2(\data_out_frame[15] [4]), 
            .I3(byte_transmit_counter[1]), .O(n37724));
    defparam byte_transmit_counter_0__bdd_4_lut_30976.LUT_INIT = 16'he4aa;
    SB_LUT4 n37724_bdd_4_lut (.I0(n37724), .I1(\data_out_frame[13] [4]), 
            .I2(\data_out_frame[12] [4]), .I3(byte_transmit_counter[1]), 
            .O(n37727));
    defparam n37724_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i7_2_lut (.I0(n18058), .I1(\data_in_frame[5] [3]), .I2(GND_net), 
            .I3(GND_net), .O(n27_adj_4191));   // verilog/coms.v(73[16:42])
    defparam i7_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1320 (.I0(\data_in_frame[1] [5]), .I1(\data_in_frame[1] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n32769));
    defparam i1_2_lut_adj_1320.LUT_INIT = 16'h6666;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_30958 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[26] [0]), .I2(\data_out_frame[27] [0]), 
            .I3(byte_transmit_counter[1]), .O(n37718));
    defparam byte_transmit_counter_0__bdd_4_lut_30958.LUT_INIT = 16'he4aa;
    SB_LUT4 n37718_bdd_4_lut (.I0(n37718), .I1(\data_out_frame[25] [0]), 
            .I2(\data_out_frame[24] [0]), .I3(byte_transmit_counter[1]), 
            .O(n37721));
    defparam n37718_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 add_43_8_lut (.I0(n2312), .I1(\FRAME_MATCHER.i [6]), .I2(GND_net), 
            .I3(n27800), .O(n2_adj_4260)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_8_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i1_2_lut_3_lut_adj_1321 (.I0(n2_adj_4082), .I1(n2_adj_4272), 
            .I2(\FRAME_MATCHER.state_c [25]), .I3(GND_net), .O(n32215));
    defparam i1_2_lut_3_lut_adj_1321.LUT_INIT = 16'he0e0;
    SB_CARRY add_43_8 (.CI(n27800), .I0(\FRAME_MATCHER.i [6]), .I1(GND_net), 
            .CO(n27801));
    SB_LUT4 add_43_7_lut (.I0(n2312), .I1(\FRAME_MATCHER.i [5]), .I2(GND_net), 
            .I3(n27799), .O(n2_adj_4262)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_7_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i1_2_lut_3_lut_adj_1322 (.I0(n2_adj_4082), .I1(n2_adj_4272), 
            .I2(\FRAME_MATCHER.state_c [26]), .I3(GND_net), .O(n32217));
    defparam i1_2_lut_3_lut_adj_1322.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_2_lut_adj_1323 (.I0(\data_in_frame[4] [4]), .I1(\data_in_frame[4] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n18235));   // verilog/coms.v(74[16:43])
    defparam i1_2_lut_adj_1323.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1324 (.I0(\data_in_frame[0] [6]), .I1(\data_in_frame[1] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n32776));   // verilog/coms.v(70[16:27])
    defparam i1_2_lut_adj_1324.LUT_INIT = 16'h6666;
    SB_CARRY add_43_7 (.CI(n27799), .I0(\FRAME_MATCHER.i [5]), .I1(GND_net), 
            .CO(n27800));
    SB_LUT4 add_43_6_lut (.I0(n2312), .I1(\FRAME_MATCHER.i [4]), .I2(GND_net), 
            .I3(n27798), .O(n2_adj_4264)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_6_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_43_6 (.CI(n27798), .I0(\FRAME_MATCHER.i [4]), .I1(GND_net), 
            .CO(n27799));
    SB_DFF data_in_frame_0__i160 (.Q(\data_in_frame[19] [7]), .C(clk32MHz), 
           .D(n19110));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut (.I0(byte_transmit_counter[1]), 
            .I1(n36270), .I2(n36271), .I3(byte_transmit_counter[2]), .O(n37712));
    defparam byte_transmit_counter_1__bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_LUT4 n37712_bdd_4_lut (.I0(n37712), .I1(n17_adj_4076), .I2(n16_adj_4075), 
            .I3(byte_transmit_counter[2]), .O(n37715));
    defparam n37712_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_30948 (.I0(byte_transmit_counter[1]), 
            .I1(n36273), .I2(n36274), .I3(byte_transmit_counter[2]), .O(n37706));
    defparam byte_transmit_counter_1__bdd_4_lut_30948.LUT_INIT = 16'he4aa;
    SB_LUT4 n37706_bdd_4_lut (.I0(n37706), .I1(n17_adj_4074), .I2(n16_adj_4072), 
            .I3(byte_transmit_counter[2]), .O(n37709));
    defparam n37706_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_30943 (.I0(byte_transmit_counter[1]), 
            .I1(n36284), .I2(n36285), .I3(byte_transmit_counter[2]), .O(n37700));
    defparam byte_transmit_counter_1__bdd_4_lut_30943.LUT_INIT = 16'he4aa;
    SB_LUT4 n37700_bdd_4_lut (.I0(n37700), .I1(n17_adj_4068), .I2(n16_adj_4067), 
            .I3(byte_transmit_counter[2]), .O(n37703));
    defparam n37700_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF data_in_frame_0__i161 (.Q(\data_in_frame[20] [0]), .C(clk32MHz), 
           .D(n19109));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i1_2_lut_adj_1325 (.I0(\data_in_frame[3] [1]), .I1(\data_in_frame[5] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n33139));   // verilog/coms.v(85[17:70])
    defparam i1_2_lut_adj_1325.LUT_INIT = 16'h6666;
    SB_DFF data_in_frame_0__i162 (.Q(\data_in_frame[20] [1]), .C(clk32MHz), 
           .D(n19108));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1326 (.I0(n2_adj_4085), .I1(n3_adj_4084), 
            .I2(n2970), .I3(n14711), .O(n6_adj_4081));
    defparam i1_2_lut_3_lut_4_lut_adj_1326.LUT_INIT = 16'hfeee;
    SB_LUT4 i1_2_lut_adj_1327 (.I0(\data_in_frame[5] [0]), .I1(\data_in_frame[4] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n33353));
    defparam i1_2_lut_adj_1327.LUT_INIT = 16'h6666;
    SB_LUT4 add_43_5_lut (.I0(n2312), .I1(\FRAME_MATCHER.i [3]), .I2(GND_net), 
            .I3(n27797), .O(n2_adj_4266)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_5_lut.LUT_INIT = 16'h8228;
    SB_DFF data_in_frame_0__i163 (.Q(\data_in_frame[20] [2]), .C(clk32MHz), 
           .D(n19107));   // verilog/coms.v(127[12] 300[6])
    SB_CARRY add_43_5 (.CI(n27797), .I0(\FRAME_MATCHER.i [3]), .I1(GND_net), 
            .CO(n27798));
    SB_LUT4 add_43_4_lut (.I0(n2312), .I1(\FRAME_MATCHER.i [2]), .I2(GND_net), 
            .I3(n27796), .O(n2_adj_4268)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_4_lut.LUT_INIT = 16'h8228;
    SB_DFF data_in_frame_0__i164 (.Q(\data_in_frame[20] [3]), .C(clk32MHz), 
           .D(n19106));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i165 (.Q(\data_in_frame[20] [4]), .C(clk32MHz), 
           .D(n19105));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i166 (.Q(\data_in_frame[20] [5]), .C(clk32MHz), 
           .D(n19104));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i167 (.Q(\data_in_frame[20] [6]), .C(clk32MHz), 
           .D(n19103));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i168 (.Q(\data_in_frame[20] [7]), .C(clk32MHz), 
           .D(n19102));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i169 (.Q(\data_in_frame[21] [0]), .C(clk32MHz), 
           .D(n19101));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i170 (.Q(\data_in_frame[21] [1]), .C(clk32MHz), 
           .D(n19100));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i171 (.Q(\data_in_frame[21] [2]), .C(clk32MHz), 
           .D(n19099));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i172 (.Q(\data_in_frame[21] [3]), .C(clk32MHz), 
           .D(n19098));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i173 (.Q(\data_in_frame[21] [4]), .C(clk32MHz), 
           .D(n19097));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i174 (.Q(\data_in_frame[21] [5]), .C(clk32MHz), 
           .D(n19096));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i175 (.Q(\data_in_frame[21] [6]), .C(clk32MHz), 
           .D(n19095));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i176 (.Q(\data_in_frame[21] [7]), .C(clk32MHz), 
           .D(n19094));   // verilog/coms.v(127[12] 300[6])
    SB_DFF control_mode_i0_i1 (.Q(control_mode[1]), .C(clk32MHz), .D(n19093));   // verilog/coms.v(127[12] 300[6])
    SB_DFF control_mode_i0_i2 (.Q(control_mode[2]), .C(clk32MHz), .D(n19092));   // verilog/coms.v(127[12] 300[6])
    SB_DFF control_mode_i0_i3 (.Q(control_mode[3]), .C(clk32MHz), .D(n19091));   // verilog/coms.v(127[12] 300[6])
    SB_DFF control_mode_i0_i4 (.Q(control_mode[4]), .C(clk32MHz), .D(n19090));   // verilog/coms.v(127[12] 300[6])
    SB_DFF control_mode_i0_i5 (.Q(control_mode[5]), .C(clk32MHz), .D(n19089));   // verilog/coms.v(127[12] 300[6])
    SB_DFF control_mode_i0_i6 (.Q(control_mode[6]), .C(clk32MHz), .D(n19088));   // verilog/coms.v(127[12] 300[6])
    SB_DFF control_mode_i0_i7 (.Q(control_mode[7]), .C(clk32MHz), .D(n19087));   // verilog/coms.v(127[12] 300[6])
    SB_DFF PWMLimit_i0_i1 (.Q(PWMLimit[1]), .C(clk32MHz), .D(n19086));   // verilog/coms.v(127[12] 300[6])
    SB_DFF PWMLimit_i0_i2 (.Q(PWMLimit[2]), .C(clk32MHz), .D(n19085));   // verilog/coms.v(127[12] 300[6])
    SB_DFF PWMLimit_i0_i3 (.Q(PWMLimit[3]), .C(clk32MHz), .D(n19084));   // verilog/coms.v(127[12] 300[6])
    SB_DFF PWMLimit_i0_i4 (.Q(PWMLimit[4]), .C(clk32MHz), .D(n19083));   // verilog/coms.v(127[12] 300[6])
    SB_DFF PWMLimit_i0_i5 (.Q(PWMLimit[5]), .C(clk32MHz), .D(n19082));   // verilog/coms.v(127[12] 300[6])
    SB_DFF PWMLimit_i0_i6 (.Q(PWMLimit[6]), .C(clk32MHz), .D(n19081));   // verilog/coms.v(127[12] 300[6])
    SB_DFF PWMLimit_i0_i7 (.Q(PWMLimit[7]), .C(clk32MHz), .D(n19080));   // verilog/coms.v(127[12] 300[6])
    SB_DFF PWMLimit_i0_i8 (.Q(PWMLimit[8]), .C(clk32MHz), .D(n19079));   // verilog/coms.v(127[12] 300[6])
    SB_DFF PWMLimit_i0_i9 (.Q(PWMLimit[9]), .C(clk32MHz), .D(n19078));   // verilog/coms.v(127[12] 300[6])
    SB_DFF PWMLimit_i0_i10 (.Q(PWMLimit[10]), .C(clk32MHz), .D(n19077));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE setpoint__i1 (.Q(setpoint[1]), .C(clk32MHz), .E(n18646), .D(n5456));   // verilog/coms.v(127[12] 300[6])
    SB_DFF PWMLimit_i0_i11 (.Q(PWMLimit[11]), .C(clk32MHz), .D(n19076));   // verilog/coms.v(127[12] 300[6])
    SB_CARRY add_43_4 (.CI(n27796), .I0(\FRAME_MATCHER.i [2]), .I1(GND_net), 
            .CO(n27797));
    SB_DFF PWMLimit_i0_i12 (.Q(PWMLimit[12]), .C(clk32MHz), .D(n19075));   // verilog/coms.v(127[12] 300[6])
    SB_DFF PWMLimit_i0_i13 (.Q(PWMLimit[13]), .C(clk32MHz), .D(n19074));   // verilog/coms.v(127[12] 300[6])
    SB_DFF PWMLimit_i0_i14 (.Q(PWMLimit[14]), .C(clk32MHz), .D(n19073));   // verilog/coms.v(127[12] 300[6])
    SB_DFF PWMLimit_i0_i15 (.Q(PWMLimit[15]), .C(clk32MHz), .D(n19072));   // verilog/coms.v(127[12] 300[6])
    SB_DFF PWMLimit_i0_i16 (.Q(PWMLimit[16]), .C(clk32MHz), .D(n19071));   // verilog/coms.v(127[12] 300[6])
    SB_DFF PWMLimit_i0_i17 (.Q(PWMLimit[17]), .C(clk32MHz), .D(n19070));   // verilog/coms.v(127[12] 300[6])
    SB_DFF PWMLimit_i0_i18 (.Q(PWMLimit[18]), .C(clk32MHz), .D(n19069));   // verilog/coms.v(127[12] 300[6])
    SB_DFF PWMLimit_i0_i19 (.Q(PWMLimit[19]), .C(clk32MHz), .D(n19068));   // verilog/coms.v(127[12] 300[6])
    SB_DFF PWMLimit_i0_i20 (.Q(PWMLimit[20]), .C(clk32MHz), .D(n19067));   // verilog/coms.v(127[12] 300[6])
    SB_DFF PWMLimit_i0_i21 (.Q(PWMLimit[21]), .C(clk32MHz), .D(n19066));   // verilog/coms.v(127[12] 300[6])
    SB_DFF PWMLimit_i0_i22 (.Q(PWMLimit[22]), .C(clk32MHz), .D(n19065));   // verilog/coms.v(127[12] 300[6])
    SB_DFF PWMLimit_i0_i23 (.Q(PWMLimit[23]), .C(clk32MHz), .D(n19064));   // verilog/coms.v(127[12] 300[6])
    SB_DFF \FRAME_MATCHER.state_i1  (.Q(\FRAME_MATCHER.state_c [1]), .C(clk32MHz), 
           .D(n38205));   // verilog/coms.v(127[12] 300[6])
    SB_DFF \FRAME_MATCHER.state_i2  (.Q(\FRAME_MATCHER.state_c [2]), .C(clk32MHz), 
           .D(n38206));   // verilog/coms.v(127[12] 300[6])
    SB_DFF \FRAME_MATCHER.state_i0  (.Q(\FRAME_MATCHER.state[0] ), .C(clk32MHz), 
           .D(n32009));   // verilog/coms.v(127[12] 300[6])
    SB_DFF PWMLimit_i0_i0 (.Q(PWMLimit[0]), .C(clk32MHz), .D(n19047));   // verilog/coms.v(127[12] 300[6])
    SB_DFF control_mode_i0_i0 (.Q(control_mode[0]), .C(clk32MHz), .D(n19046));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE setpoint__i2 (.Q(setpoint[2]), .C(clk32MHz), .E(n18646), .D(n5457));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 add_43_3_lut (.I0(n2312), .I1(\FRAME_MATCHER.i [1]), .I2(GND_net), 
            .I3(n27795), .O(n2_adj_4270)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_3_lut.LUT_INIT = 16'h8228;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_30938 (.I0(byte_transmit_counter[1]), 
            .I1(n36291), .I2(n36292), .I3(byte_transmit_counter[2]), .O(n37694));
    defparam byte_transmit_counter_1__bdd_4_lut_30938.LUT_INIT = 16'he4aa;
    SB_CARRY add_43_3 (.CI(n27795), .I0(\FRAME_MATCHER.i [1]), .I1(GND_net), 
            .CO(n27796));
    SB_LUT4 i1_2_lut_3_lut_adj_1328 (.I0(n2_adj_4082), .I1(n2_adj_4272), 
            .I2(\FRAME_MATCHER.state_c [27]), .I3(GND_net), .O(n32219));
    defparam i1_2_lut_3_lut_adj_1328.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_2_lut_adj_1329 (.I0(n17794), .I1(\data_in_frame[4] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n32784));   // verilog/coms.v(75[16:43])
    defparam i1_2_lut_adj_1329.LUT_INIT = 16'h6666;
    SB_DFFE setpoint__i3 (.Q(setpoint[3]), .C(clk32MHz), .E(n18646), .D(n5458));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE setpoint__i4 (.Q(setpoint[4]), .C(clk32MHz), .E(n18646), .D(n5459));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE setpoint__i5 (.Q(setpoint[5]), .C(clk32MHz), .E(n18646), .D(n5460));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE setpoint__i6 (.Q(setpoint[6]), .C(clk32MHz), .E(n18646), .D(n5461));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE setpoint__i7 (.Q(setpoint[7]), .C(clk32MHz), .E(n18646), .D(n5462));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE setpoint__i8 (.Q(setpoint[8]), .C(clk32MHz), .E(n18646), .D(n5463));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE setpoint__i9 (.Q(setpoint[9]), .C(clk32MHz), .E(n18646), .D(n5464));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE setpoint__i10 (.Q(setpoint[10]), .C(clk32MHz), .E(n18646), 
            .D(n5465));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE setpoint__i11 (.Q(setpoint[11]), .C(clk32MHz), .E(n18646), 
            .D(n5466));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE setpoint__i12 (.Q(setpoint[12]), .C(clk32MHz), .E(n18646), 
            .D(n5467));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE setpoint__i13 (.Q(setpoint[13]), .C(clk32MHz), .E(n18646), 
            .D(n5468));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE setpoint__i14 (.Q(setpoint[14]), .C(clk32MHz), .E(n18646), 
            .D(n5469));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE setpoint__i15 (.Q(setpoint[15]), .C(clk32MHz), .E(n18646), 
            .D(n5470));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE setpoint__i16 (.Q(setpoint[16]), .C(clk32MHz), .E(n18646), 
            .D(n5471));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE setpoint__i17 (.Q(setpoint[17]), .C(clk32MHz), .E(n18646), 
            .D(n5472));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE setpoint__i18 (.Q(setpoint[18]), .C(clk32MHz), .E(n18646), 
            .D(n5473));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE setpoint__i19 (.Q(setpoint[19]), .C(clk32MHz), .E(n18646), 
            .D(n5474));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE setpoint__i20 (.Q(setpoint[20]), .C(clk32MHz), .E(n18646), 
            .D(n5475));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE setpoint__i21 (.Q(setpoint[21]), .C(clk32MHz), .E(n18646), 
            .D(n5476));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE setpoint__i22 (.Q(setpoint[22]), .C(clk32MHz), .E(n18646), 
            .D(n5477));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE setpoint__i23 (.Q(setpoint[23]), .C(clk32MHz), .E(n18646), 
            .D(n5478));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i2_3_lut_adj_1330 (.I0(\data_in_frame[0] [2]), .I1(\data_in_frame[0] [1]), 
            .I2(\data_in_frame[2] [3]), .I3(GND_net), .O(n18264));   // verilog/coms.v(75[16:43])
    defparam i2_3_lut_adj_1330.LUT_INIT = 16'h9696;
    SB_LUT4 i3_3_lut_adj_1331 (.I0(n32794), .I1(\data_in_frame[1] [4]), 
            .I2(\data_in_frame[1] [3]), .I3(GND_net), .O(n23_adj_4292));   // verilog/coms.v(73[16:42])
    defparam i3_3_lut_adj_1331.LUT_INIT = 16'h9696;
    SB_LUT4 i11_4_lut_adj_1332 (.I0(n33139), .I1(n32776), .I2(n18235), 
            .I3(n18506), .O(n31_adj_4293));   // verilog/coms.v(73[16:42])
    defparam i11_4_lut_adj_1332.LUT_INIT = 16'h6996;
    SB_DFF data_in_frame_0__i1 (.Q(\data_in_frame[0] [0]), .C(clk32MHz), 
           .D(n19045));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i1_2_lut_3_lut_adj_1333 (.I0(n2_adj_4082), .I1(n2_adj_4272), 
            .I2(\FRAME_MATCHER.state_c [28]), .I3(GND_net), .O(n32221));
    defparam i1_2_lut_3_lut_adj_1333.LUT_INIT = 16'he0e0;
    SB_LUT4 i16_4_lut_adj_1334 (.I0(n31_adj_4293), .I1(n23_adj_4292), .I2(\data_in_frame[4] [2]), 
            .I3(n33293), .O(n36));   // verilog/coms.v(73[16:42])
    defparam i16_4_lut_adj_1334.LUT_INIT = 16'h6996;
    SB_DFF neopxl_color_i0_i0 (.Q(neopxl_color[0]), .C(clk32MHz), .D(n19044));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i14120_3_lut_4_lut (.I0(n8_adj_4090), .I1(n32657), .I2(rx_data[7]), 
            .I3(\data_in_frame[0] [7]), .O(n19262));
    defparam i14120_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFFESR LED_3874 (.Q(LED_c), .C(clk32MHz), .E(n32597), .D(n18858), 
            .R(n33587));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Ki_i0 (.Q(\Ki[0] ), .C(clk32MHz), .D(n19043));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Kp_i0 (.Q(\Kp[0] ), .C(clk32MHz), .D(n19042));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i1 (.Q(\data_in[0] [0]), .C(clk32MHz), .D(n19041));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i14121_3_lut_4_lut (.I0(n8_adj_4090), .I1(n32657), .I2(rx_data[6]), 
            .I3(\data_in_frame[0] [6]), .O(n19263));
    defparam i14121_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i14122_3_lut_4_lut (.I0(n8_adj_4090), .I1(n32657), .I2(rx_data[5]), 
            .I3(\data_in_frame[0] [5]), .O(n19264));
    defparam i14122_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i14123_3_lut_4_lut (.I0(n8_adj_4090), .I1(n32657), .I2(rx_data[4]), 
            .I3(\data_in_frame[0] [4]), .O(n19265));
    defparam i14123_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i14124_3_lut_4_lut (.I0(n8_adj_4090), .I1(n32657), .I2(rx_data[3]), 
            .I3(\data_in_frame[0] [3]), .O(n19266));
    defparam i14124_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i14125_3_lut_4_lut (.I0(n8_adj_4090), .I1(n32657), .I2(rx_data[2]), 
            .I3(\data_in_frame[0] [2]), .O(n19267));
    defparam i14125_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_3_lut_adj_1335 (.I0(n2_adj_4082), .I1(n2_adj_4272), 
            .I2(\FRAME_MATCHER.state_c [29]), .I3(GND_net), .O(n32223));
    defparam i1_2_lut_3_lut_adj_1335.LUT_INIT = 16'he0e0;
    SB_LUT4 i14126_3_lut_4_lut (.I0(n8_adj_4090), .I1(n32657), .I2(rx_data[1]), 
            .I3(\data_in_frame[0] [1]), .O(n19268));
    defparam i14126_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13903_3_lut_4_lut (.I0(n8_adj_4090), .I1(n32657), .I2(rx_data[0]), 
            .I3(\data_in_frame[0] [0]), .O(n19045));
    defparam i13903_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 add_43_2_lut (.I0(n2312), .I1(\FRAME_MATCHER.i [0]), .I2(n161), 
            .I3(GND_net), .O(n2_adj_4022)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_2_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_43_2 (.CI(GND_net), .I0(\FRAME_MATCHER.i [0]), .I1(n161), 
            .CO(n27795));
    SB_LUT4 i1_2_lut_3_lut_adj_1336 (.I0(n2_adj_4082), .I1(n2_adj_4272), 
            .I2(\FRAME_MATCHER.state_c [30]), .I3(GND_net), .O(n32225));
    defparam i1_2_lut_3_lut_adj_1336.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_2_lut_3_lut_adj_1337 (.I0(n2_adj_4082), .I1(n2_adj_4272), 
            .I2(\FRAME_MATCHER.state_c [31]), .I3(GND_net), .O(n32227));
    defparam i1_2_lut_3_lut_adj_1337.LUT_INIT = 16'he0e0;
    SB_LUT4 i15_4_lut_adj_1338 (.I0(n17749), .I1(\data_in_frame[1] [5]), 
            .I2(n32934), .I3(Kp_23__N_843), .O(n35));   // verilog/coms.v(73[16:42])
    defparam i15_4_lut_adj_1338.LUT_INIT = 16'h6996;
    SB_LUT4 i13_4_lut_adj_1339 (.I0(n32916), .I1(n32753), .I2(n32781), 
            .I3(\data_in_frame[4] [6]), .O(n33_adj_4294));   // verilog/coms.v(73[16:42])
    defparam i13_4_lut_adj_1339.LUT_INIT = 16'h6996;
    SB_LUT4 i19_4_lut_adj_1340 (.I0(n33_adj_4294), .I1(n35), .I2(n34_adj_4295), 
            .I3(n36), .O(n30031));   // verilog/coms.v(73[16:42])
    defparam i19_4_lut_adj_1340.LUT_INIT = 16'h6996;
    SB_LUT4 i3_3_lut_adj_1341 (.I0(n30031), .I1(n18264), .I2(n32784), 
            .I3(GND_net), .O(n8_adj_4042));   // verilog/coms.v(73[16:42])
    defparam i3_3_lut_adj_1341.LUT_INIT = 16'h9696;
    SB_LUT4 equal_1577_i7_2_lut (.I0(Kp_23__N_1069), .I1(\data_in_frame[8] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n7_adj_4147));   // verilog/coms.v(236[9:81])
    defparam equal_1577_i7_2_lut.LUT_INIT = 16'h6666;
    SB_DFF driver_enable_3875 (.Q(DE_c), .C(clk32MHz), .D(n32173));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i1_2_lut_3_lut_adj_1342 (.I0(n4452), .I1(n14711), .I2(\FRAME_MATCHER.state[0] ), 
            .I3(GND_net), .O(n4_adj_4083));   // verilog/coms.v(259[6] 261[9])
    defparam i1_2_lut_3_lut_adj_1342.LUT_INIT = 16'h4040;
    SB_DFF IntegralLimit_i0_i1 (.Q(IntegralLimit[1]), .C(clk32MHz), .D(n19581));   // verilog/coms.v(127[12] 300[6])
    SB_DFF IntegralLimit_i0_i2 (.Q(IntegralLimit[2]), .C(clk32MHz), .D(n19580));   // verilog/coms.v(127[12] 300[6])
    SB_DFF IntegralLimit_i0_i3 (.Q(IntegralLimit[3]), .C(clk32MHz), .D(n19579));   // verilog/coms.v(127[12] 300[6])
    SB_DFF IntegralLimit_i0_i4 (.Q(IntegralLimit[4]), .C(clk32MHz), .D(n19578));   // verilog/coms.v(127[12] 300[6])
    SB_DFF IntegralLimit_i0_i5 (.Q(IntegralLimit[5]), .C(clk32MHz), .D(n19577));   // verilog/coms.v(127[12] 300[6])
    SB_DFF IntegralLimit_i0_i6 (.Q(IntegralLimit[6]), .C(clk32MHz), .D(n19576));   // verilog/coms.v(127[12] 300[6])
    SB_DFF IntegralLimit_i0_i7 (.Q(IntegralLimit[7]), .C(clk32MHz), .D(n19575));   // verilog/coms.v(127[12] 300[6])
    SB_DFF IntegralLimit_i0_i8 (.Q(IntegralLimit[8]), .C(clk32MHz), .D(n19574));   // verilog/coms.v(127[12] 300[6])
    SB_DFF IntegralLimit_i0_i9 (.Q(IntegralLimit[9]), .C(clk32MHz), .D(n19573));   // verilog/coms.v(127[12] 300[6])
    SB_DFF IntegralLimit_i0_i10 (.Q(IntegralLimit[10]), .C(clk32MHz), .D(n19572));   // verilog/coms.v(127[12] 300[6])
    SB_DFF IntegralLimit_i0_i11 (.Q(IntegralLimit[11]), .C(clk32MHz), .D(n19571));   // verilog/coms.v(127[12] 300[6])
    SB_DFF IntegralLimit_i0_i12 (.Q(IntegralLimit[12]), .C(clk32MHz), .D(n19570));   // verilog/coms.v(127[12] 300[6])
    SB_DFF IntegralLimit_i0_i13 (.Q(IntegralLimit[13]), .C(clk32MHz), .D(n19569));   // verilog/coms.v(127[12] 300[6])
    SB_DFF IntegralLimit_i0_i14 (.Q(IntegralLimit[14]), .C(clk32MHz), .D(n19568));   // verilog/coms.v(127[12] 300[6])
    SB_DFF IntegralLimit_i0_i15 (.Q(IntegralLimit[15]), .C(clk32MHz), .D(n19567));   // verilog/coms.v(127[12] 300[6])
    SB_DFF IntegralLimit_i0_i16 (.Q(IntegralLimit[16]), .C(clk32MHz), .D(n19566));   // verilog/coms.v(127[12] 300[6])
    SB_DFF IntegralLimit_i0_i17 (.Q(IntegralLimit[17]), .C(clk32MHz), .D(n19565));   // verilog/coms.v(127[12] 300[6])
    SB_DFF IntegralLimit_i0_i18 (.Q(IntegralLimit[18]), .C(clk32MHz), .D(n19564));   // verilog/coms.v(127[12] 300[6])
    SB_DFF IntegralLimit_i0_i19 (.Q(IntegralLimit[19]), .C(clk32MHz), .D(n19563));   // verilog/coms.v(127[12] 300[6])
    SB_DFF IntegralLimit_i0_i20 (.Q(IntegralLimit[20]), .C(clk32MHz), .D(n19562));   // verilog/coms.v(127[12] 300[6])
    SB_DFF IntegralLimit_i0_i21 (.Q(IntegralLimit[21]), .C(clk32MHz), .D(n19561));   // verilog/coms.v(127[12] 300[6])
    SB_DFF IntegralLimit_i0_i22 (.Q(IntegralLimit[22]), .C(clk32MHz), .D(n19560));   // verilog/coms.v(127[12] 300[6])
    SB_DFF IntegralLimit_i0_i23 (.Q(IntegralLimit[23]), .C(clk32MHz), .D(n19559));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i2 (.Q(\data_in[0] [1]), .C(clk32MHz), .D(n19520));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i3 (.Q(\data_in[0] [2]), .C(clk32MHz), .D(n19519));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i4 (.Q(\data_in[0] [3]), .C(clk32MHz), .D(n19518));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i5 (.Q(\data_in[0] [4]), .C(clk32MHz), .D(n19517));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i6 (.Q(\data_in[0] [5]), .C(clk32MHz), .D(n19516));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i7 (.Q(\data_in[0] [6]), .C(clk32MHz), .D(n19515));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i8 (.Q(\data_in[0] [7]), .C(clk32MHz), .D(n19514));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i9 (.Q(\data_in[1] [0]), .C(clk32MHz), .D(n19513));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i10 (.Q(\data_in[1] [1]), .C(clk32MHz), .D(n19512));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i11 (.Q(\data_in[1] [2]), .C(clk32MHz), .D(n19511));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i12 (.Q(\data_in[1] [3]), .C(clk32MHz), .D(n19510));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i13 (.Q(\data_in[1] [4]), .C(clk32MHz), .D(n19509));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i14 (.Q(\data_in[1] [5]), .C(clk32MHz), .D(n19508));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i15 (.Q(\data_in[1] [6]), .C(clk32MHz), .D(n19507));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i16 (.Q(\data_in[1] [7]), .C(clk32MHz), .D(n19506));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i17 (.Q(\data_in[2] [0]), .C(clk32MHz), .D(n19505));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i18 (.Q(\data_in[2] [1]), .C(clk32MHz), .D(n19504));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i19 (.Q(\data_in[2] [2]), .C(clk32MHz), .D(n19503));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i20 (.Q(\data_in[2] [3]), .C(clk32MHz), .D(n19502));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i21 (.Q(\data_in[2] [4]), .C(clk32MHz), .D(n19501));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i22 (.Q(\data_in[2] [5]), .C(clk32MHz), .D(n19500));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i23 (.Q(\data_in[2] [6]), .C(clk32MHz), .D(n19499));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i24 (.Q(\data_in[2] [7]), .C(clk32MHz), .D(n19498));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i25 (.Q(\data_in[3] [0]), .C(clk32MHz), .D(n19497));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i26 (.Q(\data_in[3] [1]), .C(clk32MHz), .D(n19496));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i27 (.Q(\data_in[3] [2]), .C(clk32MHz), .D(n19495));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i28 (.Q(\data_in[3] [3]), .C(clk32MHz), .D(n19494));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i29 (.Q(\data_in[3] [4]), .C(clk32MHz), .D(n19493));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i30 (.Q(\data_in[3] [5]), .C(clk32MHz), .D(n19492));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i31 (.Q(\data_in[3] [6]), .C(clk32MHz), .D(n19491));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i32 (.Q(\data_in[3] [7]), .C(clk32MHz), .D(n19490));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Kp_i1 (.Q(\Kp[1] ), .C(clk32MHz), .D(n19489));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Kp_i2 (.Q(\Kp[2] ), .C(clk32MHz), .D(n19488));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Kp_i3 (.Q(\Kp[3] ), .C(clk32MHz), .D(n19487));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Kp_i4 (.Q(\Kp[4] ), .C(clk32MHz), .D(n19486));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Kp_i5 (.Q(\Kp[5] ), .C(clk32MHz), .D(n19485));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Kp_i6 (.Q(\Kp[6] ), .C(clk32MHz), .D(n19484));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Kp_i7 (.Q(\Kp[7] ), .C(clk32MHz), .D(n19483));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Kp_i8 (.Q(\Kp[8] ), .C(clk32MHz), .D(n19482));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Kp_i9 (.Q(\Kp[9] ), .C(clk32MHz), .D(n19481));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Kp_i10 (.Q(\Kp[10] ), .C(clk32MHz), .D(n19480));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Kp_i11 (.Q(\Kp[11] ), .C(clk32MHz), .D(n19479));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Kp_i12 (.Q(\Kp[12] ), .C(clk32MHz), .D(n19478));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Kp_i13 (.Q(\Kp[13] ), .C(clk32MHz), .D(n19477));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 n37694_bdd_4_lut (.I0(n37694), .I1(n17_adj_4296), .I2(n16_adj_4297), 
            .I3(byte_transmit_counter[2]), .O(n37697));
    defparam n37694_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF Kp_i14 (.Q(\Kp[14] ), .C(clk32MHz), .D(n19476));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Kp_i15 (.Q(\Kp[15] ), .C(clk32MHz), .D(n19475));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Ki_i1 (.Q(\Ki[1] ), .C(clk32MHz), .D(n19474));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Ki_i2 (.Q(\Ki[2] ), .C(clk32MHz), .D(n19473));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Ki_i3 (.Q(\Ki[3] ), .C(clk32MHz), .D(n19472));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Ki_i4 (.Q(\Ki[4] ), .C(clk32MHz), .D(n19471));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1343 (.I0(\data_in_frame[2] [4]), .I1(\data_in_frame[0] [2]), 
            .I2(\data_in_frame[0] [3]), .I3(n18264), .O(Kp_23__N_894));   // verilog/coms.v(75[16:43])
    defparam i1_2_lut_3_lut_4_lut_adj_1343.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1344 (.I0(n63_adj_4106), .I1(n63_adj_4103), 
            .I2(\FRAME_MATCHER.state_c [1]), .I3(GND_net), .O(n123));   // verilog/coms.v(136[7:86])
    defparam i1_2_lut_3_lut_adj_1344.LUT_INIT = 16'h8080;
    SB_DFF Ki_i5 (.Q(\Ki[5] ), .C(clk32MHz), .D(n19470));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Ki_i6 (.Q(\Ki[6] ), .C(clk32MHz), .D(n19469));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Ki_i7 (.Q(\Ki[7] ), .C(clk32MHz), .D(n19468));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Ki_i8 (.Q(\Ki[8] ), .C(clk32MHz), .D(n19467));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Ki_i9 (.Q(\Ki[9] ), .C(clk32MHz), .D(n19466));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Ki_i10 (.Q(\Ki[10] ), .C(clk32MHz), .D(n19465));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1345 (.I0(n4452), .I1(n14711), .I2(\FRAME_MATCHER.state[0] ), 
            .I3(n17551), .O(n2_adj_4272));   // verilog/coms.v(259[6] 261[9])
    defparam i1_2_lut_3_lut_4_lut_adj_1345.LUT_INIT = 16'h0040;
    SB_DFF Ki_i11 (.Q(\Ki[11] ), .C(clk32MHz), .D(n19464));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_30933 (.I0(byte_transmit_counter[1]), 
            .I1(n36296), .I2(n36297), .I3(byte_transmit_counter[2]), .O(n37688));
    defparam byte_transmit_counter_1__bdd_4_lut_30933.LUT_INIT = 16'he4aa;
    SB_LUT4 n37688_bdd_4_lut (.I0(n37688), .I1(n17_adj_4298), .I2(n16_adj_4299), 
            .I3(byte_transmit_counter[2]), .O(n37691));
    defparam n37688_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF Ki_i12 (.Q(\Ki[12] ), .C(clk32MHz), .D(n19463));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Ki_i13 (.Q(\Ki[13] ), .C(clk32MHz), .D(n19462));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Ki_i14 (.Q(\Ki[14] ), .C(clk32MHz), .D(n19461));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Ki_i15 (.Q(\Ki[15] ), .C(clk32MHz), .D(n19452));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i33 (.Q(\data_out_frame[4] [0]), .C(clk32MHz), 
           .D(n19451));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i34 (.Q(\data_out_frame[4] [1]), .C(clk32MHz), 
           .D(n19450));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i35 (.Q(\data_out_frame[4] [2]), .C(clk32MHz), 
           .D(n19449));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i36 (.Q(\data_out_frame[4] [3]), .C(clk32MHz), 
           .D(n19448));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i37 (.Q(\data_out_frame[4] [4]), .C(clk32MHz), 
           .D(n19447));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i38 (.Q(\data_out_frame[4] [5]), .C(clk32MHz), 
           .D(n19446));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i39 (.Q(\data_out_frame[4] [6]), .C(clk32MHz), 
           .D(n19445));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i40 (.Q(\data_out_frame[4] [7]), .C(clk32MHz), 
           .D(n19444));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i41 (.Q(\data_out_frame[5] [0]), .C(clk32MHz), 
           .D(n19443));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i42 (.Q(\data_out_frame[5] [1]), .C(clk32MHz), 
           .D(n19442));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i43 (.Q(\data_out_frame[5] [2]), .C(clk32MHz), 
           .D(n19441));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i44 (.Q(\data_out_frame[5] [3]), .C(clk32MHz), 
           .D(n19440));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i45 (.Q(\data_out_frame[5] [4]), .C(clk32MHz), 
           .D(n19439));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i46 (.Q(\data_out_frame[5] [5]), .C(clk32MHz), 
           .D(n19438));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i47 (.Q(\data_out_frame[5] [6]), .C(clk32MHz), 
           .D(n19437));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i48 (.Q(\data_out_frame[5] [7]), .C(clk32MHz), 
           .D(n19436));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i49 (.Q(\data_out_frame[6] [0]), .C(clk32MHz), 
           .D(n19435));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i50 (.Q(\data_out_frame[6] [1]), .C(clk32MHz), 
           .D(n19434));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i51 (.Q(\data_out_frame[6] [2]), .C(clk32MHz), 
           .D(n19433));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i52 (.Q(\data_out_frame[6] [3]), .C(clk32MHz), 
           .D(n19432));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i53 (.Q(\data_out_frame[6] [4]), .C(clk32MHz), 
           .D(n19431));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i54 (.Q(\data_out_frame[6] [5]), .C(clk32MHz), 
           .D(n19430));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i55 (.Q(\data_out_frame[6] [6]), .C(clk32MHz), 
           .D(n19429));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i56 (.Q(\data_out_frame[6] [7]), .C(clk32MHz), 
           .D(n19428));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i57 (.Q(\data_out_frame[7] [0]), .C(clk32MHz), 
           .D(n19427));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i58 (.Q(\data_out_frame[7] [1]), .C(clk32MHz), 
           .D(n19426));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i59 (.Q(\data_out_frame[7] [2]), .C(clk32MHz), 
           .D(n19425));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i60 (.Q(\data_out_frame[7] [3]), .C(clk32MHz), 
           .D(n19424));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i61 (.Q(\data_out_frame[7] [4]), .C(clk32MHz), 
           .D(n19423));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i62 (.Q(\data_out_frame[7] [5]), .C(clk32MHz), 
           .D(n19422));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i63 (.Q(\data_out_frame[7] [6]), .C(clk32MHz), 
           .D(n19421));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i64 (.Q(\data_out_frame[7] [7]), .C(clk32MHz), 
           .D(n19420));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i65 (.Q(\data_out_frame[8] [0]), .C(clk32MHz), 
           .D(n19419));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i66 (.Q(\data_out_frame[8] [1]), .C(clk32MHz), 
           .D(n19418));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i1_2_lut_3_lut_adj_1346 (.I0(\data_in_frame[2] [4]), .I1(\data_in_frame[0] [2]), 
            .I2(\data_in_frame[0] [3]), .I3(GND_net), .O(n17794));   // verilog/coms.v(166[9:87])
    defparam i1_2_lut_3_lut_adj_1346.LUT_INIT = 16'h9696;
    SB_DFF data_out_frame_0___i67 (.Q(\data_out_frame[8] [2]), .C(clk32MHz), 
           .D(n19417));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i68 (.Q(\data_out_frame[8] [3]), .C(clk32MHz), 
           .D(n19416));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i69 (.Q(\data_out_frame[8] [4]), .C(clk32MHz), 
           .D(n19415));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i70 (.Q(\data_out_frame[8] [5]), .C(clk32MHz), 
           .D(n19414));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i71 (.Q(\data_out_frame[8] [6]), .C(clk32MHz), 
           .D(n19413));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i72 (.Q(\data_out_frame[8] [7]), .C(clk32MHz), 
           .D(n19412));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i73 (.Q(\data_out_frame[9] [0]), .C(clk32MHz), 
           .D(n19411));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i74 (.Q(\data_out_frame[9] [1]), .C(clk32MHz), 
           .D(n19410));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i75 (.Q(\data_out_frame[9] [2]), .C(clk32MHz), 
           .D(n19409));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i76 (.Q(\data_out_frame[9] [3]), .C(clk32MHz), 
           .D(n19408));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i77 (.Q(\data_out_frame[9] [4]), .C(clk32MHz), 
           .D(n19407));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i78 (.Q(\data_out_frame[9] [5]), .C(clk32MHz), 
           .D(n19406));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i79 (.Q(\data_out_frame[9] [6]), .C(clk32MHz), 
           .D(n19405));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i80 (.Q(\data_out_frame[9] [7]), .C(clk32MHz), 
           .D(n19404));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i81 (.Q(\data_out_frame[10] [0]), .C(clk32MHz), 
           .D(n19403));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i82 (.Q(\data_out_frame[10] [1]), .C(clk32MHz), 
           .D(n19402));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i83 (.Q(\data_out_frame[10] [2]), .C(clk32MHz), 
           .D(n19401));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i84 (.Q(\data_out_frame[10] [3]), .C(clk32MHz), 
           .D(n19400));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i85 (.Q(\data_out_frame[10] [4]), .C(clk32MHz), 
           .D(n19399));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i86 (.Q(\data_out_frame[10] [5]), .C(clk32MHz), 
           .D(n19398));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i87 (.Q(\data_out_frame[10] [6]), .C(clk32MHz), 
           .D(n19397));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i88 (.Q(\data_out_frame[10] [7]), .C(clk32MHz), 
           .D(n19396));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i89 (.Q(\data_out_frame[11] [0]), .C(clk32MHz), 
           .D(n19395));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i90 (.Q(\data_out_frame[11] [1]), .C(clk32MHz), 
           .D(n19394));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i91 (.Q(\data_out_frame[11] [2]), .C(clk32MHz), 
           .D(n19393));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i92 (.Q(\data_out_frame[11] [3]), .C(clk32MHz), 
           .D(n19392));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i93 (.Q(\data_out_frame[11] [4]), .C(clk32MHz), 
           .D(n19391));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i94 (.Q(\data_out_frame[11] [5]), .C(clk32MHz), 
           .D(n19390));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i95 (.Q(\data_out_frame[11] [6]), .C(clk32MHz), 
           .D(n19389));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i96 (.Q(\data_out_frame[11] [7]), .C(clk32MHz), 
           .D(n19388));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i97 (.Q(\data_out_frame[12] [0]), .C(clk32MHz), 
           .D(n19387));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i98 (.Q(\data_out_frame[12] [1]), .C(clk32MHz), 
           .D(n19386));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i99 (.Q(\data_out_frame[12] [2]), .C(clk32MHz), 
           .D(n19385));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i100 (.Q(\data_out_frame[12] [3]), .C(clk32MHz), 
           .D(n19384));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i101 (.Q(\data_out_frame[12] [4]), .C(clk32MHz), 
           .D(n19383));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i1_2_lut_4_lut_adj_1347 (.I0(\data_in_frame[2] [4]), .I1(n32710), 
            .I2(n18264), .I3(n33353), .O(n32794));   // verilog/coms.v(70[16:27])
    defparam i1_2_lut_4_lut_adj_1347.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_1348 (.I0(\data_in_frame[5] [6]), .I1(\data_in_frame[1] [5]), 
            .I2(\data_in_frame[1] [4]), .I3(\data_in_frame[5] [7]), .O(n18506));
    defparam i2_3_lut_4_lut_adj_1348.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_1349 (.I0(\data_out_frame[15] [5]), .I1(n33218), 
            .I2(\data_out_frame[13] [1]), .I3(n17086), .O(n33034));
    defparam i2_3_lut_4_lut_adj_1349.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1350 (.I0(n63_adj_4106), .I1(n63_adj_4103), 
            .I2(n63), .I3(GND_net), .O(n14711));   // verilog/coms.v(136[7:86])
    defparam i1_2_lut_3_lut_adj_1350.LUT_INIT = 16'h8080;
    SB_LUT4 i1_2_lut_3_lut_adj_1351 (.I0(n18086), .I1(n32816), .I2(n30139), 
            .I3(GND_net), .O(n30170));
    defparam i1_2_lut_3_lut_adj_1351.LUT_INIT = 16'h9696;
    SB_LUT4 i30507_3_lut_4_lut (.I0(n17559), .I1(n63_adj_8), .I2(tx_active), 
            .I3(r_SM_Main_2__N_3490[0]), .O(n18619));
    defparam i30507_3_lut_4_lut.LUT_INIT = 16'h3337;
    SB_LUT4 i13984_3_lut_4_lut (.I0(n8_adj_4300), .I1(n32678), .I2(rx_data[7]), 
            .I3(\data_in_frame[17] [7]), .O(n19126));
    defparam i13984_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13985_3_lut_4_lut (.I0(n8_adj_4300), .I1(n32678), .I2(rx_data[6]), 
            .I3(\data_in_frame[17] [6]), .O(n19127));
    defparam i13985_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_3_lut_adj_1352 (.I0(\state[0] ), .I1(\state[2] ), .I2(\state[3] ), 
            .I3(GND_net), .O(n5690));
    defparam i1_2_lut_3_lut_adj_1352.LUT_INIT = 16'h0202;
    SB_DFF data_out_frame_0___i102 (.Q(\data_out_frame[12] [5]), .C(clk32MHz), 
           .D(n19382));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i13986_3_lut_4_lut (.I0(n8_adj_4300), .I1(n32678), .I2(rx_data[5]), 
            .I3(\data_in_frame[17] [5]), .O(n19128));
    defparam i13986_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF data_out_frame_0___i103 (.Q(\data_out_frame[12] [6]), .C(clk32MHz), 
           .D(n19381));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i13987_3_lut_4_lut (.I0(n8_adj_4300), .I1(n32678), .I2(rx_data[4]), 
            .I3(\data_in_frame[17] [4]), .O(n19129));
    defparam i13987_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_3_lut_4_lut_adj_1353 (.I0(tx_transmit_N_3387), .I1(n23740), 
            .I2(n14711), .I3(n17559), .O(n2_adj_4082));   // verilog/coms.v(213[6] 220[9])
    defparam i1_3_lut_4_lut_adj_1353.LUT_INIT = 16'h00e0;
    SB_LUT4 i2_2_lut_4_lut (.I0(\FRAME_MATCHER.state_c [2]), .I1(\FRAME_MATCHER.state_c [1]), 
            .I2(\FRAME_MATCHER.state[0] ), .I3(n32655), .O(n5592));
    defparam i2_2_lut_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_3_lut_adj_1354 (.I0(tx_transmit_N_3387), .I1(n23740), 
            .I2(n17559), .I3(GND_net), .O(n32));   // verilog/coms.v(213[6] 220[9])
    defparam i1_2_lut_3_lut_adj_1354.LUT_INIT = 16'h0e0e;
    SB_LUT4 i13988_3_lut_4_lut (.I0(n8_adj_4300), .I1(n32678), .I2(rx_data[3]), 
            .I3(\data_in_frame[17] [3]), .O(n19130));
    defparam i13988_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF data_out_frame_0___i104 (.Q(\data_out_frame[12] [7]), .C(clk32MHz), 
           .D(n19380));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i105 (.Q(\data_out_frame[13] [0]), .C(clk32MHz), 
           .D(n19379));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i13989_3_lut_4_lut (.I0(n8_adj_4300), .I1(n32678), .I2(rx_data[2]), 
            .I3(\data_in_frame[17] [2]), .O(n19131));
    defparam i13989_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF data_out_frame_0___i106 (.Q(\data_out_frame[13] [1]), .C(clk32MHz), 
           .D(n19378));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i107 (.Q(\data_out_frame[13] [2]), .C(clk32MHz), 
           .D(n19377));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i13990_3_lut_4_lut (.I0(n8_adj_4300), .I1(n32678), .I2(rx_data[1]), 
            .I3(\data_in_frame[17] [1]), .O(n19132));
    defparam i13990_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i18661_2_lut_3_lut (.I0(n24499), .I1(rx_data_ready), .I2(\FRAME_MATCHER.rx_data_ready_prev ), 
            .I3(GND_net), .O(n23788));
    defparam i18661_2_lut_3_lut.LUT_INIT = 16'h0404;
    SB_LUT4 i1_2_lut_3_lut_adj_1355 (.I0(n2_adj_4085), .I1(n3_adj_4084), 
            .I2(n2_adj_4082), .I3(GND_net), .O(n32677));
    defparam i1_2_lut_3_lut_adj_1355.LUT_INIT = 16'hfefe;
    SB_LUT4 i13991_3_lut_4_lut (.I0(n8_adj_4300), .I1(n32678), .I2(rx_data[0]), 
            .I3(\data_in_frame[17] [0]), .O(n19133));
    defparam i13991_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13976_3_lut_4_lut (.I0(n8_adj_4302), .I1(n32678), .I2(rx_data[7]), 
            .I3(\data_in_frame[18] [7]), .O(n19118));
    defparam i13976_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13977_3_lut_4_lut (.I0(n8_adj_4302), .I1(n32678), .I2(rx_data[6]), 
            .I3(\data_in_frame[18] [6]), .O(n19119));
    defparam i13977_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13978_3_lut_4_lut (.I0(n8_adj_4302), .I1(n32678), .I2(rx_data[5]), 
            .I3(\data_in_frame[18] [5]), .O(n19120));
    defparam i13978_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13979_3_lut_4_lut (.I0(n8_adj_4302), .I1(n32678), .I2(rx_data[4]), 
            .I3(\data_in_frame[18] [4]), .O(n19121));
    defparam i13979_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13980_3_lut_4_lut (.I0(n8_adj_4302), .I1(n32678), .I2(rx_data[3]), 
            .I3(\data_in_frame[18] [3]), .O(n19122));
    defparam i13980_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13981_3_lut_4_lut (.I0(n8_adj_4302), .I1(n32678), .I2(rx_data[2]), 
            .I3(\data_in_frame[18] [2]), .O(n19123));
    defparam i13981_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13982_3_lut_4_lut (.I0(n8_adj_4302), .I1(n32678), .I2(rx_data[1]), 
            .I3(\data_in_frame[18] [1]), .O(n19124));
    defparam i13982_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13983_3_lut_4_lut (.I0(n8_adj_4302), .I1(n32678), .I2(rx_data[0]), 
            .I3(\data_in_frame[18] [0]), .O(n19125));
    defparam i13983_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 equal_134_i8_2_lut_3_lut (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(\FRAME_MATCHER.i [0]), .I3(GND_net), .O(n8_adj_4302));   // verilog/coms.v(154[7:23])
    defparam equal_134_i8_2_lut_3_lut.LUT_INIT = 16'hfdfd;
    SB_LUT4 equal_125_i8_2_lut_3_lut (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(\FRAME_MATCHER.i [0]), .I3(GND_net), .O(n8_adj_4303));   // verilog/coms.v(154[7:23])
    defparam equal_125_i8_2_lut_3_lut.LUT_INIT = 16'hdfdf;
    SB_LUT4 i13968_3_lut_4_lut (.I0(n8_adj_4303), .I1(n32678), .I2(rx_data[7]), 
            .I3(\data_in_frame[19] [7]), .O(n19110));
    defparam i13968_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13969_3_lut_4_lut (.I0(n8_adj_4303), .I1(n32678), .I2(rx_data[6]), 
            .I3(\data_in_frame[19] [6]), .O(n19111));
    defparam i13969_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13970_3_lut_4_lut (.I0(n8_adj_4303), .I1(n32678), .I2(rx_data[5]), 
            .I3(\data_in_frame[19] [5]), .O(n19112));
    defparam i13970_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13971_3_lut_4_lut (.I0(n8_adj_4303), .I1(n32678), .I2(rx_data[4]), 
            .I3(\data_in_frame[19] [4]), .O(n19113));
    defparam i13971_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_3_lut_adj_1356 (.I0(\data_in_frame[0] [1]), .I1(\data_in_frame[0] [6]), 
            .I2(\data_in_frame[0] [5]), .I3(GND_net), .O(n6_adj_4229));   // verilog/coms.v(70[16:27])
    defparam i1_2_lut_3_lut_adj_1356.LUT_INIT = 16'h9696;
    SB_DFF data_out_frame_0___i108 (.Q(\data_out_frame[13] [3]), .C(clk32MHz), 
           .D(n19376));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i109 (.Q(\data_out_frame[13] [4]), .C(clk32MHz), 
           .D(n19375));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i2_2_lut_3_lut (.I0(\data_in_frame[3] [1]), .I1(\data_in_frame[5] [1]), 
            .I2(\data_in_frame[4] [7]), .I3(GND_net), .O(n10_adj_4228));   // verilog/coms.v(71[16:69])
    defparam i2_2_lut_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 i13972_3_lut_4_lut (.I0(n8_adj_4303), .I1(n32678), .I2(rx_data[3]), 
            .I3(\data_in_frame[19] [3]), .O(n19114));
    defparam i13972_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_3_lut_adj_1357 (.I0(\data_in_frame[1] [2]), .I1(\data_in_frame[3] [4]), 
            .I2(\data_in_frame[1] [4]), .I3(GND_net), .O(n6_adj_4226));
    defparam i1_2_lut_3_lut_adj_1357.LUT_INIT = 16'h9696;
    SB_DFF data_out_frame_0___i110 (.Q(\data_out_frame[13] [5]), .C(clk32MHz), 
           .D(n19374));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i111 (.Q(\data_out_frame[13] [6]), .C(clk32MHz), 
           .D(n19373));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i112 (.Q(\data_out_frame[13] [7]), .C(clk32MHz), 
           .D(n19372));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i13973_3_lut_4_lut (.I0(n8_adj_4303), .I1(n32678), .I2(rx_data[2]), 
            .I3(\data_in_frame[19] [2]), .O(n19115));
    defparam i13973_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF data_out_frame_0___i113 (.Q(\data_out_frame[14] [0]), .C(clk32MHz), 
           .D(n19371));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i114 (.Q(\data_out_frame[14] [1]), .C(clk32MHz), 
           .D(n19370));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i115 (.Q(\data_out_frame[14] [2]), .C(clk32MHz), 
           .D(n19369));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i19369_2_lut_4_lut (.I0(n2_adj_4085), .I1(n3_adj_4084), .I2(n1), 
            .I3(\FRAME_MATCHER.state_c [8]), .O(n24506));
    defparam i19369_2_lut_4_lut.LUT_INIT = 16'hfe00;
    SB_DFF data_out_frame_0___i116 (.Q(\data_out_frame[14] [3]), .C(clk32MHz), 
           .D(n19368));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i1_2_lut_4_lut_adj_1358 (.I0(\data_in_frame[6] [7]), .I1(\data_in_frame[6] [2]), 
            .I2(n10_adj_4194), .I3(\data_in_frame[6] [5]), .O(Kp_23__N_804));   // verilog/coms.v(85[17:28])
    defparam i1_2_lut_4_lut_adj_1358.LUT_INIT = 16'h6996;
    SB_DFF data_out_frame_0___i117 (.Q(\data_out_frame[14] [4]), .C(clk32MHz), 
           .D(n19367));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i2_3_lut_4_lut_adj_1359 (.I0(n18268), .I1(\data_in_frame[2] [4]), 
            .I2(n32710), .I3(\data_in_frame[4] [6]), .O(n32791));   // verilog/coms.v(74[16:43])
    defparam i2_3_lut_4_lut_adj_1359.LUT_INIT = 16'h6996;
    SB_DFF data_out_frame_0___i118 (.Q(\data_out_frame[14] [5]), .C(clk32MHz), 
           .D(n19366));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i119 (.Q(\data_out_frame[14] [6]), .C(clk32MHz), 
           .D(n19365));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i120 (.Q(\data_out_frame[14] [7]), .C(clk32MHz), 
           .D(n19364));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i2_2_lut_3_lut_adj_1360 (.I0(\data_in_frame[5] [4]), .I1(n33057), 
            .I2(n4_adj_4179), .I3(GND_net), .O(n32781));
    defparam i2_2_lut_3_lut_adj_1360.LUT_INIT = 16'h9696;
    SB_DFF data_out_frame_0___i121 (.Q(\data_out_frame[15] [0]), .C(clk32MHz), 
           .D(n19363));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i122 (.Q(\data_out_frame[15] [1]), .C(clk32MHz), 
           .D(n19362));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i123 (.Q(\data_out_frame[15] [2]), .C(clk32MHz), 
           .D(n19361));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i124 (.Q(\data_out_frame[15] [3]), .C(clk32MHz), 
           .D(n19360));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i125 (.Q(\data_out_frame[15] [4]), .C(clk32MHz), 
           .D(n19359));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i126 (.Q(\data_out_frame[15] [5]), .C(clk32MHz), 
           .D(n19358));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i127 (.Q(\data_out_frame[15] [6]), .C(clk32MHz), 
           .D(n19357));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i128 (.Q(\data_out_frame[15] [7]), .C(clk32MHz), 
           .D(n19356));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i129 (.Q(\data_out_frame[16] [0]), .C(clk32MHz), 
           .D(n19355));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i130 (.Q(\data_out_frame[16] [1]), .C(clk32MHz), 
           .D(n19354));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i131 (.Q(\data_out_frame[16] [2]), .C(clk32MHz), 
           .D(n19353));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i132 (.Q(\data_out_frame[16] [3]), .C(clk32MHz), 
           .D(n19352));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i133 (.Q(\data_out_frame[16] [4]), .C(clk32MHz), 
           .D(n19351));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i134 (.Q(\data_out_frame[16] [5]), .C(clk32MHz), 
           .D(n19350));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i135 (.Q(\data_out_frame[16] [6]), .C(clk32MHz), 
           .D(n19349));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i136 (.Q(\data_out_frame[16] [7]), .C(clk32MHz), 
           .D(n19348));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i137 (.Q(\data_out_frame[17] [0]), .C(clk32MHz), 
           .D(n19347));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i138 (.Q(\data_out_frame[17] [1]), .C(clk32MHz), 
           .D(n19346));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i139 (.Q(\data_out_frame[17] [2]), .C(clk32MHz), 
           .D(n19345));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i140 (.Q(\data_out_frame[17] [3]), .C(clk32MHz), 
           .D(n19344));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i141 (.Q(\data_out_frame[17] [4]), .C(clk32MHz), 
           .D(n19343));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i142 (.Q(\data_out_frame[17] [5]), .C(clk32MHz), 
           .D(n19342));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i143 (.Q(\data_out_frame[17] [6]), .C(clk32MHz), 
           .D(n19341));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i144 (.Q(\data_out_frame[17] [7]), .C(clk32MHz), 
           .D(n19340));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i145 (.Q(\data_out_frame[18] [0]), .C(clk32MHz), 
           .D(n19339));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i146 (.Q(\data_out_frame[18] [1]), .C(clk32MHz), 
           .D(n19338));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i147 (.Q(\data_out_frame[18] [2]), .C(clk32MHz), 
           .D(n19337));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i148 (.Q(\data_out_frame[18] [3]), .C(clk32MHz), 
           .D(n19336));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i149 (.Q(\data_out_frame[18] [4]), .C(clk32MHz), 
           .D(n19335));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i150 (.Q(\data_out_frame[18] [5]), .C(clk32MHz), 
           .D(n19334));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i151 (.Q(\data_out_frame[18] [6]), .C(clk32MHz), 
           .D(n19333));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i1_2_lut_4_lut_adj_1361 (.I0(n2_adj_4085), .I1(n3_adj_4084), 
            .I2(n1), .I3(\FRAME_MATCHER.state_c [12]), .O(n31999));
    defparam i1_2_lut_4_lut_adj_1361.LUT_INIT = 16'hfe00;
    SB_DFF data_out_frame_0___i152 (.Q(\data_out_frame[18] [7]), .C(clk32MHz), 
           .D(n19332));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i153 (.Q(\data_out_frame[19] [0]), .C(clk32MHz), 
           .D(n19331));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i154 (.Q(\data_out_frame[19] [1]), .C(clk32MHz), 
           .D(n19330));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i155 (.Q(\data_out_frame[19] [2]), .C(clk32MHz), 
           .D(n19329));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i156 (.Q(\data_out_frame[19] [3]), .C(clk32MHz), 
           .D(n19328));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i157 (.Q(\data_out_frame[19] [4]), .C(clk32MHz), 
           .D(n19327));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i158 (.Q(\data_out_frame[19] [5]), .C(clk32MHz), 
           .D(n19326));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i159 (.Q(\data_out_frame[19] [6]), .C(clk32MHz), 
           .D(n19325));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i13974_3_lut_4_lut (.I0(n8_adj_4303), .I1(n32678), .I2(rx_data[1]), 
            .I3(\data_in_frame[19] [1]), .O(n19116));
    defparam i13974_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF data_out_frame_0___i160 (.Q(\data_out_frame[19] [7]), .C(clk32MHz), 
           .D(n19324));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i161 (.Q(\data_out_frame[20] [0]), .C(clk32MHz), 
           .D(n19323));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i162 (.Q(\data_out_frame[20] [1]), .C(clk32MHz), 
           .D(n19322));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i163 (.Q(\data_out_frame[20] [2]), .C(clk32MHz), 
           .D(n19321));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i164 (.Q(\data_out_frame[20] [3]), .C(clk32MHz), 
           .D(n19320));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i165 (.Q(\data_out_frame[20] [4]), .C(clk32MHz), 
           .D(n19319));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i2_2_lut_3_lut_adj_1362 (.I0(\data_in_frame[3] [6]), .I1(\data_in_frame[6] [2]), 
            .I2(\data_in_frame[2] [0]), .I3(GND_net), .O(n10_adj_4188));   // verilog/coms.v(75[16:27])
    defparam i2_2_lut_3_lut_adj_1362.LUT_INIT = 16'h9696;
    SB_DFF data_out_frame_0___i166 (.Q(\data_out_frame[20] [5]), .C(clk32MHz), 
           .D(n19318));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i2_2_lut_4_lut_adj_1363 (.I0(n18460), .I1(\data_in_frame[13] [2]), 
            .I2(n30624), .I3(\data_in_frame[10] [6]), .O(n10_adj_4184));
    defparam i2_2_lut_4_lut_adj_1363.LUT_INIT = 16'h6996;
    SB_DFF data_out_frame_0___i167 (.Q(\data_out_frame[20] [6]), .C(clk32MHz), 
           .D(n19317));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i13975_3_lut_4_lut (.I0(n8_adj_4303), .I1(n32678), .I2(rx_data[0]), 
            .I3(\data_in_frame[19] [0]), .O(n19117));
    defparam i13975_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF data_out_frame_0___i168 (.Q(\data_out_frame[20] [7]), .C(clk32MHz), 
           .D(n19316));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i185 (.Q(\data_out_frame[23] [0]), .C(clk32MHz), 
           .D(n19315));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i5_3_lut_4_lut (.I0(n18285), .I1(\data_in_frame[7] [6]), .I2(n32781), 
            .I3(Kp_23__N_1063), .O(n14_adj_4181));
    defparam i5_3_lut_4_lut.LUT_INIT = 16'h6996;
    SB_DFF data_out_frame_0___i186 (.Q(\data_out_frame[23] [1]), .C(clk32MHz), 
           .D(n19314));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i187 (.Q(\data_out_frame[23] [2]), .C(clk32MHz), 
           .D(n19313));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i188 (.Q(\data_out_frame[23] [3]), .C(clk32MHz), 
           .D(n19312));   // verilog/coms.v(127[12] 300[6])
    SB_DFF IntegralLimit_i0_i0 (.Q(IntegralLimit[0]), .C(clk32MHz), .D(n19023));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i189 (.Q(\data_out_frame[23] [4]), .C(clk32MHz), 
           .D(n19311));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i190 (.Q(\data_out_frame[23] [5]), .C(clk32MHz), 
           .D(n19310));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i191 (.Q(\data_out_frame[23] [6]), .C(clk32MHz), 
           .D(n19309));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i192 (.Q(\data_out_frame[23] [7]), .C(clk32MHz), 
           .D(n19308));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i193 (.Q(\data_out_frame[24] [0]), .C(clk32MHz), 
           .D(n19307));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i194 (.Q(\data_out_frame[24] [1]), .C(clk32MHz), 
           .D(n19306));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i195 (.Q(\data_out_frame[24] [2]), .C(clk32MHz), 
           .D(n19305));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i196 (.Q(\data_out_frame[24] [3]), .C(clk32MHz), 
           .D(n19304));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i197 (.Q(\data_out_frame[24] [4]), .C(clk32MHz), 
           .D(n19303));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i198 (.Q(\data_out_frame[24] [5]), .C(clk32MHz), 
           .D(n19302));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i199 (.Q(\data_out_frame[24] [6]), .C(clk32MHz), 
           .D(n19301));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i200 (.Q(\data_out_frame[24] [7]), .C(clk32MHz), 
           .D(n19300));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i201 (.Q(\data_out_frame[25] [0]), .C(clk32MHz), 
           .D(n19299));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i202 (.Q(\data_out_frame[25] [1]), .C(clk32MHz), 
           .D(n19298));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i203 (.Q(\data_out_frame[25] [2]), .C(clk32MHz), 
           .D(n19297));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i204 (.Q(\data_out_frame[25] [3]), .C(clk32MHz), 
           .D(n19296));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i205 (.Q(\data_out_frame[25] [4]), .C(clk32MHz), 
           .D(n19295));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i206 (.Q(\data_out_frame[25] [5]), .C(clk32MHz), 
           .D(n19294));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i207 (.Q(\data_out_frame[25] [6]), .C(clk32MHz), 
           .D(n19293));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i208 (.Q(\data_out_frame[25] [7]), .C(clk32MHz), 
           .D(n19292));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i1 (.Q(neopxl_color[1]), .C(clk32MHz), .D(n19291));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i2 (.Q(neopxl_color[2]), .C(clk32MHz), .D(n19290));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i3 (.Q(neopxl_color[3]), .C(clk32MHz), .D(n19289));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i4 (.Q(neopxl_color[4]), .C(clk32MHz), .D(n19288));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i5 (.Q(neopxl_color[5]), .C(clk32MHz), .D(n19287));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i6 (.Q(neopxl_color[6]), .C(clk32MHz), .D(n19286));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i7 (.Q(neopxl_color[7]), .C(clk32MHz), .D(n19285));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i8 (.Q(neopxl_color[8]), .C(clk32MHz), .D(n19284));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i9 (.Q(neopxl_color[9]), .C(clk32MHz), .D(n19283));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i10 (.Q(neopxl_color[10]), .C(clk32MHz), .D(n19282));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i11 (.Q(neopxl_color[11]), .C(clk32MHz), .D(n19281));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i12 (.Q(neopxl_color[12]), .C(clk32MHz), .D(n19280));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i13 (.Q(neopxl_color[13]), .C(clk32MHz), .D(n19279));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i14 (.Q(neopxl_color[14]), .C(clk32MHz), .D(n19278));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i15 (.Q(neopxl_color[15]), .C(clk32MHz), .D(n19277));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i28577_2_lut (.I0(\FRAME_MATCHER.state [3]), .I1(\FRAME_MATCHER.state_c [2]), 
            .I2(GND_net), .I3(GND_net), .O(n35330));
    defparam i28577_2_lut.LUT_INIT = 16'heeee;
    SB_DFF neopxl_color_i0_i16 (.Q(neopxl_color[16]), .C(clk32MHz), .D(n19276));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i17 (.Q(neopxl_color[17]), .C(clk32MHz), .D(n19275));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i1_4_lut_adj_1364 (.I0(\FRAME_MATCHER.state_c [1]), .I1(n32564), 
            .I2(n35330), .I3(\FRAME_MATCHER.state[0] ), .O(n14557));
    defparam i1_4_lut_adj_1364.LUT_INIT = 16'hccce;
    SB_DFF neopxl_color_i0_i18 (.Q(neopxl_color[18]), .C(clk32MHz), .D(n19274));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i3_4_lut_adj_1365 (.I0(n14557), .I1(n32655), .I2(\FRAME_MATCHER.state_c [1]), 
            .I3(\FRAME_MATCHER.state_31__N_2598 [3]), .O(n14867));   // verilog/coms.v(127[12] 300[6])
    defparam i3_4_lut_adj_1365.LUT_INIT = 16'h2000;
    SB_DFF neopxl_color_i0_i19 (.Q(neopxl_color[19]), .C(clk32MHz), .D(n19273));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i1_3_lut_4_lut_adj_1366 (.I0(\data_in_frame[1] [3]), .I1(\data_in_frame[5] [5]), 
            .I2(\data_in_frame[1] [2]), .I3(\data_in_frame[3] [4]), .O(n4_adj_4179));
    defparam i1_3_lut_4_lut_adj_1366.LUT_INIT = 16'h6996;
    SB_DFF neopxl_color_i0_i20 (.Q(neopxl_color[20]), .C(clk32MHz), .D(n19272));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i21 (.Q(neopxl_color[21]), .C(clk32MHz), .D(n19271));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i22 (.Q(neopxl_color[22]), .C(clk32MHz), .D(n19270));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i23 (.Q(neopxl_color[23]), .C(clk32MHz), .D(n19269));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i2 (.Q(\data_in_frame[0] [1]), .C(clk32MHz), 
           .D(n19268));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i3 (.Q(\data_in_frame[0] [2]), .C(clk32MHz), 
           .D(n19267));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i4 (.Q(\data_in_frame[0] [3]), .C(clk32MHz), 
           .D(n19266));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i5 (.Q(\data_in_frame[0] [4]), .C(clk32MHz), 
           .D(n19265));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i6 (.Q(\data_in_frame[0] [5]), .C(clk32MHz), 
           .D(n19264));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i7 (.Q(\data_in_frame[0] [6]), .C(clk32MHz), 
           .D(n19263));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i8 (.Q(\data_in_frame[0] [7]), .C(clk32MHz), 
           .D(n19262));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i9 (.Q(\data_in_frame[1] [0]), .C(clk32MHz), 
           .D(n19261));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i10 (.Q(\data_in_frame[1] [1]), .C(clk32MHz), 
           .D(n19260));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i11 (.Q(\data_in_frame[1] [2]), .C(clk32MHz), 
           .D(n19259));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i12 (.Q(\data_in_frame[1] [3]), .C(clk32MHz), 
           .D(n19258));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i13 (.Q(\data_in_frame[1] [4]), .C(clk32MHz), 
           .D(n19257));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i2_3_lut_4_lut_adj_1367 (.I0(\data_in_frame[9] [5]), .I1(n30545), 
            .I2(n17885), .I3(n30872), .O(n15920));
    defparam i2_3_lut_4_lut_adj_1367.LUT_INIT = 16'h6996;
    SB_DFF data_in_frame_0__i14 (.Q(\data_in_frame[1] [5]), .C(clk32MHz), 
           .D(n19256));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i15 (.Q(\data_in_frame[1] [6]), .C(clk32MHz), 
           .D(n19255));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i16 (.Q(\data_in_frame[1] [7]), .C(clk32MHz), 
           .D(n19254));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i17 (.Q(\data_in_frame[2] [0]), .C(clk32MHz), 
           .D(n19253));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i1_2_lut_3_lut_adj_1368 (.I0(\data_in_frame[9] [2]), .I1(n17827), 
            .I2(n17846), .I3(GND_net), .O(n32824));   // verilog/coms.v(73[16:42])
    defparam i1_2_lut_3_lut_adj_1368.LUT_INIT = 16'h9696;
    SB_DFF data_in_frame_0__i18 (.Q(\data_in_frame[2] [1]), .C(clk32MHz), 
           .D(n19252));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i19 (.Q(\data_in_frame[2] [2]), .C(clk32MHz), 
           .D(n19251));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i2_3_lut_4_lut_adj_1369 (.I0(\data_in_frame[0] [6]), .I1(\data_in_frame[1] [0]), 
            .I2(\data_in_frame[3] [2]), .I3(\data_in_frame[1] [1]), .O(n33057));   // verilog/coms.v(70[16:27])
    defparam i2_3_lut_4_lut_adj_1369.LUT_INIT = 16'h6996;
    SB_DFF data_in_frame_0__i20 (.Q(\data_in_frame[2] [3]), .C(clk32MHz), 
           .D(n19250));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i21 (.Q(\data_in_frame[2] [4]), .C(clk32MHz), 
           .D(n19249));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i22 (.Q(\data_in_frame[2] [5]), .C(clk32MHz), 
           .D(n19248));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i1_2_lut_4_lut_adj_1370 (.I0(\data_in_frame[9] [2]), .I1(\data_in_frame[9] [3]), 
            .I2(\data_in_frame[9] [4]), .I3(\data_in_frame[9] [1]), .O(n18168));   // verilog/coms.v(75[16:43])
    defparam i1_2_lut_4_lut_adj_1370.LUT_INIT = 16'h6996;
    SB_DFF data_in_frame_0__i23 (.Q(\data_in_frame[2] [6]), .C(clk32MHz), 
           .D(n19247));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i24 (.Q(\data_in_frame[2] [7]), .C(clk32MHz), 
           .D(n19246));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i25 (.Q(\data_in_frame[3] [0]), .C(clk32MHz), 
           .D(n19245));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i26 (.Q(\data_in_frame[3] [1]), .C(clk32MHz), 
           .D(n19244));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i27 (.Q(\data_in_frame[3] [2]), .C(clk32MHz), 
           .D(n19243));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i28 (.Q(\data_in_frame[3] [3]), .C(clk32MHz), 
           .D(n19242));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i29 (.Q(\data_in_frame[3] [4]), .C(clk32MHz), 
           .D(n19241));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i30 (.Q(\data_in_frame[3] [5]), .C(clk32MHz), 
           .D(n19240));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i31 (.Q(\data_in_frame[3] [6]), .C(clk32MHz), 
           .D(n19239));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i32 (.Q(\data_in_frame[3] [7]), .C(clk32MHz), 
           .D(n19238));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i33 (.Q(\data_in_frame[4] [0]), .C(clk32MHz), 
           .D(n19237));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i34 (.Q(\data_in_frame[4] [1]), .C(clk32MHz), 
           .D(n19236));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i35 (.Q(\data_in_frame[4] [2]), .C(clk32MHz), 
           .D(n19235));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i36 (.Q(\data_in_frame[4] [3]), .C(clk32MHz), 
           .D(n19234));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i37 (.Q(\data_in_frame[4] [4]), .C(clk32MHz), 
           .D(n19233));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i19370_2_lut_4_lut (.I0(n2_adj_4085), .I1(n3_adj_4084), .I2(n1), 
            .I3(\FRAME_MATCHER.state_c [13]), .O(n24508));
    defparam i19370_2_lut_4_lut.LUT_INIT = 16'hfe00;
    SB_DFF data_in_frame_0__i38 (.Q(\data_in_frame[4] [5]), .C(clk32MHz), 
           .D(n19232));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i39 (.Q(\data_in_frame[4] [6]), .C(clk32MHz), 
           .D(n19231));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i40 (.Q(\data_in_frame[4] [7]), .C(clk32MHz), 
           .D(n19230));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i41 (.Q(\data_in_frame[5] [0]), .C(clk32MHz), 
           .D(n19229));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i42 (.Q(\data_in_frame[5] [1]), .C(clk32MHz), 
           .D(n19228));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i43 (.Q(\data_in_frame[5] [2]), .C(clk32MHz), 
           .D(n19227));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i44 (.Q(\data_in_frame[5] [3]), .C(clk32MHz), 
           .D(n19226));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i45 (.Q(\data_in_frame[5] [4]), .C(clk32MHz), 
           .D(n19225));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i46 (.Q(\data_in_frame[5] [5]), .C(clk32MHz), 
           .D(n19224));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i47 (.Q(\data_in_frame[5] [6]), .C(clk32MHz), 
           .D(n19223));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i48 (.Q(\data_in_frame[5] [7]), .C(clk32MHz), 
           .D(n19222));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i49 (.Q(\data_in_frame[6] [0]), .C(clk32MHz), 
           .D(n19221));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i50 (.Q(\data_in_frame[6] [1]), .C(clk32MHz), 
           .D(n19220));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i51 (.Q(\data_in_frame[6] [2]), .C(clk32MHz), 
           .D(n19219));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i52 (.Q(\data_in_frame[6] [3]), .C(clk32MHz), 
           .D(n19218));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i53 (.Q(\data_in_frame[6] [4]), .C(clk32MHz), 
           .D(n19217));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i54 (.Q(\data_in_frame[6] [5]), .C(clk32MHz), 
           .D(n19216));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i55 (.Q(\data_in_frame[6] [6]), .C(clk32MHz), 
           .D(n19215));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i56 (.Q(\data_in_frame[6] [7]), .C(clk32MHz), 
           .D(n19214));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i57 (.Q(\data_in_frame[7] [0]), .C(clk32MHz), 
           .D(n19213));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i58 (.Q(\data_in_frame[7] [1]), .C(clk32MHz), 
           .D(n19212));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_3_i16_3_lut (.I0(\data_out_frame[16] [3]), 
            .I1(\data_out_frame[17] [3]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n16_adj_4299));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_3_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF data_in_frame_0__i59 (.Q(\data_in_frame[7] [2]), .C(clk32MHz), 
           .D(n19211));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i1_2_lut_3_lut_adj_1371 (.I0(\data_in_frame[15] [7]), .I1(\data_in_frame[9] [4]), 
            .I2(\data_in_frame[13] [6]), .I3(GND_net), .O(n33299));
    defparam i1_2_lut_3_lut_adj_1371.LUT_INIT = 16'h9696;
    SB_DFF data_in_frame_0__i60 (.Q(\data_in_frame[7] [3]), .C(clk32MHz), 
           .D(n19210));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i1_2_lut_4_lut_adj_1372 (.I0(\data_in_frame[1] [5]), .I1(\data_in_frame[3] [6]), 
            .I2(n33114), .I3(\data_in_frame[8] [1]), .O(n32732));
    defparam i1_2_lut_4_lut_adj_1372.LUT_INIT = 16'h6996;
    SB_DFF data_in_frame_0__i61 (.Q(\data_in_frame[7] [4]), .C(clk32MHz), 
           .D(n19209));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i62 (.Q(\data_in_frame[7] [5]), .C(clk32MHz), 
           .D(n19208));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i63 (.Q(\data_in_frame[7] [6]), .C(clk32MHz), 
           .D(n19207));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i64 (.Q(\data_in_frame[7] [7]), .C(clk32MHz), 
           .D(n19206));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i65 (.Q(\data_in_frame[8] [0]), .C(clk32MHz), 
           .D(n19205));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i66 (.Q(\data_in_frame[8] [1]), .C(clk32MHz), 
           .D(n19204));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i67 (.Q(\data_in_frame[8] [2]), .C(clk32MHz), 
           .D(n19203));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i68 (.Q(\data_in_frame[8] [3]), .C(clk32MHz), 
           .D(n19202));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i69 (.Q(\data_in_frame[8] [4]), .C(clk32MHz), 
           .D(n19201));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i70 (.Q(\data_in_frame[8] [5]), .C(clk32MHz), 
           .D(n19200));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i71 (.Q(\data_in_frame[8] [6]), .C(clk32MHz), 
           .D(n19199));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i72 (.Q(\data_in_frame[8] [7]), .C(clk32MHz), 
           .D(n19198));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i73 (.Q(\data_in_frame[9] [0]), .C(clk32MHz), 
           .D(n19197));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i74 (.Q(\data_in_frame[9] [1]), .C(clk32MHz), 
           .D(n19196));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i75 (.Q(\data_in_frame[9] [2]), .C(clk32MHz), 
           .D(n19195));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i76 (.Q(\data_in_frame[9] [3]), .C(clk32MHz), 
           .D(n19194));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_3_i17_3_lut (.I0(\data_out_frame[18] [3]), 
            .I1(\data_out_frame[19] [3]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n17_adj_4298));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_3_i17_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF data_in_frame_0__i77 (.Q(\data_in_frame[9] [4]), .C(clk32MHz), 
           .D(n19193));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i29817_2_lut (.I0(\data_out_frame[23] [3]), .I1(byte_transmit_counter[0]), 
            .I2(GND_net), .I3(GND_net), .O(n36297));
    defparam i29817_2_lut.LUT_INIT = 16'h8888;
    SB_DFF data_in_frame_0__i78 (.Q(\data_in_frame[9] [5]), .C(clk32MHz), 
           .D(n19192));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i79 (.Q(\data_in_frame[9] [6]), .C(clk32MHz), 
           .D(n19191));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i80 (.Q(\data_in_frame[9] [7]), .C(clk32MHz), 
           .D(n19190));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i29838_2_lut (.I0(\data_out_frame[20] [3]), .I1(byte_transmit_counter[0]), 
            .I2(GND_net), .I3(GND_net), .O(n36296));
    defparam i29838_2_lut.LUT_INIT = 16'h2222;
    SB_DFF data_in_frame_0__i81 (.Q(\data_in_frame[10] [0]), .C(clk32MHz), 
           .D(n19189));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i82 (.Q(\data_in_frame[10] [1]), .C(clk32MHz), 
           .D(n19188));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i83 (.Q(\data_in_frame[10] [2]), .C(clk32MHz), 
           .D(n19187));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i84 (.Q(\data_in_frame[10] [3]), .C(clk32MHz), 
           .D(n19186));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i85 (.Q(\data_in_frame[10] [4]), .C(clk32MHz), 
           .D(n19185));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i86 (.Q(\data_in_frame[10] [5]), .C(clk32MHz), 
           .D(n19184));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i87 (.Q(\data_in_frame[10] [6]), .C(clk32MHz), 
           .D(n19183));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i88 (.Q(\data_in_frame[10] [7]), .C(clk32MHz), 
           .D(n19182));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i89 (.Q(\data_in_frame[11] [0]), .C(clk32MHz), 
           .D(n19181));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i90 (.Q(\data_in_frame[11] [1]), .C(clk32MHz), 
           .D(n19180));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i91 (.Q(\data_in_frame[11] [2]), .C(clk32MHz), 
           .D(n19179));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i5_3_lut_4_lut_adj_1373 (.I0(n18440), .I1(n18460), .I2(n10_adj_4169), 
            .I3(\data_in_frame[15] [6]), .O(n15965));   // verilog/coms.v(72[16:41])
    defparam i5_3_lut_4_lut_adj_1373.LUT_INIT = 16'h6996;
    SB_LUT4 i19371_2_lut_4_lut (.I0(n2_adj_4085), .I1(n3_adj_4084), .I2(n1), 
            .I3(\FRAME_MATCHER.state_c [14]), .O(n24510));
    defparam i19371_2_lut_4_lut.LUT_INIT = 16'hfe00;
    SB_LUT4 i1_2_lut_3_lut_adj_1374 (.I0(\data_in_frame[1] [3]), .I1(\data_in_frame[3] [5]), 
            .I2(\data_in_frame[5] [7]), .I3(GND_net), .O(n33114));   // verilog/coms.v(75[16:27])
    defparam i1_2_lut_3_lut_adj_1374.LUT_INIT = 16'h9696;
    SB_DFF data_in_frame_0__i92 (.Q(\data_in_frame[11] [3]), .C(clk32MHz), 
           .D(n19178));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i93 (.Q(\data_in_frame[11] [4]), .C(clk32MHz), 
           .D(n19177));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i94 (.Q(\data_in_frame[11] [5]), .C(clk32MHz), 
           .D(n19176));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i95 (.Q(\data_in_frame[11] [6]), .C(clk32MHz), 
           .D(n19175));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i96 (.Q(\data_in_frame[11] [7]), .C(clk32MHz), 
           .D(n19174));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i97 (.Q(\data_in_frame[12] [0]), .C(clk32MHz), 
           .D(n19173));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i1_2_lut_4_lut_adj_1375 (.I0(\data_in_frame[11] [6]), .I1(\data_in_frame[9] [5]), 
            .I2(n30848), .I3(n30872), .O(n18440));   // verilog/coms.v(74[16:43])
    defparam i1_2_lut_4_lut_adj_1375.LUT_INIT = 16'h6996;
    SB_LUT4 i14013_3_lut_4_lut (.I0(n8_adj_4304), .I1(n32666), .I2(rx_data[2]), 
            .I3(\data_in_frame[14] [2]), .O(n19155));
    defparam i14013_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF data_in_frame_0__i98 (.Q(\data_in_frame[12] [1]), .C(clk32MHz), 
           .D(n19172));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i99 (.Q(\data_in_frame[12] [2]), .C(clk32MHz), 
           .D(n19171));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i100 (.Q(\data_in_frame[12] [3]), .C(clk32MHz), 
           .D(n19170));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 add_43_33_lut (.I0(n2312), .I1(\FRAME_MATCHER.i [31]), .I2(GND_net), 
            .I3(n27825), .O(n2_adj_4212)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_33_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1376 (.I0(\data_out_frame[17] [0]), .I1(n18450), 
            .I2(n33228), .I3(\data_out_frame[17] [1]), .O(n6_adj_4031));
    defparam i1_2_lut_3_lut_4_lut_adj_1376.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_3_lut_adj_1377 (.I0(Kp_23__N_862), .I1(\data_in_frame[0] [6]), 
            .I2(\data_in_frame[1] [0]), .I3(GND_net), .O(n16400));   // verilog/coms.v(77[16:27])
    defparam i1_2_lut_3_lut_adj_1377.LUT_INIT = 16'h9696;
    SB_DFF data_in_frame_0__i101 (.Q(\data_in_frame[12] [4]), .C(clk32MHz), 
           .D(n19169));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i102 (.Q(\data_in_frame[12] [5]), .C(clk32MHz), 
           .D(n19168));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i103 (.Q(\data_in_frame[12] [6]), .C(clk32MHz), 
           .D(n19167));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 add_43_32_lut (.I0(n2312), .I1(\FRAME_MATCHER.i [30]), .I2(GND_net), 
            .I3(n27824), .O(n2_adj_4216)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_32_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_43_32 (.CI(n27824), .I0(\FRAME_MATCHER.i [30]), .I1(GND_net), 
            .CO(n27825));
    SB_DFF data_in_frame_0__i104 (.Q(\data_in_frame[12] [7]), .C(clk32MHz), 
           .D(n19166));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i105 (.Q(\data_in_frame[13] [0]), .C(clk32MHz), 
           .D(n19165));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i106 (.Q(\data_in_frame[13] [1]), .C(clk32MHz), 
           .D(n19164));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i107 (.Q(\data_in_frame[13] [2]), .C(clk32MHz), 
           .D(n19163));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i108 (.Q(\data_in_frame[13] [3]), .C(clk32MHz), 
           .D(n19162));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i109 (.Q(\data_in_frame[13] [4]), .C(clk32MHz), 
           .D(n19161));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 add_43_31_lut (.I0(n2312), .I1(\FRAME_MATCHER.i [29]), .I2(GND_net), 
            .I3(n27823), .O(n2_adj_4218)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_31_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i14014_3_lut_4_lut (.I0(n8_adj_4304), .I1(n32666), .I2(rx_data[1]), 
            .I3(\data_in_frame[14] [1]), .O(n19156));
    defparam i14014_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF data_in_frame_0__i110 (.Q(\data_in_frame[13] [5]), .C(clk32MHz), 
           .D(n19160));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i111 (.Q(\data_in_frame[13] [6]), .C(clk32MHz), 
           .D(n19159));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i112 (.Q(\data_in_frame[13] [7]), .C(clk32MHz), 
           .D(n19158));   // verilog/coms.v(127[12] 300[6])
    SB_CARRY add_43_31 (.CI(n27823), .I0(\FRAME_MATCHER.i [29]), .I1(GND_net), 
            .CO(n27824));
    SB_DFF data_in_frame_0__i113 (.Q(\data_in_frame[14] [0]), .C(clk32MHz), 
           .D(n19157));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i114 (.Q(\data_in_frame[14] [1]), .C(clk32MHz), 
           .D(n19156));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i115 (.Q(\data_in_frame[14] [2]), .C(clk32MHz), 
           .D(n19155));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i14015_3_lut_4_lut (.I0(n8_adj_4304), .I1(n32666), .I2(rx_data[0]), 
            .I3(\data_in_frame[14] [0]), .O(n19157));
    defparam i14015_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 add_43_30_lut (.I0(n2312), .I1(\FRAME_MATCHER.i [28]), .I2(GND_net), 
            .I3(n27822), .O(n2_adj_4220)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_30_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i14008_3_lut_4_lut (.I0(n8_adj_4304), .I1(n32666), .I2(rx_data[7]), 
            .I3(\data_in_frame[14] [7]), .O(n19150));
    defparam i14008_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_3_lut_adj_1378 (.I0(n17738), .I1(\data_in_frame[1] [2]), 
            .I2(\data_in_frame[3] [4]), .I3(GND_net), .O(n6_adj_4155));
    defparam i1_2_lut_3_lut_adj_1378.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1379 (.I0(\data_out_frame[17] [0]), .I1(n18450), 
            .I2(\data_out_frame[16] [5]), .I3(GND_net), .O(n6_adj_4071));
    defparam i1_2_lut_3_lut_adj_1379.LUT_INIT = 16'h9696;
    SB_LUT4 i14009_3_lut_4_lut (.I0(n8_adj_4304), .I1(n32666), .I2(rx_data[6]), 
            .I3(\data_in_frame[14] [6]), .O(n19151));
    defparam i14009_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_3_lut_adj_1380 (.I0(\data_out_frame[7] [7]), .I1(\data_out_frame[7] [6]), 
            .I2(\data_out_frame[8] [0]), .I3(GND_net), .O(n18431));   // verilog/coms.v(85[17:70])
    defparam i1_2_lut_3_lut_adj_1380.LUT_INIT = 16'h9696;
    SB_LUT4 i14010_3_lut_4_lut (.I0(n8_adj_4304), .I1(n32666), .I2(rx_data[5]), 
            .I3(\data_in_frame[14] [5]), .O(n19152));
    defparam i14010_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i14011_3_lut_4_lut (.I0(n8_adj_4304), .I1(n32666), .I2(rx_data[4]), 
            .I3(\data_in_frame[14] [4]), .O(n19153));
    defparam i14011_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i14012_3_lut_4_lut (.I0(n8_adj_4304), .I1(n32666), .I2(rx_data[3]), 
            .I3(\data_in_frame[14] [3]), .O(n19154));
    defparam i14012_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_CARRY add_43_30 (.CI(n27822), .I0(\FRAME_MATCHER.i [28]), .I1(GND_net), 
            .CO(n27823));
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1381 (.I0(\data_out_frame[23] [4]), .I1(n18363), 
            .I2(n17126), .I3(\data_out_frame[19] [2]), .O(n33256));
    defparam i1_2_lut_3_lut_4_lut_adj_1381.LUT_INIT = 16'h6996;
    SB_LUT4 i14_3_lut_4_lut (.I0(\data_in_frame[2] [6]), .I1(n17784), .I2(n17794), 
            .I3(n27_adj_4191), .O(n34_adj_4295));   // verilog/coms.v(73[16:42])
    defparam i14_3_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 add_43_29_lut (.I0(n2312), .I1(\FRAME_MATCHER.i [27]), .I2(GND_net), 
            .I3(n27821), .O(n2_adj_4222)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_29_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i1_2_lut_3_lut_adj_1382 (.I0(\data_in_frame[2] [6]), .I1(n17784), 
            .I2(\data_in_frame[4] [5]), .I3(GND_net), .O(n6_adj_4045));   // verilog/coms.v(73[16:42])
    defparam i1_2_lut_3_lut_adj_1382.LUT_INIT = 16'h9696;
    SB_CARRY add_43_29 (.CI(n27821), .I0(\FRAME_MATCHER.i [27]), .I1(GND_net), 
            .CO(n27822));
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_4_i16_3_lut (.I0(\data_out_frame[16] [4]), 
            .I1(\data_out_frame[17] [4]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n16_adj_4297));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_4_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_4_i17_3_lut (.I0(\data_out_frame[18] [4]), 
            .I1(\data_out_frame[19] [4]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n17_adj_4296));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_4_i17_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3_4_lut_4_lut (.I0(Kp_23__N_735), .I1(n17652), .I2(n30093), 
            .I3(GND_net), .O(n32702));
    defparam i3_4_lut_4_lut.LUT_INIT = 16'h6969;
    SB_LUT4 i1_2_lut_3_lut_adj_1383 (.I0(\data_out_frame[23] [4]), .I1(n18363), 
            .I2(\data_out_frame[23] [5]), .I3(GND_net), .O(n32861));
    defparam i1_2_lut_3_lut_adj_1383.LUT_INIT = 16'h9696;
    SB_LUT4 i14000_3_lut_4_lut (.I0(n24559), .I1(n32666), .I2(rx_data[7]), 
            .I3(\data_in_frame[15] [7]), .O(n19142));
    defparam i14000_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i13960_3_lut_4_lut (.I0(n8_adj_4066), .I1(n32678), .I2(rx_data[7]), 
            .I3(\data_in_frame[20] [7]), .O(n19102));
    defparam i13960_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13961_3_lut_4_lut (.I0(n8_adj_4066), .I1(n32678), .I2(rx_data[6]), 
            .I3(\data_in_frame[20] [6]), .O(n19103));
    defparam i13961_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_3_lut_4_lut_adj_1384 (.I0(\data_in_frame[16] [7]), .I1(\data_in_frame[16] [6]), 
            .I2(\data_in_frame[17] [0]), .I3(n33236), .O(n30093));
    defparam i1_3_lut_4_lut_adj_1384.LUT_INIT = 16'h9669;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_30928 (.I0(byte_transmit_counter[1]), 
            .I1(n36299), .I2(n36300), .I3(byte_transmit_counter[2]), .O(n37682));
    defparam byte_transmit_counter_1__bdd_4_lut_30928.LUT_INIT = 16'he4aa;
    SB_LUT4 i1_2_lut_4_lut_adj_1385 (.I0(n17863), .I1(\data_in_frame[10] [2]), 
            .I2(n29957), .I3(\data_in_frame[12] [4]), .O(n6_adj_4151));
    defparam i1_2_lut_4_lut_adj_1385.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_adj_1386 (.I0(\data_in_frame[0] [7]), .I1(\data_in_frame[1] [1]), 
            .I2(\data_in_frame[1] [2]), .I3(\data_in_frame[3] [3]), .O(n33212));
    defparam i1_2_lut_4_lut_adj_1386.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1387 (.I0(\data_in_frame[10] [2]), .I1(n29957), 
            .I2(\data_in_frame[12] [4]), .I3(GND_net), .O(n33302));
    defparam i1_2_lut_3_lut_adj_1387.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_4_lut_adj_1388 (.I0(Kp_23__N_1069), .I1(\data_in_frame[11] [0]), 
            .I2(\data_in_frame[8] [6]), .I3(\data_in_frame[10] [7]), .O(n33329));
    defparam i2_3_lut_4_lut_adj_1388.LUT_INIT = 16'h6996;
    SB_LUT4 i5_3_lut_4_lut_adj_1389 (.I0(\data_in_frame[11] [4]), .I1(\data_in_frame[14] [1]), 
            .I2(n10_adj_4126), .I3(n30114), .O(n33284));   // verilog/coms.v(74[16:43])
    defparam i5_3_lut_4_lut_adj_1389.LUT_INIT = 16'h6996;
    SB_LUT4 i2_2_lut_3_lut_adj_1390 (.I0(\data_in_frame[12] [7]), .I1(\data_in_frame[13] [1]), 
            .I2(\data_in_frame[10] [3]), .I3(GND_net), .O(n10_adj_4122));
    defparam i2_2_lut_3_lut_adj_1390.LUT_INIT = 16'h9696;
    SB_LUT4 i14001_3_lut_4_lut (.I0(n24559), .I1(n32666), .I2(rx_data[6]), 
            .I3(\data_in_frame[15] [6]), .O(n19143));
    defparam i14001_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1_2_lut_3_lut_adj_1391 (.I0(\data_in_frame[16] [3]), .I1(n30114), 
            .I2(\data_in_frame[14] [1]), .I3(GND_net), .O(n6_adj_4120));
    defparam i1_2_lut_3_lut_adj_1391.LUT_INIT = 16'h9696;
    SB_LUT4 i13962_3_lut_4_lut (.I0(n8_adj_4066), .I1(n32678), .I2(rx_data[5]), 
            .I3(\data_in_frame[20] [5]), .O(n19104));
    defparam i13962_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i14002_3_lut_4_lut (.I0(n24559), .I1(n32666), .I2(rx_data[5]), 
            .I3(\data_in_frame[15] [5]), .O(n19144));
    defparam i14002_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4_2_lut_4_lut (.I0(\data_in[3] [4]), .I1(n10_adj_4107), .I2(\data_in[2] [7]), 
            .I3(\data_in[3] [0]), .O(n15_adj_4102));
    defparam i4_2_lut_4_lut.LUT_INIT = 16'hffdf;
    SB_LUT4 i1_3_lut_4_lut_adj_1392 (.I0(n771), .I1(\FRAME_MATCHER.state[0] ), 
            .I2(n32653), .I3(n14711), .O(n2_adj_4085));
    defparam i1_3_lut_4_lut_adj_1392.LUT_INIT = 16'h0400;
    SB_LUT4 i1_3_lut_4_lut_adj_1393 (.I0(\FRAME_MATCHER.i [0]), .I1(\FRAME_MATCHER.i [4]), 
            .I2(n17471), .I3(\FRAME_MATCHER.i [1]), .O(n5_adj_4086));
    defparam i1_3_lut_4_lut_adj_1393.LUT_INIT = 16'hfefc;
    SB_LUT4 i1_3_lut_4_lut_adj_1394 (.I0(\FRAME_MATCHER.state [3]), .I1(n2970), 
            .I2(n14711), .I3(n2_adj_4272), .O(n32017));
    defparam i1_3_lut_4_lut_adj_1394.LUT_INIT = 16'haa80;
    SB_LUT4 i5_3_lut_4_lut_adj_1395 (.I0(Kp_23__N_843), .I1(n4_adj_4116), 
            .I2(\data_in_frame[1] [7]), .I3(\data_in_frame[0] [0]), .O(n22));
    defparam i5_3_lut_4_lut_adj_1395.LUT_INIT = 16'h2112;
    SB_LUT4 i2_3_lut_4_lut_adj_1396 (.I0(\FRAME_MATCHER.state_c [1]), .I1(n32655), 
            .I2(\FRAME_MATCHER.state [3]), .I3(n33453), .O(n18682));   // verilog/coms.v(127[12] 300[6])
    defparam i2_3_lut_4_lut_adj_1396.LUT_INIT = 16'h0010;
    SB_LUT4 i2_2_lut_4_lut_adj_1397 (.I0(\data_out_frame[8] [1]), .I1(\data_out_frame[7] [7]), 
            .I2(\data_out_frame[8] [3]), .I3(n18431), .O(n10_adj_4070));   // verilog/coms.v(85[17:70])
    defparam i2_2_lut_4_lut_adj_1397.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1398 (.I0(\data_out_frame[4] [1]), .I1(\data_out_frame[4] [0]), 
            .I2(\data_out_frame[6] [2]), .I3(GND_net), .O(n17569));   // verilog/coms.v(74[16:43])
    defparam i1_2_lut_3_lut_adj_1398.LUT_INIT = 16'h9696;
    SB_LUT4 i2_2_lut_3_lut_adj_1399 (.I0(\data_out_frame[18] [6]), .I1(n32960), 
            .I2(\data_out_frame[16] [4]), .I3(GND_net), .O(n6_adj_4065));
    defparam i2_2_lut_3_lut_adj_1399.LUT_INIT = 16'h9696;
    SB_LUT4 i13963_3_lut_4_lut (.I0(n8_adj_4066), .I1(n32678), .I2(rx_data[4]), 
            .I3(\data_in_frame[20] [4]), .O(n19105));
    defparam i13963_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i14003_3_lut_4_lut (.I0(n24559), .I1(n32666), .I2(rx_data[4]), 
            .I3(\data_in_frame[15] [4]), .O(n19145));
    defparam i14003_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i13964_3_lut_4_lut (.I0(n8_adj_4066), .I1(n32678), .I2(rx_data[3]), 
            .I3(\data_in_frame[20] [3]), .O(n19106));
    defparam i13964_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i14004_3_lut_4_lut (.I0(n24559), .I1(n32666), .I2(rx_data[3]), 
            .I3(\data_in_frame[15] [3]), .O(n19146));
    defparam i14004_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i13965_3_lut_4_lut (.I0(n8_adj_4066), .I1(n32678), .I2(rx_data[2]), 
            .I3(\data_in_frame[20] [2]), .O(n19107));
    defparam i13965_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i14005_3_lut_4_lut (.I0(n24559), .I1(n32666), .I2(rx_data[2]), 
            .I3(\data_in_frame[15] [2]), .O(n19147));
    defparam i14005_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1_2_lut_4_lut_adj_1400 (.I0(\data_out_frame[5] [1]), .I1(\data_out_frame[5] [0]), 
            .I2(\data_out_frame[7] [2]), .I3(\data_out_frame[4] [6]), .O(n32912));
    defparam i1_2_lut_4_lut_adj_1400.LUT_INIT = 16'h6996;
    SB_LUT4 i14006_3_lut_4_lut (.I0(n24559), .I1(n32666), .I2(rx_data[1]), 
            .I3(\data_in_frame[15] [1]), .O(n19148));
    defparam i14006_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i14007_3_lut_4_lut (.I0(n24559), .I1(n32666), .I2(rx_data[0]), 
            .I3(\data_in_frame[15] [0]), .O(n19149));
    defparam i14007_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i26705_2_lut_3_lut (.I0(\FRAME_MATCHER.state_c [1]), .I1(\FRAME_MATCHER.state[0] ), 
            .I2(\FRAME_MATCHER.state_c [2]), .I3(GND_net), .O(n33453));
    defparam i26705_2_lut_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i1_2_lut_4_lut_adj_1401 (.I0(\data_out_frame[4] [7]), .I1(\data_out_frame[7] [3]), 
            .I2(\data_out_frame[5] [2]), .I3(\data_out_frame[5] [1]), .O(n18333));
    defparam i1_2_lut_4_lut_adj_1401.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1402 (.I0(\FRAME_MATCHER.state_c [1]), .I1(\FRAME_MATCHER.state[0] ), 
            .I2(n32655), .I3(GND_net), .O(n4_adj_4305));
    defparam i1_2_lut_3_lut_adj_1402.LUT_INIT = 16'hfefe;
    SB_LUT4 i2_3_lut_4_lut_adj_1403 (.I0(\FRAME_MATCHER.i [4]), .I1(\FRAME_MATCHER.i [5]), 
            .I2(\FRAME_MATCHER.i [3]), .I3(n23788), .O(n32657));   // verilog/coms.v(154[7:23])
    defparam i2_3_lut_4_lut_adj_1403.LUT_INIT = 16'hfeff;
    SB_LUT4 i2_3_lut_4_lut_adj_1404 (.I0(\FRAME_MATCHER.i [4]), .I1(\FRAME_MATCHER.i [5]), 
            .I2(\FRAME_MATCHER.i [3]), .I3(n23788), .O(n32666));   // verilog/coms.v(154[7:23])
    defparam i2_3_lut_4_lut_adj_1404.LUT_INIT = 16'hefff;
    SB_LUT4 i13966_3_lut_4_lut (.I0(n8_adj_4066), .I1(n32678), .I2(rx_data[1]), 
            .I3(\data_in_frame[20] [1]), .O(n19108));
    defparam i13966_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13967_3_lut_4_lut (.I0(n8_adj_4066), .I1(n32678), .I2(rx_data[0]), 
            .I3(\data_in_frame[20] [0]), .O(n19109));
    defparam i13967_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_3_lut_adj_1405 (.I0(\data_in_frame[1] [1]), .I1(\data_in_frame[1] [2]), 
            .I2(\data_in_frame[3] [3]), .I3(GND_net), .O(n32916));   // verilog/coms.v(73[16:34])
    defparam i1_2_lut_3_lut_adj_1405.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1406 (.I0(\data_in_frame[1] [1]), .I1(\data_in_frame[1] [2]), 
            .I2(n33142), .I3(GND_net), .O(Kp_23__N_862));   // verilog/coms.v(73[16:34])
    defparam i1_2_lut_3_lut_adj_1406.LUT_INIT = 16'h9696;
    SB_LUT4 equal_132_i8_2_lut_3_lut (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(\FRAME_MATCHER.i [0]), .I3(GND_net), .O(n8_adj_4066));   // verilog/coms.v(154[7:23])
    defparam equal_132_i8_2_lut_3_lut.LUT_INIT = 16'hfbfb;
    SB_LUT4 n37682_bdd_4_lut (.I0(n37682), .I1(n17_adj_4152), .I2(n16_adj_4150), 
            .I3(byte_transmit_counter[2]), .O(n37685));
    defparam n37682_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i2_2_lut_4_lut_adj_1407 (.I0(\data_out_frame[25] [7]), .I1(n30870), 
            .I2(n30174), .I3(\data_out_frame[23] [7]), .O(n7_c));
    defparam i2_2_lut_4_lut_adj_1407.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_3_lut_adj_1408 (.I0(\data_out_frame[7] [3]), .I1(\data_out_frame[5] [2]), 
            .I2(\data_out_frame[5] [1]), .I3(GND_net), .O(n33093));
    defparam i1_2_lut_3_lut_adj_1408.LUT_INIT = 16'h9696;
    SB_LUT4 i3_4_lut_3_lut (.I0(n30870), .I1(n30174), .I2(\data_out_frame[23] [7]), 
            .I3(GND_net), .O(n32931));
    defparam i3_4_lut_3_lut.LUT_INIT = 16'h6969;
    SB_LUT4 i2_3_lut_4_lut_adj_1409 (.I0(n30870), .I1(n33028), .I2(n33000), 
            .I3(\data_out_frame[24] [2]), .O(n33784));
    defparam i2_3_lut_4_lut_adj_1409.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1410 (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(n32666), .I3(\FRAME_MATCHER.i [0]), .O(n32667));   // verilog/coms.v(154[7:23])
    defparam i1_2_lut_3_lut_4_lut_adj_1410.LUT_INIT = 16'hfbff;
    SB_LUT4 i1_2_lut_3_lut_adj_1411 (.I0(\data_out_frame[7] [5]), .I1(\data_out_frame[8] [5]), 
            .I2(\data_out_frame[7] [6]), .I3(GND_net), .O(n33265));
    defparam i1_2_lut_3_lut_adj_1411.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1412 (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(n32678), .I3(\FRAME_MATCHER.i [0]), .O(n32679));   // verilog/coms.v(154[7:23])
    defparam i1_2_lut_3_lut_4_lut_adj_1412.LUT_INIT = 16'hfbff;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_30923 (.I0(byte_transmit_counter[1]), 
            .I1(n36305), .I2(n36306), .I3(byte_transmit_counter[2]), .O(n37676));
    defparam byte_transmit_counter_1__bdd_4_lut_30923.LUT_INIT = 16'he4aa;
    SB_LUT4 i19093_2_lut_3_lut (.I0(\FRAME_MATCHER.state_c [2]), .I1(\FRAME_MATCHER.state[0] ), 
            .I2(\FRAME_MATCHER.state_c [1]), .I3(GND_net), .O(n24226));
    defparam i19093_2_lut_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 i1_2_lut_3_lut_adj_1413 (.I0(\FRAME_MATCHER.state_c [2]), .I1(\FRAME_MATCHER.state[0] ), 
            .I2(n17548), .I3(GND_net), .O(n39));
    defparam i1_2_lut_3_lut_adj_1413.LUT_INIT = 16'hf7f7;
    SB_LUT4 i5_3_lut_4_lut_adj_1414 (.I0(n30908), .I1(n30957), .I2(\data_out_frame[16] [7]), 
            .I3(\data_out_frame[16] [6]), .O(n14_adj_4060));
    defparam i5_3_lut_4_lut_adj_1414.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1415 (.I0(\FRAME_MATCHER.state [3]), .I1(n32655), 
            .I2(\FRAME_MATCHER.state_c [1]), .I3(GND_net), .O(n17548));   // verilog/coms.v(212[5:16])
    defparam i1_2_lut_3_lut_adj_1415.LUT_INIT = 16'hfefe;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1416 (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(n32657), .I3(\FRAME_MATCHER.i [0]), .O(n32660));   // verilog/coms.v(154[7:23])
    defparam i1_2_lut_3_lut_4_lut_adj_1416.LUT_INIT = 16'hfbff;
    SB_LUT4 i2_3_lut_4_lut_adj_1417 (.I0(n1247), .I1(\data_out_frame[10] [6]), 
            .I2(n34545), .I3(n33206), .O(n30018));   // verilog/coms.v(85[17:63])
    defparam i2_3_lut_4_lut_adj_1417.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_3_lut_adj_1418 (.I0(\FRAME_MATCHER.state [3]), .I1(n32655), 
            .I2(n24226), .I3(GND_net), .O(n17559));   // verilog/coms.v(212[5:16])
    defparam i1_2_lut_3_lut_adj_1418.LUT_INIT = 16'hefef;
    SB_LUT4 i3_3_lut_4_lut (.I0(\FRAME_MATCHER.state [3]), .I1(n32655), 
            .I2(\FRAME_MATCHER.state_c [2]), .I3(n5534), .O(n63_adj_4087));   // verilog/coms.v(212[5:16])
    defparam i3_3_lut_4_lut.LUT_INIT = 16'hffef;
    SB_LUT4 n37676_bdd_4_lut (.I0(n37676), .I1(n17_adj_4149), .I2(n16_adj_4145), 
            .I3(byte_transmit_counter[2]), .O(n37679));
    defparam n37676_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i2_3_lut_4_lut_adj_1419 (.I0(\FRAME_MATCHER.state [3]), .I1(n32655), 
            .I2(\FRAME_MATCHER.state_c [2]), .I3(\FRAME_MATCHER.state_c [1]), 
            .O(n17551));   // verilog/coms.v(212[5:16])
    defparam i2_3_lut_4_lut_adj_1419.LUT_INIT = 16'hfeff;
    SB_LUT4 i2123_2_lut_3_lut (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(\FRAME_MATCHER.i [3]), .I3(GND_net), .O(n8_adj_4114));
    defparam i2123_2_lut_3_lut.LUT_INIT = 16'hf8f8;
    SB_LUT4 i2_3_lut_4_lut_adj_1420 (.I0(\data_out_frame[4] [6]), .I1(\data_out_frame[5] [0]), 
            .I2(n1168), .I3(\data_out_frame[7] [0]), .O(n18496));   // verilog/coms.v(85[17:70])
    defparam i2_3_lut_4_lut_adj_1420.LUT_INIT = 16'h6996;
    SB_LUT4 i19420_2_lut_3_lut (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(\FRAME_MATCHER.i [0]), .I3(GND_net), .O(n24559));
    defparam i19420_2_lut_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 i2_3_lut_4_lut_adj_1421 (.I0(\data_out_frame[14] [2]), .I1(n30860), 
            .I2(n17232), .I3(\data_out_frame[14] [1]), .O(n30957));
    defparam i2_3_lut_4_lut_adj_1421.LUT_INIT = 16'h6996;
    SB_LUT4 select_422_Select_1_i3_2_lut (.I0(\FRAME_MATCHER.i [1]), .I1(n2994), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_4271));
    defparam select_422_Select_1_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_3_lut_adj_1422 (.I0(\data_out_frame[14] [2]), .I1(n30860), 
            .I2(n33889), .I3(GND_net), .O(n32939));
    defparam i1_2_lut_3_lut_adj_1422.LUT_INIT = 16'h6969;
    SB_LUT4 equal_122_i8_2_lut_3_lut (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(\FRAME_MATCHER.i [0]), .I3(GND_net), .O(n8_adj_4304));
    defparam equal_122_i8_2_lut_3_lut.LUT_INIT = 16'hf7f7;
    SB_LUT4 i13992_3_lut_4_lut (.I0(n8_adj_4090), .I1(n32678), .I2(rx_data[7]), 
            .I3(\data_in_frame[16] [7]), .O(n19134));
    defparam i13992_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 select_422_Select_2_i3_2_lut (.I0(\FRAME_MATCHER.i [2]), .I1(n2994), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_4269));
    defparam select_422_Select_2_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i13993_3_lut_4_lut (.I0(n8_adj_4090), .I1(n32678), .I2(rx_data[6]), 
            .I3(\data_in_frame[16] [6]), .O(n19135));
    defparam i13993_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 select_422_Select_3_i3_2_lut (.I0(\FRAME_MATCHER.i [3]), .I1(n2994), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_4267));
    defparam select_422_Select_3_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 select_422_Select_4_i3_2_lut (.I0(\FRAME_MATCHER.i [4]), .I1(n2994), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_4265));
    defparam select_422_Select_4_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 select_422_Select_5_i3_2_lut (.I0(\FRAME_MATCHER.i [5]), .I1(n2994), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_4263));
    defparam select_422_Select_5_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 select_422_Select_6_i3_2_lut (.I0(\FRAME_MATCHER.i [6]), .I1(n2994), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_4261));
    defparam select_422_Select_6_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 select_422_Select_7_i3_2_lut (.I0(\FRAME_MATCHER.i [7]), .I1(n2994), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_4259));
    defparam select_422_Select_7_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 select_422_Select_8_i3_2_lut (.I0(\FRAME_MATCHER.i [8]), .I1(n2994), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_4257));
    defparam select_422_Select_8_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 select_422_Select_9_i3_2_lut (.I0(\FRAME_MATCHER.i [9]), .I1(n2994), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_4255));
    defparam select_422_Select_9_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 select_422_Select_10_i3_2_lut (.I0(\FRAME_MATCHER.i [10]), .I1(n2994), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_4253));
    defparam select_422_Select_10_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 select_422_Select_11_i3_2_lut (.I0(\FRAME_MATCHER.i [11]), .I1(n2994), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_4251));
    defparam select_422_Select_11_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 select_422_Select_12_i3_2_lut (.I0(\FRAME_MATCHER.i [12]), .I1(n2994), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_4249));
    defparam select_422_Select_12_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i13994_3_lut_4_lut (.I0(n8_adj_4090), .I1(n32678), .I2(rx_data[5]), 
            .I3(\data_in_frame[16] [5]), .O(n19136));
    defparam i13994_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13995_3_lut_4_lut (.I0(n8_adj_4090), .I1(n32678), .I2(rx_data[4]), 
            .I3(\data_in_frame[16] [4]), .O(n19137));
    defparam i13995_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 select_422_Select_13_i3_2_lut (.I0(\FRAME_MATCHER.i [13]), .I1(n2994), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_4247));
    defparam select_422_Select_13_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i2_3_lut_4_lut_adj_1423 (.I0(\data_out_frame[5] [0]), .I1(n1168), 
            .I2(\data_out_frame[6] [7]), .I3(\data_out_frame[4] [5]), .O(n32844));   // verilog/coms.v(85[17:70])
    defparam i2_3_lut_4_lut_adj_1423.LUT_INIT = 16'h6996;
    SB_LUT4 i13996_3_lut_4_lut (.I0(n8_adj_4090), .I1(n32678), .I2(rx_data[3]), 
            .I3(\data_in_frame[16] [3]), .O(n19138));
    defparam i13996_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 select_422_Select_14_i3_2_lut (.I0(\FRAME_MATCHER.i [14]), .I1(n2994), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_4245));
    defparam select_422_Select_14_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i13997_3_lut_4_lut (.I0(n8_adj_4090), .I1(n32678), .I2(rx_data[2]), 
            .I3(\data_in_frame[16] [2]), .O(n19139));
    defparam i13997_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 select_422_Select_15_i3_2_lut (.I0(\FRAME_MATCHER.i [15]), .I1(n2994), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_4243));
    defparam select_422_Select_15_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 select_422_Select_16_i3_2_lut (.I0(\FRAME_MATCHER.i [16]), .I1(n2994), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_4241));
    defparam select_422_Select_16_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 select_422_Select_17_i3_2_lut (.I0(\FRAME_MATCHER.i [17]), .I1(n2994), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_4240));
    defparam select_422_Select_17_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i13998_3_lut_4_lut (.I0(n8_adj_4090), .I1(n32678), .I2(rx_data[1]), 
            .I3(\data_in_frame[16] [1]), .O(n19140));
    defparam i13998_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13999_3_lut_4_lut (.I0(n8_adj_4090), .I1(n32678), .I2(rx_data[0]), 
            .I3(\data_in_frame[16] [0]), .O(n19141));
    defparam i13999_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_3_lut_adj_1424 (.I0(n29786), .I1(\data_in_frame[10] [0]), 
            .I2(\data_in_frame[12] [2]), .I3(GND_net), .O(n33341));
    defparam i1_2_lut_3_lut_adj_1424.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_4_lut_adj_1425 (.I0(\data_in_frame[1] [7]), .I1(\data_in_frame[1] [6]), 
            .I2(\data_in_frame[1] [3]), .I3(n32769), .O(n33142));   // verilog/coms.v(78[16:27])
    defparam i2_3_lut_4_lut_adj_1425.LUT_INIT = 16'h6996;
    SB_LUT4 select_422_Select_18_i3_2_lut (.I0(\FRAME_MATCHER.i [18]), .I1(n2994), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_4239));
    defparam select_422_Select_18_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 select_422_Select_19_i3_2_lut (.I0(\FRAME_MATCHER.i [19]), .I1(n2994), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_4238));
    defparam select_422_Select_19_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 select_422_Select_20_i3_2_lut (.I0(\FRAME_MATCHER.i [20]), .I1(n2994), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_4237));
    defparam select_422_Select_20_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 select_422_Select_21_i3_2_lut (.I0(\FRAME_MATCHER.i [21]), .I1(n2994), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_4235));
    defparam select_422_Select_21_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 select_422_Select_22_i3_2_lut (.I0(\FRAME_MATCHER.i [22]), .I1(n2994), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_4234));
    defparam select_422_Select_22_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 select_422_Select_23_i3_2_lut (.I0(\FRAME_MATCHER.i [23]), .I1(n2994), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_4233));
    defparam select_422_Select_23_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 select_422_Select_24_i3_2_lut (.I0(\FRAME_MATCHER.i [24]), .I1(n2994), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_4231));
    defparam select_422_Select_24_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_30918 (.I0(byte_transmit_counter[1]), 
            .I1(n36302), .I2(n36303), .I3(byte_transmit_counter[2]), .O(n37670));
    defparam byte_transmit_counter_1__bdd_4_lut_30918.LUT_INIT = 16'he4aa;
    SB_LUT4 i1_2_lut_3_lut_adj_1426 (.I0(\data_in_frame[1] [7]), .I1(\data_in_frame[1] [6]), 
            .I2(\data_in_frame[4] [2]), .I3(GND_net), .O(n17714));   // verilog/coms.v(78[16:27])
    defparam i1_2_lut_3_lut_adj_1426.LUT_INIT = 16'h9696;
    SB_LUT4 i14112_3_lut_4_lut (.I0(n8_adj_4300), .I1(n32657), .I2(rx_data[7]), 
            .I3(\data_in_frame[1] [7]), .O(n19254));
    defparam i14112_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 select_422_Select_25_i3_2_lut (.I0(\FRAME_MATCHER.i [25]), .I1(n2994), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_4225));
    defparam select_422_Select_25_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 select_422_Select_26_i3_2_lut (.I0(\FRAME_MATCHER.i [26]), .I1(n2994), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_4224));
    defparam select_422_Select_26_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 select_422_Select_27_i3_2_lut (.I0(\FRAME_MATCHER.i [27]), .I1(n2994), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_4223));
    defparam select_422_Select_27_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 select_422_Select_28_i3_2_lut (.I0(\FRAME_MATCHER.i [28]), .I1(n2994), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_4221));
    defparam select_422_Select_28_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 select_422_Select_29_i3_2_lut (.I0(\FRAME_MATCHER.i [29]), .I1(n2994), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_4219));
    defparam select_422_Select_29_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 select_422_Select_30_i3_2_lut (.I0(\FRAME_MATCHER.i [30]), .I1(n2994), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_4217));
    defparam select_422_Select_30_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_4_lut_adj_1427 (.I0(\data_out_frame[8] [4]), .I1(\data_out_frame[8] [2]), 
            .I2(\data_out_frame[5] [7]), .I3(\data_out_frame[5] [6]), .O(n32735));   // verilog/coms.v(76[16:43])
    defparam i1_2_lut_4_lut_adj_1427.LUT_INIT = 16'h6996;
    SB_LUT4 i14113_3_lut_4_lut (.I0(n8_adj_4300), .I1(n32657), .I2(rx_data[6]), 
            .I3(\data_in_frame[1] [6]), .O(n19255));
    defparam i14113_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_3_lut_adj_1428 (.I0(\data_out_frame[8] [2]), .I1(\data_out_frame[5] [7]), 
            .I2(\data_out_frame[5] [6]), .I3(GND_net), .O(n33356));
    defparam i1_2_lut_3_lut_adj_1428.LUT_INIT = 16'h9696;
    SB_LUT4 i14114_3_lut_4_lut (.I0(n8_adj_4300), .I1(n32657), .I2(rx_data[5]), 
            .I3(\data_in_frame[1] [5]), .O(n19256));
    defparam i14114_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i14115_3_lut_4_lut (.I0(n8_adj_4300), .I1(n32657), .I2(rx_data[4]), 
            .I3(\data_in_frame[1] [4]), .O(n19257));
    defparam i14115_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_3_lut_4_lut_adj_1429 (.I0(\data_out_frame[4] [1]), .I1(\data_out_frame[4] [3]), 
            .I2(\data_out_frame[6] [4]), .I3(\data_out_frame[6] [3]), .O(n1247));   // verilog/coms.v(75[16:43])
    defparam i2_3_lut_4_lut_adj_1429.LUT_INIT = 16'h6996;
    SB_LUT4 i14116_3_lut_4_lut (.I0(n8_adj_4300), .I1(n32657), .I2(rx_data[3]), 
            .I3(\data_in_frame[1] [3]), .O(n19258));
    defparam i14116_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i14117_3_lut_4_lut (.I0(n8_adj_4300), .I1(n32657), .I2(rx_data[2]), 
            .I3(\data_in_frame[1] [2]), .O(n19259));
    defparam i14117_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i5_3_lut_4_lut_adj_1430 (.I0(\data_out_frame[12] [5]), .I1(\data_out_frame[12] [4]), 
            .I2(n10_adj_4039), .I3(\data_out_frame[12] [2]), .O(n33308));
    defparam i5_3_lut_4_lut_adj_1430.LUT_INIT = 16'h6996;
    SB_LUT4 i14118_3_lut_4_lut (.I0(n8_adj_4300), .I1(n32657), .I2(rx_data[1]), 
            .I3(\data_in_frame[1] [1]), .O(n19260));
    defparam i14118_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_4_lut_adj_1431 (.I0(\data_out_frame[8] [6]), .I1(\data_out_frame[4] [2]), 
            .I2(\data_out_frame[4] [3]), .I3(\data_out_frame[6] [4]), .O(n18503));   // verilog/coms.v(75[16:43])
    defparam i1_2_lut_4_lut_adj_1431.LUT_INIT = 16'h6996;
    SB_LUT4 n37670_bdd_4_lut (.I0(n37670), .I1(n17_adj_4144), .I2(n16_adj_4142), 
            .I3(byte_transmit_counter[2]), .O(n37673));
    defparam n37670_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i14119_3_lut_4_lut (.I0(n8_adj_4300), .I1(n32657), .I2(rx_data[0]), 
            .I3(\data_in_frame[1] [0]), .O(n19261));
    defparam i14119_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_3_lut_adj_1432 (.I0(\data_out_frame[4] [2]), .I1(\data_out_frame[4] [3]), 
            .I2(\data_out_frame[6] [4]), .I3(GND_net), .O(n33148));   // verilog/coms.v(75[16:43])
    defparam i1_2_lut_3_lut_adj_1432.LUT_INIT = 16'h9696;
    SB_LUT4 equal_119_i8_2_lut_3_lut (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(\FRAME_MATCHER.i [0]), .I3(GND_net), .O(n8_adj_4300));   // verilog/coms.v(154[7:23])
    defparam equal_119_i8_2_lut_3_lut.LUT_INIT = 16'hefef;
    SB_LUT4 select_422_Select_31_i3_2_lut (.I0(\FRAME_MATCHER.i [31]), .I1(n2994), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_4213));
    defparam select_422_Select_31_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i4_4_lut_adj_1433 (.I0(n30116), .I1(\data_out_frame[25] [6]), 
            .I2(\data_out_frame[25] [7]), .I3(n6_adj_4306), .O(n34053));
    defparam i4_4_lut_adj_1433.LUT_INIT = 16'h9669;
    SB_LUT4 equal_120_i8_2_lut_3_lut (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(\FRAME_MATCHER.i [0]), .I3(GND_net), .O(n8_adj_4090));   // verilog/coms.v(154[7:23])
    defparam equal_120_i8_2_lut_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i14104_3_lut_4_lut (.I0(n8_adj_4302), .I1(n32657), .I2(rx_data[7]), 
            .I3(\data_in_frame[2] [7]), .O(n19246));
    defparam i14104_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i14105_3_lut_4_lut (.I0(n8_adj_4302), .I1(n32657), .I2(rx_data[6]), 
            .I3(\data_in_frame[2] [6]), .O(n19247));
    defparam i14105_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i14106_3_lut_4_lut (.I0(n8_adj_4302), .I1(n32657), .I2(rx_data[5]), 
            .I3(\data_in_frame[2] [5]), .O(n19248));
    defparam i14106_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i14107_3_lut_4_lut (.I0(n8_adj_4302), .I1(n32657), .I2(rx_data[4]), 
            .I3(\data_in_frame[2] [4]), .O(n19249));
    defparam i14107_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i14108_3_lut_4_lut (.I0(n8_adj_4302), .I1(n32657), .I2(rx_data[3]), 
            .I3(\data_in_frame[2] [3]), .O(n19250));
    defparam i14108_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i14109_3_lut_4_lut (.I0(n8_adj_4302), .I1(n32657), .I2(rx_data[2]), 
            .I3(\data_in_frame[2] [2]), .O(n19251));
    defparam i14109_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_3_lut_4_lut_adj_1434 (.I0(\data_out_frame[9] [4]), .I1(n18333), 
            .I2(n32844), .I3(n33181), .O(n17243));
    defparam i2_3_lut_4_lut_adj_1434.LUT_INIT = 16'h6996;
    SB_LUT4 i14110_3_lut_4_lut (.I0(n8_adj_4302), .I1(n32657), .I2(rx_data[1]), 
            .I3(\data_in_frame[2] [1]), .O(n19252));
    defparam i14110_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i14111_3_lut_4_lut (.I0(n8_adj_4302), .I1(n32657), .I2(rx_data[0]), 
            .I3(\data_in_frame[2] [0]), .O(n19253));
    defparam i14111_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i14096_3_lut_4_lut (.I0(n8_adj_4303), .I1(n32657), .I2(rx_data[7]), 
            .I3(\data_in_frame[3] [7]), .O(n19238));
    defparam i14096_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i14097_3_lut_4_lut (.I0(n8_adj_4303), .I1(n32657), .I2(rx_data[6]), 
            .I3(\data_in_frame[3] [6]), .O(n19239));
    defparam i14097_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i14098_3_lut_4_lut (.I0(n8_adj_4303), .I1(n32657), .I2(rx_data[5]), 
            .I3(\data_in_frame[3] [5]), .O(n19240));
    defparam i14098_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i14099_3_lut_4_lut (.I0(n8_adj_4303), .I1(n32657), .I2(rx_data[4]), 
            .I3(\data_in_frame[3] [4]), .O(n19241));
    defparam i14099_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i14100_3_lut_4_lut (.I0(n8_adj_4303), .I1(n32657), .I2(rx_data[3]), 
            .I3(\data_in_frame[3] [3]), .O(n19242));
    defparam i14100_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_3_lut_4_lut_adj_1435 (.I0(\data_out_frame[9] [4]), .I1(n18333), 
            .I2(n32912), .I3(\data_out_frame[11] [6]), .O(n33074));
    defparam i2_3_lut_4_lut_adj_1435.LUT_INIT = 16'h6996;
    SB_LUT4 i14101_3_lut_4_lut (.I0(n8_adj_4303), .I1(n32657), .I2(rx_data[2]), 
            .I3(\data_in_frame[3] [2]), .O(n19243));
    defparam i14101_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i14102_3_lut_4_lut (.I0(n8_adj_4303), .I1(n32657), .I2(rx_data[1]), 
            .I3(\data_in_frame[3] [1]), .O(n19244));
    defparam i14102_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i5_3_lut_4_lut_adj_1436 (.I0(\data_out_frame[5] [2]), .I1(\data_out_frame[7] [4]), 
            .I2(n10_adj_4062), .I3(n33096), .O(n30860));
    defparam i5_3_lut_4_lut_adj_1436.LUT_INIT = 16'h6996;
    SB_LUT4 i2_2_lut_3_lut_adj_1437 (.I0(\data_out_frame[8] [7]), .I1(\data_out_frame[8] [6]), 
            .I2(\data_out_frame[6] [6]), .I3(GND_net), .O(n10_adj_4036));   // verilog/coms.v(85[17:28])
    defparam i2_2_lut_3_lut_adj_1437.LUT_INIT = 16'h9696;
    SB_LUT4 i14103_3_lut_4_lut (.I0(n8_adj_4303), .I1(n32657), .I2(rx_data[0]), 
            .I3(\data_in_frame[3] [0]), .O(n19245));
    defparam i14103_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_30953 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[26] [1]), .I2(\data_out_frame[27] [1]), 
            .I3(byte_transmit_counter[1]), .O(n37658));
    defparam byte_transmit_counter_0__bdd_4_lut_30953.LUT_INIT = 16'he4aa;
    SB_LUT4 i14088_3_lut_4_lut (.I0(n8_adj_4066), .I1(n32657), .I2(rx_data[7]), 
            .I3(\data_in_frame[4] [7]), .O(n19230));
    defparam i14088_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i14089_3_lut_4_lut (.I0(n8_adj_4066), .I1(n32657), .I2(rx_data[6]), 
            .I3(\data_in_frame[4] [6]), .O(n19231));
    defparam i14089_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_3_lut_4_lut_adj_1438 (.I0(\data_out_frame[5] [2]), .I1(\data_out_frame[7] [4]), 
            .I2(n18333), .I3(n33197), .O(n17768));
    defparam i2_3_lut_4_lut_adj_1438.LUT_INIT = 16'h6996;
    SB_LUT4 i14090_3_lut_4_lut (.I0(n8_adj_4066), .I1(n32657), .I2(rx_data[5]), 
            .I3(\data_in_frame[4] [5]), .O(n19232));
    defparam i14090_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i14091_3_lut_4_lut (.I0(n8_adj_4066), .I1(n32657), .I2(rx_data[4]), 
            .I3(\data_in_frame[4] [4]), .O(n19233));
    defparam i14091_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i14092_3_lut_4_lut (.I0(n8_adj_4066), .I1(n32657), .I2(rx_data[3]), 
            .I3(\data_in_frame[4] [3]), .O(n19234));
    defparam i14092_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_3_lut_4_lut_adj_1439 (.I0(n18431), .I1(n32878), .I2(\data_out_frame[14] [3]), 
            .I3(n33096), .O(n33889));   // verilog/coms.v(74[16:27])
    defparam i2_3_lut_4_lut_adj_1439.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_adj_1440 (.I0(\data_out_frame[19] [4]), .I1(n30895), 
            .I2(n32963), .I3(n33256), .O(n6_adj_4306));
    defparam i1_2_lut_4_lut_adj_1440.LUT_INIT = 16'h9669;
    SB_LUT4 i14093_3_lut_4_lut (.I0(n8_adj_4066), .I1(n32657), .I2(rx_data[2]), 
            .I3(\data_in_frame[4] [2]), .O(n19235));
    defparam i14093_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 n37658_bdd_4_lut (.I0(n37658), .I1(\data_out_frame[25] [1]), 
            .I2(\data_out_frame[24] [1]), .I3(byte_transmit_counter[1]), 
            .O(n37661));
    defparam n37658_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i14094_3_lut_4_lut (.I0(n8_adj_4066), .I1(n32657), .I2(rx_data[1]), 
            .I3(\data_in_frame[4] [1]), .O(n19236));
    defparam i14094_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_3_lut_adj_1441 (.I0(n18431), .I1(n32878), .I2(\data_out_frame[14] [4]), 
            .I3(GND_net), .O(n33172));   // verilog/coms.v(74[16:27])
    defparam i1_2_lut_3_lut_adj_1441.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1442 (.I0(\data_out_frame[4] [3]), .I1(\data_out_frame[4] [4]), 
            .I2(\data_out_frame[6] [5]), .I3(GND_net), .O(n18075));
    defparam i1_2_lut_3_lut_adj_1442.LUT_INIT = 16'h9696;
    SB_LUT4 i14095_3_lut_4_lut (.I0(n8_adj_4066), .I1(n32657), .I2(rx_data[0]), 
            .I3(\data_in_frame[4] [0]), .O(n19237));
    defparam i14095_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_3_lut_adj_1443 (.I0(\data_out_frame[13] [1]), .I1(n17086), 
            .I2(n32949), .I3(GND_net), .O(n33230));
    defparam i1_2_lut_3_lut_adj_1443.LUT_INIT = 16'h9696;
    SB_LUT4 i2_2_lut_3_lut_adj_1444 (.I0(\data_in_frame[0] [3]), .I1(\data_in_frame[2] [5]), 
            .I2(\data_in_frame[0] [4]), .I3(GND_net), .O(n18268));   // verilog/coms.v(74[16:43])
    defparam i2_2_lut_3_lut_adj_1444.LUT_INIT = 16'h9696;
    SB_LUT4 i5_3_lut_4_lut_adj_1445 (.I0(\data_out_frame[19] [2]), .I1(n17126), 
            .I2(n18330), .I3(n10_adj_4073), .O(n32713));
    defparam i5_3_lut_4_lut_adj_1445.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_3_lut_adj_1446 (.I0(\data_in_frame[0] [3]), .I1(\data_in_frame[2] [5]), 
            .I2(\data_in_frame[0] [5]), .I3(GND_net), .O(n17784));   // verilog/coms.v(74[16:43])
    defparam i1_2_lut_3_lut_adj_1446.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1447 (.I0(\data_in_frame[0] [1]), .I1(\data_in_frame[0] [0]), 
            .I2(\data_in_frame[2] [2]), .I3(GND_net), .O(n4_adj_4116));   // verilog/coms.v(72[16:27])
    defparam i1_2_lut_3_lut_adj_1447.LUT_INIT = 16'h9696;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_30905 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[26] [3]), .I2(\data_out_frame[27] [3]), 
            .I3(byte_transmit_counter[1]), .O(n37652));
    defparam byte_transmit_counter_0__bdd_4_lut_30905.LUT_INIT = 16'he4aa;
    SB_LUT4 i2_3_lut_4_lut_adj_1448 (.I0(\data_in_frame[0] [1]), .I1(\data_in_frame[0] [0]), 
            .I2(\data_in_frame[4] [4]), .I3(\data_in_frame[2] [2]), .O(n33127));   // verilog/coms.v(72[16:27])
    defparam i2_3_lut_4_lut_adj_1448.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_1449 (.I0(\data_out_frame[10] [2]), .I1(\data_out_frame[10] [1]), 
            .I2(n33350), .I3(n32908), .O(n33206));   // verilog/coms.v(75[16:27])
    defparam i2_3_lut_4_lut_adj_1449.LUT_INIT = 16'h6996;
    SB_LUT4 i14072_3_lut_4_lut (.I0(n8_adj_4304), .I1(n32657), .I2(rx_data[7]), 
            .I3(\data_in_frame[6] [7]), .O(n19214));
    defparam i14072_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i14073_3_lut_4_lut (.I0(n8_adj_4304), .I1(n32657), .I2(rx_data[6]), 
            .I3(\data_in_frame[6] [6]), .O(n19215));
    defparam i14073_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i14074_3_lut_4_lut (.I0(n8_adj_4304), .I1(n32657), .I2(rx_data[5]), 
            .I3(\data_in_frame[6] [5]), .O(n19216));
    defparam i14074_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_4_lut_adj_1450 (.I0(\FRAME_MATCHER.state_c [2]), .I1(n17503), 
            .I2(\FRAME_MATCHER.state_c [1]), .I3(n4_adj_4305), .O(n17504));
    defparam i1_4_lut_adj_1450.LUT_INIT = 16'hfeee;
    SB_LUT4 i2_3_lut_4_lut_adj_1451 (.I0(\data_out_frame[10] [2]), .I1(\data_out_frame[10] [1]), 
            .I2(\data_out_frame[6] [0]), .I3(\data_out_frame[12] [3]), .O(n33069));   // verilog/coms.v(75[16:27])
    defparam i2_3_lut_4_lut_adj_1451.LUT_INIT = 16'h6996;
    SB_LUT4 i14075_3_lut_4_lut (.I0(n8_adj_4304), .I1(n32657), .I2(rx_data[4]), 
            .I3(\data_in_frame[6] [4]), .O(n19217));
    defparam i14075_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 n37652_bdd_4_lut (.I0(n37652), .I1(\data_out_frame[25] [3]), 
            .I2(\data_out_frame[24] [3]), .I3(byte_transmit_counter[1]), 
            .O(n37655));
    defparam n37652_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i14076_3_lut_4_lut (.I0(n8_adj_4304), .I1(n32657), .I2(rx_data[3]), 
            .I3(\data_in_frame[6] [3]), .O(n19218));
    defparam i14076_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i14077_3_lut_4_lut (.I0(n8_adj_4304), .I1(n32657), .I2(rx_data[2]), 
            .I3(\data_in_frame[6] [2]), .O(n19219));
    defparam i14077_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_4_lut_adj_1452 (.I0(\data_out_frame[20] [5]), .I1(\data_out_frame[20] [6]), 
            .I2(n30073), .I3(n30986), .O(n33086));
    defparam i1_2_lut_4_lut_adj_1452.LUT_INIT = 16'h9669;
    SB_LUT4 i14078_3_lut_4_lut (.I0(n8_adj_4304), .I1(n32657), .I2(rx_data[1]), 
            .I3(\data_in_frame[6] [1]), .O(n19220));
    defparam i14078_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i14079_3_lut_4_lut (.I0(n8_adj_4304), .I1(n32657), .I2(rx_data[0]), 
            .I3(\data_in_frame[6] [0]), .O(n19221));
    defparam i14079_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i14064_3_lut_4_lut (.I0(n24559), .I1(n32657), .I2(rx_data[7]), 
            .I3(\data_in_frame[7] [7]), .O(n19206));
    defparam i14064_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i14065_3_lut_4_lut (.I0(n24559), .I1(n32657), .I2(rx_data[6]), 
            .I3(\data_in_frame[7] [6]), .O(n19207));
    defparam i14065_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i14066_3_lut_4_lut (.I0(n24559), .I1(n32657), .I2(rx_data[5]), 
            .I3(\data_in_frame[7] [5]), .O(n19208));
    defparam i14066_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i14067_3_lut_4_lut (.I0(n24559), .I1(n32657), .I2(rx_data[4]), 
            .I3(\data_in_frame[7] [4]), .O(n19209));
    defparam i14067_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i14068_3_lut_4_lut (.I0(n24559), .I1(n32657), .I2(rx_data[3]), 
            .I3(\data_in_frame[7] [3]), .O(n19210));
    defparam i14068_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1_2_lut_4_lut_adj_1453 (.I0(\data_out_frame[14] [0]), .I1(n33074), 
            .I2(n17768), .I3(n30108), .O(n4_c));
    defparam i1_2_lut_4_lut_adj_1453.LUT_INIT = 16'h6996;
    SB_LUT4 i14069_3_lut_4_lut (.I0(n24559), .I1(n32657), .I2(rx_data[2]), 
            .I3(\data_in_frame[7] [2]), .O(n19211));
    defparam i14069_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i14070_3_lut_4_lut (.I0(n24559), .I1(n32657), .I2(rx_data[1]), 
            .I3(\data_in_frame[7] [1]), .O(n19212));
    defparam i14070_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i13_3_lut_4_lut (.I0(\data_out_frame[15] [0]), .I1(n17676), 
            .I2(n33172), .I3(n32881), .O(n38));
    defparam i13_3_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i14071_3_lut_4_lut (.I0(n24559), .I1(n32657), .I2(rx_data[0]), 
            .I3(\data_in_frame[7] [0]), .O(n19213));
    defparam i14071_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1_2_lut_3_lut_adj_1454 (.I0(\data_out_frame[20] [6]), .I1(n30073), 
            .I2(n30986), .I3(GND_net), .O(n33085));
    defparam i1_2_lut_3_lut_adj_1454.LUT_INIT = 16'h6969;
    SB_LUT4 i14056_3_lut_4_lut (.I0(n8_adj_4090), .I1(n32666), .I2(rx_data[7]), 
            .I3(\data_in_frame[8] [7]), .O(n19198));
    defparam i14056_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_3_lut_4_lut_adj_1455 (.I0(n30885), .I1(n30874), .I2(n33086), 
            .I3(n31000), .O(n17112));
    defparam i2_3_lut_4_lut_adj_1455.LUT_INIT = 16'h9669;
    SB_LUT4 i5_3_lut_4_lut_adj_1456 (.I0(\data_out_frame[15] [7]), .I1(\data_out_frame[15] [6]), 
            .I2(n10_adj_4028), .I3(n33193), .O(n32984));
    defparam i5_3_lut_4_lut_adj_1456.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_1457 (.I0(\data_out_frame[15] [0]), .I1(n17676), 
            .I2(n17084), .I3(n32949), .O(n33227));
    defparam i2_3_lut_4_lut_adj_1457.LUT_INIT = 16'h6996;
    SB_LUT4 i14057_3_lut_4_lut (.I0(n8_adj_4090), .I1(n32666), .I2(rx_data[6]), 
            .I3(\data_in_frame[8] [6]), .O(n19199));
    defparam i14057_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_30900 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[26] [2]), .I2(\data_out_frame[27] [2]), 
            .I3(byte_transmit_counter[1]), .O(n37646));
    defparam byte_transmit_counter_0__bdd_4_lut_30900.LUT_INIT = 16'he4aa;
    SB_LUT4 i14058_3_lut_4_lut (.I0(n8_adj_4090), .I1(n32666), .I2(rx_data[5]), 
            .I3(\data_in_frame[8] [5]), .O(n19200));
    defparam i14058_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 n37646_bdd_4_lut (.I0(n37646), .I1(\data_out_frame[25] [2]), 
            .I2(\data_out_frame[24] [2]), .I3(byte_transmit_counter[1]), 
            .O(n37649));
    defparam n37646_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i14059_3_lut_4_lut (.I0(n8_adj_4090), .I1(n32666), .I2(rx_data[4]), 
            .I3(\data_in_frame[8] [4]), .O(n19201));
    defparam i14059_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i14060_3_lut_4_lut (.I0(n8_adj_4090), .I1(n32666), .I2(rx_data[3]), 
            .I3(\data_in_frame[8] [3]), .O(n19202));
    defparam i14060_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_3_lut_4_lut_adj_1458 (.I0(n30049), .I1(n30866), .I2(\data_out_frame[23] [0]), 
            .I3(n30986), .O(n33130));
    defparam i2_3_lut_4_lut_adj_1458.LUT_INIT = 16'h6996;
    SB_LUT4 i14061_3_lut_4_lut (.I0(n8_adj_4090), .I1(n32666), .I2(rx_data[2]), 
            .I3(\data_in_frame[8] [2]), .O(n19203));
    defparam i14061_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i14062_3_lut_4_lut (.I0(n8_adj_4090), .I1(n32666), .I2(rx_data[1]), 
            .I3(\data_in_frame[8] [1]), .O(n19204));
    defparam i14062_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i14063_3_lut_4_lut (.I0(n8_adj_4090), .I1(n32666), .I2(rx_data[0]), 
            .I3(\data_in_frame[8] [0]), .O(n19205));
    defparam i14063_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_4_lut_adj_1459 (.I0(\data_out_frame[24] [7]), .I1(n30885), 
            .I2(n30995), .I3(n31000), .O(n30058));
    defparam i1_2_lut_4_lut_adj_1459.LUT_INIT = 16'h6996;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_7_i7_3_lut_4_lut (.I0(byte_transmit_counter[2]), 
            .I1(byte_transmit_counter[1]), .I2(n35440), .I3(n35438), .O(n7_adj_4291));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_7_i7_3_lut_4_lut.LUT_INIT = 16'hf2d0;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_6_i7_3_lut_4_lut (.I0(byte_transmit_counter[2]), 
            .I1(byte_transmit_counter[1]), .I2(n35434), .I3(n35432), .O(n7_adj_4290));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_6_i7_3_lut_4_lut.LUT_INIT = 16'hf2d0;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_5_i7_3_lut_4_lut (.I0(byte_transmit_counter[2]), 
            .I1(byte_transmit_counter[1]), .I2(n35428), .I3(n35426), .O(n7_adj_4289));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_5_i7_3_lut_4_lut.LUT_INIT = 16'hf2d0;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_4_i7_3_lut_4_lut (.I0(byte_transmit_counter[2]), 
            .I1(byte_transmit_counter[1]), .I2(n35422), .I3(n35420), .O(n7_adj_4288));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_4_i7_3_lut_4_lut.LUT_INIT = 16'hf2d0;
    SB_LUT4 i30425_3_lut (.I0(n32655), .I1(n33453), .I2(n17503), .I3(GND_net), 
            .O(n33587));
    defparam i30425_3_lut.LUT_INIT = 16'h0101;
    SB_LUT4 i1_2_lut_4_lut_adj_1460 (.I0(n17704), .I1(\data_in_frame[9] [2]), 
            .I2(n17827), .I3(n17846), .O(n17595));   // verilog/coms.v(73[16:42])
    defparam i1_2_lut_4_lut_adj_1460.LUT_INIT = 16'h6996;
    SB_LUT4 i2_2_lut_4_lut_adj_1461 (.I0(\data_out_frame[18] [1]), .I1(n32902), 
            .I2(n10_adj_4026), .I3(GND_net), .O(n6_adj_4027));
    defparam i2_2_lut_4_lut_adj_1461.LUT_INIT = 16'h6969;
    SB_LUT4 i2_3_lut_4_lut_adj_1462 (.I0(n33057), .I1(n18058), .I2(\data_in_frame[5] [3]), 
            .I3(\data_in_frame[7] [4]), .O(n33338));
    defparam i2_3_lut_4_lut_adj_1462.LUT_INIT = 16'h6996;
    SB_LUT4 i30833_4_lut (.I0(n17503), .I1(n5592), .I2(n5_adj_4282), .I3(n6_adj_4283), 
            .O(n32597));
    defparam i30833_4_lut.LUT_INIT = 16'h1115;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_3_i7_3_lut_4_lut (.I0(byte_transmit_counter[2]), 
            .I1(byte_transmit_counter[1]), .I2(n35416), .I3(n35414), .O(n7_adj_4287));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_3_i7_3_lut_4_lut.LUT_INIT = 16'hf2d0;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1463 (.I0(n17885), .I1(n18168), .I2(n32923), 
            .I3(n30876), .O(n30950));
    defparam i1_2_lut_3_lut_4_lut_adj_1463.LUT_INIT = 16'h6996;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_1_i7_3_lut_4_lut (.I0(byte_transmit_counter[2]), 
            .I1(byte_transmit_counter[1]), .I2(n35404), .I3(n35402), .O(n7_adj_4284));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_1_i7_3_lut_4_lut.LUT_INIT = 16'hf2d0;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_0_i7_3_lut_4_lut (.I0(byte_transmit_counter[2]), 
            .I1(byte_transmit_counter[1]), .I2(n35401), .I3(n35399), .O(n7_adj_4285));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_0_i7_3_lut_4_lut.LUT_INIT = 16'hf2d0;
    SB_LUT4 i2_3_lut_4_lut_adj_1464 (.I0(n30866), .I1(n32816), .I2(n33133), 
            .I3(\data_out_frame[24] [6]), .O(n33020));
    defparam i2_3_lut_4_lut_adj_1464.LUT_INIT = 16'h6996;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_2_i7_3_lut_4_lut (.I0(byte_transmit_counter[2]), 
            .I1(byte_transmit_counter[1]), .I2(n35410), .I3(n35408), .O(n7_adj_4286));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_2_i7_3_lut_4_lut.LUT_INIT = 16'hf2d0;
    SB_LUT4 i2_3_lut_4_lut_adj_1465 (.I0(\data_out_frame[17] [7]), .I1(\data_out_frame[15] [6]), 
            .I2(n30108), .I3(\data_out_frame[15] [4]), .O(n33218));   // verilog/coms.v(74[16:43])
    defparam i2_3_lut_4_lut_adj_1465.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_adj_1466 (.I0(n30858), .I1(n33130), .I2(n30058), 
            .I3(n30948), .O(n30823));
    defparam i1_2_lut_4_lut_adj_1466.LUT_INIT = 16'h9669;
    SB_LUT4 mux_1387_i24_3_lut (.I0(\data_in_frame[17] [7]), .I1(\data_in_frame[1] [7]), 
            .I2(n5454), .I3(GND_net), .O(n5478));
    defparam mux_1387_i24_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_1387_i23_3_lut (.I0(\data_in_frame[17] [6]), .I1(\data_in_frame[1] [6]), 
            .I2(n5454), .I3(GND_net), .O(n5477));
    defparam mux_1387_i23_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_1387_i22_3_lut (.I0(\data_in_frame[17] [5]), .I1(\data_in_frame[1] [5]), 
            .I2(n5454), .I3(GND_net), .O(n5476));
    defparam mux_1387_i22_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_1387_i21_3_lut (.I0(\data_in_frame[17] [4]), .I1(\data_in_frame[1] [4]), 
            .I2(n5454), .I3(GND_net), .O(n5475));
    defparam mux_1387_i21_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_1387_i20_3_lut (.I0(\data_in_frame[17] [3]), .I1(\data_in_frame[1] [3]), 
            .I2(n5454), .I3(GND_net), .O(n5474));
    defparam mux_1387_i20_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_1387_i19_3_lut (.I0(\data_in_frame[17] [2]), .I1(\data_in_frame[1] [2]), 
            .I2(n5454), .I3(GND_net), .O(n5473));
    defparam mux_1387_i19_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_1387_i18_3_lut (.I0(\data_in_frame[17] [1]), .I1(\data_in_frame[1] [1]), 
            .I2(n5454), .I3(GND_net), .O(n5472));
    defparam mux_1387_i18_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_1387_i17_3_lut (.I0(\data_in_frame[17] [0]), .I1(\data_in_frame[1] [0]), 
            .I2(n5454), .I3(GND_net), .O(n5471));
    defparam mux_1387_i17_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_1387_i16_3_lut (.I0(\data_in_frame[18] [7]), .I1(\data_in_frame[2] [7]), 
            .I2(n5454), .I3(GND_net), .O(n5470));
    defparam mux_1387_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_1387_i15_3_lut (.I0(\data_in_frame[18] [6]), .I1(\data_in_frame[2] [6]), 
            .I2(n5454), .I3(GND_net), .O(n5469));
    defparam mux_1387_i15_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_1387_i14_3_lut (.I0(\data_in_frame[18] [5]), .I1(\data_in_frame[2] [5]), 
            .I2(n5454), .I3(GND_net), .O(n5468));
    defparam mux_1387_i14_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_1387_i13_3_lut (.I0(\data_in_frame[18] [4]), .I1(\data_in_frame[2] [4]), 
            .I2(n5454), .I3(GND_net), .O(n5467));
    defparam mux_1387_i13_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_1387_i12_3_lut (.I0(\data_in_frame[18] [3]), .I1(\data_in_frame[2] [3]), 
            .I2(n5454), .I3(GND_net), .O(n5466));
    defparam mux_1387_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_1387_i11_3_lut (.I0(\data_in_frame[18] [2]), .I1(\data_in_frame[2] [2]), 
            .I2(n5454), .I3(GND_net), .O(n5465));
    defparam mux_1387_i11_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_1387_i10_3_lut (.I0(\data_in_frame[18] [1]), .I1(\data_in_frame[2] [1]), 
            .I2(n5454), .I3(GND_net), .O(n5464));
    defparam mux_1387_i10_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_1387_i9_3_lut (.I0(\data_in_frame[18] [0]), .I1(\data_in_frame[2] [0]), 
            .I2(n5454), .I3(GND_net), .O(n5463));
    defparam mux_1387_i9_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_1387_i8_3_lut (.I0(\data_in_frame[19] [7]), .I1(\data_in_frame[3] [7]), 
            .I2(n5454), .I3(GND_net), .O(n5462));
    defparam mux_1387_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_1387_i7_3_lut (.I0(\data_in_frame[19] [6]), .I1(\data_in_frame[3] [6]), 
            .I2(n5454), .I3(GND_net), .O(n5461));
    defparam mux_1387_i7_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_1387_i6_3_lut (.I0(\data_in_frame[19] [5]), .I1(\data_in_frame[3] [5]), 
            .I2(n5454), .I3(GND_net), .O(n5460));
    defparam mux_1387_i6_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_1387_i5_3_lut (.I0(\data_in_frame[19] [4]), .I1(\data_in_frame[3] [4]), 
            .I2(n5454), .I3(GND_net), .O(n5459));
    defparam mux_1387_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i5_3_lut_4_lut_adj_1467 (.I0(\data_out_frame[18] [0]), .I1(\data_out_frame[15] [3]), 
            .I2(n10_adj_4023), .I3(\data_out_frame[17] [5]), .O(n30139));
    defparam i5_3_lut_4_lut_adj_1467.LUT_INIT = 16'h6996;
    SB_LUT4 i14048_3_lut_4_lut (.I0(n8_adj_4300), .I1(n32666), .I2(rx_data[7]), 
            .I3(\data_in_frame[9] [7]), .O(n19190));
    defparam i14048_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 mux_1387_i4_3_lut (.I0(\data_in_frame[19] [3]), .I1(\data_in_frame[3] [3]), 
            .I2(n5454), .I3(GND_net), .O(n5458));
    defparam mux_1387_i4_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_4_lut_adj_1468 (.I0(n18086), .I1(n32816), .I2(n30139), 
            .I3(n32981), .O(n32982));
    defparam i1_2_lut_4_lut_adj_1468.LUT_INIT = 16'h9669;
    SB_LUT4 i14049_3_lut_4_lut (.I0(n8_adj_4300), .I1(n32666), .I2(rx_data[6]), 
            .I3(\data_in_frame[9] [6]), .O(n19191));
    defparam i14049_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i14050_3_lut_4_lut (.I0(n8_adj_4300), .I1(n32666), .I2(rx_data[5]), 
            .I3(\data_in_frame[9] [5]), .O(n19192));
    defparam i14050_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i29820_2_lut (.I0(\data_out_frame[23] [4]), .I1(byte_transmit_counter[0]), 
            .I2(GND_net), .I3(GND_net), .O(n36292));
    defparam i29820_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i29822_2_lut (.I0(\data_out_frame[20] [4]), .I1(byte_transmit_counter[0]), 
            .I2(GND_net), .I3(GND_net), .O(n36291));
    defparam i29822_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i14051_3_lut_4_lut (.I0(n8_adj_4300), .I1(n32666), .I2(rx_data[4]), 
            .I3(\data_in_frame[9] [4]), .O(n19193));
    defparam i14051_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i14052_3_lut_4_lut (.I0(n8_adj_4300), .I1(n32666), .I2(rx_data[3]), 
            .I3(\data_in_frame[9] [3]), .O(n19194));
    defparam i14052_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 mux_1387_i3_3_lut (.I0(\data_in_frame[19] [2]), .I1(\data_in_frame[3] [2]), 
            .I2(n5454), .I3(GND_net), .O(n5457));
    defparam mux_1387_i3_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14053_3_lut_4_lut (.I0(n8_adj_4300), .I1(n32666), .I2(rx_data[2]), 
            .I3(\data_in_frame[9] [2]), .O(n19195));
    defparam i14053_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i14054_3_lut_4_lut (.I0(n8_adj_4300), .I1(n32666), .I2(rx_data[1]), 
            .I3(\data_in_frame[9] [1]), .O(n19196));
    defparam i14054_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_4_lut_adj_1469 (.I0(\data_out_frame[24] [3]), .I1(n32991), 
            .I2(n10_adj_4021), .I3(n30870), .O(n33000));
    defparam i1_2_lut_4_lut_adj_1469.LUT_INIT = 16'h9669;
    SB_LUT4 i14055_3_lut_4_lut (.I0(n8_adj_4300), .I1(n32666), .I2(rx_data[0]), 
            .I3(\data_in_frame[9] [0]), .O(n19197));
    defparam i14055_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_3_lut_4_lut_adj_1470 (.I0(\data_in_frame[2] [0]), .I1(\data_in_frame[0] [0]), 
            .I2(Kp_23__N_843), .I3(\data_in_frame[1] [6]), .O(n19_adj_4079));   // verilog/coms.v(73[16:42])
    defparam i2_3_lut_4_lut_adj_1470.LUT_INIT = 16'h6900;
    SB_LUT4 i1_2_lut_3_lut_adj_1471 (.I0(\data_out_frame[19] [7]), .I1(\data_out_frame[19] [6]), 
            .I2(n17098), .I3(GND_net), .O(n32975));   // verilog/coms.v(71[16:27])
    defparam i1_2_lut_3_lut_adj_1471.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1472 (.I0(\data_in_frame[2] [0]), .I1(\data_in_frame[0] [0]), 
            .I2(n32749), .I3(GND_net), .O(n33117));   // verilog/coms.v(73[16:42])
    defparam i1_2_lut_3_lut_adj_1472.LUT_INIT = 16'h9696;
    SB_LUT4 i14040_3_lut_4_lut (.I0(n8_adj_4302), .I1(n32666), .I2(rx_data[7]), 
            .I3(\data_in_frame[10] [7]), .O(n19182));
    defparam i14040_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i6_3_lut_4_lut (.I0(n17569), .I1(n32926), .I2(n18241), .I3(n17676), 
            .O(n17_adj_4051));
    defparam i6_3_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i14041_3_lut_4_lut (.I0(n8_adj_4302), .I1(n32666), .I2(rx_data[6]), 
            .I3(\data_in_frame[10] [6]), .O(n19183));
    defparam i14041_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i14042_3_lut_4_lut (.I0(n8_adj_4302), .I1(n32666), .I2(rx_data[5]), 
            .I3(\data_in_frame[10] [5]), .O(n19184));
    defparam i14042_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_3_lut_4_lut_adj_1473 (.I0(\data_out_frame[19] [7]), .I1(\data_out_frame[19] [6]), 
            .I2(\data_out_frame[18] [0]), .I3(\data_out_frame[17] [4]), 
            .O(n33007));   // verilog/coms.v(71[16:27])
    defparam i2_3_lut_4_lut_adj_1473.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_adj_1474 (.I0(\data_in_frame[4] [2]), .I1(\data_in_frame[2] [0]), 
            .I2(\data_in_frame[0] [0]), .I3(n32749), .O(n6));   // verilog/coms.v(78[16:27])
    defparam i1_2_lut_4_lut_adj_1474.LUT_INIT = 16'h6996;
    SB_LUT4 i14043_3_lut_4_lut (.I0(n8_adj_4302), .I1(n32666), .I2(rx_data[4]), 
            .I3(\data_in_frame[10] [4]), .O(n19185));
    defparam i14043_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i14044_3_lut_4_lut (.I0(n8_adj_4302), .I1(n32666), .I2(rx_data[3]), 
            .I3(\data_in_frame[10] [3]), .O(n19186));
    defparam i14044_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i14045_3_lut_4_lut (.I0(n8_adj_4302), .I1(n32666), .I2(rx_data[2]), 
            .I3(\data_in_frame[10] [2]), .O(n19187));
    defparam i14045_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i14046_3_lut_4_lut (.I0(n8_adj_4302), .I1(n32666), .I2(rx_data[1]), 
            .I3(\data_in_frame[10] [1]), .O(n19188));
    defparam i14046_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i14047_3_lut_4_lut (.I0(n8_adj_4302), .I1(n32666), .I2(rx_data[0]), 
            .I3(\data_in_frame[10] [0]), .O(n19189));
    defparam i14047_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i14032_3_lut_4_lut (.I0(n8_adj_4303), .I1(n32666), .I2(rx_data[7]), 
            .I3(\data_in_frame[11] [7]), .O(n19174));
    defparam i14032_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i14033_3_lut_4_lut (.I0(n8_adj_4303), .I1(n32666), .I2(rx_data[6]), 
            .I3(\data_in_frame[11] [6]), .O(n19175));
    defparam i14033_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i14034_3_lut_4_lut (.I0(n8_adj_4303), .I1(n32666), .I2(rx_data[5]), 
            .I3(\data_in_frame[11] [5]), .O(n19176));
    defparam i14034_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i14035_3_lut_4_lut (.I0(n8_adj_4303), .I1(n32666), .I2(rx_data[4]), 
            .I3(\data_in_frame[11] [4]), .O(n19177));
    defparam i14035_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i14036_3_lut_4_lut (.I0(n8_adj_4303), .I1(n32666), .I2(rx_data[3]), 
            .I3(\data_in_frame[11] [3]), .O(n19178));
    defparam i14036_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i14037_3_lut_4_lut (.I0(n8_adj_4303), .I1(n32666), .I2(rx_data[2]), 
            .I3(\data_in_frame[11] [2]), .O(n19179));
    defparam i14037_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i14038_3_lut_4_lut (.I0(n8_adj_4303), .I1(n32666), .I2(rx_data[1]), 
            .I3(\data_in_frame[11] [1]), .O(n19180));
    defparam i14038_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i14039_3_lut_4_lut (.I0(n8_adj_4303), .I1(n32666), .I2(rx_data[0]), 
            .I3(\data_in_frame[11] [0]), .O(n19181));
    defparam i14039_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_3_lut_4_lut_adj_1475 (.I0(\data_in_frame[8] [6]), .I1(n8), 
            .I2(n33344), .I3(Kp_23__N_1069), .O(n18460));   // verilog/coms.v(77[16:43])
    defparam i2_3_lut_4_lut_adj_1475.LUT_INIT = 16'h6996;
    SB_LUT4 i2_2_lut_3_lut_adj_1476 (.I0(\data_out_frame[17] [6]), .I1(\data_out_frame[20] [0]), 
            .I2(\data_out_frame[24] [0]), .I3(GND_net), .O(n10_c));
    defparam i2_2_lut_3_lut_adj_1476.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_4_lut_adj_1477 (.I0(\data_in_frame[8] [6]), .I1(n8), 
            .I2(\data_in_frame[8] [0]), .I3(n17730), .O(n33108));   // verilog/coms.v(77[16:43])
    defparam i2_3_lut_4_lut_adj_1477.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_1478 (.I0(\data_in_frame[9] [7]), .I1(\data_in_frame[9] [6]), 
            .I2(n17894), .I3(n17885), .O(n29786));   // verilog/coms.v(85[17:28])
    defparam i2_3_lut_4_lut_adj_1478.LUT_INIT = 16'h6996;
    SB_LUT4 i2_2_lut_4_lut_adj_1479 (.I0(n17126), .I1(n33865), .I2(n30908), 
            .I3(n18363), .O(n7_adj_4029));
    defparam i2_2_lut_4_lut_adj_1479.LUT_INIT = 16'h6996;
    SB_LUT4 i5_3_lut_4_lut_adj_1480 (.I0(\data_in_frame[9] [7]), .I1(\data_in_frame[9] [6]), 
            .I2(n10_adj_4182), .I3(n15920), .O(n33268));   // verilog/coms.v(85[17:28])
    defparam i5_3_lut_4_lut_adj_1480.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1481 (.I0(\data_in_frame[9] [7]), .I1(\data_in_frame[9] [6]), 
            .I2(\data_in_frame[9] [5]), .I3(GND_net), .O(n32923));   // verilog/coms.v(85[17:28])
    defparam i1_2_lut_3_lut_adj_1481.LUT_INIT = 16'h9696;
    SB_LUT4 i1_3_lut_adj_1482 (.I0(\FRAME_MATCHER.state_c [2]), .I1(n63_adj_4103), 
            .I2(n63_adj_4106), .I3(GND_net), .O(n20830));   // verilog/coms.v(112[11:16])
    defparam i1_3_lut_adj_1482.LUT_INIT = 16'hb3b3;
    SB_LUT4 select_450_Select_2_i5_4_lut (.I0(n3303), .I1(n39), .I2(n63), 
            .I3(n20830), .O(n5));
    defparam select_450_Select_2_i5_4_lut.LUT_INIT = 16'h3222;
    SB_LUT4 i1_rep_297_2_lut (.I0(n63), .I1(n20830), .I2(GND_net), .I3(GND_net), 
            .O(n38579));   // verilog/coms.v(112[11:16])
    defparam i1_rep_297_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_3_lut_adj_1483 (.I0(n30545), .I1(n18285), .I2(\data_in_frame[11] [5]), 
            .I3(GND_net), .O(n30880));
    defparam i1_2_lut_3_lut_adj_1483.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1484 (.I0(n30545), .I1(n18285), .I2(\data_in_frame[9] [4]), 
            .I3(GND_net), .O(n30872));
    defparam i1_2_lut_3_lut_adj_1484.LUT_INIT = 16'h9696;
    uart_tx tx (.clk32MHz(clk32MHz), .n18738(n18738), .n18956(n18956), 
            .tx_o(tx_o), .tx_data({tx_data}), .r_SM_Main({r_SM_Main}), 
            .GND_net(GND_net), .VCC_net(VCC_net), .\r_SM_Main_2__N_3490[0] (r_SM_Main_2__N_3490[0]), 
            .\r_SM_Main_2__N_3487[1] (\r_SM_Main_2__N_3487[1] ), .n4(n4), 
            .\r_Bit_Index[0] (\r_Bit_Index[0] ), .n19052(n19052), .tx_active(tx_active), 
            .n19460(n19460), .n38214(n38214), .tx_enable(tx_enable), .n10524(n10524)) /* synthesis syn_module_defined=1 */ ;   // verilog/coms.v(107[10:70])
    uart_rx rx (.n18732(n18732), .clk32MHz(clk32MHz), .n18954(n18954), 
            .GND_net(GND_net), .r_Rx_Data(r_Rx_Data), .RX_N_10(RX_N_10), 
            .VCC_net(VCC_net), .\r_Bit_Index[0] (\r_Bit_Index[0]_adj_9 ), 
            .n23879(n23879), .n4(n4_adj_10), .n4_adj_6(n4_adj_11), .n17539(n17539), 
            .n19524(n19524), .rx_data_ready(rx_data_ready), .n19583(n19583), 
            .rx_data({rx_data}), .n19035(n19035), .n19034(n19034), .n19033(n19033), 
            .n19032(n19032), .n19031(n19031), .n19030(n19030), .n19029(n19029), 
            .n17534(n17534), .n4_adj_7(n4_adj_12)) /* synthesis syn_module_defined=1 */ ;   // verilog/coms.v(93[10:44])
    
endmodule
//
// Verilog Description of module uart_tx
//

module uart_tx (clk32MHz, n18738, n18956, tx_o, tx_data, r_SM_Main, 
            GND_net, VCC_net, \r_SM_Main_2__N_3490[0] , \r_SM_Main_2__N_3487[1] , 
            n4, \r_Bit_Index[0] , n19052, tx_active, n19460, n38214, 
            tx_enable, n10524) /* synthesis syn_module_defined=1 */ ;
    input clk32MHz;
    output n18738;
    output n18956;
    output tx_o;
    input [7:0]tx_data;
    output [2:0]r_SM_Main;
    input GND_net;
    input VCC_net;
    input \r_SM_Main_2__N_3490[0] ;
    output \r_SM_Main_2__N_3487[1] ;
    output n4;
    output \r_Bit_Index[0] ;
    input n19052;
    output tx_active;
    input n19460;
    input n38214;
    output tx_enable;
    output n10524;
    
    wire clk32MHz /* synthesis SET_AS_NETWORK=clk32MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(33[6:14])
    wire [8:0]n41;
    
    wire n1;
    wire [8:0]r_Clock_Count;   // verilog/uart_tx.v(32[16:29])
    
    wire n18920;
    wire [2:0]n307;
    wire [2:0]r_Bit_Index;   // verilog/uart_tx.v(33[16:27])
    
    wire n3, n14784;
    wire [7:0]r_Tx_Data;   // verilog/uart_tx.v(34[16:25])
    
    wire n12453, n28612, n28611, n28610, n28609, n28608, n28607, 
        n28606, n28605, n24300, n12452, n37895, n37739, o_Tx_Serial_N_3518, 
        n10, n34484, n37892, n37736, n3_adj_4020;
    
    SB_DFFESR r_Clock_Count_1584__i8 (.Q(r_Clock_Count[8]), .C(clk32MHz), 
            .E(n1), .D(n41[8]), .R(n18920));   // verilog/uart_tx.v(118[34:51])
    SB_DFFESR r_Clock_Count_1584__i7 (.Q(r_Clock_Count[7]), .C(clk32MHz), 
            .E(n1), .D(n41[7]), .R(n18920));   // verilog/uart_tx.v(118[34:51])
    SB_DFFESR r_Clock_Count_1584__i6 (.Q(r_Clock_Count[6]), .C(clk32MHz), 
            .E(n1), .D(n41[6]), .R(n18920));   // verilog/uart_tx.v(118[34:51])
    SB_DFFESR r_Clock_Count_1584__i5 (.Q(r_Clock_Count[5]), .C(clk32MHz), 
            .E(n1), .D(n41[5]), .R(n18920));   // verilog/uart_tx.v(118[34:51])
    SB_DFFESR r_Clock_Count_1584__i4 (.Q(r_Clock_Count[4]), .C(clk32MHz), 
            .E(n1), .D(n41[4]), .R(n18920));   // verilog/uart_tx.v(118[34:51])
    SB_DFFESR r_Clock_Count_1584__i3 (.Q(r_Clock_Count[3]), .C(clk32MHz), 
            .E(n1), .D(n41[3]), .R(n18920));   // verilog/uart_tx.v(118[34:51])
    SB_DFFESR r_Bit_Index_i2 (.Q(r_Bit_Index[2]), .C(clk32MHz), .E(n18738), 
            .D(n307[2]), .R(n18956));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFESR r_Bit_Index_i1 (.Q(r_Bit_Index[1]), .C(clk32MHz), .E(n18738), 
            .D(n307[1]), .R(n18956));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFESR r_Clock_Count_1584__i2 (.Q(r_Clock_Count[2]), .C(clk32MHz), 
            .E(n1), .D(n41[2]), .R(n18920));   // verilog/uart_tx.v(118[34:51])
    SB_DFFESR r_Clock_Count_1584__i1 (.Q(r_Clock_Count[1]), .C(clk32MHz), 
            .E(n1), .D(n41[1]), .R(n18920));   // verilog/uart_tx.v(118[34:51])
    SB_DFFESR r_Clock_Count_1584__i0 (.Q(r_Clock_Count[0]), .C(clk32MHz), 
            .E(n1), .D(n41[0]), .R(n18920));   // verilog/uart_tx.v(118[34:51])
    SB_DFFE o_Tx_Serial_45 (.Q(tx_o), .C(clk32MHz), .E(n1), .D(n3));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFE r_Tx_Data_i0 (.Q(r_Tx_Data[0]), .C(clk32MHz), .E(n14784), 
            .D(tx_data[0]));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFSR r_SM_Main_i0 (.Q(r_SM_Main[0]), .C(clk32MHz), .D(n12453), 
            .R(r_SM_Main[2]));   // verilog/uart_tx.v(40[10] 143[8])
    SB_LUT4 r_Clock_Count_1584_add_4_10_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[8]), .I3(n28612), .O(n41[8])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1584_add_4_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 r_Clock_Count_1584_add_4_9_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[7]), .I3(n28611), .O(n41[7])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1584_add_4_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_1584_add_4_9 (.CI(n28611), .I0(GND_net), .I1(r_Clock_Count[7]), 
            .CO(n28612));
    SB_LUT4 r_Clock_Count_1584_add_4_8_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[6]), .I3(n28610), .O(n41[6])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1584_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_1584_add_4_8 (.CI(n28610), .I0(GND_net), .I1(r_Clock_Count[6]), 
            .CO(n28611));
    SB_LUT4 r_Clock_Count_1584_add_4_7_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[5]), .I3(n28609), .O(n41[5])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1584_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_1584_add_4_7 (.CI(n28609), .I0(GND_net), .I1(r_Clock_Count[5]), 
            .CO(n28610));
    SB_LUT4 r_Clock_Count_1584_add_4_6_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[4]), .I3(n28608), .O(n41[4])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1584_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_1584_add_4_6 (.CI(n28608), .I0(GND_net), .I1(r_Clock_Count[4]), 
            .CO(n28609));
    SB_LUT4 r_Clock_Count_1584_add_4_5_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[3]), .I3(n28607), .O(n41[3])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1584_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_1584_add_4_5 (.CI(n28607), .I0(GND_net), .I1(r_Clock_Count[3]), 
            .CO(n28608));
    SB_LUT4 r_Clock_Count_1584_add_4_4_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[2]), .I3(n28606), .O(n41[2])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1584_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_1584_add_4_4 (.CI(n28606), .I0(GND_net), .I1(r_Clock_Count[2]), 
            .CO(n28607));
    SB_LUT4 r_Clock_Count_1584_add_4_3_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[1]), .I3(n28605), .O(n41[1])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1584_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_1584_add_4_3 (.CI(n28605), .I0(GND_net), .I1(r_Clock_Count[1]), 
            .CO(n28606));
    SB_LUT4 r_Clock_Count_1584_add_4_2_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[0]), .I3(VCC_net), .O(n41[0])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1584_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_1584_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(r_Clock_Count[0]), 
            .CO(n28605));
    SB_LUT4 i7391_4_lut (.I0(\r_SM_Main_2__N_3490[0] ), .I1(n24300), .I2(r_SM_Main[1]), 
            .I3(\r_SM_Main_2__N_3487[1] ), .O(n12452));   // verilog/uart_tx.v(43[7] 142[14])
    defparam i7391_4_lut.LUT_INIT = 16'hca0a;
    SB_LUT4 i7392_3_lut (.I0(n12452), .I1(\r_SM_Main_2__N_3487[1] ), .I2(r_SM_Main[0]), 
            .I3(GND_net), .O(n12453));   // verilog/uart_tx.v(43[7] 142[14])
    defparam i7392_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i1986372_i1_3_lut (.I0(n37895), .I1(n37739), .I2(r_Bit_Index[2]), 
            .I3(GND_net), .O(o_Tx_Serial_N_3518));
    defparam i1986372_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 r_SM_Main_2__I_0_56_i3_3_lut (.I0(r_SM_Main[0]), .I1(o_Tx_Serial_N_3518), 
            .I2(r_SM_Main[1]), .I3(GND_net), .O(n3));   // verilog/uart_tx.v(43[7] 142[14])
    defparam r_SM_Main_2__I_0_56_i3_3_lut.LUT_INIT = 16'he5e5;
    SB_LUT4 i1_3_lut_4_lut_4_lut (.I0(\r_SM_Main_2__N_3487[1] ), .I1(r_SM_Main[0]), 
            .I2(r_SM_Main[1]), .I3(r_SM_Main[2]), .O(n4));   // verilog/uart_tx.v(43[7] 142[14])
    defparam i1_3_lut_4_lut_4_lut.LUT_INIT = 16'h008f;
    SB_LUT4 i1684_2_lut (.I0(r_Bit_Index[1]), .I1(\r_Bit_Index[0] ), .I2(GND_net), 
            .I3(GND_net), .O(n307[1]));   // verilog/uart_tx.v(98[36:51])
    defparam i1684_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[2]), .I2(\r_Bit_Index[0] ), 
            .I3(GND_net), .O(n24300));
    defparam i2_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 i13814_3_lut (.I0(n18738), .I1(n24300), .I2(r_SM_Main[1]), 
            .I3(GND_net), .O(n18956));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i13814_3_lut.LUT_INIT = 16'h8a8a;
    SB_LUT4 i1691_3_lut (.I0(r_Bit_Index[2]), .I1(r_Bit_Index[1]), .I2(\r_Bit_Index[0] ), 
            .I3(GND_net), .O(n307[2]));   // verilog/uart_tx.v(98[36:51])
    defparam i1691_3_lut.LUT_INIT = 16'h6a6a;
    SB_LUT4 i4_4_lut (.I0(r_Clock_Count[1]), .I1(r_Clock_Count[5]), .I2(r_Clock_Count[0]), 
            .I3(r_Clock_Count[2]), .O(n10));
    defparam i4_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i5_3_lut (.I0(r_Clock_Count[3]), .I1(n10), .I2(r_Clock_Count[4]), 
            .I3(GND_net), .O(n34484));
    defparam i5_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 i3_4_lut (.I0(n34484), .I1(r_Clock_Count[8]), .I2(r_Clock_Count[6]), 
            .I3(r_Clock_Count[7]), .O(\r_SM_Main_2__N_3487[1] ));
    defparam i3_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i30393_4_lut (.I0(r_SM_Main[2]), .I1(\r_SM_Main_2__N_3487[1] ), 
            .I2(r_SM_Main[1]), .I3(r_SM_Main[0]), .O(n18920));
    defparam i30393_4_lut.LUT_INIT = 16'h4445;
    SB_LUT4 i1_1_lut (.I0(r_SM_Main[2]), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n1));
    defparam i1_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 r_Bit_Index_0__bdd_4_lut (.I0(\r_Bit_Index[0] ), .I1(r_Tx_Data[2]), 
            .I2(r_Tx_Data[3]), .I3(r_Bit_Index[1]), .O(n37892));
    defparam r_Bit_Index_0__bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_LUT4 n37892_bdd_4_lut (.I0(n37892), .I1(r_Tx_Data[1]), .I2(r_Tx_Data[0]), 
            .I3(r_Bit_Index[1]), .O(n37895));
    defparam n37892_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 r_Bit_Index_0__bdd_4_lut_31095 (.I0(\r_Bit_Index[0] ), .I1(r_Tx_Data[6]), 
            .I2(r_Tx_Data[7]), .I3(r_Bit_Index[1]), .O(n37736));
    defparam r_Bit_Index_0__bdd_4_lut_31095.LUT_INIT = 16'he4aa;
    SB_LUT4 n37736_bdd_4_lut (.I0(n37736), .I1(r_Tx_Data[5]), .I2(r_Tx_Data[4]), 
            .I3(r_Bit_Index[1]), .O(n37739));
    defparam n37736_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFFE r_Tx_Data_i1 (.Q(r_Tx_Data[1]), .C(clk32MHz), .E(n14784), 
            .D(tx_data[1]));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFE r_Tx_Data_i2 (.Q(r_Tx_Data[2]), .C(clk32MHz), .E(n14784), 
            .D(tx_data[2]));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFE r_Tx_Data_i3 (.Q(r_Tx_Data[3]), .C(clk32MHz), .E(n14784), 
            .D(tx_data[3]));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFE r_Tx_Data_i4 (.Q(r_Tx_Data[4]), .C(clk32MHz), .E(n14784), 
            .D(tx_data[4]));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFE r_Tx_Data_i5 (.Q(r_Tx_Data[5]), .C(clk32MHz), .E(n14784), 
            .D(tx_data[5]));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFE r_Tx_Data_i6 (.Q(r_Tx_Data[6]), .C(clk32MHz), .E(n14784), 
            .D(tx_data[6]));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFE r_Tx_Data_i7 (.Q(r_Tx_Data[7]), .C(clk32MHz), .E(n14784), 
            .D(tx_data[7]));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFSR r_SM_Main_i1 (.Q(r_SM_Main[1]), .C(clk32MHz), .D(n3_adj_4020), 
            .R(r_SM_Main[2]));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFF r_Tx_Active_47 (.Q(tx_active), .C(clk32MHz), .D(n19052));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFF r_Bit_Index_i0 (.Q(\r_Bit_Index[0] ), .C(clk32MHz), .D(n19460));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFF r_SM_Main_i2 (.Q(r_SM_Main[2]), .C(clk32MHz), .D(n38214));   // verilog/uart_tx.v(40[10] 143[8])
    SB_LUT4 i2_3_lut_4_lut (.I0(r_SM_Main[2]), .I1(r_SM_Main[0]), .I2(\r_SM_Main_2__N_3490[0] ), 
            .I3(r_SM_Main[1]), .O(n14784));
    defparam i2_3_lut_4_lut.LUT_INIT = 16'h0010;
    SB_LUT4 i1_3_lut_4_lut (.I0(r_SM_Main[2]), .I1(r_SM_Main[0]), .I2(r_SM_Main[1]), 
            .I3(\r_SM_Main_2__N_3487[1] ), .O(n18738));
    defparam i1_3_lut_4_lut.LUT_INIT = 16'h1101;
    SB_LUT4 i9460_2_lut_3_lut (.I0(\r_SM_Main_2__N_3487[1] ), .I1(r_SM_Main[0]), 
            .I2(r_SM_Main[1]), .I3(GND_net), .O(n3_adj_4020));   // verilog/uart_tx.v(43[7] 142[14])
    defparam i9460_2_lut_3_lut.LUT_INIT = 16'h7878;
    SB_LUT4 o_Tx_Serial_I_0_1_lut (.I0(tx_o), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(tx_enable));   // verilog/uart_tx.v(38[24:36])
    defparam o_Tx_Serial_I_0_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i5471_2_lut (.I0(\r_SM_Main_2__N_3490[0] ), .I1(r_SM_Main[0]), 
            .I2(GND_net), .I3(GND_net), .O(n10524));   // verilog/uart_tx.v(43[7] 142[14])
    defparam i5471_2_lut.LUT_INIT = 16'h2222;
    
endmodule
//
// Verilog Description of module uart_rx
//

module uart_rx (n18732, clk32MHz, n18954, GND_net, r_Rx_Data, RX_N_10, 
            VCC_net, \r_Bit_Index[0] , n23879, n4, n4_adj_6, n17539, 
            n19524, rx_data_ready, n19583, rx_data, n19035, n19034, 
            n19033, n19032, n19031, n19030, n19029, n17534, n4_adj_7) /* synthesis syn_module_defined=1 */ ;
    output n18732;
    input clk32MHz;
    output n18954;
    input GND_net;
    output r_Rx_Data;
    input RX_N_10;
    input VCC_net;
    output \r_Bit_Index[0] ;
    output n23879;
    output n4;
    output n4_adj_6;
    output n17539;
    input n19524;
    output rx_data_ready;
    input n19583;
    output [7:0]rx_data;
    input n19035;
    input n19034;
    input n19033;
    input n19032;
    input n19031;
    input n19030;
    input n19029;
    output n17534;
    output n4_adj_7;
    
    wire clk32MHz /* synthesis SET_AS_NETWORK=clk32MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(33[6:14])
    wire [2:0]n326;
    wire [2:0]r_Bit_Index;   // verilog/uart_rx.v(33[17:28])
    wire [7:0]n37;
    
    wire n18687;
    wire [7:0]r_Clock_Count;   // verilog/uart_rx.v(32[17:30])
    
    wire n18918;
    wire [2:0]r_SM_Main_2__N_3416;
    wire [2:0]r_SM_Main;   // verilog/uart_rx.v(36[17:26])
    
    wire n32642, n24649, n21649, n3, n21655, r_Rx_Data_R, n28604, 
        n28603, n28602, n28601, n28600, n28599, n28598, n21641, 
        n24291, n24591, n21654, n31, n5, n8, n6, n17343, n32269, 
        n18626;
    
    SB_DFFESR r_Bit_Index_i2 (.Q(r_Bit_Index[2]), .C(clk32MHz), .E(n18732), 
            .D(n326[2]), .R(n18954));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFFESR r_Bit_Index_i1 (.Q(r_Bit_Index[1]), .C(clk32MHz), .E(n18732), 
            .D(n326[1]), .R(n18954));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFFESR r_Clock_Count_1582__i7 (.Q(r_Clock_Count[7]), .C(clk32MHz), 
            .E(n18687), .D(n37[7]), .R(n18918));   // verilog/uart_rx.v(120[34:51])
    SB_DFFESR r_Clock_Count_1582__i6 (.Q(r_Clock_Count[6]), .C(clk32MHz), 
            .E(n18687), .D(n37[6]), .R(n18918));   // verilog/uart_rx.v(120[34:51])
    SB_DFFESR r_Clock_Count_1582__i5 (.Q(r_Clock_Count[5]), .C(clk32MHz), 
            .E(n18687), .D(n37[5]), .R(n18918));   // verilog/uart_rx.v(120[34:51])
    SB_DFFESR r_Clock_Count_1582__i4 (.Q(r_Clock_Count[4]), .C(clk32MHz), 
            .E(n18687), .D(n37[4]), .R(n18918));   // verilog/uart_rx.v(120[34:51])
    SB_DFFESR r_Clock_Count_1582__i3 (.Q(r_Clock_Count[3]), .C(clk32MHz), 
            .E(n18687), .D(n37[3]), .R(n18918));   // verilog/uart_rx.v(120[34:51])
    SB_DFFSR r_SM_Main_i2 (.Q(r_SM_Main[2]), .C(clk32MHz), .D(r_SM_Main_2__N_3416[2]), 
            .R(n32642));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFFESR r_Clock_Count_1582__i0 (.Q(r_Clock_Count[0]), .C(clk32MHz), 
            .E(n18687), .D(n37[0]), .R(n18918));   // verilog/uart_rx.v(120[34:51])
    SB_DFFESR r_Clock_Count_1582__i2 (.Q(r_Clock_Count[2]), .C(clk32MHz), 
            .E(n18687), .D(n37[2]), .R(n18918));   // verilog/uart_rx.v(120[34:51])
    SB_DFFESR r_Clock_Count_1582__i1 (.Q(r_Clock_Count[1]), .C(clk32MHz), 
            .E(n18687), .D(n37[1]), .R(n18918));   // verilog/uart_rx.v(120[34:51])
    SB_LUT4 i19506_2_lut (.I0(r_SM_Main_2__N_3416[2]), .I1(r_SM_Main[0]), 
            .I2(GND_net), .I3(GND_net), .O(n24649));
    defparam i19506_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i16517_4_lut (.I0(r_Rx_Data), .I1(n24649), .I2(r_SM_Main[1]), 
            .I3(n21649), .O(n3));   // verilog/uart_rx.v(36[17:26])
    defparam i16517_4_lut.LUT_INIT = 16'h3530;
    SB_DFFSR r_SM_Main_i0 (.Q(r_SM_Main[0]), .C(clk32MHz), .D(n21655), 
            .R(r_SM_Main[2]));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_Data_50 (.Q(r_Rx_Data), .C(clk32MHz), .D(r_Rx_Data_R));   // verilog/uart_rx.v(41[10] 45[8])
    SB_DFF r_Rx_Data_R_49 (.Q(r_Rx_Data_R), .C(clk32MHz), .D(RX_N_10));   // verilog/uart_rx.v(41[10] 45[8])
    SB_LUT4 r_Clock_Count_1582_add_4_9_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[7]), .I3(n28604), .O(n37[7])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1582_add_4_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 r_Clock_Count_1582_add_4_8_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[6]), .I3(n28603), .O(n37[6])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1582_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_1582_add_4_8 (.CI(n28603), .I0(GND_net), .I1(r_Clock_Count[6]), 
            .CO(n28604));
    SB_LUT4 r_Clock_Count_1582_add_4_7_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[5]), .I3(n28602), .O(n37[5])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1582_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_1582_add_4_7 (.CI(n28602), .I0(GND_net), .I1(r_Clock_Count[5]), 
            .CO(n28603));
    SB_LUT4 r_Clock_Count_1582_add_4_6_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[4]), .I3(n28601), .O(n37[4])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1582_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_1582_add_4_6 (.CI(n28601), .I0(GND_net), .I1(r_Clock_Count[4]), 
            .CO(n28602));
    SB_LUT4 r_Clock_Count_1582_add_4_5_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[3]), .I3(n28600), .O(n37[3])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1582_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_1582_add_4_5 (.CI(n28600), .I0(GND_net), .I1(r_Clock_Count[3]), 
            .CO(n28601));
    SB_LUT4 r_Clock_Count_1582_add_4_4_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[2]), .I3(n28599), .O(n37[2])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1582_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_1582_add_4_4 (.CI(n28599), .I0(GND_net), .I1(r_Clock_Count[2]), 
            .CO(n28600));
    SB_LUT4 r_Clock_Count_1582_add_4_3_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[1]), .I3(n28598), .O(n37[1])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1582_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_1582_add_4_3 (.CI(n28598), .I0(GND_net), .I1(r_Clock_Count[1]), 
            .CO(n28599));
    SB_LUT4 r_Clock_Count_1582_add_4_2_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[0]), .I3(VCC_net), .O(n37[0])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1582_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_1582_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(r_Clock_Count[0]), 
            .CO(n28598));
    SB_LUT4 i1_2_lut (.I0(r_SM_Main[0]), .I1(n21641), .I2(GND_net), .I3(GND_net), 
            .O(n21649));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i1_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 r_SM_Main_2__I_0_56_Mux_0_i2_3_lut (.I0(n24291), .I1(r_SM_Main_2__N_3416[2]), 
            .I2(r_SM_Main[0]), .I3(GND_net), .O(n24591));   // verilog/uart_rx.v(52[7] 143[14])
    defparam r_SM_Main_2__I_0_56_Mux_0_i2_3_lut.LUT_INIT = 16'hc7c7;
    SB_LUT4 i16521_3_lut (.I0(n21654), .I1(n24591), .I2(r_SM_Main[1]), 
            .I3(GND_net), .O(n21655));   // verilog/uart_rx.v(36[17:26])
    defparam i16521_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i3_4_lut (.I0(r_Clock_Count[2]), .I1(r_Clock_Count[5]), .I2(n31), 
            .I3(n5), .O(n21641));
    defparam i3_4_lut.LUT_INIT = 16'hfdff;
    SB_LUT4 i13776_3_lut (.I0(n18687), .I1(r_SM_Main[2]), .I2(n8), .I3(GND_net), 
            .O(n18918));   // verilog/uart_rx.v(120[34:51])
    defparam i13776_3_lut.LUT_INIT = 16'h8a8a;
    SB_LUT4 i2_2_lut (.I0(n21641), .I1(r_SM_Main[0]), .I2(GND_net), .I3(GND_net), 
            .O(n6));   // verilog/uart_rx.v(36[17:26])
    defparam i2_2_lut.LUT_INIT = 16'hbbbb;
    SB_LUT4 i1_4_lut (.I0(r_SM_Main[1]), .I1(r_SM_Main[2]), .I2(n6), .I3(r_Rx_Data), 
            .O(n18687));   // verilog/uart_rx.v(36[17:26])
    defparam i1_4_lut.LUT_INIT = 16'h3233;
    SB_LUT4 i1662_2_lut (.I0(r_Bit_Index[1]), .I1(\r_Bit_Index[0] ), .I2(GND_net), 
            .I3(GND_net), .O(n326[1]));   // verilog/uart_rx.v(102[36:51])
    defparam i1662_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_841 (.I0(r_Clock_Count[1]), .I1(r_Clock_Count[0]), 
            .I2(r_Clock_Count[4]), .I3(r_Clock_Count[3]), .O(n5));
    defparam i3_4_lut_adj_841.LUT_INIT = 16'h8000;
    SB_LUT4 i1_2_lut_adj_842 (.I0(r_Clock_Count[7]), .I1(r_Clock_Count[6]), 
            .I2(GND_net), .I3(GND_net), .O(n31));   // verilog/uart_rx.v(120[34:51])
    defparam i1_2_lut_adj_842.LUT_INIT = 16'heeee;
    SB_LUT4 i19160_4_lut (.I0(r_Clock_Count[5]), .I1(n31), .I2(r_Clock_Count[2]), 
            .I3(n5), .O(r_SM_Main_2__N_3416[2]));
    defparam i19160_4_lut.LUT_INIT = 16'heccc;
    SB_LUT4 i2_3_lut (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[2]), .I2(\r_Bit_Index[0] ), 
            .I3(GND_net), .O(n24291));
    defparam i2_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 i13812_3_lut (.I0(n18732), .I1(n24291), .I2(r_SM_Main[1]), 
            .I3(GND_net), .O(n18954));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i13812_3_lut.LUT_INIT = 16'h8a8a;
    SB_LUT4 i2_4_lut (.I0(r_SM_Main[2]), .I1(r_SM_Main_2__N_3416[2]), .I2(r_SM_Main[0]), 
            .I3(r_SM_Main[1]), .O(n18732));
    defparam i2_4_lut.LUT_INIT = 16'h0405;
    SB_LUT4 i1669_3_lut (.I0(r_Bit_Index[2]), .I1(r_Bit_Index[1]), .I2(\r_Bit_Index[0] ), 
            .I3(GND_net), .O(n326[2]));   // verilog/uart_rx.v(102[36:51])
    defparam i1669_3_lut.LUT_INIT = 16'h6a6a;
    SB_LUT4 i16520_3_lut_4_lut_3_lut (.I0(r_SM_Main[0]), .I1(n21641), .I2(r_Rx_Data), 
            .I3(GND_net), .O(n21654));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i16520_3_lut_4_lut_3_lut.LUT_INIT = 16'h8d8d;
    SB_LUT4 i18752_2_lut (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[2]), .I2(GND_net), 
            .I3(GND_net), .O(n23879));
    defparam i18752_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 equal_148_i4_2_lut (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[2]), 
            .I2(GND_net), .I3(GND_net), .O(n4));   // verilog/uart_rx.v(97[17:39])
    defparam equal_148_i4_2_lut.LUT_INIT = 16'hbbbb;
    SB_LUT4 equal_150_i4_2_lut (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[2]), 
            .I2(GND_net), .I3(GND_net), .O(n4_adj_6));   // verilog/uart_rx.v(97[17:39])
    defparam equal_150_i4_2_lut.LUT_INIT = 16'hdddd;
    SB_LUT4 i1_2_lut_adj_843 (.I0(n17343), .I1(\r_Bit_Index[0] ), .I2(GND_net), 
            .I3(GND_net), .O(n17539));   // verilog/uart_rx.v(52[7] 143[14])
    defparam i1_2_lut_adj_843.LUT_INIT = 16'hbbbb;
    SB_DFFSR r_SM_Main_i1 (.Q(r_SM_Main[1]), .C(clk32MHz), .D(n3), .R(r_SM_Main[2]));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Bit_Index_i0 (.Q(\r_Bit_Index[0] ), .C(clk32MHz), .D(n19524));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_DV_52 (.Q(rx_data_ready), .C(clk32MHz), .D(n32269));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_Byte_i0 (.Q(rx_data[0]), .C(clk32MHz), .D(n19583));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_Byte_i1 (.Q(rx_data[1]), .C(clk32MHz), .D(n19035));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_Byte_i2 (.Q(rx_data[2]), .C(clk32MHz), .D(n19034));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_Byte_i3 (.Q(rx_data[3]), .C(clk32MHz), .D(n19033));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_Byte_i4 (.Q(rx_data[4]), .C(clk32MHz), .D(n19032));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_Byte_i5 (.Q(rx_data[5]), .C(clk32MHz), .D(n19031));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_Byte_i6 (.Q(rx_data[6]), .C(clk32MHz), .D(n19030));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_Byte_i7 (.Q(rx_data[7]), .C(clk32MHz), .D(n19029));   // verilog/uart_rx.v(49[10] 144[8])
    SB_LUT4 i19_3_lut_4_lut (.I0(r_SM_Main[0]), .I1(n21641), .I2(r_SM_Main[1]), 
            .I3(r_SM_Main_2__N_3416[2]), .O(n8));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i19_3_lut_4_lut.LUT_INIT = 16'h08f8;
    SB_LUT4 i21_4_lut_4_lut (.I0(r_SM_Main[1]), .I1(r_SM_Main[2]), .I2(r_SM_Main_2__N_3416[2]), 
            .I3(r_SM_Main[0]), .O(n18626));   // verilog/uart_rx.v(52[7] 143[14])
    defparam i21_4_lut_4_lut.LUT_INIT = 16'h2055;
    SB_LUT4 i12_3_lut_4_lut (.I0(r_SM_Main[1]), .I1(r_SM_Main[2]), .I2(n18626), 
            .I3(rx_data_ready), .O(n32269));   // verilog/uart_rx.v(52[7] 143[14])
    defparam i12_3_lut_4_lut.LUT_INIT = 16'h2f20;
    SB_LUT4 i30539_2_lut_3_lut (.I0(r_SM_Main[1]), .I1(r_SM_Main[2]), .I2(r_SM_Main[0]), 
            .I3(GND_net), .O(n32642));   // verilog/uart_rx.v(52[7] 143[14])
    defparam i30539_2_lut_3_lut.LUT_INIT = 16'hdfdf;
    SB_LUT4 i3_4_lut_adj_844 (.I0(r_SM_Main[2]), .I1(r_SM_Main[0]), .I2(r_SM_Main[1]), 
            .I3(r_SM_Main_2__N_3416[2]), .O(n17343));   // verilog/uart_rx.v(52[7] 143[14])
    defparam i3_4_lut_adj_844.LUT_INIT = 16'hefff;
    SB_LUT4 i1_2_lut_adj_845 (.I0(\r_Bit_Index[0] ), .I1(n17343), .I2(GND_net), 
            .I3(GND_net), .O(n17534));   // verilog/uart_rx.v(52[7] 143[14])
    defparam i1_2_lut_adj_845.LUT_INIT = 16'heeee;
    SB_LUT4 equal_151_i4_2_lut (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[2]), 
            .I2(GND_net), .I3(GND_net), .O(n4_adj_7));   // verilog/uart_rx.v(97[17:39])
    defparam equal_151_i4_2_lut.LUT_INIT = 16'heeee;
    
endmodule
//
// Verilog Description of module pwm
//

module pwm (n36951, VCC_net, INHA_c, clk32MHz, n17362, GND_net, 
            pwm_counter, n17360) /* synthesis syn_module_defined=1 */ ;
    input n36951;
    input VCC_net;
    output INHA_c;
    input clk32MHz;
    input n17362;
    input GND_net;
    output [31:0]pwm_counter;
    input n17360;
    
    wire clk32MHz /* synthesis SET_AS_NETWORK=clk32MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(33[6:14])
    wire [31:0]n133;
    
    wire n28597, n28596, n28595, n28594, n28593, n28592, n28591, 
        n28590, n28589, n28588, n28587, n28586, n28585, n28584, 
        n28583, n28582, n28581, n28580, n28579, n28578, n28577, 
        n28576, n28575, n28574, n28573, n28572, n28571, n28570, 
        n28569, n28568, n28567, n34838, n18, n24, n22, n26, 
        n21, pwm_counter_31__N_685;
    
    SB_DFFESR pwm_out_12 (.Q(INHA_c), .C(clk32MHz), .E(VCC_net), .D(n36951), 
            .R(n17362));   // verilog/pwm.v(16[12] 26[6])
    SB_LUT4 pwm_counter_1580_add_4_33_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[31]), 
            .I3(n28597), .O(n133[31])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1580_add_4_33_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 pwm_counter_1580_add_4_32_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[30]), 
            .I3(n28596), .O(n133[30])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1580_add_4_32_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_1580_add_4_32 (.CI(n28596), .I0(GND_net), .I1(pwm_counter[30]), 
            .CO(n28597));
    SB_LUT4 pwm_counter_1580_add_4_31_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[29]), 
            .I3(n28595), .O(n133[29])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1580_add_4_31_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_1580_add_4_31 (.CI(n28595), .I0(GND_net), .I1(pwm_counter[29]), 
            .CO(n28596));
    SB_LUT4 pwm_counter_1580_add_4_30_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[28]), 
            .I3(n28594), .O(n133[28])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1580_add_4_30_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_1580_add_4_30 (.CI(n28594), .I0(GND_net), .I1(pwm_counter[28]), 
            .CO(n28595));
    SB_LUT4 pwm_counter_1580_add_4_29_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[27]), 
            .I3(n28593), .O(n133[27])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1580_add_4_29_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_1580_add_4_29 (.CI(n28593), .I0(GND_net), .I1(pwm_counter[27]), 
            .CO(n28594));
    SB_LUT4 pwm_counter_1580_add_4_28_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[26]), 
            .I3(n28592), .O(n133[26])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1580_add_4_28_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_1580_add_4_28 (.CI(n28592), .I0(GND_net), .I1(pwm_counter[26]), 
            .CO(n28593));
    SB_LUT4 pwm_counter_1580_add_4_27_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[25]), 
            .I3(n28591), .O(n133[25])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1580_add_4_27_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_1580_add_4_27 (.CI(n28591), .I0(GND_net), .I1(pwm_counter[25]), 
            .CO(n28592));
    SB_LUT4 pwm_counter_1580_add_4_26_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[24]), 
            .I3(n28590), .O(n133[24])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1580_add_4_26_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_1580_add_4_26 (.CI(n28590), .I0(GND_net), .I1(pwm_counter[24]), 
            .CO(n28591));
    SB_LUT4 pwm_counter_1580_add_4_25_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[23]), 
            .I3(n28589), .O(n133[23])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1580_add_4_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_1580_add_4_25 (.CI(n28589), .I0(GND_net), .I1(pwm_counter[23]), 
            .CO(n28590));
    SB_LUT4 pwm_counter_1580_add_4_24_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[22]), 
            .I3(n28588), .O(n133[22])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1580_add_4_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_1580_add_4_24 (.CI(n28588), .I0(GND_net), .I1(pwm_counter[22]), 
            .CO(n28589));
    SB_LUT4 pwm_counter_1580_add_4_23_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[21]), 
            .I3(n28587), .O(n133[21])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1580_add_4_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_1580_add_4_23 (.CI(n28587), .I0(GND_net), .I1(pwm_counter[21]), 
            .CO(n28588));
    SB_LUT4 pwm_counter_1580_add_4_22_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[20]), 
            .I3(n28586), .O(n133[20])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1580_add_4_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_1580_add_4_22 (.CI(n28586), .I0(GND_net), .I1(pwm_counter[20]), 
            .CO(n28587));
    SB_LUT4 pwm_counter_1580_add_4_21_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[19]), 
            .I3(n28585), .O(n133[19])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1580_add_4_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_1580_add_4_21 (.CI(n28585), .I0(GND_net), .I1(pwm_counter[19]), 
            .CO(n28586));
    SB_LUT4 pwm_counter_1580_add_4_20_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[18]), 
            .I3(n28584), .O(n133[18])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1580_add_4_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_1580_add_4_20 (.CI(n28584), .I0(GND_net), .I1(pwm_counter[18]), 
            .CO(n28585));
    SB_LUT4 pwm_counter_1580_add_4_19_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[17]), 
            .I3(n28583), .O(n133[17])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1580_add_4_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_1580_add_4_19 (.CI(n28583), .I0(GND_net), .I1(pwm_counter[17]), 
            .CO(n28584));
    SB_LUT4 pwm_counter_1580_add_4_18_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[16]), 
            .I3(n28582), .O(n133[16])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1580_add_4_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_1580_add_4_18 (.CI(n28582), .I0(GND_net), .I1(pwm_counter[16]), 
            .CO(n28583));
    SB_LUT4 pwm_counter_1580_add_4_17_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[15]), 
            .I3(n28581), .O(n133[15])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1580_add_4_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_1580_add_4_17 (.CI(n28581), .I0(GND_net), .I1(pwm_counter[15]), 
            .CO(n28582));
    SB_LUT4 pwm_counter_1580_add_4_16_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[14]), 
            .I3(n28580), .O(n133[14])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1580_add_4_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_1580_add_4_16 (.CI(n28580), .I0(GND_net), .I1(pwm_counter[14]), 
            .CO(n28581));
    SB_LUT4 pwm_counter_1580_add_4_15_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[13]), 
            .I3(n28579), .O(n133[13])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1580_add_4_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_1580_add_4_15 (.CI(n28579), .I0(GND_net), .I1(pwm_counter[13]), 
            .CO(n28580));
    SB_LUT4 pwm_counter_1580_add_4_14_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[12]), 
            .I3(n28578), .O(n133[12])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1580_add_4_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_1580_add_4_14 (.CI(n28578), .I0(GND_net), .I1(pwm_counter[12]), 
            .CO(n28579));
    SB_LUT4 pwm_counter_1580_add_4_13_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[11]), 
            .I3(n28577), .O(n133[11])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1580_add_4_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_1580_add_4_13 (.CI(n28577), .I0(GND_net), .I1(pwm_counter[11]), 
            .CO(n28578));
    SB_LUT4 pwm_counter_1580_add_4_12_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[10]), 
            .I3(n28576), .O(n133[10])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1580_add_4_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_1580_add_4_12 (.CI(n28576), .I0(GND_net), .I1(pwm_counter[10]), 
            .CO(n28577));
    SB_LUT4 pwm_counter_1580_add_4_11_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[9]), 
            .I3(n28575), .O(n133[9])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1580_add_4_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_1580_add_4_11 (.CI(n28575), .I0(GND_net), .I1(pwm_counter[9]), 
            .CO(n28576));
    SB_LUT4 pwm_counter_1580_add_4_10_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[8]), 
            .I3(n28574), .O(n133[8])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1580_add_4_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_1580_add_4_10 (.CI(n28574), .I0(GND_net), .I1(pwm_counter[8]), 
            .CO(n28575));
    SB_LUT4 pwm_counter_1580_add_4_9_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[7]), 
            .I3(n28573), .O(n133[7])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1580_add_4_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_1580_add_4_9 (.CI(n28573), .I0(GND_net), .I1(pwm_counter[7]), 
            .CO(n28574));
    SB_LUT4 pwm_counter_1580_add_4_8_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[6]), 
            .I3(n28572), .O(n133[6])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1580_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_1580_add_4_8 (.CI(n28572), .I0(GND_net), .I1(pwm_counter[6]), 
            .CO(n28573));
    SB_LUT4 pwm_counter_1580_add_4_7_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[5]), 
            .I3(n28571), .O(n133[5])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1580_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_1580_add_4_7 (.CI(n28571), .I0(GND_net), .I1(pwm_counter[5]), 
            .CO(n28572));
    SB_LUT4 pwm_counter_1580_add_4_6_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[4]), 
            .I3(n28570), .O(n133[4])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1580_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_1580_add_4_6 (.CI(n28570), .I0(GND_net), .I1(pwm_counter[4]), 
            .CO(n28571));
    SB_LUT4 pwm_counter_1580_add_4_5_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[3]), 
            .I3(n28569), .O(n133[3])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1580_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_1580_add_4_5 (.CI(n28569), .I0(GND_net), .I1(pwm_counter[3]), 
            .CO(n28570));
    SB_LUT4 pwm_counter_1580_add_4_4_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[2]), 
            .I3(n28568), .O(n133[2])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1580_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_1580_add_4_4 (.CI(n28568), .I0(GND_net), .I1(pwm_counter[2]), 
            .CO(n28569));
    SB_LUT4 pwm_counter_1580_add_4_3_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[1]), 
            .I3(n28567), .O(n133[1])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1580_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_1580_add_4_3 (.CI(n28567), .I0(GND_net), .I1(pwm_counter[1]), 
            .CO(n28568));
    SB_LUT4 pwm_counter_1580_add_4_2_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[0]), 
            .I3(VCC_net), .O(n133[0])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1580_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_1580_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(pwm_counter[0]), 
            .CO(n28567));
    SB_LUT4 i2_3_lut (.I0(pwm_counter[6]), .I1(pwm_counter[8]), .I2(pwm_counter[7]), 
            .I3(GND_net), .O(n34838));
    defparam i2_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i4_4_lut (.I0(n34838), .I1(pwm_counter[13]), .I2(pwm_counter[10]), 
            .I3(pwm_counter[9]), .O(n18));
    defparam i4_4_lut.LUT_INIT = 16'heccc;
    SB_LUT4 i10_4_lut (.I0(pwm_counter[17]), .I1(pwm_counter[22]), .I2(pwm_counter[14]), 
            .I3(pwm_counter[18]), .O(n24));
    defparam i10_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i8_4_lut (.I0(pwm_counter[21]), .I1(n17360), .I2(pwm_counter[16]), 
            .I3(pwm_counter[12]), .O(n22));
    defparam i8_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i12_4_lut (.I0(pwm_counter[15]), .I1(n24), .I2(n18), .I3(pwm_counter[19]), 
            .O(n26));
    defparam i12_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i7_2_lut (.I0(pwm_counter[11]), .I1(pwm_counter[20]), .I2(GND_net), 
            .I3(GND_net), .O(n21));
    defparam i7_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i18782_4_lut (.I0(n21), .I1(pwm_counter[31]), .I2(n26), .I3(n22), 
            .O(pwm_counter_31__N_685));   // verilog/pwm.v(18[8:40])
    defparam i18782_4_lut.LUT_INIT = 16'h3332;
    SB_DFFSR pwm_counter_1580__i0 (.Q(pwm_counter[0]), .C(clk32MHz), .D(n133[0]), 
            .R(pwm_counter_31__N_685));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_1580__i1 (.Q(pwm_counter[1]), .C(clk32MHz), .D(n133[1]), 
            .R(pwm_counter_31__N_685));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_1580__i2 (.Q(pwm_counter[2]), .C(clk32MHz), .D(n133[2]), 
            .R(pwm_counter_31__N_685));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_1580__i3 (.Q(pwm_counter[3]), .C(clk32MHz), .D(n133[3]), 
            .R(pwm_counter_31__N_685));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_1580__i4 (.Q(pwm_counter[4]), .C(clk32MHz), .D(n133[4]), 
            .R(pwm_counter_31__N_685));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_1580__i5 (.Q(pwm_counter[5]), .C(clk32MHz), .D(n133[5]), 
            .R(pwm_counter_31__N_685));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_1580__i6 (.Q(pwm_counter[6]), .C(clk32MHz), .D(n133[6]), 
            .R(pwm_counter_31__N_685));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_1580__i7 (.Q(pwm_counter[7]), .C(clk32MHz), .D(n133[7]), 
            .R(pwm_counter_31__N_685));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_1580__i8 (.Q(pwm_counter[8]), .C(clk32MHz), .D(n133[8]), 
            .R(pwm_counter_31__N_685));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_1580__i9 (.Q(pwm_counter[9]), .C(clk32MHz), .D(n133[9]), 
            .R(pwm_counter_31__N_685));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_1580__i10 (.Q(pwm_counter[10]), .C(clk32MHz), .D(n133[10]), 
            .R(pwm_counter_31__N_685));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_1580__i11 (.Q(pwm_counter[11]), .C(clk32MHz), .D(n133[11]), 
            .R(pwm_counter_31__N_685));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_1580__i12 (.Q(pwm_counter[12]), .C(clk32MHz), .D(n133[12]), 
            .R(pwm_counter_31__N_685));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_1580__i13 (.Q(pwm_counter[13]), .C(clk32MHz), .D(n133[13]), 
            .R(pwm_counter_31__N_685));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_1580__i14 (.Q(pwm_counter[14]), .C(clk32MHz), .D(n133[14]), 
            .R(pwm_counter_31__N_685));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_1580__i15 (.Q(pwm_counter[15]), .C(clk32MHz), .D(n133[15]), 
            .R(pwm_counter_31__N_685));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_1580__i16 (.Q(pwm_counter[16]), .C(clk32MHz), .D(n133[16]), 
            .R(pwm_counter_31__N_685));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_1580__i17 (.Q(pwm_counter[17]), .C(clk32MHz), .D(n133[17]), 
            .R(pwm_counter_31__N_685));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_1580__i18 (.Q(pwm_counter[18]), .C(clk32MHz), .D(n133[18]), 
            .R(pwm_counter_31__N_685));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_1580__i19 (.Q(pwm_counter[19]), .C(clk32MHz), .D(n133[19]), 
            .R(pwm_counter_31__N_685));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_1580__i20 (.Q(pwm_counter[20]), .C(clk32MHz), .D(n133[20]), 
            .R(pwm_counter_31__N_685));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_1580__i21 (.Q(pwm_counter[21]), .C(clk32MHz), .D(n133[21]), 
            .R(pwm_counter_31__N_685));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_1580__i22 (.Q(pwm_counter[22]), .C(clk32MHz), .D(n133[22]), 
            .R(pwm_counter_31__N_685));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_1580__i23 (.Q(pwm_counter[23]), .C(clk32MHz), .D(n133[23]), 
            .R(pwm_counter_31__N_685));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_1580__i24 (.Q(pwm_counter[24]), .C(clk32MHz), .D(n133[24]), 
            .R(pwm_counter_31__N_685));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_1580__i25 (.Q(pwm_counter[25]), .C(clk32MHz), .D(n133[25]), 
            .R(pwm_counter_31__N_685));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_1580__i26 (.Q(pwm_counter[26]), .C(clk32MHz), .D(n133[26]), 
            .R(pwm_counter_31__N_685));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_1580__i27 (.Q(pwm_counter[27]), .C(clk32MHz), .D(n133[27]), 
            .R(pwm_counter_31__N_685));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_1580__i28 (.Q(pwm_counter[28]), .C(clk32MHz), .D(n133[28]), 
            .R(pwm_counter_31__N_685));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_1580__i29 (.Q(pwm_counter[29]), .C(clk32MHz), .D(n133[29]), 
            .R(pwm_counter_31__N_685));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_1580__i30 (.Q(pwm_counter[30]), .C(clk32MHz), .D(n133[30]), 
            .R(pwm_counter_31__N_685));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_1580__i31 (.Q(pwm_counter[31]), .C(clk32MHz), .D(n133[31]), 
            .R(pwm_counter_31__N_685));   // verilog/pwm.v(17[20:33])
    
endmodule
//
// Verilog Description of module EEPROM
//

module EEPROM (CLK_c, n3646, \state[1] , enable_slow_N_4001, GND_net, 
            read, \state[0] , \state[2] , n7, n19051, rw, n32425, 
            data_ready, n24036, n33471, n33535, n32331, n32323, 
            \state[3] , n6, n5212, \state_7__N_3914[3] , \saved_addr[0] , 
            \state[0]_adj_3 , \state_7__N_3898[0] , n10, scl_enable, 
            VCC_net, sda_enable, n23736, n10_adj_4, n5690, n19061, 
            data, n19060, n19056, n19055, n19054, n19592, n19584, 
            n19582, n19558, n8, scl, sda_out, n36289, n4, n23836, 
            n17518, n4_adj_5, n17513) /* synthesis syn_noprune=1, syn_module_defined=1 */ ;
    input CLK_c;
    output [0:0]n3646;
    output \state[1] ;
    output enable_slow_N_4001;
    input GND_net;
    input read;
    output \state[0] ;
    output \state[2] ;
    output n7;
    input n19051;
    output rw;
    input n32425;
    output data_ready;
    output n24036;
    input n33471;
    output n33535;
    input n32331;
    input n32323;
    output \state[3] ;
    output n6;
    output n5212;
    input \state_7__N_3914[3] ;
    output \saved_addr[0] ;
    output \state[0]_adj_3 ;
    output \state_7__N_3898[0] ;
    output n10;
    output scl_enable;
    input VCC_net;
    output sda_enable;
    output n23736;
    input n10_adj_4;
    input n5690;
    input n19061;
    output [7:0]data;
    input n19060;
    input n19056;
    input n19055;
    input n19054;
    input n19592;
    input n19584;
    input n19582;
    input n19558;
    input n8;
    output scl;
    output sda_out;
    output n36289;
    output n4;
    output n23836;
    output n17518;
    output n4_adj_5;
    output n17513;
    
    wire CLK_c /* synthesis SET_AS_NETWORK=CLK_c, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(3[9:12])
    wire [15:0]delay_counter_15__N_3800;
    
    wire n18717;
    wire [15:0]delay_counter;   // verilog/eeprom.v(24[12:25])
    
    wire n18923, enable, n17332;
    wire [15:0]n3338;
    
    wire n28, n26, n27, n25;
    wire [7:0]state;   // verilog/i2c_controller.v(33[12:17])
    
    wire n27897, n27896, n27895, n27894, n27893, n27892, n27891, 
        n27890, n27889, n27888, n27887, n27886, n27885, n27884, 
        n27883;
    
    SB_DFFESR delay_counter_i0_i15 (.Q(delay_counter[15]), .C(CLK_c), .E(n18717), 
            .D(delay_counter_15__N_3800[15]), .R(n18923));   // verilog/eeprom.v(26[8] 58[4])
    SB_DFFESR delay_counter_i0_i14 (.Q(delay_counter[14]), .C(CLK_c), .E(n18717), 
            .D(delay_counter_15__N_3800[14]), .R(n18923));   // verilog/eeprom.v(26[8] 58[4])
    SB_DFFESR delay_counter_i0_i13 (.Q(delay_counter[13]), .C(CLK_c), .E(n18717), 
            .D(delay_counter_15__N_3800[13]), .R(n18923));   // verilog/eeprom.v(26[8] 58[4])
    SB_DFFESR delay_counter_i0_i12 (.Q(delay_counter[12]), .C(CLK_c), .E(n18717), 
            .D(delay_counter_15__N_3800[12]), .R(n18923));   // verilog/eeprom.v(26[8] 58[4])
    SB_DFFESR delay_counter_i0_i11 (.Q(delay_counter[11]), .C(CLK_c), .E(n18717), 
            .D(delay_counter_15__N_3800[11]), .R(n18923));   // verilog/eeprom.v(26[8] 58[4])
    SB_DFFESS delay_counter_i0_i10 (.Q(delay_counter[10]), .C(CLK_c), .E(n18717), 
            .D(delay_counter_15__N_3800[10]), .S(n18923));   // verilog/eeprom.v(26[8] 58[4])
    SB_DFFESS delay_counter_i0_i9 (.Q(delay_counter[9]), .C(CLK_c), .E(n18717), 
            .D(delay_counter_15__N_3800[9]), .S(n18923));   // verilog/eeprom.v(26[8] 58[4])
    SB_DFFESS delay_counter_i0_i8 (.Q(delay_counter[8]), .C(CLK_c), .E(n18717), 
            .D(delay_counter_15__N_3800[8]), .S(n18923));   // verilog/eeprom.v(26[8] 58[4])
    SB_DFFESS delay_counter_i0_i7 (.Q(delay_counter[7]), .C(CLK_c), .E(n18717), 
            .D(delay_counter_15__N_3800[7]), .S(n18923));   // verilog/eeprom.v(26[8] 58[4])
    SB_DFFESS delay_counter_i0_i6 (.Q(delay_counter[6]), .C(CLK_c), .E(n18717), 
            .D(delay_counter_15__N_3800[6]), .S(n18923));   // verilog/eeprom.v(26[8] 58[4])
    SB_DFFESR delay_counter_i0_i5 (.Q(delay_counter[5]), .C(CLK_c), .E(n18717), 
            .D(delay_counter_15__N_3800[5]), .R(n18923));   // verilog/eeprom.v(26[8] 58[4])
    SB_DFFESS delay_counter_i0_i4 (.Q(delay_counter[4]), .C(CLK_c), .E(n18717), 
            .D(delay_counter_15__N_3800[4]), .S(n18923));   // verilog/eeprom.v(26[8] 58[4])
    SB_DFFESR delay_counter_i0_i3 (.Q(delay_counter[3]), .C(CLK_c), .E(n18717), 
            .D(delay_counter_15__N_3800[3]), .R(n18923));   // verilog/eeprom.v(26[8] 58[4])
    SB_DFFESR delay_counter_i0_i2 (.Q(delay_counter[2]), .C(CLK_c), .E(n18717), 
            .D(delay_counter_15__N_3800[2]), .R(n18923));   // verilog/eeprom.v(26[8] 58[4])
    SB_DFFESR delay_counter_i0_i1 (.Q(delay_counter[1]), .C(CLK_c), .E(n18717), 
            .D(delay_counter_15__N_3800[1]), .R(n18923));   // verilog/eeprom.v(26[8] 58[4])
    SB_DFFSR enable_39 (.Q(enable), .C(CLK_c), .D(n3646[0]), .R(\state[1] ));   // verilog/eeprom.v(26[8] 58[4])
    SB_LUT4 i30413_2_lut (.I0(n17332), .I1(enable_slow_N_4001), .I2(GND_net), 
            .I3(GND_net), .O(n3338[14]));   // verilog/eeprom.v(46[18] 48[12])
    defparam i30413_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i12_4_lut (.I0(delay_counter[6]), .I1(delay_counter[10]), .I2(delay_counter[12]), 
            .I3(delay_counter[8]), .O(n28));   // verilog/eeprom.v(42[12:28])
    defparam i12_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i10_4_lut (.I0(delay_counter[11]), .I1(delay_counter[2]), .I2(delay_counter[7]), 
            .I3(delay_counter[5]), .O(n26));   // verilog/eeprom.v(42[12:28])
    defparam i10_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i11_4_lut (.I0(delay_counter[15]), .I1(delay_counter[3]), .I2(delay_counter[14]), 
            .I3(delay_counter[1]), .O(n27));   // verilog/eeprom.v(42[12:28])
    defparam i11_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i9_4_lut (.I0(delay_counter[4]), .I1(delay_counter[9]), .I2(delay_counter[13]), 
            .I3(delay_counter[0]), .O(n25));   // verilog/eeprom.v(42[12:28])
    defparam i9_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i15_4_lut (.I0(n25), .I1(n27), .I2(n26), .I3(n28), .O(n17332));   // verilog/eeprom.v(42[12:28])
    defparam i15_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 mux_937_Mux_0_i1_4_lut (.I0(read), .I1(n17332), .I2(\state[0] ), 
            .I3(enable_slow_N_4001), .O(n3646[0]));   // verilog/eeprom.v(29[3] 57[10])
    defparam mux_937_Mux_0_i1_4_lut.LUT_INIT = 16'h0a3a;
    SB_LUT4 i2_2_lut (.I0(state[1]), .I1(\state[2] ), .I2(GND_net), .I3(GND_net), 
            .O(n7));   // verilog/eeprom.v(42[12:28])
    defparam i2_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i13794_2_lut (.I0(n18717), .I1(\state[0] ), .I2(GND_net), 
            .I3(GND_net), .O(n18923));   // verilog/eeprom.v(26[8] 58[4])
    defparam i13794_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i1_3_lut (.I0(read), .I1(\state[1] ), .I2(\state[0] ), .I3(GND_net), 
            .O(n18717));
    defparam i1_3_lut.LUT_INIT = 16'h3232;
    SB_LUT4 add_755_17_lut (.I0(GND_net), .I1(delay_counter[15]), .I2(n3338[14]), 
            .I3(n27897), .O(delay_counter_15__N_3800[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_755_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_755_16_lut (.I0(GND_net), .I1(delay_counter[14]), .I2(n3338[14]), 
            .I3(n27896), .O(delay_counter_15__N_3800[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_755_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_755_16 (.CI(n27896), .I0(delay_counter[14]), .I1(n3338[14]), 
            .CO(n27897));
    SB_LUT4 add_755_15_lut (.I0(GND_net), .I1(delay_counter[13]), .I2(n3338[14]), 
            .I3(n27895), .O(delay_counter_15__N_3800[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_755_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_755_15 (.CI(n27895), .I0(delay_counter[13]), .I1(n3338[14]), 
            .CO(n27896));
    SB_LUT4 add_755_14_lut (.I0(GND_net), .I1(delay_counter[12]), .I2(n3338[14]), 
            .I3(n27894), .O(delay_counter_15__N_3800[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_755_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_755_14 (.CI(n27894), .I0(delay_counter[12]), .I1(n3338[14]), 
            .CO(n27895));
    SB_LUT4 add_755_13_lut (.I0(GND_net), .I1(delay_counter[11]), .I2(n3338[14]), 
            .I3(n27893), .O(delay_counter_15__N_3800[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_755_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_755_13 (.CI(n27893), .I0(delay_counter[11]), .I1(n3338[14]), 
            .CO(n27894));
    SB_LUT4 add_755_12_lut (.I0(GND_net), .I1(delay_counter[10]), .I2(n3338[14]), 
            .I3(n27892), .O(delay_counter_15__N_3800[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_755_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_755_12 (.CI(n27892), .I0(delay_counter[10]), .I1(n3338[14]), 
            .CO(n27893));
    SB_LUT4 add_755_11_lut (.I0(GND_net), .I1(delay_counter[9]), .I2(n3338[14]), 
            .I3(n27891), .O(delay_counter_15__N_3800[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_755_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_755_11 (.CI(n27891), .I0(delay_counter[9]), .I1(n3338[14]), 
            .CO(n27892));
    SB_LUT4 add_755_10_lut (.I0(GND_net), .I1(delay_counter[8]), .I2(n3338[14]), 
            .I3(n27890), .O(delay_counter_15__N_3800[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_755_10_lut.LUT_INIT = 16'hC33C;
    SB_DFFESR delay_counter_i0_i0 (.Q(delay_counter[0]), .C(CLK_c), .E(n18717), 
            .D(delay_counter_15__N_3800[0]), .R(n18923));   // verilog/eeprom.v(26[8] 58[4])
    SB_CARRY add_755_10 (.CI(n27890), .I0(delay_counter[8]), .I1(n3338[14]), 
            .CO(n27891));
    SB_LUT4 add_755_9_lut (.I0(GND_net), .I1(delay_counter[7]), .I2(n3338[14]), 
            .I3(n27889), .O(delay_counter_15__N_3800[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_755_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_755_9 (.CI(n27889), .I0(delay_counter[7]), .I1(n3338[14]), 
            .CO(n27890));
    SB_LUT4 add_755_8_lut (.I0(GND_net), .I1(delay_counter[6]), .I2(n3338[14]), 
            .I3(n27888), .O(delay_counter_15__N_3800[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_755_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_755_8 (.CI(n27888), .I0(delay_counter[6]), .I1(n3338[14]), 
            .CO(n27889));
    SB_LUT4 add_755_7_lut (.I0(GND_net), .I1(delay_counter[5]), .I2(n3338[14]), 
            .I3(n27887), .O(delay_counter_15__N_3800[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_755_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_755_7 (.CI(n27887), .I0(delay_counter[5]), .I1(n3338[14]), 
            .CO(n27888));
    SB_LUT4 add_755_6_lut (.I0(GND_net), .I1(delay_counter[4]), .I2(n3338[14]), 
            .I3(n27886), .O(delay_counter_15__N_3800[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_755_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_755_6 (.CI(n27886), .I0(delay_counter[4]), .I1(n3338[14]), 
            .CO(n27887));
    SB_LUT4 add_755_5_lut (.I0(GND_net), .I1(delay_counter[3]), .I2(n3338[14]), 
            .I3(n27885), .O(delay_counter_15__N_3800[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_755_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_755_5 (.CI(n27885), .I0(delay_counter[3]), .I1(n3338[14]), 
            .CO(n27886));
    SB_DFF rw_43 (.Q(rw), .C(CLK_c), .D(n19051));   // verilog/eeprom.v(26[8] 58[4])
    SB_DFF data_ready_42 (.Q(data_ready), .C(CLK_c), .D(n32425));   // verilog/eeprom.v(26[8] 58[4])
    SB_LUT4 add_755_4_lut (.I0(GND_net), .I1(delay_counter[2]), .I2(n3338[14]), 
            .I3(n27884), .O(delay_counter_15__N_3800[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_755_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_755_4 (.CI(n27884), .I0(delay_counter[2]), .I1(n3338[14]), 
            .CO(n27885));
    SB_LUT4 i18903_2_lut_3_lut (.I0(\state[0] ), .I1(\state[1] ), .I2(enable_slow_N_4001), 
            .I3(GND_net), .O(n24036));   // verilog/eeprom.v(51[5:9])
    defparam i18903_2_lut_3_lut.LUT_INIT = 16'hfbfb;
    SB_LUT4 i26785_4_lut_4_lut (.I0(\state[0] ), .I1(\state[1] ), .I2(n33471), 
            .I3(enable_slow_N_4001), .O(n33535));   // verilog/eeprom.v(51[5:9])
    defparam i26785_4_lut_4_lut.LUT_INIT = 16'hfcf8;
    SB_LUT4 add_755_3_lut (.I0(GND_net), .I1(delay_counter[1]), .I2(n3338[14]), 
            .I3(n27883), .O(delay_counter_15__N_3800[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_755_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_755_3 (.CI(n27883), .I0(delay_counter[1]), .I1(n3338[14]), 
            .CO(n27884));
    SB_DFF state__i1 (.Q(\state[1] ), .C(CLK_c), .D(n32331));   // verilog/eeprom.v(26[8] 58[4])
    SB_DFF state__i0 (.Q(\state[0] ), .C(CLK_c), .D(n32323));   // verilog/eeprom.v(26[8] 58[4])
    SB_LUT4 add_755_2_lut (.I0(GND_net), .I1(delay_counter[0]), .I2(n3338[14]), 
            .I3(GND_net), .O(delay_counter_15__N_3800[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_755_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_755_2 (.CI(GND_net), .I0(delay_counter[0]), .I1(n3338[14]), 
            .CO(n27883));
    SB_LUT4 i2_2_lut_adj_840 (.I0(\state[3] ), .I1(n17332), .I2(GND_net), 
            .I3(GND_net), .O(n6));   // verilog/eeprom.v(42[12:28])
    defparam i2_2_lut_adj_840.LUT_INIT = 16'heeee;
    i2c_controller i2c (.n5212(n5212), .\state[3] (\state[3] ), .\state[2] (\state[2] ), 
            .\state[1] (state[1]), .GND_net(GND_net), .CLK_c(CLK_c), .\state_7__N_3914[3] (\state_7__N_3914[3] ), 
            .\saved_addr[0] (\saved_addr[0] ), .\state[0] (\state[0]_adj_3 ), 
            .\state_7__N_3898[0] (\state_7__N_3898[0] ), .enable_slow_N_4001(enable_slow_N_4001), 
            .n10(n10), .scl_enable(scl_enable), .VCC_net(VCC_net), .sda_enable(sda_enable), 
            .n23736(n23736), .n10_adj_1(n10_adj_4), .enable(enable), .n5690(n5690), 
            .n19061(n19061), .data({data}), .n19060(n19060), .n19056(n19056), 
            .n19055(n19055), .n19054(n19054), .n19592(n19592), .n19584(n19584), 
            .n19582(n19582), .n19558(n19558), .n8(n8), .scl(scl), .sda_out(sda_out), 
            .n36289(n36289), .n4(n4), .n23836(n23836), .n17518(n17518), 
            .n4_adj_2(n4_adj_5), .n17513(n17513)) /* synthesis syn_noprune=1, syn_module_defined=1 */ ;   // verilog/eeprom.v(60[16] 74[4])
    
endmodule
//
// Verilog Description of module i2c_controller
//

module i2c_controller (n5212, \state[3] , \state[2] , \state[1] , GND_net, 
            CLK_c, \state_7__N_3914[3] , \saved_addr[0] , \state[0] , 
            \state_7__N_3898[0] , enable_slow_N_4001, n10, scl_enable, 
            VCC_net, sda_enable, n23736, n10_adj_1, enable, n5690, 
            n19061, data, n19060, n19056, n19055, n19054, n19592, 
            n19584, n19582, n19558, n8, scl, sda_out, n36289, 
            n4, n23836, n17518, n4_adj_2, n17513) /* synthesis syn_noprune=1, syn_module_defined=1 */ ;
    output n5212;
    output \state[3] ;
    output \state[2] ;
    output \state[1] ;
    input GND_net;
    input CLK_c;
    input \state_7__N_3914[3] ;
    output \saved_addr[0] ;
    output \state[0] ;
    output \state_7__N_3898[0] ;
    output enable_slow_N_4001;
    output n10;
    output scl_enable;
    input VCC_net;
    output sda_enable;
    output n23736;
    input n10_adj_1;
    input enable;
    input n5690;
    input n19061;
    output [7:0]data;
    input n19060;
    input n19056;
    input n19055;
    input n19054;
    input n19592;
    input n19584;
    input n19582;
    input n19558;
    input n8;
    output scl;
    output sda_out;
    output n36289;
    output n4;
    output n23836;
    output n17518;
    output n4_adj_2;
    output n17513;
    
    wire i2c_clk /* synthesis is_clock=1, SET_AS_NETWORK=\eeprom/i2c/i2c_clk */ ;   // verilog/i2c_controller.v(41[6:13])
    wire CLK_c /* synthesis SET_AS_NETWORK=CLK_c, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(3[9:12])
    
    wire n32481, n34096, n24009, n24285, n5, n24595, n15, n11;
    wire [5:0]n29;
    wire [7:0]counter2;   // verilog/i2c_controller.v(37[12:20])
    
    wire n18921;
    wire [7:0]n119;
    
    wire n18768;
    wire [7:0]counter;   // verilog/i2c_controller.v(36[12:19])
    
    wire n19001, n11_adj_4002, n36282, n36214, n11_adj_4003, n36320, 
        n33, n37, n18884, n34, n39, n7, i2c_clk_N_3987, enable_slow_N_4000, 
        n18648, scl_enable_N_3988, n12, n28629, n28628, n28627, 
        n28626, n28625, n10595, n5574, n32365, sda_out_adj_4006, 
        n5205, n28112, n28111, n28110, n28109, n28108, n28107, 
        n28106, n10_adj_4007, n18565, n11_adj_4008, n36307, n15_adj_4010, 
        n33475, n10_adj_4011, n11_adj_4012;
    
    SB_DFFESS state_i0_i3 (.Q(\state[3] ), .C(i2c_clk), .E(n5212), .D(n32481), 
            .S(n34096));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFFESS state_i0_i2 (.Q(\state[2] ), .C(i2c_clk), .E(n5212), .D(n24009), 
            .S(n24285));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFFESS state_i0_i1 (.Q(\state[1] ), .C(i2c_clk), .E(n5212), .D(n5), 
            .S(n24595));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_LUT4 i30563_3_lut (.I0(n5212), .I1(n15), .I2(n11), .I3(GND_net), 
            .O(n24285));
    defparam i30563_3_lut.LUT_INIT = 16'h2a2a;
    SB_DFFSR counter2_1587_1588__i1 (.Q(counter2[0]), .C(CLK_c), .D(n29[0]), 
            .R(n18921));   // verilog/i2c_controller.v(69[20:35])
    SB_DFFESR counter_i7 (.Q(counter[7]), .C(i2c_clk), .E(n18768), .D(n119[7]), 
            .R(n19001));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFFESR counter_i6 (.Q(counter[6]), .C(i2c_clk), .E(n18768), .D(n119[6]), 
            .R(n19001));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFFESR counter_i5 (.Q(counter[5]), .C(i2c_clk), .E(n18768), .D(n119[5]), 
            .R(n19001));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_LUT4 i30501_2_lut (.I0(\state_7__N_3914[3] ), .I1(n11_adj_4002), 
            .I2(GND_net), .I3(GND_net), .O(n24009));
    defparam i30501_2_lut.LUT_INIT = 16'h1111;
    SB_DFFESR counter_i4 (.Q(counter[4]), .C(i2c_clk), .E(n18768), .D(n119[4]), 
            .R(n19001));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFFESR counter_i3 (.Q(counter[3]), .C(i2c_clk), .E(n18768), .D(n119[3]), 
            .R(n19001));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFFESS counter_i2 (.Q(counter[2]), .C(i2c_clk), .E(n18768), .D(n119[2]), 
            .S(n19001));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFFESS counter_i1 (.Q(counter[1]), .C(i2c_clk), .E(n18768), .D(n119[1]), 
            .S(n19001));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_LUT4 i29842_2_lut (.I0(counter[1]), .I1(\saved_addr[0] ), .I2(GND_net), 
            .I3(GND_net), .O(n36282));   // verilog/i2c_controller.v(198[28:35])
    defparam i29842_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i29833_4_lut (.I0(n36282), .I1(\state[1] ), .I2(counter[0]), 
            .I3(counter[2]), .O(n36214));   // verilog/i2c_controller.v(181[4] 214[11])
    defparam i29833_4_lut.LUT_INIT = 16'hc008;
    SB_LUT4 i29850_4_lut (.I0(n36214), .I1(\state[2] ), .I2(\state[0] ), 
            .I3(n11_adj_4003), .O(n36320));   // verilog/i2c_controller.v(181[4] 214[11])
    defparam i29850_4_lut.LUT_INIT = 16'h0322;
    SB_LUT4 i1_3_lut (.I0(\state[1] ), .I1(n33), .I2(n37), .I3(GND_net), 
            .O(n18884));
    defparam i1_3_lut.LUT_INIT = 16'h5454;
    SB_LUT4 i1_2_lut (.I0(n34), .I1(n37), .I2(GND_net), .I3(GND_net), 
            .O(n39));
    defparam i1_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i1_2_lut_adj_835 (.I0(\state[2] ), .I1(\state[3] ), .I2(GND_net), 
            .I3(GND_net), .O(n7));
    defparam i1_2_lut_adj_835.LUT_INIT = 16'h4444;
    SB_LUT4 i1_2_lut_adj_836 (.I0(i2c_clk), .I1(n18921), .I2(GND_net), 
            .I3(GND_net), .O(i2c_clk_N_3987));
    defparam i1_2_lut_adj_836.LUT_INIT = 16'h6666;
    SB_LUT4 i30386_2_lut (.I0(\state_7__N_3898[0] ), .I1(enable_slow_N_4001), 
            .I2(GND_net), .I3(GND_net), .O(enable_slow_N_4000));   // verilog/i2c_controller.v(62[6:32])
    defparam i30386_2_lut.LUT_INIT = 16'h7777;
    SB_LUT4 i2_2_lut (.I0(counter[2]), .I1(counter[1]), .I2(GND_net), 
            .I3(GND_net), .O(n10));   // verilog/i2c_controller.v(110[10:22])
    defparam i2_2_lut.LUT_INIT = 16'heeee;
    SB_DFFE enable_slow_120 (.Q(\state_7__N_3898[0] ), .C(CLK_c), .E(n18648), 
            .D(enable_slow_N_4000));   // verilog/i2c_controller.v(58[9] 71[5])
    SB_DFF i2c_clk_121 (.Q(i2c_clk), .C(CLK_c), .D(i2c_clk_N_3987));   // verilog/i2c_controller.v(58[9] 71[5])
    SB_DFFN i2c_scl_enable_123 (.Q(scl_enable), .C(i2c_clk), .D(scl_enable_N_3988));   // verilog/i2c_controller.v(76[12] 82[6])
    SB_LUT4 i5_4_lut (.I0(counter[0]), .I1(counter[3]), .I2(counter[6]), 
            .I3(counter[5]), .O(n12));   // verilog/i2c_controller.v(110[10:22])
    defparam i5_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 counter2_1587_1588_add_4_7_lut (.I0(GND_net), .I1(GND_net), 
            .I2(counter2[5]), .I3(n28629), .O(n29[5])) /* synthesis syn_instantiated=1 */ ;
    defparam counter2_1587_1588_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 counter2_1587_1588_add_4_6_lut (.I0(GND_net), .I1(GND_net), 
            .I2(counter2[4]), .I3(n28628), .O(n29[4])) /* synthesis syn_instantiated=1 */ ;
    defparam counter2_1587_1588_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter2_1587_1588_add_4_6 (.CI(n28628), .I0(GND_net), .I1(counter2[4]), 
            .CO(n28629));
    SB_LUT4 counter2_1587_1588_add_4_5_lut (.I0(GND_net), .I1(GND_net), 
            .I2(counter2[3]), .I3(n28627), .O(n29[3])) /* synthesis syn_instantiated=1 */ ;
    defparam counter2_1587_1588_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter2_1587_1588_add_4_5 (.CI(n28627), .I0(GND_net), .I1(counter2[3]), 
            .CO(n28628));
    SB_LUT4 counter2_1587_1588_add_4_4_lut (.I0(GND_net), .I1(GND_net), 
            .I2(counter2[2]), .I3(n28626), .O(n29[2])) /* synthesis syn_instantiated=1 */ ;
    defparam counter2_1587_1588_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter2_1587_1588_add_4_4 (.CI(n28626), .I0(GND_net), .I1(counter2[2]), 
            .CO(n28627));
    SB_LUT4 counter2_1587_1588_add_4_3_lut (.I0(GND_net), .I1(GND_net), 
            .I2(counter2[1]), .I3(n28625), .O(n29[1])) /* synthesis syn_instantiated=1 */ ;
    defparam counter2_1587_1588_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter2_1587_1588_add_4_3 (.CI(n28625), .I0(GND_net), .I1(counter2[1]), 
            .CO(n28626));
    SB_LUT4 counter2_1587_1588_add_4_2_lut (.I0(GND_net), .I1(GND_net), 
            .I2(counter2[0]), .I3(VCC_net), .O(n29[0])) /* synthesis syn_instantiated=1 */ ;
    defparam counter2_1587_1588_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter2_1587_1588_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(counter2[0]), 
            .CO(n28625));
    SB_DFFNESS write_enable_131 (.Q(sda_enable), .C(i2c_clk), .E(n5574), 
            .D(n10595), .S(n18884));   // verilog/i2c_controller.v(180[12] 215[6])
    SB_DFFNE sda_out_132 (.Q(sda_out_adj_4006), .C(i2c_clk), .E(n32365), 
            .D(n36320));   // verilog/i2c_controller.v(180[12] 215[6])
    SB_DFFESS counter_i0 (.Q(counter[0]), .C(i2c_clk), .E(n18768), .D(n119[0]), 
            .S(n19001));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_LUT4 i6_4_lut (.I0(counter[4]), .I1(n12), .I2(counter[7]), .I3(n10), 
            .O(n5205));   // verilog/i2c_controller.v(110[10:22])
    defparam i6_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 sub_39_add_2_9_lut (.I0(GND_net), .I1(counter[7]), .I2(VCC_net), 
            .I3(n28112), .O(n119[7])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_39_add_2_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_39_add_2_8_lut (.I0(GND_net), .I1(counter[6]), .I2(VCC_net), 
            .I3(n28111), .O(n119[6])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_39_add_2_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_39_add_2_8 (.CI(n28111), .I0(counter[6]), .I1(VCC_net), 
            .CO(n28112));
    SB_LUT4 sub_39_add_2_7_lut (.I0(GND_net), .I1(counter[5]), .I2(VCC_net), 
            .I3(n28110), .O(n119[5])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_39_add_2_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_39_add_2_7 (.CI(n28110), .I0(counter[5]), .I1(VCC_net), 
            .CO(n28111));
    SB_LUT4 sub_39_add_2_6_lut (.I0(GND_net), .I1(counter[4]), .I2(VCC_net), 
            .I3(n28109), .O(n119[4])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_39_add_2_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_39_add_2_6 (.CI(n28109), .I0(counter[4]), .I1(VCC_net), 
            .CO(n28110));
    SB_LUT4 sub_39_add_2_5_lut (.I0(GND_net), .I1(counter[3]), .I2(VCC_net), 
            .I3(n28108), .O(n119[3])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_39_add_2_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_39_add_2_5 (.CI(n28108), .I0(counter[3]), .I1(VCC_net), 
            .CO(n28109));
    SB_LUT4 sub_39_add_2_4_lut (.I0(GND_net), .I1(counter[2]), .I2(VCC_net), 
            .I3(n28107), .O(n119[2])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_39_add_2_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_39_add_2_4 (.CI(n28107), .I0(counter[2]), .I1(VCC_net), 
            .CO(n28108));
    SB_LUT4 sub_39_add_2_3_lut (.I0(GND_net), .I1(counter[1]), .I2(VCC_net), 
            .I3(n28106), .O(n119[1])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_39_add_2_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_39_add_2_3 (.CI(n28106), .I0(counter[1]), .I1(VCC_net), 
            .CO(n28107));
    SB_LUT4 sub_39_add_2_2_lut (.I0(GND_net), .I1(counter[0]), .I2(GND_net), 
            .I3(VCC_net), .O(n119[0])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_39_add_2_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_39_add_2_2 (.CI(VCC_net), .I0(counter[0]), .I1(GND_net), 
            .CO(n28106));
    SB_LUT4 i30420_4_lut_4_lut (.I0(\state[2] ), .I1(n11_adj_4003), .I2(\state[1] ), 
            .I3(n39), .O(n5574));
    defparam i30420_4_lut_4_lut.LUT_INIT = 16'hef00;
    SB_LUT4 i30449_2_lut_3_lut (.I0(\state[2] ), .I1(n11_adj_4003), .I2(\state[0] ), 
            .I3(GND_net), .O(n10595));
    defparam i30449_2_lut_3_lut.LUT_INIT = 16'h0404;
    SB_LUT4 state_7__I_0_143_i10_2_lut (.I0(\state[2] ), .I1(\state[3] ), 
            .I2(GND_net), .I3(GND_net), .O(n10_adj_4007));   // verilog/i2c_controller.v(151[5:14])
    defparam state_7__I_0_143_i10_2_lut.LUT_INIT = 16'hdddd;
    SB_LUT4 i30399_4_lut (.I0(n18565), .I1(n5205), .I2(n11_adj_4008), 
            .I3(n23736), .O(n5212));
    defparam i30399_4_lut.LUT_INIT = 16'h5111;
    SB_LUT4 i29773_4_lut (.I0(n10_adj_1), .I1(n10_adj_4007), .I2(\state_7__N_3914[3] ), 
            .I3(enable), .O(n36307));   // verilog/i2c_controller.v(92[4] 172[11])
    defparam i29773_4_lut.LUT_INIT = 16'h7073;
    SB_LUT4 i1_4_lut (.I0(\state[1] ), .I1(n7), .I2(n36307), .I3(\state[0] ), 
            .O(n32481));   // verilog/i2c_controller.v(92[4] 172[11])
    defparam i1_4_lut.LUT_INIT = 16'ha088;
    SB_LUT4 state_7__I_0_139_i11_2_lut_3_lut_4_lut (.I0(\state[0] ), .I1(\state[1] ), 
            .I2(\state[2] ), .I3(\state[3] ), .O(n11_adj_4002));
    defparam state_7__I_0_139_i11_2_lut_3_lut_4_lut.LUT_INIT = 16'hfff7;
    SB_LUT4 i26727_2_lut (.I0(\state_7__N_3914[3] ), .I1(n15_adj_4010), 
            .I2(GND_net), .I3(GND_net), .O(n33475));
    defparam i26727_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i17_4_lut (.I0(n5205), .I1(n33475), .I2(n5690), .I3(n37), 
            .O(n18768));
    defparam i17_4_lut.LUT_INIT = 16'h3a30;
    SB_LUT4 i4_4_lut (.I0(counter2[3]), .I1(counter2[5]), .I2(counter2[2]), 
            .I3(counter2[4]), .O(n10_adj_4011));
    defparam i4_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i5_3_lut (.I0(counter2[1]), .I1(n10_adj_4011), .I2(counter2[0]), 
            .I3(GND_net), .O(n18921));
    defparam i5_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 equal_1573_i19_2_lut_3_lut_4_lut (.I0(\state[1] ), .I1(\state[0] ), 
            .I2(\state[2] ), .I3(\state[3] ), .O(enable_slow_N_4001));
    defparam equal_1573_i19_2_lut_3_lut_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_4_lut_4_lut (.I0(\state[1] ), .I1(\state[2] ), .I2(\state[3] ), 
            .I3(\state[0] ), .O(n34));
    defparam i1_2_lut_4_lut_4_lut.LUT_INIT = 16'h0510;
    SB_LUT4 equal_100_i11_2_lut_3_lut_4_lut (.I0(\state[0] ), .I1(\state[1] ), 
            .I2(\state[2] ), .I3(\state[3] ), .O(n15_adj_4010));   // verilog/i2c_controller.v(77[27:43])
    defparam equal_100_i11_2_lut_3_lut_4_lut.LUT_INIT = 16'hfffd;
    SB_LUT4 state_7__I_0_144_i11_2_lut_3_lut_4_lut (.I0(\state[0] ), .I1(\state[1] ), 
            .I2(\state[2] ), .I3(\state[3] ), .O(n11_adj_4012));   // verilog/i2c_controller.v(77[27:43])
    defparam state_7__I_0_144_i11_2_lut_3_lut_4_lut.LUT_INIT = 16'hffdf;
    SB_LUT4 i1_4_lut_adj_837 (.I0(n11_adj_4012), .I1(n11_adj_4002), .I2(\state_7__N_3914[3] ), 
            .I3(\saved_addr[0] ), .O(n5));   // verilog/i2c_controller.v(92[4] 172[11])
    defparam i1_4_lut_adj_837.LUT_INIT = 16'h5755;
    SB_DFF data_out_i0_i0 (.Q(data[0]), .C(i2c_clk), .D(n19061));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFF data_out_i0_i5 (.Q(data[5]), .C(i2c_clk), .D(n19060));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFF saved_addr__i1 (.Q(\saved_addr[0] ), .C(i2c_clk), .D(n19056));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFF data_out_i0_i6 (.Q(data[6]), .C(i2c_clk), .D(n19055));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFF data_out_i0_i7 (.Q(data[7]), .C(i2c_clk), .D(n19054));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFF data_out_i0_i1 (.Q(data[1]), .C(i2c_clk), .D(n19592));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFF data_out_i0_i2 (.Q(data[2]), .C(i2c_clk), .D(n19584));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFF data_out_i0_i3 (.Q(data[3]), .C(i2c_clk), .D(n19582));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFF data_out_i0_i4 (.Q(data[4]), .C(i2c_clk), .D(n19558));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFFE state_i0_i0 (.Q(\state[0] ), .C(i2c_clk), .E(VCC_net), .D(n8));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_LUT4 i18699_2_lut (.I0(i2c_clk), .I1(scl_enable), .I2(GND_net), 
            .I3(GND_net), .O(scl));   // verilog/i2c_controller.v(45[19:61])
    defparam i18699_2_lut.LUT_INIT = 16'hbbbb;
    SB_LUT4 i1844_2_lut (.I0(sda_out_adj_4006), .I1(sda_enable), .I2(GND_net), 
            .I3(GND_net), .O(sda_out));   // verilog/i2c_controller.v(46[9:20])
    defparam i1844_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i26696_2_lut_4_lut (.I0(\state[0] ), .I1(\state[2] ), .I2(\state[3] ), 
            .I3(n33475), .O(n19001));   // verilog/i2c_controller.v(91[8] 173[6])
    defparam i26696_2_lut_4_lut.LUT_INIT = 16'h0002;
    SB_LUT4 i1_2_lut_4_lut (.I0(\state[3] ), .I1(\state[1] ), .I2(\state[2] ), 
            .I3(\state[0] ), .O(n37));
    defparam i1_2_lut_4_lut.LUT_INIT = 16'h0554;
    SB_LUT4 i30566_3_lut_4_lut (.I0(\state[2] ), .I1(\state[3] ), .I2(\state[1] ), 
            .I3(n5212), .O(n34096));
    defparam i30566_3_lut_4_lut.LUT_INIT = 16'h0200;
    SB_DFFSR counter2_1587_1588__i2 (.Q(counter2[1]), .C(CLK_c), .D(n29[1]), 
            .R(n18921));   // verilog/i2c_controller.v(69[20:35])
    SB_DFFSR counter2_1587_1588__i3 (.Q(counter2[2]), .C(CLK_c), .D(n29[2]), 
            .R(n18921));   // verilog/i2c_controller.v(69[20:35])
    SB_DFFSR counter2_1587_1588__i4 (.Q(counter2[3]), .C(CLK_c), .D(n29[3]), 
            .R(n18921));   // verilog/i2c_controller.v(69[20:35])
    SB_DFFSR counter2_1587_1588__i5 (.Q(counter2[4]), .C(CLK_c), .D(n29[4]), 
            .R(n18921));   // verilog/i2c_controller.v(69[20:35])
    SB_DFFSR counter2_1587_1588__i6 (.Q(counter2[5]), .C(CLK_c), .D(n29[5]), 
            .R(n18921));   // verilog/i2c_controller.v(69[20:35])
    SB_LUT4 i19164_2_lut_3_lut (.I0(\state[2] ), .I1(\state[3] ), .I2(\state[0] ), 
            .I3(GND_net), .O(n23736));
    defparam i19164_2_lut_3_lut.LUT_INIT = 16'hfdfd;
    SB_LUT4 i2_3_lut_4_lut (.I0(\state[0] ), .I1(\state[1] ), .I2(\state[2] ), 
            .I3(\state[3] ), .O(n11));   // verilog/i2c_controller.v(77[27:43])
    defparam i2_3_lut_4_lut.LUT_INIT = 16'hfdff;
    SB_LUT4 i29805_3_lut_4_lut (.I0(n11_adj_4008), .I1(n11), .I2(enable_slow_N_4001), 
            .I3(\state_7__N_3898[0] ), .O(n36289));
    defparam i29805_3_lut_4_lut.LUT_INIT = 16'h8088;
    SB_LUT4 i30561_3_lut_4_lut (.I0(n11_adj_4008), .I1(n11), .I2(n15_adj_4010), 
            .I3(n5212), .O(n24595));
    defparam i30561_3_lut_4_lut.LUT_INIT = 16'h7f00;
    SB_LUT4 state_7__I_0_143_i11_2_lut_3_lut_4_lut (.I0(\state[0] ), .I1(\state[1] ), 
            .I2(\state[2] ), .I3(\state[3] ), .O(n15));   // verilog/i2c_controller.v(151[5:14])
    defparam state_7__I_0_143_i11_2_lut_3_lut_4_lut.LUT_INIT = 16'hffbf;
    SB_LUT4 state_7__I_0_138_i11_2_lut_3_lut_4_lut (.I0(\state[0] ), .I1(\state[1] ), 
            .I2(\state[2] ), .I3(\state[3] ), .O(n11_adj_4008));   // verilog/i2c_controller.v(151[5:14])
    defparam state_7__I_0_138_i11_2_lut_3_lut_4_lut.LUT_INIT = 16'hfffb;
    SB_LUT4 i1_2_lut_3_lut (.I0(enable), .I1(\state_7__N_3898[0] ), .I2(enable_slow_N_4001), 
            .I3(GND_net), .O(n18648));
    defparam i1_2_lut_3_lut.LUT_INIT = 16'heaea;
    SB_LUT4 i56_3_lut_3_lut (.I0(\state[2] ), .I1(\state[3] ), .I2(\state[0] ), 
            .I3(GND_net), .O(n33));
    defparam i56_3_lut_3_lut.LUT_INIT = 16'h3434;
    SB_LUT4 i22_3_lut_3_lut (.I0(\state[1] ), .I1(\state[0] ), .I2(\state[3] ), 
            .I3(GND_net), .O(n11_adj_4003));
    defparam i22_3_lut_3_lut.LUT_INIT = 16'h1c1c;
    SB_LUT4 i19558_3_lut_4_lut (.I0(\state[1] ), .I1(\state[0] ), .I2(\state[2] ), 
            .I3(n15_adj_4010), .O(scl_enable_N_3988));
    defparam i19558_3_lut_4_lut.LUT_INIT = 16'hfe00;
    SB_LUT4 i1_3_lut_4_lut (.I0(\state[0] ), .I1(\state[1] ), .I2(\state[2] ), 
            .I3(\state[3] ), .O(n18565));
    defparam i1_3_lut_4_lut.LUT_INIT = 16'hf800;
    SB_LUT4 equal_158_i4_2_lut (.I0(counter[1]), .I1(counter[2]), .I2(GND_net), 
            .I3(GND_net), .O(n4));   // verilog/i2c_controller.v(153[6:23])
    defparam equal_158_i4_2_lut.LUT_INIT = 16'hdddd;
    SB_LUT4 i30418_4_lut_4_lut (.I0(\state[1] ), .I1(\state[2] ), .I2(\state[0] ), 
            .I3(\state[3] ), .O(n32365));
    defparam i30418_4_lut_4_lut.LUT_INIT = 16'h0156;
    SB_LUT4 i18709_2_lut (.I0(counter[1]), .I1(counter[2]), .I2(GND_net), 
            .I3(GND_net), .O(n23836));
    defparam i18709_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_838 (.I0(n15), .I1(counter[0]), .I2(GND_net), 
            .I3(GND_net), .O(n17518));   // verilog/i2c_controller.v(91[8] 173[6])
    defparam i1_2_lut_adj_838.LUT_INIT = 16'hbbbb;
    SB_LUT4 equal_155_i4_2_lut (.I0(counter[1]), .I1(counter[2]), .I2(GND_net), 
            .I3(GND_net), .O(n4_adj_2));   // verilog/i2c_controller.v(153[6:23])
    defparam equal_155_i4_2_lut.LUT_INIT = 16'hbbbb;
    SB_LUT4 i1_2_lut_adj_839 (.I0(counter[0]), .I1(n15), .I2(GND_net), 
            .I3(GND_net), .O(n17513));   // verilog/i2c_controller.v(91[8] 173[6])
    defparam i1_2_lut_adj_839.LUT_INIT = 16'heeee;
    
endmodule
//
// Verilog Description of module \quad(DEBOUNCE_TICKS=100) 
//

module \quad(DEBOUNCE_TICKS=100)  (encoder1_position, clk32MHz, data_o, 
            GND_net, ENCODER1_A_c_1, reg_B, VCC_net, n35209, n19053, 
            ENCODER1_B_c_0, n19593) /* synthesis syn_module_defined=1 */ ;
    output [23:0]encoder1_position;
    input clk32MHz;
    output [1:0]data_o;
    input GND_net;
    input ENCODER1_A_c_1;
    output [1:0]reg_B;
    input VCC_net;
    output n35209;
    input n19053;
    input ENCODER1_B_c_0;
    input n19593;
    
    wire clk32MHz /* synthesis SET_AS_NETWORK=clk32MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(33[6:14])
    wire [23:0]n3153;
    
    wire count_enable, B_delayed, A_delayed, count_direction, n3142, 
        n28073, n28072, n28071, n28070, n28069, n28068, n28067, 
        n28066, n28065, n28064, n28063, n28062, n28061, n28060, 
        n28059, n28058, n28057, n28056, n28055, n28054, n28053, 
        n28052, n28051, n28050;
    
    SB_DFFE count_i0_i0 (.Q(encoder1_position[0]), .C(clk32MHz), .E(count_enable), 
            .D(n3153[0]));   // quad.v(35[10] 41[6])
    SB_DFF B_delayed_16 (.Q(B_delayed), .C(clk32MHz), .D(data_o[0]));   // quad.v(23[10:54])
    SB_DFF A_delayed_15 (.Q(A_delayed), .C(clk32MHz), .D(data_o[1]));   // quad.v(22[10:54])
    SB_LUT4 quadA_debounced_I_0_2_lut (.I0(data_o[1]), .I1(B_delayed), .I2(GND_net), 
            .I3(GND_net), .O(count_direction));   // quad.v(26[26:53])
    defparam quadA_debounced_I_0_2_lut.LUT_INIT = 16'h6666;
    SB_DFFE count_i0_i23 (.Q(encoder1_position[23]), .C(clk32MHz), .E(count_enable), 
            .D(n3153[23]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i22 (.Q(encoder1_position[22]), .C(clk32MHz), .E(count_enable), 
            .D(n3153[22]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i21 (.Q(encoder1_position[21]), .C(clk32MHz), .E(count_enable), 
            .D(n3153[21]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i20 (.Q(encoder1_position[20]), .C(clk32MHz), .E(count_enable), 
            .D(n3153[20]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i19 (.Q(encoder1_position[19]), .C(clk32MHz), .E(count_enable), 
            .D(n3153[19]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i18 (.Q(encoder1_position[18]), .C(clk32MHz), .E(count_enable), 
            .D(n3153[18]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i17 (.Q(encoder1_position[17]), .C(clk32MHz), .E(count_enable), 
            .D(n3153[17]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i16 (.Q(encoder1_position[16]), .C(clk32MHz), .E(count_enable), 
            .D(n3153[16]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i15 (.Q(encoder1_position[15]), .C(clk32MHz), .E(count_enable), 
            .D(n3153[15]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i14 (.Q(encoder1_position[14]), .C(clk32MHz), .E(count_enable), 
            .D(n3153[14]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i13 (.Q(encoder1_position[13]), .C(clk32MHz), .E(count_enable), 
            .D(n3153[13]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i12 (.Q(encoder1_position[12]), .C(clk32MHz), .E(count_enable), 
            .D(n3153[12]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i11 (.Q(encoder1_position[11]), .C(clk32MHz), .E(count_enable), 
            .D(n3153[11]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i10 (.Q(encoder1_position[10]), .C(clk32MHz), .E(count_enable), 
            .D(n3153[10]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i9 (.Q(encoder1_position[9]), .C(clk32MHz), .E(count_enable), 
            .D(n3153[9]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i8 (.Q(encoder1_position[8]), .C(clk32MHz), .E(count_enable), 
            .D(n3153[8]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i7 (.Q(encoder1_position[7]), .C(clk32MHz), .E(count_enable), 
            .D(n3153[7]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i6 (.Q(encoder1_position[6]), .C(clk32MHz), .E(count_enable), 
            .D(n3153[6]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i5 (.Q(encoder1_position[5]), .C(clk32MHz), .E(count_enable), 
            .D(n3153[5]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i4 (.Q(encoder1_position[4]), .C(clk32MHz), .E(count_enable), 
            .D(n3153[4]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i3 (.Q(encoder1_position[3]), .C(clk32MHz), .E(count_enable), 
            .D(n3153[3]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i2 (.Q(encoder1_position[2]), .C(clk32MHz), .E(count_enable), 
            .D(n3153[2]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i1 (.Q(encoder1_position[1]), .C(clk32MHz), .E(count_enable), 
            .D(n3153[1]));   // quad.v(35[10] 41[6])
    SB_LUT4 i3_4_lut (.I0(data_o[1]), .I1(A_delayed), .I2(B_delayed), 
            .I3(data_o[0]), .O(count_enable));   // quad.v(25[23:80])
    defparam i3_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 add_715_25_lut (.I0(GND_net), .I1(encoder1_position[23]), .I2(n3142), 
            .I3(n28073), .O(n3153[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_715_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_715_24_lut (.I0(GND_net), .I1(encoder1_position[22]), .I2(n3142), 
            .I3(n28072), .O(n3153[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_715_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_715_24 (.CI(n28072), .I0(encoder1_position[22]), .I1(n3142), 
            .CO(n28073));
    SB_LUT4 add_715_23_lut (.I0(GND_net), .I1(encoder1_position[21]), .I2(n3142), 
            .I3(n28071), .O(n3153[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_715_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_715_23 (.CI(n28071), .I0(encoder1_position[21]), .I1(n3142), 
            .CO(n28072));
    SB_LUT4 add_715_22_lut (.I0(GND_net), .I1(encoder1_position[20]), .I2(n3142), 
            .I3(n28070), .O(n3153[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_715_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_715_22 (.CI(n28070), .I0(encoder1_position[20]), .I1(n3142), 
            .CO(n28071));
    SB_LUT4 add_715_21_lut (.I0(GND_net), .I1(encoder1_position[19]), .I2(n3142), 
            .I3(n28069), .O(n3153[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_715_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_715_21 (.CI(n28069), .I0(encoder1_position[19]), .I1(n3142), 
            .CO(n28070));
    SB_LUT4 add_715_20_lut (.I0(GND_net), .I1(encoder1_position[18]), .I2(n3142), 
            .I3(n28068), .O(n3153[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_715_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_715_20 (.CI(n28068), .I0(encoder1_position[18]), .I1(n3142), 
            .CO(n28069));
    SB_LUT4 add_715_19_lut (.I0(GND_net), .I1(encoder1_position[17]), .I2(n3142), 
            .I3(n28067), .O(n3153[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_715_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_715_19 (.CI(n28067), .I0(encoder1_position[17]), .I1(n3142), 
            .CO(n28068));
    SB_LUT4 add_715_18_lut (.I0(GND_net), .I1(encoder1_position[16]), .I2(n3142), 
            .I3(n28066), .O(n3153[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_715_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_715_18 (.CI(n28066), .I0(encoder1_position[16]), .I1(n3142), 
            .CO(n28067));
    SB_LUT4 add_715_17_lut (.I0(GND_net), .I1(encoder1_position[15]), .I2(n3142), 
            .I3(n28065), .O(n3153[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_715_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_715_17 (.CI(n28065), .I0(encoder1_position[15]), .I1(n3142), 
            .CO(n28066));
    SB_LUT4 add_715_16_lut (.I0(GND_net), .I1(encoder1_position[14]), .I2(n3142), 
            .I3(n28064), .O(n3153[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_715_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_715_16 (.CI(n28064), .I0(encoder1_position[14]), .I1(n3142), 
            .CO(n28065));
    SB_LUT4 add_715_15_lut (.I0(GND_net), .I1(encoder1_position[13]), .I2(n3142), 
            .I3(n28063), .O(n3153[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_715_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_715_15 (.CI(n28063), .I0(encoder1_position[13]), .I1(n3142), 
            .CO(n28064));
    SB_LUT4 add_715_14_lut (.I0(GND_net), .I1(encoder1_position[12]), .I2(n3142), 
            .I3(n28062), .O(n3153[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_715_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_715_14 (.CI(n28062), .I0(encoder1_position[12]), .I1(n3142), 
            .CO(n28063));
    SB_LUT4 add_715_13_lut (.I0(GND_net), .I1(encoder1_position[11]), .I2(n3142), 
            .I3(n28061), .O(n3153[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_715_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_715_13 (.CI(n28061), .I0(encoder1_position[11]), .I1(n3142), 
            .CO(n28062));
    SB_LUT4 add_715_12_lut (.I0(GND_net), .I1(encoder1_position[10]), .I2(n3142), 
            .I3(n28060), .O(n3153[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_715_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_715_12 (.CI(n28060), .I0(encoder1_position[10]), .I1(n3142), 
            .CO(n28061));
    SB_LUT4 add_715_11_lut (.I0(GND_net), .I1(encoder1_position[9]), .I2(n3142), 
            .I3(n28059), .O(n3153[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_715_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_715_11 (.CI(n28059), .I0(encoder1_position[9]), .I1(n3142), 
            .CO(n28060));
    SB_LUT4 add_715_10_lut (.I0(GND_net), .I1(encoder1_position[8]), .I2(n3142), 
            .I3(n28058), .O(n3153[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_715_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_715_10 (.CI(n28058), .I0(encoder1_position[8]), .I1(n3142), 
            .CO(n28059));
    SB_LUT4 add_715_9_lut (.I0(GND_net), .I1(encoder1_position[7]), .I2(n3142), 
            .I3(n28057), .O(n3153[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_715_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_715_9 (.CI(n28057), .I0(encoder1_position[7]), .I1(n3142), 
            .CO(n28058));
    SB_LUT4 add_715_8_lut (.I0(GND_net), .I1(encoder1_position[6]), .I2(n3142), 
            .I3(n28056), .O(n3153[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_715_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_715_8 (.CI(n28056), .I0(encoder1_position[6]), .I1(n3142), 
            .CO(n28057));
    SB_LUT4 add_715_7_lut (.I0(GND_net), .I1(encoder1_position[5]), .I2(n3142), 
            .I3(n28055), .O(n3153[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_715_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_715_7 (.CI(n28055), .I0(encoder1_position[5]), .I1(n3142), 
            .CO(n28056));
    SB_LUT4 add_715_6_lut (.I0(GND_net), .I1(encoder1_position[4]), .I2(n3142), 
            .I3(n28054), .O(n3153[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_715_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_715_6 (.CI(n28054), .I0(encoder1_position[4]), .I1(n3142), 
            .CO(n28055));
    SB_LUT4 add_715_5_lut (.I0(GND_net), .I1(encoder1_position[3]), .I2(n3142), 
            .I3(n28053), .O(n3153[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_715_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_715_5 (.CI(n28053), .I0(encoder1_position[3]), .I1(n3142), 
            .CO(n28054));
    SB_LUT4 add_715_4_lut (.I0(GND_net), .I1(encoder1_position[2]), .I2(n3142), 
            .I3(n28052), .O(n3153[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_715_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_715_4 (.CI(n28052), .I0(encoder1_position[2]), .I1(n3142), 
            .CO(n28053));
    SB_LUT4 add_715_3_lut (.I0(GND_net), .I1(encoder1_position[1]), .I2(n3142), 
            .I3(n28051), .O(n3153[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_715_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_715_3 (.CI(n28051), .I0(encoder1_position[1]), .I1(n3142), 
            .CO(n28052));
    SB_LUT4 add_715_2_lut (.I0(GND_net), .I1(encoder1_position[0]), .I2(count_direction), 
            .I3(n28050), .O(n3153[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_715_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_715_2 (.CI(n28050), .I0(encoder1_position[0]), .I1(count_direction), 
            .CO(n28051));
    SB_CARRY add_715_1 (.CI(GND_net), .I0(n3142), .I1(n3142), .CO(n28050));
    SB_LUT4 i1191_1_lut_2_lut (.I0(data_o[1]), .I1(B_delayed), .I2(GND_net), 
            .I3(GND_net), .O(n3142));   // quad.v(37[5] 40[8])
    defparam i1191_1_lut_2_lut.LUT_INIT = 16'h9999;
    \grp_debouncer(2,100)  debounce (.ENCODER1_A_c_1(ENCODER1_A_c_1), .clk32MHz(clk32MHz), 
            .reg_B({reg_B}), .GND_net(GND_net), .VCC_net(VCC_net), .n35209(n35209), 
            .n19053(n19053), .data_o({data_o}), .ENCODER1_B_c_0(ENCODER1_B_c_0), 
            .n19593(n19593));   // quad.v(15[37] 19[4])
    
endmodule
//
// Verilog Description of module \grp_debouncer(2,100) 
//

module \grp_debouncer(2,100)  (ENCODER1_A_c_1, clk32MHz, reg_B, GND_net, 
            VCC_net, n35209, n19053, data_o, ENCODER1_B_c_0, n19593);
    input ENCODER1_A_c_1;
    input clk32MHz;
    output [1:0]reg_B;
    input GND_net;
    input VCC_net;
    output n35209;
    input n19053;
    output [1:0]data_o;
    input ENCODER1_B_c_0;
    input n19593;
    
    wire clk32MHz /* synthesis SET_AS_NETWORK=clk32MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(33[6:14])
    wire [1:0]reg_A;   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(142[12:17])
    wire [6:0]n33;
    wire [6:0]cnt_reg;   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(149[12:19])
    
    wire n28624, n28623, n28622, n28621, n28620, n28619, n12, 
        n2, cnt_next_6__N_3730;
    
    SB_DFF reg_A_i1 (.Q(reg_A[1]), .C(clk32MHz), .D(ENCODER1_A_c_1));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(178[9] 184[16])
    SB_DFF reg_B_i0 (.Q(reg_B[0]), .C(clk32MHz), .D(reg_A[0]));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(178[9] 184[16])
    SB_LUT4 cnt_reg_1586_add_4_8_lut (.I0(GND_net), .I1(GND_net), .I2(cnt_reg[6]), 
            .I3(n28624), .O(n33[6])) /* synthesis syn_instantiated=1 */ ;
    defparam cnt_reg_1586_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 cnt_reg_1586_add_4_7_lut (.I0(GND_net), .I1(GND_net), .I2(cnt_reg[5]), 
            .I3(n28623), .O(n33[5])) /* synthesis syn_instantiated=1 */ ;
    defparam cnt_reg_1586_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY cnt_reg_1586_add_4_7 (.CI(n28623), .I0(GND_net), .I1(cnt_reg[5]), 
            .CO(n28624));
    SB_LUT4 cnt_reg_1586_add_4_6_lut (.I0(GND_net), .I1(GND_net), .I2(cnt_reg[4]), 
            .I3(n28622), .O(n33[4])) /* synthesis syn_instantiated=1 */ ;
    defparam cnt_reg_1586_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY cnt_reg_1586_add_4_6 (.CI(n28622), .I0(GND_net), .I1(cnt_reg[4]), 
            .CO(n28623));
    SB_LUT4 cnt_reg_1586_add_4_5_lut (.I0(GND_net), .I1(GND_net), .I2(cnt_reg[3]), 
            .I3(n28621), .O(n33[3])) /* synthesis syn_instantiated=1 */ ;
    defparam cnt_reg_1586_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY cnt_reg_1586_add_4_5 (.CI(n28621), .I0(GND_net), .I1(cnt_reg[3]), 
            .CO(n28622));
    SB_LUT4 cnt_reg_1586_add_4_4_lut (.I0(GND_net), .I1(GND_net), .I2(cnt_reg[2]), 
            .I3(n28620), .O(n33[2])) /* synthesis syn_instantiated=1 */ ;
    defparam cnt_reg_1586_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY cnt_reg_1586_add_4_4 (.CI(n28620), .I0(GND_net), .I1(cnt_reg[2]), 
            .CO(n28621));
    SB_LUT4 cnt_reg_1586_add_4_3_lut (.I0(GND_net), .I1(GND_net), .I2(cnt_reg[1]), 
            .I3(n28619), .O(n33[1])) /* synthesis syn_instantiated=1 */ ;
    defparam cnt_reg_1586_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY cnt_reg_1586_add_4_3 (.CI(n28619), .I0(GND_net), .I1(cnt_reg[1]), 
            .CO(n28620));
    SB_LUT4 cnt_reg_1586_add_4_2_lut (.I0(GND_net), .I1(GND_net), .I2(cnt_reg[0]), 
            .I3(VCC_net), .O(n33[0])) /* synthesis syn_instantiated=1 */ ;
    defparam cnt_reg_1586_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY cnt_reg_1586_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(cnt_reg[0]), 
            .CO(n28619));
    SB_LUT4 i5_4_lut (.I0(cnt_reg[1]), .I1(cnt_reg[4]), .I2(cnt_reg[3]), 
            .I3(cnt_reg[6]), .O(n12));
    defparam i5_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i6_4_lut (.I0(cnt_reg[5]), .I1(n12), .I2(cnt_reg[0]), .I3(cnt_reg[2]), 
            .O(n35209));
    defparam i6_4_lut.LUT_INIT = 16'hfdff;
    SB_LUT4 reg_B_1__I_0_i2_2_lut (.I0(reg_B[1]), .I1(reg_A[1]), .I2(GND_net), 
            .I3(GND_net), .O(n2));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(193[46:60])
    defparam reg_B_1__I_0_i2_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i2_4_lut (.I0(reg_B[0]), .I1(n35209), .I2(reg_A[0]), .I3(n2), 
            .O(cnt_next_6__N_3730));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[40:72])
    defparam i2_4_lut.LUT_INIT = 16'hff7b;
    SB_DFFSR cnt_reg_1586__i0 (.Q(cnt_reg[0]), .C(clk32MHz), .D(n33[0]), 
            .R(cnt_next_6__N_3730));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[78:85])
    SB_DFF reg_out_i0_i0 (.Q(data_o[0]), .C(clk32MHz), .D(n19053));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(186[9] 190[16])
    SB_DFF reg_B_i1 (.Q(reg_B[1]), .C(clk32MHz), .D(reg_A[1]));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(178[9] 184[16])
    SB_DFF reg_A_i0 (.Q(reg_A[0]), .C(clk32MHz), .D(ENCODER1_B_c_0));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(178[9] 184[16])
    SB_DFF reg_out_i0_i1 (.Q(data_o[1]), .C(clk32MHz), .D(n19593));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(186[9] 190[16])
    SB_DFFSR cnt_reg_1586__i1 (.Q(cnt_reg[1]), .C(clk32MHz), .D(n33[1]), 
            .R(cnt_next_6__N_3730));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[78:85])
    SB_DFFSR cnt_reg_1586__i2 (.Q(cnt_reg[2]), .C(clk32MHz), .D(n33[2]), 
            .R(cnt_next_6__N_3730));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[78:85])
    SB_DFFSR cnt_reg_1586__i3 (.Q(cnt_reg[3]), .C(clk32MHz), .D(n33[3]), 
            .R(cnt_next_6__N_3730));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[78:85])
    SB_DFFSR cnt_reg_1586__i4 (.Q(cnt_reg[4]), .C(clk32MHz), .D(n33[4]), 
            .R(cnt_next_6__N_3730));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[78:85])
    SB_DFFSR cnt_reg_1586__i5 (.Q(cnt_reg[5]), .C(clk32MHz), .D(n33[5]), 
            .R(cnt_next_6__N_3730));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[78:85])
    SB_DFFSR cnt_reg_1586__i6 (.Q(cnt_reg[6]), .C(clk32MHz), .D(n33[6]), 
            .R(cnt_next_6__N_3730));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[78:85])
    
endmodule
