// Verilog netlist produced by program LSE :  version Diamond Version 0.0.0
// Netlist written on Thu Jan  2 15:12:42 2020
//
// Verilog Description of module TinyFPGA_B
//

module TinyFPGA_B (CLK, LED, USBPU, PIN_1, PIN_2, PIN_3, PIN_4, 
            PIN_5, PIN_6, PIN_7, PIN_8, PIN_9, PIN_10, PIN_11, 
            PIN_12, PIN_13, PIN_14, PIN_15, PIN_16, PIN_17, PIN_18, 
            PIN_19, PIN_20, PIN_21, PIN_22, PIN_23, PIN_24) /* synthesis syn_preserve=0, syn_noprune=0, syn_module_defined=1 */ ;   // verilog/TinyFPGA_B.v(2[8:18])
    input CLK;   // verilog/TinyFPGA_B.v(3[9:12])
    output LED;   // verilog/TinyFPGA_B.v(4[10:13])
    output USBPU;   // verilog/TinyFPGA_B.v(5[10:15])
    input PIN_1 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(6[9:14])
    input PIN_2 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(7[9:14])
    inout PIN_3 /* synthesis black_box_pad_pin=1 */ ;   // verilog/TinyFPGA_B.v(8[9:14])
    inout PIN_4 /* synthesis black_box_pad_pin=1 */ ;   // verilog/TinyFPGA_B.v(9[9:14])
    inout PIN_5 /* synthesis black_box_pad_pin=1 */ ;   // verilog/TinyFPGA_B.v(10[9:14])
    input PIN_6 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(11[9:14])
    input PIN_7 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(12[9:14])
    output PIN_8 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(13[9:14])
    input PIN_9 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(14[9:14])
    input PIN_10 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(15[9:15])
    output PIN_11 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(16[9:15])
    inout PIN_12 /* synthesis black_box_pad_pin=1 */ ;   // verilog/TinyFPGA_B.v(17[9:15])
    input PIN_13 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(18[9:15])
    input PIN_14 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(19[9:15])
    input PIN_15 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(20[9:15])
    input PIN_16 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(21[9:15])
    input PIN_17 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(22[9:15])
    input PIN_18 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(23[9:15])
    output PIN_19 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(24[9:15])
    output PIN_20 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(25[9:15])
    output PIN_21 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(26[9:15])
    output PIN_22 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(27[9:15])
    output PIN_23 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(28[9:15])
    output PIN_24 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(29[9:15])
    
    wire CLK_c /* synthesis SET_AS_NETWORK=CLK_c, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(3[9:12])
    wire LED_c /* synthesis SET_AS_NETWORK=LED_c, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(4[10:13])
    wire clk32MHz /* synthesis SET_AS_NETWORK=clk32MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(34[6:14])
    
    wire GND_net, VCC_net, PIN_1_c_1, PIN_2_c_0, PIN_8_c, PIN_9_c_1, 
        PIN_10_c_0, PIN_11_c, PIN_13_c, PIN_19_c_0, PIN_20_c, PIN_21_c, 
        PIN_22_c, PIN_23_c;
    wire [31:0]communication_counter;   // verilog/TinyFPGA_B.v(45[9:30])
    wire [23:0]color;   // verilog/TinyFPGA_B.v(46[12:17])
    
    wire blink, hall1, hall2, hall3;
    wire [22:0]pwm_setpoint;   // verilog/TinyFPGA_B.v(129[13:25])
    wire [23:0]duty;   // verilog/TinyFPGA_B.v(130[21:25])
    
    wire tx_o, tx_enable;
    wire [23:0]encoder0_position;   // verilog/TinyFPGA_B.v(167[22:39])
    wire [23:0]encoder1_position;   // verilog/TinyFPGA_B.v(168[22:39])
    wire [23:0]displacement;   // verilog/TinyFPGA_B.v(169[21:33])
    wire [23:0]setpoint;   // verilog/TinyFPGA_B.v(170[22:30])
    wire [23:0]Kp;   // verilog/TinyFPGA_B.v(171[22:24])
    wire [23:0]Ki;   // verilog/TinyFPGA_B.v(172[22:24])
    
    wire n1722, n29596, n29595, n29594;
    wire [7:0]control_mode;   // verilog/TinyFPGA_B.v(174[14:26])
    wire [23:0]PWMLimit;   // verilog/TinyFPGA_B.v(175[22:30])
    wire [23:0]IntegralLimit;   // verilog/TinyFPGA_B.v(176[22:35])
    
    wire n1522, n1517, n1481, n28577;
    wire [23:0]motor_state;   // verilog/TinyFPGA_B.v(207[22:33])
    
    wire n28576, n29593, n28575, n1458, n37363, n37362, n28425, 
        n28424, n1449, n1448, n1847, n28423;
    wire [7:0]color_23__N_209;
    wire [31:0]timer;   // verilog/neopixel.v(9[12:17])
    
    wire n29592, n28574, n1623, n28573, n1558, n28572, n28191, 
        n20, blink_N_354;
    wire [22:0]pwm_setpoint_22__N_57;
    
    wire PIN_13_N_105, n29591, n28190, n28422, n1466, n1460, n28421, 
        n28189, n28571, n1817, n28188, n29590, n3219, n29589, 
        n28420, n3218, n29588, n3217, n37361, n29587, n29586;
    wire [23:0]displacement_23__N_80;
    
    wire n1825, n1824, n28187, n28570, n1823, n29585, n1822, n1821, 
        n1619, n1618, n29584, n1819, n28419, n29583, n1818, n1816, 
        n1815, n1778, n1756, n1755, n1753, n1751, n1750, n28569, 
        n28418, n28186, n28568, n28417, n1525, n1524, n1523, n1521, 
        n1520, n1519, n1518;
    wire [3:0]state;   // verilog/neopixel.v(16[20:25])
    wire [31:0]bit_ctr;   // verilog/neopixel.v(18[12:19])
    
    wire start, \neo_pixel_transmitter.done ;
    wire [31:0]\neo_pixel_transmitter.t0 ;   // verilog/neopixel.v(28[14:16])
    
    wire n1516, n28416, n1814, n63, n28415, n1617, n29582, n29581, 
        n28185, n28414, n29580, n28413, n28567, n28184, n28566;
    wire [3:0]state_3__N_462;
    
    wire n29579, n1717, n28565, n28564, n28412, n28183, n37360, 
        n1418, n1417, n1813, n28411, n29578, n28563, n28410, n28409, 
        n28562, n28714, n28561, n28713, n28408, n28407, n28406, 
        n28712, n28711, n3216, n3215, n3214, n28710, n28709, n29577, 
        n28708, n28560, n28405, n28404, n28559, n28558, n28403, 
        n28402, n1358, n1357, n1356, n1355, n1354, n28707, n5439, 
        n3213, n3212, n28706, n28705, n28557, n1749, n3211, n37359, 
        n28704, n3210, n1353, n29576, n28401, n29575, n28703, 
        n1452, n1352, n29574, n29573, n18147, n18146, n37, n28702, 
        n3209, n3182, n3181, n3180, n3179, n1351, n1350, n1349, 
        n28701, n28700, n28699, n37358, n28698, n28400, n28182, 
        n35, n34, n28697, n28696, n28556, n28695, n3178, n33975, 
        n3177, n29572, n3176, n3175, n1324, n1715, n1752, n3174, 
        n3173, n2958, n29571, n3172, n3171, n3170, n3169, n3168, 
        n3167, n3166, n3165, n3164, n3163, n3162, n3161, n3160, 
        n28555, n28694, n3159, n28693, n32, n31, n28554, n28553, 
        n29570, n28399, n28398, n28552, n29569, n28692, n4, n37357, 
        n25, n28181, n28180, n28691, n17567, n1748, n1820, n28690, 
        n1724, n39, n1425, n31599, n1557;
    wire [9:0]half_duty_new;   // vhdl/pwm.vhd(53[12:25])
    
    wire n1554, n37_adj_4770;
    wire [9:0]\half_duty[0] ;   // vhdl/pwm.vhd(55[11:20])
    
    wire n1553, n1424, n1423, n1552, n1549, n1547, n36, n1382, 
        n12, n34_adj_4771, n33, n28551, n28689, n28550, n3, n4_adj_4772, 
        n5, n6, n7, n8, n9, n10, n11, n12_adj_4773, n13, n14, 
        n15, n16, n17, n18, n19, n20_adj_4774, n21, n22, n23, 
        n24, n25_adj_4775, rx_data_ready;
    wire [7:0]rx_data;   // verilog/coms.v(90[13:20])
    wire [7:0]\data_in[3] ;   // verilog/coms.v(94[12:19])
    wire [7:0]\data_in[2] ;   // verilog/coms.v(94[12:19])
    wire [7:0]\data_in[1] ;   // verilog/coms.v(94[12:19])
    wire [7:0]\data_in[0] ;   // verilog/coms.v(94[12:19])
    wire [7:0]\data_in_frame[17] ;   // verilog/coms.v(95[12:25])
    wire [7:0]\data_in_frame[13] ;   // verilog/coms.v(95[12:25])
    wire [7:0]\data_in_frame[12] ;   // verilog/coms.v(95[12:25])
    wire [7:0]\data_in_frame[11] ;   // verilog/coms.v(95[12:25])
    wire [7:0]\data_in_frame[10] ;   // verilog/coms.v(95[12:25])
    wire [7:0]\data_in_frame[9] ;   // verilog/coms.v(95[12:25])
    wire [7:0]\data_in_frame[8] ;   // verilog/coms.v(95[12:25])
    wire [7:0]\data_in_frame[5] ;   // verilog/coms.v(95[12:25])
    wire [7:0]\data_in_frame[4] ;   // verilog/coms.v(95[12:25])
    wire [7:0]\data_in_frame[3] ;   // verilog/coms.v(95[12:25])
    wire [7:0]\data_in_frame[2] ;   // verilog/coms.v(95[12:25])
    wire [7:0]\data_in_frame[1] ;   // verilog/coms.v(95[12:25])
    wire [7:0]\data_out_frame[23] ;   // verilog/coms.v(96[12:26])
    
    wire n27;
    wire [7:0]\data_out_frame[20] ;   // verilog/coms.v(96[12:26])
    wire [7:0]\data_out_frame[19] ;   // verilog/coms.v(96[12:26])
    wire [7:0]\data_out_frame[18] ;   // verilog/coms.v(96[12:26])
    wire [7:0]\data_out_frame[17] ;   // verilog/coms.v(96[12:26])
    wire [7:0]\data_out_frame[16] ;   // verilog/coms.v(96[12:26])
    wire [7:0]\data_out_frame[15] ;   // verilog/coms.v(96[12:26])
    wire [7:0]\data_out_frame[14] ;   // verilog/coms.v(96[12:26])
    wire [7:0]\data_out_frame[13] ;   // verilog/coms.v(96[12:26])
    wire [7:0]\data_out_frame[12] ;   // verilog/coms.v(96[12:26])
    wire [7:0]\data_out_frame[11] ;   // verilog/coms.v(96[12:26])
    wire [7:0]\data_out_frame[10] ;   // verilog/coms.v(96[12:26])
    wire [7:0]\data_out_frame[9] ;   // verilog/coms.v(96[12:26])
    wire [7:0]\data_out_frame[8] ;   // verilog/coms.v(96[12:26])
    wire [7:0]\data_out_frame[7] ;   // verilog/coms.v(96[12:26])
    wire [7:0]\data_out_frame[6] ;   // verilog/coms.v(96[12:26])
    wire [7:0]\data_out_frame[5] ;   // verilog/coms.v(96[12:26])
    
    wire n22_adj_4776;
    wire [7:0]byte_transmit_counter;   // verilog/coms.v(101[12:33])
    
    wire tx_active, n28688, n40, n39_adj_4777, n38, n37_adj_4778, 
        n28549, n28548, n28547, n28546, n28545, n28544, n35_adj_4779, 
        n31583;
    wire [31:0]\FRAME_MATCHER.state_31__N_2566 ;
    
    wire n34_adj_4780, n1757, n1747, n1746, n1745, n28, n28543, 
        n28397, n28179, n28542, n28178, n28687, n28177, n28396, 
        n28541, n28395, n28394, n28540, n28176, n28175, n28174, 
        n28173, n28686, n28172, n28539, n28685, n28393, n28538, 
        n28392, n33879, n4_adj_4781, n28171, n1758, n1754, n28684, 
        n34531, n33944, n10_adj_4782, n33228, n737, n28391, n28390, 
        n28389, n28388, n28387, n30, n29, n28_adj_4783, n27_adj_4784, 
        n28537, n18_adj_4785, n28170, n28169, n28168, n28167, n28386, 
        n13724, n28683, n28536, n28682, n28535, n28534, n28681, 
        n28533, n28532, n1, n37356, n37355, n36489, n28680, n28679, 
        n37713, n28531, n32849, n37354, n37353, n37369, n5_adj_4786, 
        n16159, n31527, n16154, n28385, n28678, n36654, n37711, 
        tx_transmit_N_3355, n1422, n37368, n28677, n31521, n28384, 
        n3007, n28383, n28382, n28381, n28380, n28379, n28378, 
        n28377, n17534, n16143, n17527, n37364, n37365, n1421, 
        n1420, n3893, n28676, n28675, n28674, n28673, n28672, 
        n28671, n42, n41, n40_adj_4787, n39_adj_4788, n37_adj_4789, 
        n36_adj_4790, n30_adj_4791, n44, n43, n42_adj_4792, n41_adj_4793, 
        n40_adj_4794, n13_adj_4795, n36485, n11_adj_4796, n37352, 
        n37351, n38_adj_4797, n38232, n37350, n37349, n28670, n28530, 
        n28376, n28166, n28085, n28084, n28165, n28083, n28082, 
        n34029, n28375, n28164, n28081, n28080, n28163, n34037, 
        n28079, n33985, n33873, n33917, n1457, n1456, n1455, n1454, 
        n1453, n1451, n1450, n37348, n28529, n28528, n28527, n28526, 
        n28078, n28077, n28669, n1719, n28525, n28374, n28162, 
        n24786, n28076, n28075, n28161, n28074, n28073, n18278, 
        n18275, n18274, n18273, n18272, n18271, n18270, n18268, 
        n18267, n18266, n18265, n1419, n18264, n18261, n18260, 
        n18256, n18255, n18254, n18253, n18252, n18251, n18250, 
        n18249, n18248, n28373, n18247, n18246, n18245, n1718, 
        n4_adj_4798, n18244, n18243, n18242, n18241, n18240, n18239, 
        n18238, n18237, n18236, n18235, n18234, n18231, n18230, 
        n18229, n18025, n18024, n18023, n18022, n18021, n18020, 
        n18019, n18018, n18010, n18009, n18008, n18007, n18006, 
        n18005, n18004, n18003, n18002, n18001, n18000, n17999, 
        n17998, n17997, n17996, n17995, n17994, n17993, n17992, 
        n17991, n17990, n17989, n17988, n17987, n17986, n17985, 
        n17984, n17983, n17982, n17981, n17980, n17979, n17978, 
        n17977, n17976, n17975, n17974, n17973, n17972, n17971, 
        n17970, n17969, n17968, n17967, n17966, n17965, n17964, 
        n17963, n17962, n17961, n17960, n17959, n17958, n17957, 
        n17956, n17955, n17954, n17953, n17952, n17951, n17950, 
        n17949, n17948, n17947, n17946, n17945, n17944, n17943, 
        n17942, n17941, n17940, n17939, n17938, n17937, n17936, 
        n17935, n17934, n17933, n17932, n17931, n17930, n17929, 
        n17928, n17927, n17926, n17925, n17924, n17923, n17922, 
        n17921, n17920, n17919, n17918, n17917, n17916, n17915, 
        n17914, n17913, n17912, n17911, n17910, n17909, n17908, 
        n17907, n17906, n17905, n17904, n17903, n17902, n17901, 
        n17900, n17899, n17898, n17897, n17896, n17895, n17894, 
        n17893, n17892, n17891, n17890, n17889, n17888, n17887, 
        n17886, n17885, n17884, n17883, n17882, n17881, n17880, 
        n17879, n17878, n17877, n17876, n17875, n17874, n17873, 
        n17872, n17871, n17870, n17869, n17868, n17867, n17866, 
        n17865, n17864, n17863, n17862, n17861, n17860, n17859, 
        n17858, n17857, n17856, n17855, n17854, n17853, n17852, 
        n17851, n17850, n17849, n17848, n17847, n17846, n17845, 
        n17844, n17843, n17842, n17841, n17840, n17839, n17838, 
        n17837, n17836, n17835, n18228, n18227, n18226, n18225, 
        n18224, n18223, n18222, n28160, n16157, n16158, n18221, 
        n18220, n18219, n18218, n18217, n18216, n18215, n18214, 
        n18213, n18212, n18211, n18210, n18209, n17834, n17833, 
        n17832, n17831, n17830, n17829, n17828, n17827, n17826, 
        n17825, n17824, n17823, n17822, n17821, n17820, n17818, 
        n17816, n17814, n17813, n17812, n17810, n17808, n17806, 
        n17805, n17804, n17803, n17802, n18208, n18207, n18206, 
        n18205, n18204, n18203, n18202, n18201, n18200, n18199, 
        n18198, n18197, n18196, n18195, n18194, n1655, n18193, 
        n18192, n18191, n18190, n18189, n18188, n18187, n18186, 
        n28072, n28372, n30_adj_4799, n28071, n17801, n28159, n28070, 
        n17800, n17799, n17798, n28668, n17500, n17362, n1580, 
        n28524, n28371, n17797, n54, n5578, n17796, n17795, n17794, 
        n26, n28158, n26_adj_4800, n24_adj_4801, n36481, n22_adj_4802, 
        n28667, n28523, n7_adj_4803, n28370, n37347, n37346, n37345, 
        n17793, n37344, n37343, n17791, n8014, n18_adj_4804, n28157, 
        n28522, quadA_debounced, quadB_debounced, count_enable, n28069, 
        n28666, n5600, n28521, n28068, n18148, n28156, n28369, 
        n37342, n28067, n37341, n1647, quadA_debounced_adj_4805, quadB_debounced_adj_4806, 
        count_enable_adj_4807, n28066, n37340, n37339, n28065, n28665, 
        n3232, n3231, n3230, n3229, n3228, n3227, n3226, n3225, 
        n17308, n17790, n37338, n17789, n28064, n17788, n17787, 
        n1550, n37337, n17786, n17785, n17784, n17783, n17782, 
        n17781, n17780, n17779, n17778, n17777, n17776, n17775, 
        n37336, n17774, n17773, n17772, n28368, n17771, n17770, 
        n4_adj_4808, n17769, n28664, n28520, n17768, n47, n28063, 
        n17767, n17766, n46, n1556, n17765, n17764, n17763, n17762, 
        n17761, n1720, n17760, n17759, n17758, n17757, n1846, 
        n1844, n1624, n1616, n17756, n37335, n17755, n37333, n17754, 
        n17753, n17752, n10_adj_4809, n28062, n17751, n37332, n28061, 
        n1621, n1615, n17750, n28519, n17749, n3224, n3223, n3222, 
        n3221, n3220, n17748, n17747, n17746, n17745, n17744, 
        n17743, n17742, n17741, n17740, n17739, n17738, n17737, 
        n24193, n17735, n34002, n17229, n17731, n17728, n43_adj_4810, 
        n31529, n42_adj_4811, r_Rx_Data;
    wire [2:0]r_Bit_Index;   // verilog/uart_rx.v(33[17:28])
    wire [2:0]r_SM_Main;   // verilog/uart_rx.v(36[17:26])
    
    wire n9_adj_4812, n31531, n31533, n31535, n17713, n17710, n17708, 
        n40_adj_4813, n1548, n39_adj_4814, n28060, n28059, n33949, 
        n17705, n17701, n17700, n17699, n28058, n38238, n17697, 
        n17696, n17694, n17693, n17692, n17691, n17690, n17689;
    wire [2:0]r_SM_Main_adj_5047;   // verilog/uart_tx.v(31[16:25])
    wire [8:0]r_Clock_Count_adj_5048;   // verilog/uart_tx.v(32[16:29])
    wire [2:0]r_Bit_Index_adj_5049;   // verilog/uart_tx.v(33[16:27])
    
    wire n28367, n37330, n5019, n5018;
    wire [2:0]r_SM_Main_2__N_3458;
    
    wire n5017, n313, n314, n315, n5016, n5015, n28366, n38_adj_4819, 
        n17688, n17687, n17686, n17685, n17684, n17683, n17682, 
        n17681, n5014, n5013, n28518, n17679, n5478, n17676, n17674, 
        n17673, n17671, n316, n318, n321, n18152;
    wire [1:0]reg_B;   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(142[19:24])
    
    wire n17670, n17668, n17667, n17665;
    wire [1:0]reg_B_adj_5056;   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(142[19:24])
    
    wire n17664, n17662, n17661, n17659, n5012, n5011, n5010, 
        n5009, n5008, n5007, n5006, n5005, n5004, n5003, n5002, 
        n5001, n5000, n4999, n4998, n4997, n4996, n17658, n17656, 
        n17655, n1646, n1625, n4_adj_4822, n18153, n17652, n1649, 
        n8_adj_4823, n28517, n1622, n31537, n1620, n7_adj_4824, 
        n31539, n31541, n31543, n1658, n6_adj_4825, n28365, n31545, 
        n1648, n1657, n31547, n1650, n31549, n32_adj_4826, n31551, 
        n5_adj_4827, n1654, n17559, n34_adj_4828, n1716, n33_adj_4829, 
        n28364, n1714, n1656, n28057, n28056, n4_adj_4830, n32_adj_4831, 
        n31_adj_4832, n30_adj_4833, n28663, n28662, n1725, n1653, 
        n28661, n3_adj_4834, n1652, n28516, n1723, n1651, n28363, 
        n28055, n28054, n1721, n31553, n2, n1845, n1555, n31555, 
        n1551, n11_adj_4835, n12_adj_4836, n13_adj_4837, n14_adj_4838, 
        n15_adj_4839, n16_adj_4840, n17_adj_4841, n18_adj_4842, n19_adj_4843, 
        n20_adj_4844, n21_adj_4845, n22_adj_4846, n23_adj_4847, n24_adj_4848, 
        n25_adj_4849, n31557, n15_adj_4850, n31559, n33_adj_4851, 
        n32_adj_4852, n31_adj_4853, n30_adj_4854, n29_adj_4855, n28_adj_4856, 
        n27_adj_4857, n26_adj_4858, n25_adj_4859, n24_adj_4860, n23_adj_4861, 
        n22_adj_4862, n21_adj_4863, n20_adj_4864, n19_adj_4865, n18_adj_4866, 
        n17_adj_4867, n16_adj_4868, n15_adj_4869, n14_adj_4870, n13_adj_4871, 
        n12_adj_4872, n1325, n28515, n1323, n1322, n28514, n1321, 
        n28660, n1320, n1319, n1318, n28513, n28512, n28659, n28511, 
        n28510, n28658, n28509, n28508, n28657, n1283, n28053, 
        n28507, n28506, n28656, n1258, n1257, n1256, n1255, n28362, 
        n1254, n28052, n1253, n1252, n1251, n28505, n1250, n28504, 
        n28655, n28503, n28051, n28050, n1225, n1224, n1223, n1222, 
        n1221, n1220, n1219, n27896, n27895, n27894, n1184, n27893, 
        n28247, n37310, n1158, n1157, n1156, n1155, n1154, n28502, 
        n1153, n28501, n28500, n1152, n33925, n1151, n37309, n11_adj_4873, 
        n10_adj_4874, n9_adj_4875, n8_adj_4876, n7_adj_4877, n6_adj_4878, 
        n5_adj_4879, n4_adj_4880, n3_adj_4881, n1021, n1053, n1022, 
        n1054, n1023, n1055, n1024, n1056, n1025, n1057, n1058, 
        n37308, n1052, n134, n135, n136, n137, n138, n139, n140, 
        n141, n142, n143, n144, n145, n146, n147, n148, n149, 
        n150, n151, n152, n153, n154, n155, n156, n157, n158, 
        n159, n160, n161, n162, n163, n164, n165, n986, n37304, 
        n953, n954, n955, n956, n957, n958, n1125, n1679, n1124, 
        n1123, n1122, n1121, n1120, n852, n855, n746, n748, 
        n749, n17553, n17550, n17549, n31561, n31563, n31565, 
        n31567, n36301, n28246, n36297, n31569, n31571, n31573, 
        n31575, n31577, n31585, n31587, n31589, n28654, n1085, 
        n28653, n31591, n28499, n1848, n1849, n1850, n1851, n1852, 
        n1853, n1854, n1855, n1856, n1857, n1858, n1877, n1912, 
        n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, 
        n1921, n1922, n1923, n1924, n1925, n1943, n1944, n1945, 
        n1946, n1947, n1948, n1949, n1950, n1951, n1952, n1953, 
        n1954, n1955, n1956, n1957, n1958, n28652, n28245, n1976, 
        n2011, n2012, n2013, n2014, n2015, n2016, n2017, n2018, 
        n2019, n2020, n2021, n2022, n2023, n2024, n2025, n2042, 
        n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, 
        n2051, n2052, n2053, n2054, n2055, n2056, n2057, n2058, 
        n2075, n2110, n2111, n2112, n2113, n2114, n2115, n2116, 
        n2117, n2118, n2119, n2120, n2121, n2122, n2123, n2124, 
        n2125, n2141, n2142, n2143, n2144, n2145, n2146, n2147, 
        n2148, n2149, n2150, n2151, n2152, n2153, n2154, n2155, 
        n2156, n2157, n2158, n2174, n2209, n2210, n2211, n2212, 
        n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220, 
        n2221, n2222, n2223, n2224, n2225, n2240, n2241, n2242, 
        n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250, 
        n2251, n2252, n2253, n2254, n2255, n2256, n2257, n2258, 
        n2273, n2308, n2309, n2310, n2311, n2312, n2313, n2314, 
        n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322, 
        n2323, n2324, n2325, n2339, n2340, n2341, n2342, n2343, 
        n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351, 
        n2352, n2353, n2354, n2355, n2356, n2357, n2358, n2372, 
        n2407, n2408, n2409, n2410, n2411, n2412, n2413, n2414, 
        n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422, 
        n2423, n2424, n2425, n2438, n2439, n2440, n2441, n2442, 
        n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450, 
        n2451, n2452, n2453, n2454, n2455, n2456, n2457, n2458, 
        n2471, n2506, n2507, n2508, n2509, n2510, n2511, n2512, 
        n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520, 
        n2521, n2522, n2523, n2524, n2525, n2537, n2538, n2539, 
        n2540, n2541, n2542, n2543, n2544, n2545, n2546, n2547, 
        n2548, n2549, n2550, n2551, n2552, n2553, n2554, n2555, 
        n2556, n2557, n2558, n2570, n2605, n2606, n2607, n2608, 
        n2609, n2610, n2611, n2612, n2613, n2614, n2615, n2616, 
        n2617, n2618, n2619, n2620, n2621, n2622, n2623, n2624, 
        n2625, n2636, n2637, n2638, n2639, n2640, n2641, n2642, 
        n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650, 
        n2651, n2652, n2653, n2654, n2655, n2656, n2657, n2658, 
        n2669, n2735, n2736, n2737, n2738, n2739, n2740, n2741, 
        n2742, n2743, n2744, n2745, n2746, n2747, n2748, n2749, 
        n2750, n2751, n2752, n2753, n2754, n2755, n2756, n2757, 
        n2758, n2759, n2768, n2803, n2804, n2805, n2806, n2807, 
        n2808, n2809, n2810, n2811, n2812, n2813, n2814, n2815, 
        n2816, n2817, n2818, n2819, n2820, n2821, n2822, n2823, 
        n2824, n2825, n2834, n2835, n2836, n2837, n2838, n2839, 
        n2840, n2841, n2842, n2843, n2844, n2845, n2846, n2847, 
        n2848, n2849, n2850, n2851, n2852, n2853, n2854, n2855, 
        n2856, n2857, n2865, n2867, n2902, n2903, n2904, n2905, 
        n2906, n2907, n2908, n2909, n2910, n2911, n2912, n2913, 
        n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921, 
        n2922, n2923, n2924, n2925, n2933, n2934, n2935, n2936, 
        n2937, n2938, n2939, n2940, n2941, n2942, n2943, n2944, 
        n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952, 
        n2953, n2954, n2955, n2956, n2957, n2958_adj_4882, n2966, 
        n3001, n3002, n3003, n3004, n3005, n3006, n3007_adj_4883, 
        n3008, n3009, n3010, n3011, n3012, n3013, n3014, n3015, 
        n3016, n3017, n3018, n3019, n3020, n3021, n3022, n3023, 
        n3024, n3025, n3032, n3033, n3034, n3035, n3036, n3037, 
        n3038, n3039, n3040, n3041, n3042, n3043, n3044, n3045, 
        n3046, n3047, n3048, n3049, n3050, n3051, n3052, n3053, 
        n3054, n3055, n3056, n3057, n3058, n3065, n3100, n3101, 
        n3102, n3103, n3104, n3105, n3106, n3107, n3108, n3109, 
        n3110, n3111, n3112, n3113, n3114, n3115, n3116, n3117, 
        n3118, n3119, n3120, n3121, n3122, n3123, n3124, n3125, 
        n3131, n3132, n3133, n3134, n3135, n3136, n3137, n3138, 
        n3139, n3140, n3141, n3142, n3143, n3144, n3145, n3146, 
        n3147, n3148, n3149, n3150, n3151, n3152, n3153, n3154, 
        n3155, n3156, n3157, n3158, n3164_adj_4884, n3199, n3200, 
        n3201, n3202, n3203, n3204, n3205, n3206, n3207, n3208, 
        n3209_adj_4885, n3210_adj_4886, n3211_adj_4887, n3212_adj_4888, 
        n3213_adj_4889, n3214_adj_4890, n3215_adj_4891, n3216_adj_4892, 
        n3217_adj_4893, n3218_adj_4894, n3219_adj_4895, n3220_adj_4896, 
        n3221_adj_4897, n3222_adj_4898, n3223_adj_4899, n3224_adj_4900, 
        n3225_adj_4901, n3230_adj_4902, n3231_adj_4903, n3232_adj_4904, 
        n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240, 
        n3241, n3242, n3243, n3244, n3245, n3246, n3247, n3248, 
        n3249, n3250, n3251, n3252, n3253, n3254, n3255, n3256, 
        n3257, n3258, n3263, n3298, n3299, n3300, n3301, n3302, 
        n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310, 
        n3311, n3312, n3313, n3314, n3315, n3316, n3317, n3318, 
        n3319, n3320, n3321, n3322, n3323, n3324, n3325, n3330, 
        n3331, n3342, n3343, n3344, n3345, n3346, n3348, n3353, 
        n3354, n3355, n3356, n3357, n3358, n3362, n28361, n3452, 
        n3453, n3454, n3455, n3456, n3457, n3458, n38182, n38185, 
        n38188, n38191, n38194, n38197, n28049, n28244, n28651, 
        n28650, n28649, n18082, n28648, n28048, n28243, n28242, 
        n28241, n27892, n28047, n28046, n27891, n28_adj_4905, n27_adj_4906, 
        n26_adj_4907, n25_adj_4908, n28240, n28360, n28045, n28239, 
        n28044, n28647, n28359, n28358, n28238, n28043, n28646, 
        n28357, n28237, n28236, n28645, n28356, n28355, n28644, 
        n34021, n36177, n4_adj_4909, n28235, n27890, n28042, n28643, 
        n28041, n28642, n27889, n28354, n28353, n28352, n27888, 
        n28641, n10395, n10394, n10393, n10392, n10391, n10390, 
        n28040, n28640, n28639, n24_adj_4910, n22_adj_4911, n20_adj_4912, 
        n27887, n28638, n32957, n27886, n28637, n16_adj_4913, n28636, 
        n32941, n28635, n28351, n28234, n28233, n28232, n28634, 
        n28633, n33769, n28632, n32962, n28350, n28349, n28631, 
        n28231, n33930, n28630, n28230, n28629, n28348, n28347, 
        n28229, n28628, n34970, n28346, n28345, n28228, n33960, 
        n28344, n28627, n28343, n36067, n28342, n28341, n28340, 
        n28626, n27885, n33901, n28339, n28227, n28625, n28624, 
        n28623, n33701, n28226, n28225, n22_adj_4914, n28224, n28622, 
        n37263, n37262, n19_adj_4915, n37261, n37260, n18_adj_4916, 
        n28338, n28337, n28336, n27884, n28621, n33657, n15_adj_4917, 
        n28223, n28620, n34_adj_4918, n28222, n31_adj_4919, n30_adj_4920, 
        n28_adj_4921, n28619, n36011, n22_adj_4922, n1_adj_4923, n21_adj_4924, 
        n28618, n18089, n28221, n25050, n1_adj_4925, n13_adj_4926, 
        n11_adj_4927, n28617, n27883, n33970, n27882, n28616, n27881, 
        n28335, n28334, n27880, n28220, n27879, n28615, n28614, 
        n28613, n28612, n27878, n28611, n37252, n33898, n28333, 
        n28610, n28332, n28609, n28219, n27877, n27876, n18088, 
        n28331, n35933, n28218, n1_adj_4928, n1_adj_4929, n1_adj_4930, 
        n1_adj_4931, n1_adj_4932, n1_adj_4933, n1_adj_4934, n1_adj_4935, 
        n1_adj_4936, n1_adj_4937, n1_adj_4938, n1_adj_4939, n1_adj_4940, 
        n1_adj_4941, n1_adj_4942, n1_adj_4943, n1_adj_4944, n1_adj_4945, 
        n1_adj_4946, n1_adj_4947, n1_adj_4948, n1_adj_4949, n1_adj_4950, 
        n18150, n35917, n35913, n28608, n28607, n2_adj_4951, n3_adj_4952, 
        n4_adj_4953, n5_adj_4954, n6_adj_4955, n7_adj_4956, n8_adj_4957, 
        n9_adj_4958, n10_adj_4959, n11_adj_4960, n12_adj_4961, n13_adj_4962, 
        n14_adj_4963, n15_adj_4964, n16_adj_4965, n17_adj_4966, n18_adj_4967, 
        n19_adj_4968, n20_adj_4969, n21_adj_4970, n22_adj_4971, n23_adj_4972, 
        n24_adj_4973, n25_adj_4974, n26_adj_4975, n27_adj_4976, n28_adj_4977, 
        n29_adj_4978, n30_adj_4979, n31_adj_4980, n32_adj_4981, n33_adj_4982, 
        n37251, n28330, n28606, n28329, n35869, n35867, n28217, 
        n35865, n36494, n28216, n35863, n35861, n35859, n35857, 
        n37245, n35855, n37244, n18149, n37243, n34007, n35853, 
        n35851, n28605, n12_adj_4983, n6_adj_4984, n18151, n8_adj_4985, 
        n7_adj_4986, n6_adj_4987, n18087, n28_adj_4988, n26_adj_4989, 
        n24_adj_4990, n20_adj_4991, n19_adj_4992, n37241, n16_adj_4993, 
        n18_adj_4994, n16_adj_4995, n35849, n35845, n35843, n38508, 
        n35837, n35835, n35833, n35831, n35829, n34206, n33942, 
        n34066, n36410, n18086, n28328, n28327, n28215, n28214, 
        n5_adj_4996, n33989, n18_adj_4997, n34042, n27875, n28604, 
        n16_adj_4998, n28326, n28325, n28603, n34919, n28213, n13_adj_4999, 
        n33877, n28212, n28602, n25070, n33871, n28211, n28324, 
        n28210, n28323, n28209, n28208, n28601, n28207, n28322, 
        n28321, n28206, n6_adj_5000, n37232, n28205, n28320, n28600, 
        n33867, n28599, n28319, n18085, n17546, n28318, n28317, 
        n28204, n28316, n28203, n28315, n28598, n28597, n28596, 
        n28314, n29597, n28202, n28595, n32973, n25112, n37231, 
        n29598, n28594, n34971, n29599, n37230, n37229, n28201, 
        n28593, n37228, n28200, n37227, n28199, n28592, n28198, 
        n28591, n28197, n28196, n28590, n28589, n33909, n37226, 
        n28195, n28588, n16_adj_5001, n11_adj_5002, n37225, n28587, 
        n10_adj_5003, n18084, n28434, n28433, n28432, n35088, n28194, 
        n18083, n28193, n28586, n36391, n28431, n28192, n28430, 
        n28585, n28584, n28583, n28582, n16148, n28429, n28428, 
        n28581, n35492, n28427, n28426, n28580, n28579, n28578, 
        n37224;
    
    VCC i2 (.Y(VCC_net));
    SB_DFF pwm_setpoint_i0 (.Q(pwm_setpoint[0]), .C(clk32MHz), .D(pwm_setpoint_22__N_57[0]));   // verilog/TinyFPGA_B.v(139[10] 152[6])
    SB_DFF h2_68 (.Q(PIN_21_c), .C(clk32MHz), .D(hall2));   // verilog/TinyFPGA_B.v(139[10] 152[6])
    SB_DFF displacement_i0 (.Q(displacement[0]), .C(clk32MHz), .D(displacement_23__N_80[0]));   // verilog/TinyFPGA_B.v(247[10] 249[6])
    SB_IO hall2_input (.PACKAGE_PIN(PIN_4), .LATCH_INPUT_VALUE(GND_net), 
          .INPUT_CLK(GND_net), .OUTPUT_CLK(GND_net), .OUTPUT_ENABLE(GND_net), 
          .D_OUT_1(GND_net), .D_OUT_0(GND_net), .D_IN_0(hall2)) /* synthesis lattice_noprune=1, syn_instantiated=1 */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam hall2_input.PIN_TYPE = 6'b000001;
    defparam hall2_input.PULLUP = 1'b1;
    defparam hall2_input.NEG_TRIGGER = 1'b0;
    defparam hall2_input.IO_STANDARD = "SB_LVCMOS";
    SB_IO hall3_input (.PACKAGE_PIN(PIN_5), .LATCH_INPUT_VALUE(GND_net), 
          .INPUT_CLK(GND_net), .OUTPUT_CLK(GND_net), .OUTPUT_ENABLE(GND_net), 
          .D_OUT_1(GND_net), .D_OUT_0(GND_net), .D_IN_0(hall3)) /* synthesis lattice_noprune=1, syn_instantiated=1 */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam hall3_input.PIN_TYPE = 6'b000001;
    defparam hall3_input.PULLUP = 1'b1;
    defparam hall3_input.NEG_TRIGGER = 1'b0;
    defparam hall3_input.IO_STANDARD = "SB_LVCMOS";
    SB_IO tx_output (.PACKAGE_PIN(PIN_12), .LATCH_INPUT_VALUE(GND_net), 
          .INPUT_CLK(GND_net), .OUTPUT_CLK(GND_net), .OUTPUT_ENABLE(tx_enable), 
          .D_OUT_1(GND_net), .D_OUT_0(tx_o)) /* synthesis lattice_noprune=1, syn_instantiated=1 */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam tx_output.PIN_TYPE = 6'b101001;
    defparam tx_output.PULLUP = 1'b1;
    defparam tx_output.NEG_TRIGGER = 1'b0;
    defparam tx_output.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 i13439_3_lut (.I0(\half_duty[0] [4]), .I1(half_duty_new[4]), 
            .I2(n1466), .I3(GND_net), .O(n18268));   // vhdl/pwm.vhd(59[5] 95[12])
    defparam i13439_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF h3_69 (.Q(PIN_22_c), .C(clk32MHz), .D(hall3));   // verilog/TinyFPGA_B.v(139[10] 152[6])
    SB_DFF dir_73 (.Q(PIN_23_c), .C(clk32MHz), .D(duty[23]));   // verilog/TinyFPGA_B.v(139[10] 152[6])
    neopixel nx (.\neo_pixel_transmitter.done (\neo_pixel_transmitter.done ), 
            .clk32MHz(clk32MHz), .n31521(n31521), .VCC_net(VCC_net), .bit_ctr({bit_ctr}), 
            .\neo_pixel_transmitter.t0 ({\neo_pixel_transmitter.t0 }), .GND_net(GND_net), 
            .timer({timer}), .n37232(n37232), .n1(n1), .n37224(n37224), 
            .\state[0] (state[0]), .n7(n7_adj_4803), .n4(n4), .\state[1] (state[1]), 
            .n17229(n17229), .n35088(n35088), .n17500(n17500), .n17567(n17567), 
            .n37244(n37244), .n37260(n37260), .start(start), .\state_3__N_462[1] (state_3__N_462[1]), 
            .n5(n5_adj_4996), .n1460(n1460), .n33701(n33701), .n37261(n37261), 
            .n37225(n37225), .n37262(n37262), .n20(n20), .n37226(n37226), 
            .n37263(n37263), .n37304(n37304), .\color[10] (color[10]), 
            .\color[11] (color[11]), .\color[12] (color[12]), .\color[9] (color[9]), 
            .n37308(n37308), .n37309(n37309), .n37330(n37330), .PIN_8_c(PIN_8_c), 
            .n37251(n37251), .n17546(n17546), .n17767(n17767), .n17766(n17766), 
            .n17765(n17765), .n17764(n17764), .n17763(n17763), .n17762(n17762), 
            .n17761(n17761), .n17760(n17760), .n17759(n17759), .n17758(n17758), 
            .n17757(n17757), .n17756(n17756), .n17755(n17755), .n17754(n17754), 
            .n17753(n17753), .n17752(n17752), .n17751(n17751), .n17750(n17750), 
            .n17749(n17749), .n17748(n17748), .n17747(n17747), .n17746(n17746), 
            .n17745(n17745), .n17744(n17744), .n17743(n17743), .n17742(n17742), 
            .n17741(n17741), .n17740(n17740), .n17739(n17739), .n17738(n17738), 
            .n17737(n17737), .n37335(n37335), .n37227(n37227), .n37359(n37359), 
            .n37360(n37360), .n37241(n37241), .n37228(n37228), .n37361(n37361), 
            .n37362(n37362), .n37229(n37229), .n37230(n37230), .n37245(n37245), 
            .n37363(n37363), .n37364(n37364), .n31591(n31591), .n31589(n31589), 
            .n31587(n31587), .n31585(n31585), .n37252(n37252), .n31583(n31583), 
            .n31577(n31577), .n37365(n37365), .n31575(n31575), .n31573(n31573), 
            .n31571(n31571), .n31569(n31569), .n31567(n31567), .n31565(n31565), 
            .n31563(n31563), .n31561(n31561), .n31559(n31559), .n31557(n31557), 
            .n37368(n37368), .n31555(n31555), .n31553(n31553), .n31551(n31551), 
            .n31549(n31549), .n31547(n31547), .n31545(n31545), .n31543(n31543), 
            .n31541(n31541), .n31539(n31539), .n31537(n31537), .n31535(n31535), 
            .n31533(n31533), .n31531(n31531), .n31529(n31529), .n31527(n31527), 
            .n31599(n31599), .n37231(n37231), .n37369(n37369)) /* synthesis lattice_noprune=1, syn_preserve=0, syn_module_defined=1, syn_noprune=0 */ ;   // verilog/TinyFPGA_B.v(76[10] 82[2])
    SB_IO hall1_input (.PACKAGE_PIN(PIN_3), .LATCH_INPUT_VALUE(GND_net), 
          .INPUT_CLK(GND_net), .OUTPUT_CLK(GND_net), .OUTPUT_ENABLE(GND_net), 
          .D_OUT_1(GND_net), .D_OUT_0(GND_net), .D_IN_0(hall1)) /* synthesis lattice_noprune=1, syn_instantiated=1 */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam hall1_input.PIN_TYPE = 6'b000001;
    defparam hall1_input.PULLUP = 1'b1;
    defparam hall1_input.NEG_TRIGGER = 1'b0;
    defparam hall1_input.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 rem_4_add_1586_13_lut (.I0(GND_net), .I1(n2347), .I2(VCC_net), 
            .I3(n28188), .O(n2414)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1586_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1787_11 (.CI(n27883), .I0(n2649), .I1(n2669), .CO(n27884));
    SB_LUT4 rem_4_add_1720_9_lut (.I0(GND_net), .I1(n2551), .I2(VCC_net), 
            .I3(n28051), .O(n2618)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1720_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i30693_2_lut (.I0(state_3__N_462[1]), .I1(state[1]), .I2(GND_net), 
            .I3(GND_net), .O(n37243));   // verilog/neopixel.v(35[12] 117[6])
    defparam i30693_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY rem_4_add_1586_13 (.CI(n28188), .I0(n2347), .I1(VCC_net), 
            .CO(n28189));
    SB_LUT4 rem_4_add_1586_12_lut (.I0(GND_net), .I1(n2348), .I2(VCC_net), 
            .I3(n28187), .O(n2415)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1586_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1787_10_lut (.I0(n2650), .I1(n2650), .I2(n2669), 
            .I3(n27882), .O(n2749)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1787_10_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY rem_4_add_1720_9 (.CI(n28051), .I0(n2551), .I1(VCC_net), 
            .CO(n28052));
    SB_CARRY rem_4_add_1586_12 (.CI(n28187), .I0(n2348), .I1(VCC_net), 
            .CO(n28188));
    SB_LUT4 rem_4_add_1720_8_lut (.I0(GND_net), .I1(n2552), .I2(VCC_net), 
            .I3(n28050), .O(n2619)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1720_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1586_11_lut (.I0(GND_net), .I1(n2349), .I2(VCC_net), 
            .I3(n28186), .O(n2416)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1586_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1586_11 (.CI(n28186), .I0(n2349), .I1(VCC_net), 
            .CO(n28187));
    SB_LUT4 rem_4_add_1586_10_lut (.I0(GND_net), .I1(n2350), .I2(VCC_net), 
            .I3(n28185), .O(n2417)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1586_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1720_8 (.CI(n28050), .I0(n2552), .I1(VCC_net), 
            .CO(n28051));
    SB_CARRY rem_4_add_1787_10 (.CI(n27882), .I0(n2650), .I1(n2669), .CO(n27883));
    SB_CARRY rem_4_add_1586_10 (.CI(n28185), .I0(n2350), .I1(VCC_net), 
            .CO(n28186));
    SB_LUT4 rem_4_add_1720_7_lut (.I0(GND_net), .I1(n2553), .I2(VCC_net), 
            .I3(n28049), .O(n2620)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1720_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1586_9_lut (.I0(GND_net), .I1(n2351), .I2(VCC_net), 
            .I3(n28184), .O(n2418)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1586_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1720_7 (.CI(n28049), .I0(n2553), .I1(VCC_net), 
            .CO(n28050));
    SB_CARRY rem_4_add_1586_9 (.CI(n28184), .I0(n2351), .I1(VCC_net), 
            .CO(n28185));
    SB_LUT4 rem_4_add_1787_9_lut (.I0(n2651), .I1(n2651), .I2(n2669), 
            .I3(n27881), .O(n2750)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1787_9_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 rem_4_add_1586_8_lut (.I0(GND_net), .I1(n2352), .I2(VCC_net), 
            .I3(n28183), .O(n2419)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1586_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i27_4_lut (.I0(n1460), .I1(n37243), .I2(state[0]), .I3(n5_adj_4996), 
            .O(n1));   // verilog/neopixel.v(35[12] 117[6])
    defparam i27_4_lut.LUT_INIT = 16'h3505;
    SB_LUT4 i12947_3_lut (.I0(IntegralLimit[9]), .I1(\data_in_frame[12] [1]), 
            .I2(n5439), .I3(GND_net), .O(n17776));   // verilog/coms.v(126[12] 293[6])
    defparam i12947_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13016_3_lut (.I0(Ki[9]), .I1(\data_in_frame[4] [1]), .I2(n34066), 
            .I3(GND_net), .O(n17845));   // verilog/coms.v(126[12] 293[6])
    defparam i13016_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13017_3_lut (.I0(Ki[10]), .I1(\data_in_frame[4] [2]), .I2(n34066), 
            .I3(GND_net), .O(n17846));   // verilog/coms.v(126[12] 293[6])
    defparam i13017_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13018_3_lut (.I0(Ki[11]), .I1(\data_in_frame[4] [3]), .I2(n34066), 
            .I3(GND_net), .O(n17847));   // verilog/coms.v(126[12] 293[6])
    defparam i13018_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12948_3_lut (.I0(IntegralLimit[10]), .I1(\data_in_frame[12] [2]), 
            .I2(n5439), .I3(GND_net), .O(n17777));   // verilog/coms.v(126[12] 293[6])
    defparam i12948_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13019_3_lut (.I0(Ki[12]), .I1(\data_in_frame[4] [4]), .I2(n34066), 
            .I3(GND_net), .O(n17848));   // verilog/coms.v(126[12] 293[6])
    defparam i13019_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13020_3_lut (.I0(Ki[13]), .I1(\data_in_frame[4] [5]), .I2(n34066), 
            .I3(GND_net), .O(n17849));   // verilog/coms.v(126[12] 293[6])
    defparam i13020_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13021_3_lut (.I0(Ki[14]), .I1(\data_in_frame[4] [6]), .I2(n34066), 
            .I3(GND_net), .O(n17850));   // verilog/coms.v(126[12] 293[6])
    defparam i13021_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY rem_4_add_1586_8 (.CI(n28183), .I0(n2352), .I1(VCC_net), 
            .CO(n28184));
    SB_LUT4 i13022_3_lut (.I0(Ki[15]), .I1(\data_in_frame[4] [7]), .I2(n34066), 
            .I3(GND_net), .O(n17851));   // verilog/coms.v(126[12] 293[6])
    defparam i13022_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13023_3_lut (.I0(setpoint[1]), .I1(n4997), .I2(n35492), .I3(GND_net), 
            .O(n17852));   // verilog/coms.v(126[12] 293[6])
    defparam i13023_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13024_3_lut (.I0(setpoint[2]), .I1(n4998), .I2(n35492), .I3(GND_net), 
            .O(n17853));   // verilog/coms.v(126[12] 293[6])
    defparam i13024_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13025_3_lut (.I0(setpoint[3]), .I1(n4999), .I2(n35492), .I3(GND_net), 
            .O(n17854));   // verilog/coms.v(126[12] 293[6])
    defparam i13025_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13026_3_lut (.I0(setpoint[4]), .I1(n5000), .I2(n35492), .I3(GND_net), 
            .O(n17855));   // verilog/coms.v(126[12] 293[6])
    defparam i13026_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13027_3_lut (.I0(setpoint[5]), .I1(n5001), .I2(n35492), .I3(GND_net), 
            .O(n17856));   // verilog/coms.v(126[12] 293[6])
    defparam i13027_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13028_3_lut (.I0(setpoint[6]), .I1(n5002), .I2(n35492), .I3(GND_net), 
            .O(n17857));   // verilog/coms.v(126[12] 293[6])
    defparam i13028_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13029_3_lut (.I0(setpoint[7]), .I1(n5003), .I2(n35492), .I3(GND_net), 
            .O(n17858));   // verilog/coms.v(126[12] 293[6])
    defparam i13029_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 unary_minus_28_inv_0_i23_1_lut (.I0(duty[22]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n3));   // verilog/TinyFPGA_B.v(149[23:28])
    defparam unary_minus_28_inv_0_i23_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i13030_3_lut (.I0(setpoint[8]), .I1(n5004), .I2(n35492), .I3(GND_net), 
            .O(n17859));   // verilog/coms.v(126[12] 293[6])
    defparam i13030_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13031_3_lut (.I0(setpoint[9]), .I1(n5005), .I2(n35492), .I3(GND_net), 
            .O(n17860));   // verilog/coms.v(126[12] 293[6])
    defparam i13031_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13032_3_lut (.I0(setpoint[10]), .I1(n5006), .I2(n35492), 
            .I3(GND_net), .O(n17861));   // verilog/coms.v(126[12] 293[6])
    defparam i13032_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13033_3_lut (.I0(setpoint[11]), .I1(n5007), .I2(n35492), 
            .I3(GND_net), .O(n17862));   // verilog/coms.v(126[12] 293[6])
    defparam i13033_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13034_3_lut (.I0(setpoint[12]), .I1(n5008), .I2(n35492), 
            .I3(GND_net), .O(n17863));   // verilog/coms.v(126[12] 293[6])
    defparam i13034_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13035_3_lut (.I0(setpoint[13]), .I1(n5009), .I2(n35492), 
            .I3(GND_net), .O(n17864));   // verilog/coms.v(126[12] 293[6])
    defparam i13035_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13036_3_lut (.I0(setpoint[14]), .I1(n5010), .I2(n35492), 
            .I3(GND_net), .O(n17865));   // verilog/coms.v(126[12] 293[6])
    defparam i13036_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13037_3_lut (.I0(setpoint[15]), .I1(n5011), .I2(n35492), 
            .I3(GND_net), .O(n17866));   // verilog/coms.v(126[12] 293[6])
    defparam i13037_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13038_3_lut (.I0(setpoint[16]), .I1(n5012), .I2(n35492), 
            .I3(GND_net), .O(n17867));   // verilog/coms.v(126[12] 293[6])
    defparam i13038_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13039_3_lut (.I0(setpoint[17]), .I1(n5013), .I2(n35492), 
            .I3(GND_net), .O(n17868));   // verilog/coms.v(126[12] 293[6])
    defparam i13039_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13040_3_lut (.I0(setpoint[18]), .I1(n5014), .I2(n35492), 
            .I3(GND_net), .O(n17869));   // verilog/coms.v(126[12] 293[6])
    defparam i13040_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 rem_4_add_1586_7_lut (.I0(GND_net), .I1(n2353), .I2(VCC_net), 
            .I3(n28182), .O(n2420)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1586_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1720_6_lut (.I0(GND_net), .I1(n2554), .I2(GND_net), 
            .I3(n28048), .O(n2621)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1720_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i13041_3_lut (.I0(setpoint[19]), .I1(n5015), .I2(n35492), 
            .I3(GND_net), .O(n17870));   // verilog/coms.v(126[12] 293[6])
    defparam i13041_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13042_3_lut (.I0(setpoint[20]), .I1(n5016), .I2(n35492), 
            .I3(GND_net), .O(n17871));   // verilog/coms.v(126[12] 293[6])
    defparam i13042_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13043_3_lut (.I0(setpoint[21]), .I1(n5017), .I2(n35492), 
            .I3(GND_net), .O(n17872));   // verilog/coms.v(126[12] 293[6])
    defparam i13043_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13044_3_lut (.I0(setpoint[22]), .I1(n5018), .I2(n35492), 
            .I3(GND_net), .O(n17873));   // verilog/coms.v(126[12] 293[6])
    defparam i13044_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY rem_4_add_1720_6 (.CI(n28048), .I0(n2554), .I1(GND_net), 
            .CO(n28049));
    SB_CARRY rem_4_add_1586_7 (.CI(n28182), .I0(n2353), .I1(VCC_net), 
            .CO(n28183));
    SB_LUT4 i1_3_lut (.I0(start), .I1(\neo_pixel_transmitter.done ), .I2(n7_adj_4803), 
            .I3(GND_net), .O(n4));   // verilog/neopixel.v(35[12] 117[6])
    defparam i1_3_lut.LUT_INIT = 16'h4040;
    SB_LUT4 i12738_4_lut (.I0(n17500), .I1(state[1]), .I2(state_3__N_462[1]), 
            .I3(n17229), .O(n17567));   // verilog/neopixel.v(35[12] 117[6])
    defparam i12738_4_lut.LUT_INIT = 16'hfaee;
    SB_LUT4 unary_minus_28_inv_0_i1_1_lut (.I0(duty[0]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n25_adj_4775));   // verilog/TinyFPGA_B.v(149[23:28])
    defparam unary_minus_28_inv_0_i1_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i13045_3_lut (.I0(setpoint[23]), .I1(n5019), .I2(n35492), 
            .I3(GND_net), .O(n17874));   // verilog/coms.v(126[12] 293[6])
    defparam i13045_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13046_3_lut (.I0(\data_out_frame[5] [0]), .I1(control_mode[0]), 
            .I2(n13724), .I3(GND_net), .O(n17875));   // verilog/coms.v(126[12] 293[6])
    defparam i13046_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13047_3_lut (.I0(\data_out_frame[5] [1]), .I1(control_mode[1]), 
            .I2(n13724), .I3(GND_net), .O(n17876));   // verilog/coms.v(126[12] 293[6])
    defparam i13047_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13048_3_lut (.I0(\data_out_frame[5] [2]), .I1(control_mode[2]), 
            .I2(n13724), .I3(GND_net), .O(n17877));   // verilog/coms.v(126[12] 293[6])
    defparam i13048_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13049_3_lut (.I0(\data_out_frame[5] [3]), .I1(control_mode[3]), 
            .I2(n13724), .I3(GND_net), .O(n17878));   // verilog/coms.v(126[12] 293[6])
    defparam i13049_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13191_3_lut (.I0(\data_in_frame[1] [2]), .I1(rx_data[2]), .I2(n32962), 
            .I3(GND_net), .O(n18020));   // verilog/coms.v(126[12] 293[6])
    defparam i13191_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13192_3_lut (.I0(\data_in_frame[1] [3]), .I1(rx_data[3]), .I2(n32962), 
            .I3(GND_net), .O(n18021));   // verilog/coms.v(126[12] 293[6])
    defparam i13192_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13193_3_lut (.I0(\data_in_frame[1] [4]), .I1(rx_data[4]), .I2(n32962), 
            .I3(GND_net), .O(n18022));   // verilog/coms.v(126[12] 293[6])
    defparam i13193_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13194_3_lut (.I0(\data_in_frame[1] [5]), .I1(rx_data[5]), .I2(n32962), 
            .I3(GND_net), .O(n18023));   // verilog/coms.v(126[12] 293[6])
    defparam i13194_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13050_3_lut (.I0(\data_out_frame[5] [4]), .I1(control_mode[4]), 
            .I2(n13724), .I3(GND_net), .O(n17879));   // verilog/coms.v(126[12] 293[6])
    defparam i13050_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13051_3_lut (.I0(\data_out_frame[5] [5]), .I1(control_mode[5]), 
            .I2(n13724), .I3(GND_net), .O(n17880));   // verilog/coms.v(126[12] 293[6])
    defparam i13051_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 unary_minus_28_inv_0_i8_1_lut (.I0(duty[7]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n18));   // verilog/TinyFPGA_B.v(149[23:28])
    defparam unary_minus_28_inv_0_i8_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 rem_4_unary_minus_2_inv_0_i1_1_lut (.I0(communication_counter[0]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n33_adj_4982));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_unary_minus_2_inv_0_i1_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i13195_3_lut (.I0(\data_in_frame[1] [6]), .I1(rx_data[6]), .I2(n32962), 
            .I3(GND_net), .O(n18024));   // verilog/coms.v(126[12] 293[6])
    defparam i13195_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 rem_4_unary_minus_2_inv_0_i2_1_lut (.I0(communication_counter[1]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n32_adj_4981));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_unary_minus_2_inv_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i13196_3_lut (.I0(\data_in_frame[1] [7]), .I1(rx_data[7]), .I2(n32962), 
            .I3(GND_net), .O(n18025));   // verilog/coms.v(126[12] 293[6])
    defparam i13196_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 rem_4_unary_minus_2_inv_0_i3_1_lut (.I0(communication_counter[2]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n31_adj_4980));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_unary_minus_2_inv_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i13052_3_lut (.I0(\data_out_frame[5] [6]), .I1(control_mode[6]), 
            .I2(n13724), .I3(GND_net), .O(n17881));   // verilog/coms.v(126[12] 293[6])
    defparam i13052_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13053_3_lut (.I0(\data_out_frame[5] [7]), .I1(control_mode[7]), 
            .I2(n13724), .I3(GND_net), .O(n17882));   // verilog/coms.v(126[12] 293[6])
    defparam i13053_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13054_3_lut (.I0(\data_out_frame[6] [0]), .I1(encoder0_position[16]), 
            .I2(n13724), .I3(GND_net), .O(n17883));   // verilog/coms.v(126[12] 293[6])
    defparam i13054_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i30835_2_lut (.I0(displacement[0]), .I1(control_mode[0]), .I2(GND_net), 
            .I3(GND_net), .O(n37310));   // verilog/TinyFPGA_B.v(210[5] 214[10])
    defparam i30835_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 unary_minus_28_inv_0_i9_1_lut (.I0(duty[8]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n17));   // verilog/TinyFPGA_B.v(149[23:28])
    defparam unary_minus_28_inv_0_i9_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mux_843_Mux_0_i1_3_lut (.I0(encoder0_position[0]), .I1(encoder1_position[0]), 
            .I2(control_mode[0]), .I3(GND_net), .O(n1_adj_4925));   // verilog/TinyFPGA_B.v(210[5] 214[10])
    defparam mux_843_Mux_0_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13055_3_lut (.I0(\data_out_frame[6] [1]), .I1(encoder0_position[17]), 
            .I2(n13724), .I3(GND_net), .O(n17884));   // verilog/coms.v(126[12] 293[6])
    defparam i13055_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13056_3_lut (.I0(\data_out_frame[6] [2]), .I1(encoder0_position[18]), 
            .I2(n13724), .I3(GND_net), .O(n17885));   // verilog/coms.v(126[12] 293[6])
    defparam i13056_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i19339_4_lut (.I0(n1_adj_4925), .I1(n34919), .I2(n37310), 
            .I3(control_mode[1]), .O(motor_state[0]));   // verilog/TinyFPGA_B.v(210[5] 214[10])
    defparam i19339_4_lut.LUT_INIT = 16'h3022;
    SB_LUT4 unary_minus_28_inv_0_i10_1_lut (.I0(duty[9]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n16));   // verilog/TinyFPGA_B.v(149[23:28])
    defparam unary_minus_28_inv_0_i10_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_28_inv_0_i11_1_lut (.I0(duty[10]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n15));   // verilog/TinyFPGA_B.v(149[23:28])
    defparam unary_minus_28_inv_0_i11_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i30960_2_lut (.I0(displacement[1]), .I1(control_mode[0]), .I2(GND_net), 
            .I3(GND_net), .O(n37336));   // verilog/TinyFPGA_B.v(210[5] 214[10])
    defparam i30960_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 rem_4_add_1586_6_lut (.I0(GND_net), .I1(n2354), .I2(GND_net), 
            .I3(n28181), .O(n2421)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1586_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mux_843_Mux_1_i1_3_lut (.I0(encoder0_position[1]), .I1(encoder1_position[1]), 
            .I2(control_mode[0]), .I3(GND_net), .O(n1_adj_4928));   // verilog/TinyFPGA_B.v(210[5] 214[10])
    defparam mux_843_Mux_1_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i19540_4_lut (.I0(n1_adj_4928), .I1(n34919), .I2(n37336), 
            .I3(control_mode[1]), .O(motor_state[1]));   // verilog/TinyFPGA_B.v(210[5] 214[10])
    defparam i19540_4_lut.LUT_INIT = 16'h3022;
    SB_LUT4 i13057_3_lut (.I0(\data_out_frame[6] [3]), .I1(encoder0_position[19]), 
            .I2(n13724), .I3(GND_net), .O(n17886));   // verilog/coms.v(126[12] 293[6])
    defparam i13057_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 unary_minus_28_inv_0_i12_1_lut (.I0(duty[11]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n14));   // verilog/TinyFPGA_B.v(149[23:28])
    defparam unary_minus_28_inv_0_i12_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i30888_2_lut (.I0(displacement[2]), .I1(control_mode[0]), .I2(GND_net), 
            .I3(GND_net), .O(n37337));   // verilog/TinyFPGA_B.v(210[5] 214[10])
    defparam i30888_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 mux_843_Mux_2_i1_3_lut (.I0(encoder0_position[2]), .I1(encoder1_position[2]), 
            .I2(control_mode[0]), .I3(GND_net), .O(n1_adj_4929));   // verilog/TinyFPGA_B.v(210[5] 214[10])
    defparam mux_843_Mux_2_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13058_3_lut (.I0(\data_out_frame[6] [4]), .I1(encoder0_position[20]), 
            .I2(n13724), .I3(GND_net), .O(n17887));   // verilog/coms.v(126[12] 293[6])
    defparam i13058_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13059_3_lut (.I0(\data_out_frame[6] [5]), .I1(encoder0_position[21]), 
            .I2(n13724), .I3(GND_net), .O(n17888));   // verilog/coms.v(126[12] 293[6])
    defparam i13059_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i19541_4_lut (.I0(n1_adj_4929), .I1(n34919), .I2(n37337), 
            .I3(control_mode[1]), .O(motor_state[2]));   // verilog/TinyFPGA_B.v(210[5] 214[10])
    defparam i19541_4_lut.LUT_INIT = 16'h3022;
    SB_LUT4 i13060_3_lut (.I0(\data_out_frame[6] [6]), .I1(encoder0_position[22]), 
            .I2(n13724), .I3(GND_net), .O(n17889));   // verilog/coms.v(126[12] 293[6])
    defparam i13060_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13061_3_lut (.I0(\data_out_frame[6] [7]), .I1(encoder0_position[23]), 
            .I2(n13724), .I3(GND_net), .O(n17890));   // verilog/coms.v(126[12] 293[6])
    defparam i13061_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12949_3_lut (.I0(IntegralLimit[11]), .I1(\data_in_frame[12] [3]), 
            .I2(n5439), .I3(GND_net), .O(n17778));   // verilog/coms.v(126[12] 293[6])
    defparam i12949_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12950_3_lut (.I0(IntegralLimit[12]), .I1(\data_in_frame[12] [4]), 
            .I2(n5439), .I3(GND_net), .O(n17779));   // verilog/coms.v(126[12] 293[6])
    defparam i12950_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13062_3_lut (.I0(\data_out_frame[7] [0]), .I1(encoder0_position[8]), 
            .I2(n13724), .I3(GND_net), .O(n17891));   // verilog/coms.v(126[12] 293[6])
    defparam i13062_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13063_3_lut (.I0(\data_out_frame[7] [1]), .I1(encoder0_position[9]), 
            .I2(n13724), .I3(GND_net), .O(n17892));   // verilog/coms.v(126[12] 293[6])
    defparam i13063_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13064_3_lut (.I0(\data_out_frame[7] [2]), .I1(encoder0_position[10]), 
            .I2(n13724), .I3(GND_net), .O(n17893));   // verilog/coms.v(126[12] 293[6])
    defparam i13064_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13065_3_lut (.I0(\data_out_frame[7] [3]), .I1(encoder0_position[11]), 
            .I2(n13724), .I3(GND_net), .O(n17894));   // verilog/coms.v(126[12] 293[6])
    defparam i13065_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13066_3_lut (.I0(\data_out_frame[7] [4]), .I1(encoder0_position[12]), 
            .I2(n13724), .I3(GND_net), .O(n17895));   // verilog/coms.v(126[12] 293[6])
    defparam i13066_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13067_3_lut (.I0(\data_out_frame[7] [5]), .I1(encoder0_position[13]), 
            .I2(n13724), .I3(GND_net), .O(n17896));   // verilog/coms.v(126[12] 293[6])
    defparam i13067_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12951_3_lut (.I0(IntegralLimit[13]), .I1(\data_in_frame[12] [5]), 
            .I2(n5439), .I3(GND_net), .O(n17780));   // verilog/coms.v(126[12] 293[6])
    defparam i12951_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12952_3_lut (.I0(IntegralLimit[14]), .I1(\data_in_frame[12] [6]), 
            .I2(n5439), .I3(GND_net), .O(n17781));   // verilog/coms.v(126[12] 293[6])
    defparam i12952_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12953_3_lut (.I0(IntegralLimit[15]), .I1(\data_in_frame[12] [7]), 
            .I2(n5439), .I3(GND_net), .O(n17782));   // verilog/coms.v(126[12] 293[6])
    defparam i12953_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13068_3_lut (.I0(\data_out_frame[7] [6]), .I1(encoder0_position[14]), 
            .I2(n13724), .I3(GND_net), .O(n17897));   // verilog/coms.v(126[12] 293[6])
    defparam i13068_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i30895_2_lut (.I0(displacement[3]), .I1(control_mode[0]), .I2(GND_net), 
            .I3(GND_net), .O(n37338));   // verilog/TinyFPGA_B.v(210[5] 214[10])
    defparam i30895_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i13069_3_lut (.I0(\data_out_frame[7] [7]), .I1(encoder0_position[15]), 
            .I2(n13724), .I3(GND_net), .O(n17898));   // verilog/coms.v(126[12] 293[6])
    defparam i13069_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13070_3_lut (.I0(\data_out_frame[8] [0]), .I1(encoder0_position[0]), 
            .I2(n13724), .I3(GND_net), .O(n17899));   // verilog/coms.v(126[12] 293[6])
    defparam i13070_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13071_3_lut (.I0(\data_out_frame[8] [1]), .I1(encoder0_position[1]), 
            .I2(n13724), .I3(GND_net), .O(n17900));   // verilog/coms.v(126[12] 293[6])
    defparam i13071_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13072_3_lut (.I0(\data_out_frame[8] [2]), .I1(encoder0_position[2]), 
            .I2(n13724), .I3(GND_net), .O(n17901));   // verilog/coms.v(126[12] 293[6])
    defparam i13072_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_843_Mux_3_i1_3_lut (.I0(encoder0_position[3]), .I1(encoder1_position[3]), 
            .I2(control_mode[0]), .I3(GND_net), .O(n1_adj_4930));   // verilog/TinyFPGA_B.v(210[5] 214[10])
    defparam mux_843_Mux_3_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13073_3_lut (.I0(\data_out_frame[8] [3]), .I1(encoder0_position[3]), 
            .I2(n13724), .I3(GND_net), .O(n17902));   // verilog/coms.v(126[12] 293[6])
    defparam i13073_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i19542_4_lut (.I0(n1_adj_4930), .I1(n34919), .I2(n37338), 
            .I3(control_mode[1]), .O(motor_state[3]));   // verilog/TinyFPGA_B.v(210[5] 214[10])
    defparam i19542_4_lut.LUT_INIT = 16'h3022;
    SB_LUT4 i12954_3_lut (.I0(IntegralLimit[16]), .I1(\data_in_frame[11] [0]), 
            .I2(n5439), .I3(GND_net), .O(n17783));   // verilog/coms.v(126[12] 293[6])
    defparam i12954_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY rem_4_add_1586_6 (.CI(n28181), .I0(n2354), .I1(GND_net), 
            .CO(n28182));
    SB_LUT4 i12955_3_lut (.I0(IntegralLimit[17]), .I1(\data_in_frame[11] [1]), 
            .I2(n5439), .I3(GND_net), .O(n17784));   // verilog/coms.v(126[12] 293[6])
    defparam i12955_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13074_3_lut (.I0(\data_out_frame[8] [4]), .I1(encoder0_position[4]), 
            .I2(n13724), .I3(GND_net), .O(n17903));   // verilog/coms.v(126[12] 293[6])
    defparam i13074_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_add_1586_5_lut (.I0(GND_net), .I1(n2355), .I2(GND_net), 
            .I3(n28180), .O(n2422)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1586_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1586_5 (.CI(n28180), .I0(n2355), .I1(GND_net), 
            .CO(n28181));
    SB_LUT4 i13075_3_lut (.I0(\data_out_frame[8] [5]), .I1(encoder0_position[5]), 
            .I2(n13724), .I3(GND_net), .O(n17904));   // verilog/coms.v(126[12] 293[6])
    defparam i13075_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13076_3_lut (.I0(\data_out_frame[8] [6]), .I1(encoder0_position[6]), 
            .I2(n13724), .I3(GND_net), .O(n17905));   // verilog/coms.v(126[12] 293[6])
    defparam i13076_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13077_3_lut (.I0(\data_out_frame[8] [7]), .I1(encoder0_position[7]), 
            .I2(n13724), .I3(GND_net), .O(n17906));   // verilog/coms.v(126[12] 293[6])
    defparam i13077_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13078_3_lut (.I0(\data_out_frame[9] [0]), .I1(encoder1_position[16]), 
            .I2(n13724), .I3(GND_net), .O(n17907));   // verilog/coms.v(126[12] 293[6])
    defparam i13078_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13079_3_lut (.I0(\data_out_frame[9] [1]), .I1(encoder1_position[17]), 
            .I2(n13724), .I3(GND_net), .O(n17908));   // verilog/coms.v(126[12] 293[6])
    defparam i13079_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13080_3_lut (.I0(\data_out_frame[9] [2]), .I1(encoder1_position[18]), 
            .I2(n13724), .I3(GND_net), .O(n17909));   // verilog/coms.v(126[12] 293[6])
    defparam i13080_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13081_3_lut (.I0(\data_out_frame[9] [3]), .I1(encoder1_position[19]), 
            .I2(n13724), .I3(GND_net), .O(n17910));   // verilog/coms.v(126[12] 293[6])
    defparam i13081_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13082_3_lut (.I0(\data_out_frame[9] [4]), .I1(encoder1_position[20]), 
            .I2(n13724), .I3(GND_net), .O(n17911));   // verilog/coms.v(126[12] 293[6])
    defparam i13082_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13083_3_lut (.I0(\data_out_frame[9] [5]), .I1(encoder1_position[21]), 
            .I2(n13724), .I3(GND_net), .O(n17912));   // verilog/coms.v(126[12] 293[6])
    defparam i13083_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13084_3_lut (.I0(\data_out_frame[9] [6]), .I1(encoder1_position[22]), 
            .I2(n13724), .I3(GND_net), .O(n17913));   // verilog/coms.v(126[12] 293[6])
    defparam i13084_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13085_3_lut (.I0(\data_out_frame[9] [7]), .I1(encoder1_position[23]), 
            .I2(n13724), .I3(GND_net), .O(n17914));   // verilog/coms.v(126[12] 293[6])
    defparam i13085_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13086_3_lut (.I0(\data_out_frame[10] [0]), .I1(encoder1_position[8]), 
            .I2(n13724), .I3(GND_net), .O(n17915));   // verilog/coms.v(126[12] 293[6])
    defparam i13086_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13087_3_lut (.I0(\data_out_frame[10] [1]), .I1(encoder1_position[9]), 
            .I2(n13724), .I3(GND_net), .O(n17916));   // verilog/coms.v(126[12] 293[6])
    defparam i13087_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i30896_2_lut (.I0(displacement[4]), .I1(control_mode[0]), .I2(GND_net), 
            .I3(GND_net), .O(n37339));   // verilog/TinyFPGA_B.v(210[5] 214[10])
    defparam i30896_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 mux_843_Mux_4_i1_3_lut (.I0(encoder0_position[4]), .I1(encoder1_position[4]), 
            .I2(control_mode[0]), .I3(GND_net), .O(n1_adj_4931));   // verilog/TinyFPGA_B.v(210[5] 214[10])
    defparam mux_843_Mux_4_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13088_3_lut (.I0(\data_out_frame[10] [2]), .I1(encoder1_position[10]), 
            .I2(n13724), .I3(GND_net), .O(n17917));   // verilog/coms.v(126[12] 293[6])
    defparam i13088_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12956_3_lut (.I0(IntegralLimit[18]), .I1(\data_in_frame[11] [2]), 
            .I2(n5439), .I3(GND_net), .O(n17785));   // verilog/coms.v(126[12] 293[6])
    defparam i12956_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13089_3_lut (.I0(\data_out_frame[10] [3]), .I1(encoder1_position[11]), 
            .I2(n13724), .I3(GND_net), .O(n17918));   // verilog/coms.v(126[12] 293[6])
    defparam i13089_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i19543_4_lut (.I0(n1_adj_4931), .I1(n34919), .I2(n37339), 
            .I3(control_mode[1]), .O(motor_state[4]));   // verilog/TinyFPGA_B.v(210[5] 214[10])
    defparam i19543_4_lut.LUT_INIT = 16'h3022;
    SB_LUT4 i13090_3_lut (.I0(\data_out_frame[10] [4]), .I1(encoder1_position[12]), 
            .I2(n13724), .I3(GND_net), .O(n17919));   // verilog/coms.v(126[12] 293[6])
    defparam i13090_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12957_3_lut (.I0(IntegralLimit[19]), .I1(\data_in_frame[11] [3]), 
            .I2(n5439), .I3(GND_net), .O(n17786));   // verilog/coms.v(126[12] 293[6])
    defparam i12957_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13091_3_lut (.I0(\data_out_frame[10] [5]), .I1(encoder1_position[13]), 
            .I2(n13724), .I3(GND_net), .O(n17920));   // verilog/coms.v(126[12] 293[6])
    defparam i13091_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13092_3_lut (.I0(\data_out_frame[10] [6]), .I1(encoder1_position[14]), 
            .I2(n13724), .I3(GND_net), .O(n17921));   // verilog/coms.v(126[12] 293[6])
    defparam i13092_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13093_3_lut (.I0(\data_out_frame[10] [7]), .I1(encoder1_position[15]), 
            .I2(n13724), .I3(GND_net), .O(n17922));   // verilog/coms.v(126[12] 293[6])
    defparam i13093_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13094_3_lut (.I0(\data_out_frame[11] [0]), .I1(encoder1_position[0]), 
            .I2(n13724), .I3(GND_net), .O(n17923));   // verilog/coms.v(126[12] 293[6])
    defparam i13094_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i30897_2_lut (.I0(displacement[5]), .I1(control_mode[0]), .I2(GND_net), 
            .I3(GND_net), .O(n37340));   // verilog/TinyFPGA_B.v(210[5] 214[10])
    defparam i30897_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 mux_843_Mux_5_i1_3_lut (.I0(encoder0_position[5]), .I1(encoder1_position[5]), 
            .I2(control_mode[0]), .I3(GND_net), .O(n1_adj_4932));   // verilog/TinyFPGA_B.v(210[5] 214[10])
    defparam mux_843_Mux_5_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i19544_4_lut (.I0(n1_adj_4932), .I1(n34919), .I2(n37340), 
            .I3(control_mode[1]), .O(motor_state[5]));   // verilog/TinyFPGA_B.v(210[5] 214[10])
    defparam i19544_4_lut.LUT_INIT = 16'h3022;
    SB_LUT4 i12958_3_lut (.I0(IntegralLimit[20]), .I1(\data_in_frame[11] [4]), 
            .I2(n5439), .I3(GND_net), .O(n17787));   // verilog/coms.v(126[12] 293[6])
    defparam i12958_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13095_3_lut (.I0(\data_out_frame[11] [1]), .I1(encoder1_position[1]), 
            .I2(n13724), .I3(GND_net), .O(n17924));   // verilog/coms.v(126[12] 293[6])
    defparam i13095_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12959_3_lut (.I0(IntegralLimit[21]), .I1(\data_in_frame[11] [5]), 
            .I2(n5439), .I3(GND_net), .O(n17788));   // verilog/coms.v(126[12] 293[6])
    defparam i12959_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13096_3_lut (.I0(\data_out_frame[11] [2]), .I1(encoder1_position[2]), 
            .I2(n13724), .I3(GND_net), .O(n17925));   // verilog/coms.v(126[12] 293[6])
    defparam i13096_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13097_3_lut (.I0(\data_out_frame[11] [3]), .I1(encoder1_position[3]), 
            .I2(n13724), .I3(GND_net), .O(n17926));   // verilog/coms.v(126[12] 293[6])
    defparam i13097_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13098_3_lut (.I0(\data_out_frame[11] [4]), .I1(encoder1_position[4]), 
            .I2(n13724), .I3(GND_net), .O(n17927));   // verilog/coms.v(126[12] 293[6])
    defparam i13098_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12960_3_lut (.I0(IntegralLimit[22]), .I1(\data_in_frame[11] [6]), 
            .I2(n5439), .I3(GND_net), .O(n17789));   // verilog/coms.v(126[12] 293[6])
    defparam i12960_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13099_3_lut (.I0(\data_out_frame[11] [5]), .I1(encoder1_position[5]), 
            .I2(n13724), .I3(GND_net), .O(n17928));   // verilog/coms.v(126[12] 293[6])
    defparam i13099_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12961_3_lut (.I0(IntegralLimit[23]), .I1(\data_in_frame[11] [7]), 
            .I2(n5439), .I3(GND_net), .O(n17790));   // verilog/coms.v(126[12] 293[6])
    defparam i12961_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i30898_2_lut (.I0(displacement[6]), .I1(control_mode[0]), .I2(GND_net), 
            .I3(GND_net), .O(n37341));   // verilog/TinyFPGA_B.v(210[5] 214[10])
    defparam i30898_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i12962_3_lut (.I0(\data_in[0] [1]), .I1(\data_in[1] [1]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n17791));   // verilog/coms.v(126[12] 293[6])
    defparam i12962_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_843_Mux_6_i1_3_lut (.I0(encoder0_position[6]), .I1(encoder1_position[6]), 
            .I2(control_mode[0]), .I3(GND_net), .O(n1_adj_4933));   // verilog/TinyFPGA_B.v(210[5] 214[10])
    defparam mux_843_Mux_6_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12964_3_lut (.I0(\data_in[0] [3]), .I1(\data_in[1] [3]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n17793));   // verilog/coms.v(126[12] 293[6])
    defparam i12964_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13100_3_lut (.I0(\data_out_frame[11] [6]), .I1(encoder1_position[6]), 
            .I2(n13724), .I3(GND_net), .O(n17929));   // verilog/coms.v(126[12] 293[6])
    defparam i13100_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i19545_4_lut (.I0(n1_adj_4933), .I1(n34919), .I2(n37341), 
            .I3(control_mode[1]), .O(motor_state[6]));   // verilog/TinyFPGA_B.v(210[5] 214[10])
    defparam i19545_4_lut.LUT_INIT = 16'h3022;
    SB_LUT4 i13101_3_lut (.I0(\data_out_frame[11] [7]), .I1(encoder1_position[7]), 
            .I2(n13724), .I3(GND_net), .O(n17930));   // verilog/coms.v(126[12] 293[6])
    defparam i13101_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13102_3_lut (.I0(\data_out_frame[12] [0]), .I1(setpoint[16]), 
            .I2(n13724), .I3(GND_net), .O(n17931));   // verilog/coms.v(126[12] 293[6])
    defparam i13102_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13103_3_lut (.I0(\data_out_frame[12] [1]), .I1(setpoint[17]), 
            .I2(n13724), .I3(GND_net), .O(n17932));   // verilog/coms.v(126[12] 293[6])
    defparam i13103_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12965_3_lut (.I0(\data_in[0] [4]), .I1(\data_in[1] [4]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n17794));   // verilog/coms.v(126[12] 293[6])
    defparam i12965_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13104_3_lut (.I0(\data_out_frame[12] [2]), .I1(setpoint[18]), 
            .I2(n13724), .I3(GND_net), .O(n17933));   // verilog/coms.v(126[12] 293[6])
    defparam i13104_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12966_3_lut (.I0(\data_in[0] [5]), .I1(\data_in[1] [5]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n17795));   // verilog/coms.v(126[12] 293[6])
    defparam i12966_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12967_3_lut (.I0(\data_in[0] [6]), .I1(\data_in[1] [6]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n17796));   // verilog/coms.v(126[12] 293[6])
    defparam i12967_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12968_3_lut (.I0(\data_in[0] [7]), .I1(\data_in[1] [7]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n17797));   // verilog/coms.v(126[12] 293[6])
    defparam i12968_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12969_3_lut (.I0(\data_in[1] [0]), .I1(\data_in[2] [0]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n17798));   // verilog/coms.v(126[12] 293[6])
    defparam i12969_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12970_3_lut (.I0(\data_in[1] [1]), .I1(\data_in[2] [1]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n17799));   // verilog/coms.v(126[12] 293[6])
    defparam i12970_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13105_3_lut (.I0(\data_out_frame[12] [3]), .I1(setpoint[19]), 
            .I2(n13724), .I3(GND_net), .O(n17934));   // verilog/coms.v(126[12] 293[6])
    defparam i13105_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12971_3_lut (.I0(\data_in[1] [2]), .I1(\data_in[2] [2]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n17800));   // verilog/coms.v(126[12] 293[6])
    defparam i12971_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13106_3_lut (.I0(\data_out_frame[12] [4]), .I1(setpoint[20]), 
            .I2(n13724), .I3(GND_net), .O(n17935));   // verilog/coms.v(126[12] 293[6])
    defparam i13106_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13107_3_lut (.I0(\data_out_frame[12] [5]), .I1(setpoint[21]), 
            .I2(n13724), .I3(GND_net), .O(n17936));   // verilog/coms.v(126[12] 293[6])
    defparam i13107_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13108_3_lut (.I0(\data_out_frame[12] [6]), .I1(setpoint[22]), 
            .I2(n13724), .I3(GND_net), .O(n17937));   // verilog/coms.v(126[12] 293[6])
    defparam i13108_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i30899_2_lut (.I0(displacement[7]), .I1(control_mode[0]), .I2(GND_net), 
            .I3(GND_net), .O(n37342));   // verilog/TinyFPGA_B.v(210[5] 214[10])
    defparam i30899_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 mux_843_Mux_7_i1_3_lut (.I0(encoder0_position[7]), .I1(encoder1_position[7]), 
            .I2(control_mode[0]), .I3(GND_net), .O(n1_adj_4934));   // verilog/TinyFPGA_B.v(210[5] 214[10])
    defparam mux_843_Mux_7_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12972_3_lut (.I0(\data_in[1] [3]), .I1(\data_in[2] [3]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n17801));   // verilog/coms.v(126[12] 293[6])
    defparam i12972_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12973_3_lut (.I0(\data_in[1] [4]), .I1(\data_in[2] [4]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n17802));   // verilog/coms.v(126[12] 293[6])
    defparam i12973_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13109_3_lut (.I0(\data_out_frame[12] [7]), .I1(setpoint[23]), 
            .I2(n13724), .I3(GND_net), .O(n17938));   // verilog/coms.v(126[12] 293[6])
    defparam i13109_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i19546_4_lut (.I0(n1_adj_4934), .I1(n34919), .I2(n37342), 
            .I3(control_mode[1]), .O(motor_state[7]));   // verilog/TinyFPGA_B.v(210[5] 214[10])
    defparam i19546_4_lut.LUT_INIT = 16'h3022;
    SB_LUT4 i13110_3_lut (.I0(\data_out_frame[13] [0]), .I1(setpoint[8]), 
            .I2(n13724), .I3(GND_net), .O(n17939));   // verilog/coms.v(126[12] 293[6])
    defparam i13110_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12974_3_lut (.I0(\data_in[1] [5]), .I1(\data_in[2] [5]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n17803));   // verilog/coms.v(126[12] 293[6])
    defparam i12974_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13111_3_lut (.I0(\data_out_frame[13] [1]), .I1(setpoint[9]), 
            .I2(n13724), .I3(GND_net), .O(n17940));   // verilog/coms.v(126[12] 293[6])
    defparam i13111_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13112_3_lut (.I0(\data_out_frame[13] [2]), .I1(setpoint[10]), 
            .I2(n13724), .I3(GND_net), .O(n17941));   // verilog/coms.v(126[12] 293[6])
    defparam i13112_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13113_3_lut (.I0(\data_out_frame[13] [3]), .I1(setpoint[11]), 
            .I2(n13724), .I3(GND_net), .O(n17942));   // verilog/coms.v(126[12] 293[6])
    defparam i13113_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13114_3_lut (.I0(\data_out_frame[13] [4]), .I1(setpoint[12]), 
            .I2(n13724), .I3(GND_net), .O(n17943));   // verilog/coms.v(126[12] 293[6])
    defparam i13114_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13115_3_lut (.I0(\data_out_frame[13] [5]), .I1(setpoint[13]), 
            .I2(n13724), .I3(GND_net), .O(n17944));   // verilog/coms.v(126[12] 293[6])
    defparam i13115_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13116_3_lut (.I0(\data_out_frame[13] [6]), .I1(setpoint[14]), 
            .I2(n13724), .I3(GND_net), .O(n17945));   // verilog/coms.v(126[12] 293[6])
    defparam i13116_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12975_3_lut (.I0(\data_in[1] [6]), .I1(\data_in[2] [6]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n17804));   // verilog/coms.v(126[12] 293[6])
    defparam i12975_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13117_3_lut (.I0(\data_out_frame[13] [7]), .I1(setpoint[15]), 
            .I2(n13724), .I3(GND_net), .O(n17946));   // verilog/coms.v(126[12] 293[6])
    defparam i13117_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13118_3_lut (.I0(\data_out_frame[14] [0]), .I1(setpoint[0]), 
            .I2(n13724), .I3(GND_net), .O(n17947));   // verilog/coms.v(126[12] 293[6])
    defparam i13118_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13119_3_lut (.I0(\data_out_frame[14] [1]), .I1(setpoint[1]), 
            .I2(n13724), .I3(GND_net), .O(n17948));   // verilog/coms.v(126[12] 293[6])
    defparam i13119_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13120_3_lut (.I0(\data_out_frame[14] [2]), .I1(setpoint[2]), 
            .I2(n13724), .I3(GND_net), .O(n17949));   // verilog/coms.v(126[12] 293[6])
    defparam i13120_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13121_3_lut (.I0(\data_out_frame[14] [3]), .I1(setpoint[3]), 
            .I2(n13724), .I3(GND_net), .O(n17950));   // verilog/coms.v(126[12] 293[6])
    defparam i13121_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13122_3_lut (.I0(\data_out_frame[14] [4]), .I1(setpoint[4]), 
            .I2(n13724), .I3(GND_net), .O(n17951));   // verilog/coms.v(126[12] 293[6])
    defparam i13122_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13123_3_lut (.I0(\data_out_frame[14] [5]), .I1(setpoint[5]), 
            .I2(n13724), .I3(GND_net), .O(n17952));   // verilog/coms.v(126[12] 293[6])
    defparam i13123_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13124_3_lut (.I0(\data_out_frame[14] [6]), .I1(setpoint[6]), 
            .I2(n13724), .I3(GND_net), .O(n17953));   // verilog/coms.v(126[12] 293[6])
    defparam i13124_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13125_3_lut (.I0(\data_out_frame[14] [7]), .I1(setpoint[7]), 
            .I2(n13724), .I3(GND_net), .O(n17954));   // verilog/coms.v(126[12] 293[6])
    defparam i13125_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13126_3_lut (.I0(\data_out_frame[15] [0]), .I1(duty[16]), .I2(n13724), 
            .I3(GND_net), .O(n17955));   // verilog/coms.v(126[12] 293[6])
    defparam i13126_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13127_3_lut (.I0(\data_out_frame[15] [1]), .I1(duty[17]), .I2(n13724), 
            .I3(GND_net), .O(n17956));   // verilog/coms.v(126[12] 293[6])
    defparam i13127_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13128_3_lut (.I0(\data_out_frame[15] [2]), .I1(duty[18]), .I2(n13724), 
            .I3(GND_net), .O(n17957));   // verilog/coms.v(126[12] 293[6])
    defparam i13128_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13129_3_lut (.I0(\data_out_frame[15] [3]), .I1(duty[19]), .I2(n13724), 
            .I3(GND_net), .O(n17958));   // verilog/coms.v(126[12] 293[6])
    defparam i13129_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13130_3_lut (.I0(\data_out_frame[15] [4]), .I1(duty[20]), .I2(n13724), 
            .I3(GND_net), .O(n17959));   // verilog/coms.v(126[12] 293[6])
    defparam i13130_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13131_3_lut (.I0(\data_out_frame[15] [5]), .I1(duty[21]), .I2(n13724), 
            .I3(GND_net), .O(n17960));   // verilog/coms.v(126[12] 293[6])
    defparam i13131_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13132_3_lut (.I0(\data_out_frame[15] [6]), .I1(duty[22]), .I2(n13724), 
            .I3(GND_net), .O(n17961));   // verilog/coms.v(126[12] 293[6])
    defparam i13132_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_add_1586_4_lut (.I0(GND_net), .I1(n2356), .I2(VCC_net), 
            .I3(n28179), .O(n2423)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1586_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1720_5_lut (.I0(GND_net), .I1(n2555), .I2(GND_net), 
            .I3(n28047), .O(n2622)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1720_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1586_4 (.CI(n28179), .I0(n2356), .I1(VCC_net), 
            .CO(n28180));
    SB_LUT4 rem_4_add_1586_3_lut (.I0(GND_net), .I1(n2357), .I2(VCC_net), 
            .I3(n28178), .O(n2424)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1586_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i13133_3_lut (.I0(\data_out_frame[15] [7]), .I1(duty[23]), .I2(n13724), 
            .I3(GND_net), .O(n17962));   // verilog/coms.v(126[12] 293[6])
    defparam i13133_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY rem_4_add_1720_5 (.CI(n28047), .I0(n2555), .I1(GND_net), 
            .CO(n28048));
    SB_LUT4 i13134_3_lut (.I0(\data_out_frame[16] [0]), .I1(duty[8]), .I2(n13724), 
            .I3(GND_net), .O(n17963));   // verilog/coms.v(126[12] 293[6])
    defparam i13134_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13135_3_lut (.I0(\data_out_frame[16] [1]), .I1(duty[9]), .I2(n13724), 
            .I3(GND_net), .O(n17964));   // verilog/coms.v(126[12] 293[6])
    defparam i13135_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i30900_2_lut (.I0(displacement[8]), .I1(control_mode[0]), .I2(GND_net), 
            .I3(GND_net), .O(n37343));   // verilog/TinyFPGA_B.v(210[5] 214[10])
    defparam i30900_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i13136_3_lut (.I0(\data_out_frame[16] [2]), .I1(duty[10]), .I2(n13724), 
            .I3(GND_net), .O(n17965));   // verilog/coms.v(126[12] 293[6])
    defparam i13136_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_unary_minus_2_inv_0_i4_1_lut (.I0(communication_counter[3]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n30_adj_4979));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_unary_minus_2_inv_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i13137_3_lut (.I0(\data_out_frame[16] [3]), .I1(duty[11]), .I2(n13724), 
            .I3(GND_net), .O(n17966));   // verilog/coms.v(126[12] 293[6])
    defparam i13137_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13138_3_lut (.I0(\data_out_frame[16] [4]), .I1(duty[12]), .I2(n13724), 
            .I3(GND_net), .O(n17967));   // verilog/coms.v(126[12] 293[6])
    defparam i13138_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13139_3_lut (.I0(\data_out_frame[16] [5]), .I1(duty[13]), .I2(n13724), 
            .I3(GND_net), .O(n17968));   // verilog/coms.v(126[12] 293[6])
    defparam i13139_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13140_3_lut (.I0(\data_out_frame[16] [6]), .I1(duty[14]), .I2(n13724), 
            .I3(GND_net), .O(n17969));   // verilog/coms.v(126[12] 293[6])
    defparam i13140_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_843_Mux_8_i1_3_lut (.I0(encoder0_position[8]), .I1(encoder1_position[8]), 
            .I2(control_mode[0]), .I3(GND_net), .O(n1_adj_4935));   // verilog/TinyFPGA_B.v(210[5] 214[10])
    defparam mux_843_Mux_8_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13141_3_lut (.I0(\data_out_frame[16] [7]), .I1(duty[15]), .I2(n13724), 
            .I3(GND_net), .O(n17970));   // verilog/coms.v(126[12] 293[6])
    defparam i13141_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13142_3_lut (.I0(\data_out_frame[17] [0]), .I1(duty[0]), .I2(n13724), 
            .I3(GND_net), .O(n17971));   // verilog/coms.v(126[12] 293[6])
    defparam i13142_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i19547_4_lut (.I0(n1_adj_4935), .I1(n34919), .I2(n37343), 
            .I3(control_mode[1]), .O(motor_state[8]));   // verilog/TinyFPGA_B.v(210[5] 214[10])
    defparam i19547_4_lut.LUT_INIT = 16'h3022;
    SB_LUT4 i13143_3_lut (.I0(\data_out_frame[17] [1]), .I1(duty[1]), .I2(n13724), 
            .I3(GND_net), .O(n17972));   // verilog/coms.v(126[12] 293[6])
    defparam i13143_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_unary_minus_2_inv_0_i5_1_lut (.I0(communication_counter[4]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n29_adj_4978));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_unary_minus_2_inv_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i13144_3_lut (.I0(\data_out_frame[17] [2]), .I1(duty[2]), .I2(n13724), 
            .I3(GND_net), .O(n17973));   // verilog/coms.v(126[12] 293[6])
    defparam i13144_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13145_3_lut (.I0(\data_out_frame[17] [3]), .I1(duty[3]), .I2(n13724), 
            .I3(GND_net), .O(n17974));   // verilog/coms.v(126[12] 293[6])
    defparam i13145_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13146_3_lut (.I0(\data_out_frame[17] [4]), .I1(duty[4]), .I2(n13724), 
            .I3(GND_net), .O(n17975));   // verilog/coms.v(126[12] 293[6])
    defparam i13146_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i30901_2_lut (.I0(displacement[9]), .I1(control_mode[0]), .I2(GND_net), 
            .I3(GND_net), .O(n37344));   // verilog/TinyFPGA_B.v(210[5] 214[10])
    defparam i30901_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 mux_843_Mux_9_i1_3_lut (.I0(encoder0_position[9]), .I1(encoder1_position[9]), 
            .I2(control_mode[0]), .I3(GND_net), .O(n1_adj_4936));   // verilog/TinyFPGA_B.v(210[5] 214[10])
    defparam mux_843_Mux_9_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13147_3_lut (.I0(\data_out_frame[17] [5]), .I1(duty[5]), .I2(n13724), 
            .I3(GND_net), .O(n17976));   // verilog/coms.v(126[12] 293[6])
    defparam i13147_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13148_3_lut (.I0(\data_out_frame[17] [6]), .I1(duty[6]), .I2(n13724), 
            .I3(GND_net), .O(n17977));   // verilog/coms.v(126[12] 293[6])
    defparam i13148_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13149_3_lut (.I0(\data_out_frame[17] [7]), .I1(duty[7]), .I2(n13724), 
            .I3(GND_net), .O(n17978));   // verilog/coms.v(126[12] 293[6])
    defparam i13149_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13150_3_lut (.I0(\data_out_frame[18] [0]), .I1(displacement[16]), 
            .I2(n13724), .I3(GND_net), .O(n17979));   // verilog/coms.v(126[12] 293[6])
    defparam i13150_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13151_3_lut (.I0(\data_out_frame[18] [1]), .I1(displacement[17]), 
            .I2(n13724), .I3(GND_net), .O(n17980));   // verilog/coms.v(126[12] 293[6])
    defparam i13151_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i19548_4_lut (.I0(n1_adj_4936), .I1(n34919), .I2(n37344), 
            .I3(control_mode[1]), .O(motor_state[9]));   // verilog/TinyFPGA_B.v(210[5] 214[10])
    defparam i19548_4_lut.LUT_INIT = 16'h3022;
    SB_CARRY rem_4_add_1586_3 (.CI(n28178), .I0(n2357), .I1(VCC_net), 
            .CO(n28179));
    SB_LUT4 rem_4_add_1720_4_lut (.I0(GND_net), .I1(n2556), .I2(VCC_net), 
            .I3(n28046), .O(n2623)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1720_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1586_2_lut (.I0(GND_net), .I1(n2358), .I2(GND_net), 
            .I3(VCC_net), .O(n2425)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1586_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1720_4 (.CI(n28046), .I0(n2556), .I1(VCC_net), 
            .CO(n28047));
    SB_CARRY rem_4_add_1586_2 (.CI(VCC_net), .I0(n2358), .I1(GND_net), 
            .CO(n28178));
    SB_LUT4 add_582_24_lut (.I0(duty[22]), .I1(n38238), .I2(n3), .I3(n28177), 
            .O(pwm_setpoint_22__N_57[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_582_24_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 rem_4_add_1720_3_lut (.I0(GND_net), .I1(n2557), .I2(VCC_net), 
            .I3(n28045), .O(n2624)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1720_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i30902_2_lut (.I0(displacement[10]), .I1(control_mode[0]), .I2(GND_net), 
            .I3(GND_net), .O(n37345));   // verilog/TinyFPGA_B.v(210[5] 214[10])
    defparam i30902_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 mux_843_Mux_10_i1_3_lut (.I0(encoder0_position[10]), .I1(encoder1_position[10]), 
            .I2(control_mode[0]), .I3(GND_net), .O(n1_adj_4937));   // verilog/TinyFPGA_B.v(210[5] 214[10])
    defparam mux_843_Mux_10_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i19549_4_lut (.I0(n1_adj_4937), .I1(n34919), .I2(n37345), 
            .I3(control_mode[1]), .O(motor_state[10]));   // verilog/TinyFPGA_B.v(210[5] 214[10])
    defparam i19549_4_lut.LUT_INIT = 16'h3022;
    SB_LUT4 rem_4_unary_minus_2_inv_0_i6_1_lut (.I0(communication_counter[5]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n28_adj_4977));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_unary_minus_2_inv_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i12976_3_lut (.I0(\data_in[1] [7]), .I1(\data_in[2] [7]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n17805));   // verilog/coms.v(126[12] 293[6])
    defparam i12976_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_unary_minus_2_inv_0_i7_1_lut (.I0(communication_counter[6]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n27_adj_4976));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_unary_minus_2_inv_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_582_23_lut (.I0(duty[21]), .I1(n38238), .I2(n4_adj_4772), 
            .I3(n28176), .O(pwm_setpoint_22__N_57[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_582_23_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_582_23 (.CI(n28176), .I0(n38238), .I1(n4_adj_4772), .CO(n28177));
    SB_CARRY rem_4_add_1720_3 (.CI(n28045), .I0(n2557), .I1(VCC_net), 
            .CO(n28046));
    SB_LUT4 i13152_3_lut (.I0(\data_out_frame[18] [2]), .I1(displacement[18]), 
            .I2(n13724), .I3(GND_net), .O(n17981));   // verilog/coms.v(126[12] 293[6])
    defparam i13152_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i30903_2_lut (.I0(displacement[11]), .I1(control_mode[0]), .I2(GND_net), 
            .I3(GND_net), .O(n37346));   // verilog/TinyFPGA_B.v(210[5] 214[10])
    defparam i30903_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 rem_4_mux_3_i3_3_lut (.I0(communication_counter[2]), .I1(n31_adj_4853), 
            .I2(communication_counter[31]), .I3(GND_net), .O(n3358));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_mux_3_i3_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_add_1720_2_lut (.I0(GND_net), .I1(n2558), .I2(GND_net), 
            .I3(VCC_net), .O(n2625)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1720_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mux_843_Mux_11_i1_3_lut (.I0(encoder0_position[11]), .I1(encoder1_position[11]), 
            .I2(control_mode[0]), .I3(GND_net), .O(n1_adj_4938));   // verilog/TinyFPGA_B.v(210[5] 214[10])
    defparam mux_843_Mux_11_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY rem_4_add_1720_2 (.CI(VCC_net), .I0(n2558), .I1(GND_net), 
            .CO(n28045));
    SB_LUT4 i19550_4_lut (.I0(n1_adj_4938), .I1(n34919), .I2(n37346), 
            .I3(control_mode[1]), .O(motor_state[11]));   // verilog/TinyFPGA_B.v(210[5] 214[10])
    defparam i19550_4_lut.LUT_INIT = 16'h3022;
    SB_CARRY rem_4_add_1787_9 (.CI(n27881), .I0(n2651), .I1(n2669), .CO(n27882));
    SB_LUT4 i13153_3_lut (.I0(\data_out_frame[18] [3]), .I1(displacement[19]), 
            .I2(n13724), .I3(GND_net), .O(n17982));   // verilog/coms.v(126[12] 293[6])
    defparam i13153_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_add_1787_8_lut (.I0(n2652), .I1(n2652), .I2(n2669), 
            .I3(n27880), .O(n2751)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1787_8_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i30904_2_lut (.I0(displacement[12]), .I1(control_mode[0]), .I2(GND_net), 
            .I3(GND_net), .O(n37347));   // verilog/TinyFPGA_B.v(210[5] 214[10])
    defparam i30904_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 mux_843_Mux_12_i1_3_lut (.I0(encoder0_position[12]), .I1(encoder1_position[12]), 
            .I2(control_mode[0]), .I3(GND_net), .O(n1_adj_4939));   // verilog/TinyFPGA_B.v(210[5] 214[10])
    defparam mux_843_Mux_12_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i19551_4_lut (.I0(n1_adj_4939), .I1(n34919), .I2(n37347), 
            .I3(control_mode[1]), .O(motor_state[12]));   // verilog/TinyFPGA_B.v(210[5] 214[10])
    defparam i19551_4_lut.LUT_INIT = 16'h3022;
    SB_CARRY rem_4_add_1787_8 (.CI(n27880), .I0(n2652), .I1(n2669), .CO(n27881));
    SB_LUT4 add_5647_7_lut (.I0(GND_net), .I1(n3353), .I2(VCC_net), .I3(n28044), 
            .O(n10390)) /* synthesis syn_instantiated=1 */ ;
    defparam add_5647_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1787_7_lut (.I0(n2653), .I1(n2653), .I2(n2669), 
            .I3(n27879), .O(n2752)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1787_7_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 add_582_22_lut (.I0(duty[20]), .I1(n38238), .I2(n5), .I3(n28175), 
            .O(pwm_setpoint_22__N_57[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_582_22_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY rem_4_add_1787_7 (.CI(n27879), .I0(n2653), .I1(n2669), .CO(n27880));
    SB_CARRY add_582_22 (.CI(n28175), .I0(n38238), .I1(n5), .CO(n28176));
    SB_LUT4 add_582_21_lut (.I0(duty[19]), .I1(n38238), .I2(n6), .I3(n28174), 
            .O(pwm_setpoint_22__N_57[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_582_21_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 i30905_2_lut (.I0(displacement[13]), .I1(control_mode[0]), .I2(GND_net), 
            .I3(GND_net), .O(n37348));   // verilog/TinyFPGA_B.v(210[5] 214[10])
    defparam i30905_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 mux_843_Mux_13_i1_3_lut (.I0(encoder0_position[13]), .I1(encoder1_position[13]), 
            .I2(control_mode[0]), .I3(GND_net), .O(n1_adj_4940));   // verilog/TinyFPGA_B.v(210[5] 214[10])
    defparam mux_843_Mux_13_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_582_21 (.CI(n28174), .I0(n38238), .I1(n6), .CO(n28175));
    SB_LUT4 i19552_4_lut (.I0(n1_adj_4940), .I1(n34919), .I2(n37348), 
            .I3(control_mode[1]), .O(motor_state[13]));   // verilog/TinyFPGA_B.v(210[5] 214[10])
    defparam i19552_4_lut.LUT_INIT = 16'h3022;
    SB_LUT4 unary_minus_28_inv_0_i13_1_lut (.I0(duty[12]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n13));   // verilog/TinyFPGA_B.v(149[23:28])
    defparam unary_minus_28_inv_0_i13_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 rem_4_add_1787_6_lut (.I0(n2654), .I1(n2654), .I2(n38232), 
            .I3(n27878), .O(n2753)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1787_6_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY rem_4_add_1787_6 (.CI(n27878), .I0(n2654), .I1(n38232), .CO(n27879));
    SB_LUT4 i13154_3_lut (.I0(\data_out_frame[18] [4]), .I1(displacement[20]), 
            .I2(n13724), .I3(GND_net), .O(n17983));   // verilog/coms.v(126[12] 293[6])
    defparam i13154_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13443_3_lut (.I0(color[9]), .I1(n54), .I2(n15_adj_4850), 
            .I3(GND_net), .O(n18272));   // verilog/TinyFPGA_B.v(51[8] 74[4])
    defparam i13443_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13155_3_lut (.I0(\data_out_frame[18] [5]), .I1(displacement[21]), 
            .I2(n13724), .I3(GND_net), .O(n17984));   // verilog/coms.v(126[12] 293[6])
    defparam i13155_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13156_3_lut (.I0(\data_out_frame[18] [6]), .I1(displacement[22]), 
            .I2(n13724), .I3(GND_net), .O(n17985));   // verilog/coms.v(126[12] 293[6])
    defparam i13156_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13444_3_lut (.I0(color[10]), .I1(n54), .I2(n15_adj_4850), 
            .I3(GND_net), .O(n18273));   // verilog/TinyFPGA_B.v(51[8] 74[4])
    defparam i13444_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 rem_4_i2219_3_lut (.I0(n3258), .I1(n3325), .I2(n3263), .I3(GND_net), 
            .O(n3357));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i2219_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13157_3_lut (.I0(\data_out_frame[18] [7]), .I1(displacement[23]), 
            .I2(n13724), .I3(GND_net), .O(n17986));   // verilog/coms.v(126[12] 293[6])
    defparam i13157_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13158_3_lut (.I0(\data_out_frame[19] [0]), .I1(displacement[8]), 
            .I2(n13724), .I3(GND_net), .O(n17987));   // verilog/coms.v(126[12] 293[6])
    defparam i13158_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13159_3_lut (.I0(\data_out_frame[19] [1]), .I1(displacement[9]), 
            .I2(n13724), .I3(GND_net), .O(n17988));   // verilog/coms.v(126[12] 293[6])
    defparam i13159_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13364_3_lut (.I0(PWMLimit[8]), .I1(\data_in_frame[9] [0]), 
            .I2(n5439), .I3(GND_net), .O(n18193));   // verilog/coms.v(126[12] 293[6])
    defparam i13364_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13445_3_lut (.I0(color[11]), .I1(n54), .I2(n15_adj_4850), 
            .I3(GND_net), .O(n18274));   // verilog/TinyFPGA_B.v(51[8] 74[4])
    defparam i13445_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13363_3_lut (.I0(PWMLimit[7]), .I1(\data_in_frame[10] [7]), 
            .I2(n5439), .I3(GND_net), .O(n18192));   // verilog/coms.v(126[12] 293[6])
    defparam i13363_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13362_3_lut (.I0(PWMLimit[6]), .I1(\data_in_frame[10] [6]), 
            .I2(n5439), .I3(GND_net), .O(n18191));   // verilog/coms.v(126[12] 293[6])
    defparam i13362_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut (.I0(blink), .I1(n15_adj_4850), .I2(GND_net), .I3(GND_net), 
            .O(blink_N_354));
    defparam i1_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i13361_3_lut (.I0(PWMLimit[5]), .I1(\data_in_frame[10] [5]), 
            .I2(n5439), .I3(GND_net), .O(n18190));   // verilog/coms.v(126[12] 293[6])
    defparam i13361_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3_2_lut (.I0(color_23__N_209[3]), .I1(color_23__N_209[5]), 
            .I2(GND_net), .I3(GND_net), .O(n11_adj_4927));   // verilog/TinyFPGA_B.v(54[6:36])
    defparam i3_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i1_4_lut (.I0(color_23__N_209[4]), .I1(color_23__N_209[6]), 
            .I2(color_23__N_209[2]), .I3(color_23__N_209[0]), .O(n13_adj_4926));   // verilog/TinyFPGA_B.v(54[6:36])
    defparam i1_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 rem_4_unary_minus_2_inv_0_i8_1_lut (.I0(communication_counter[7]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n26_adj_4975));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_unary_minus_2_inv_0_i8_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1_4_lut_adj_1600 (.I0(color_23__N_209[7]), .I1(n13_adj_4926), 
            .I2(n11_adj_4927), .I3(color_23__N_209[1]), .O(n15_adj_4850));   // verilog/TinyFPGA_B.v(54[6:36])
    defparam i1_4_lut_adj_1600.LUT_INIT = 16'hfffe;
    SB_LUT4 rem_4_unary_minus_2_inv_0_i9_1_lut (.I0(communication_counter[8]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n25_adj_4974));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_unary_minus_2_inv_0_i9_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i13360_3_lut (.I0(PWMLimit[4]), .I1(\data_in_frame[10] [4]), 
            .I2(n5439), .I3(GND_net), .O(n18189));   // verilog/coms.v(126[12] 293[6])
    defparam i13360_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_adj_1601 (.I0(color_23__N_209[1]), .I1(blink), .I2(GND_net), 
            .I3(GND_net), .O(n35933));   // verilog/TinyFPGA_B.v(54[6:36])
    defparam i1_2_lut_adj_1601.LUT_INIT = 16'heeee;
    SB_LUT4 i1_4_lut_adj_1602 (.I0(color_23__N_209[7]), .I1(n13_adj_4926), 
            .I2(n11_adj_4927), .I3(n35933), .O(n54));   // verilog/TinyFPGA_B.v(54[6:36])
    defparam i1_4_lut_adj_1602.LUT_INIT = 16'hfffe;
    SB_LUT4 i13359_3_lut (.I0(PWMLimit[3]), .I1(\data_in_frame[10] [3]), 
            .I2(n5439), .I3(GND_net), .O(n18188));   // verilog/coms.v(126[12] 293[6])
    defparam i13359_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_unary_minus_2_inv_0_i10_1_lut (.I0(communication_counter[9]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n24_adj_4973));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_unary_minus_2_inv_0_i10_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_28_inv_0_i14_1_lut (.I0(duty[13]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n12_adj_4773));   // verilog/TinyFPGA_B.v(149[23:28])
    defparam unary_minus_28_inv_0_i14_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i13446_3_lut (.I0(color[12]), .I1(n54), .I2(n15_adj_4850), 
            .I3(GND_net), .O(n18275));   // verilog/TinyFPGA_B.v(51[8] 74[4])
    defparam i13446_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 add_582_20_lut (.I0(duty[18]), .I1(n38238), .I2(n7), .I3(n28173), 
            .O(pwm_setpoint_22__N_57[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_582_20_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_582_20 (.CI(n28173), .I0(n38238), .I1(n7), .CO(n28174));
    SB_LUT4 add_582_19_lut (.I0(duty[17]), .I1(n38238), .I2(n8), .I3(n28172), 
            .O(pwm_setpoint_22__N_57[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_582_19_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_582_19 (.CI(n28172), .I0(n38238), .I1(n8), .CO(n28173));
    SB_LUT4 i18_4_lut (.I0(n4), .I1(n35088), .I2(state[1]), .I3(start), 
            .O(n31599));   // verilog/neopixel.v(35[12] 117[6])
    defparam i18_4_lut.LUT_INIT = 16'hfa3a;
    SB_LUT4 add_582_18_lut (.I0(duty[16]), .I1(n38238), .I2(n9), .I3(n28171), 
            .O(pwm_setpoint_22__N_57[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_582_18_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 rem_4_unary_minus_2_add_3_33_lut (.I0(communication_counter[31]), 
            .I1(GND_net), .I2(n2_adj_4951), .I3(n29599), .O(n746)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_unary_minus_2_add_3_33_lut.LUT_INIT = 16'h8228;
    SB_LUT4 rem_4_unary_minus_2_inv_0_i11_1_lut (.I0(communication_counter[10]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n23_adj_4972));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_unary_minus_2_inv_0_i11_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i13160_3_lut (.I0(\data_out_frame[19] [2]), .I1(displacement[10]), 
            .I2(n13724), .I3(GND_net), .O(n17989));   // verilog/coms.v(126[12] 293[6])
    defparam i13160_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_unary_minus_2_add_3_32_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n3_adj_4952), .I3(n29598), .O(n3_adj_4881)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_unary_minus_2_add_3_32_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i30906_2_lut (.I0(displacement[14]), .I1(control_mode[0]), .I2(GND_net), 
            .I3(GND_net), .O(n37349));   // verilog/TinyFPGA_B.v(210[5] 214[10])
    defparam i30906_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 mux_843_Mux_14_i1_3_lut (.I0(encoder0_position[14]), .I1(encoder1_position[14]), 
            .I2(control_mode[0]), .I3(GND_net), .O(n1_adj_4941));   // verilog/TinyFPGA_B.v(210[5] 214[10])
    defparam mux_843_Mux_14_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i19553_4_lut (.I0(n1_adj_4941), .I1(n34919), .I2(n37349), 
            .I3(control_mode[1]), .O(motor_state[14]));   // verilog/TinyFPGA_B.v(210[5] 214[10])
    defparam i19553_4_lut.LUT_INIT = 16'h3022;
    SB_CARRY rem_4_unary_minus_2_add_3_32 (.CI(n29598), .I0(GND_net), .I1(n3_adj_4952), 
            .CO(n29599));
    SB_LUT4 rem_4_unary_minus_2_inv_0_i12_1_lut (.I0(communication_counter[11]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n22_adj_4971));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_unary_minus_2_inv_0_i12_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 rem_4_unary_minus_2_add_3_31_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n4_adj_4953), .I3(n29597), .O(n4_adj_4880)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_unary_minus_2_add_3_31_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i12724_4_lut (.I0(n5478), .I1(r_Clock_Count_adj_5048[5]), .I2(n316), 
            .I3(r_SM_Main_adj_5047[2]), .O(n17553));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i12724_4_lut.LUT_INIT = 16'h4450;
    SB_LUT4 i13358_3_lut (.I0(PWMLimit[2]), .I1(\data_in_frame[10] [2]), 
            .I2(n5439), .I3(GND_net), .O(n18187));   // verilog/coms.v(126[12] 293[6])
    defparam i13358_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_add_1787_5_lut (.I0(n2655), .I1(n2655), .I2(n38232), 
            .I3(n27877), .O(n2754)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1787_5_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY rem_4_add_1787_5 (.CI(n27877), .I0(n2655), .I1(n38232), .CO(n27878));
    SB_CARRY rem_4_unary_minus_2_add_3_31 (.CI(n29597), .I0(GND_net), .I1(n4_adj_4953), 
            .CO(n29598));
    SB_LUT4 i13357_3_lut (.I0(PWMLimit[1]), .I1(\data_in_frame[10] [1]), 
            .I2(n5439), .I3(GND_net), .O(n18186));   // verilog/coms.v(126[12] 293[6])
    defparam i13357_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_unary_minus_2_add_3_30_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n5_adj_4954), .I3(n29596), .O(n5_adj_4879)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_unary_minus_2_add_3_30_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_unary_minus_2_add_3_30 (.CI(n29596), .I0(GND_net), .I1(n5_adj_4954), 
            .CO(n29597));
    SB_LUT4 rem_4_unary_minus_2_inv_0_i13_1_lut (.I0(communication_counter[12]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n21_adj_4970));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_unary_minus_2_inv_0_i13_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_28_inv_0_i15_1_lut (.I0(duty[14]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n11));   // verilog/TinyFPGA_B.v(149[23:28])
    defparam unary_minus_28_inv_0_i15_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i30907_2_lut (.I0(displacement[15]), .I1(control_mode[0]), .I2(GND_net), 
            .I3(GND_net), .O(n37350));   // verilog/TinyFPGA_B.v(210[5] 214[10])
    defparam i30907_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 rem_4_i1462_3_lut (.I0(n2149), .I1(n2216), .I2(n2174), .I3(GND_net), 
            .O(n2248));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1462_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1529_3_lut (.I0(n2248), .I1(n2315), .I2(n2273), .I3(GND_net), 
            .O(n2347));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1529_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_unary_minus_2_add_3_29_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n6_adj_4955), .I3(n29595), .O(n6_adj_4878)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_unary_minus_2_add_3_29_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mux_843_Mux_15_i1_3_lut (.I0(encoder0_position[15]), .I1(encoder1_position[15]), 
            .I2(control_mode[0]), .I3(GND_net), .O(n1_adj_4942));   // verilog/TinyFPGA_B.v(210[5] 214[10])
    defparam mux_843_Mux_15_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY rem_4_unary_minus_2_add_3_29 (.CI(n29595), .I0(GND_net), .I1(n6_adj_4955), 
            .CO(n29596));
    SB_LUT4 i13161_3_lut (.I0(\data_out_frame[19] [3]), .I1(displacement[11]), 
            .I2(n13724), .I3(GND_net), .O(n17990));   // verilog/coms.v(126[12] 293[6])
    defparam i13161_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_582_18 (.CI(n28171), .I0(n38238), .I1(n9), .CO(n28172));
    SB_LUT4 i19554_4_lut (.I0(n1_adj_4942), .I1(n34919), .I2(n37350), 
            .I3(control_mode[1]), .O(motor_state[15]));   // verilog/TinyFPGA_B.v(210[5] 214[10])
    defparam i19554_4_lut.LUT_INIT = 16'h3022;
    SB_LUT4 i13162_3_lut (.I0(\data_out_frame[19] [4]), .I1(displacement[12]), 
            .I2(n13724), .I3(GND_net), .O(n17991));   // verilog/coms.v(126[12] 293[6])
    defparam i13162_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_unary_minus_2_add_3_28_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n7_adj_4956), .I3(n29594), .O(n7_adj_4877)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_unary_minus_2_add_3_28_lut.LUT_INIT = 16'hC33C;
    SB_IO PIN_20_pad (.PACKAGE_PIN(PIN_20), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(PIN_20_c)) /* synthesis IO_FF_OUT=TRUE */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam PIN_20_pad.PIN_TYPE = 6'b011001;
    defparam PIN_20_pad.PULLUP = 1'b0;
    defparam PIN_20_pad.NEG_TRIGGER = 1'b0;
    defparam PIN_20_pad.IO_STANDARD = "SB_LVCMOS";
    SB_CARRY rem_4_unary_minus_2_add_3_28 (.CI(n29594), .I0(GND_net), .I1(n7_adj_4956), 
            .CO(n29595));
    SB_LUT4 i13163_3_lut (.I0(\data_out_frame[19] [5]), .I1(displacement[13]), 
            .I2(n13724), .I3(GND_net), .O(n17992));   // verilog/coms.v(126[12] 293[6])
    defparam i13163_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_unary_minus_2_inv_0_i14_1_lut (.I0(communication_counter[13]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n20_adj_4969));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_unary_minus_2_inv_0_i14_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 rem_4_unary_minus_2_inv_0_i15_1_lut (.I0(communication_counter[14]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n19_adj_4968));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_unary_minus_2_inv_0_i15_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i13372_3_lut (.I0(PWMLimit[16]), .I1(\data_in_frame[8] [0]), 
            .I2(n5439), .I3(GND_net), .O(n18201));   // verilog/coms.v(126[12] 293[6])
    defparam i13372_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13371_3_lut (.I0(PWMLimit[15]), .I1(\data_in_frame[9] [7]), 
            .I2(n5439), .I3(GND_net), .O(n18200));   // verilog/coms.v(126[12] 293[6])
    defparam i13371_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13382_3_lut (.I0(encoder0_position[3]), .I1(n3229), .I2(count_enable), 
            .I3(GND_net), .O(n18211));   // quad.v(35[10] 41[6])
    defparam i13382_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_unary_minus_2_inv_0_i16_1_lut (.I0(communication_counter[15]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n18_adj_4967));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_unary_minus_2_inv_0_i16_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i13381_3_lut (.I0(encoder0_position[2]), .I1(n3230), .I2(count_enable), 
            .I3(GND_net), .O(n18210));   // quad.v(35[10] 41[6])
    defparam i13381_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13380_3_lut (.I0(encoder0_position[1]), .I1(n3231), .I2(count_enable), 
            .I3(GND_net), .O(n18209));   // quad.v(35[10] 41[6])
    defparam i13380_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i30908_2_lut (.I0(displacement[16]), .I1(control_mode[0]), .I2(GND_net), 
            .I3(GND_net), .O(n37351));   // verilog/TinyFPGA_B.v(210[5] 214[10])
    defparam i30908_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 mux_843_Mux_16_i1_3_lut (.I0(encoder0_position[16]), .I1(encoder1_position[16]), 
            .I2(control_mode[0]), .I3(GND_net), .O(n1_adj_4943));   // verilog/TinyFPGA_B.v(210[5] 214[10])
    defparam mux_843_Mux_16_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i19555_4_lut (.I0(n1_adj_4943), .I1(n34919), .I2(n37351), 
            .I3(control_mode[1]), .O(motor_state[16]));   // verilog/TinyFPGA_B.v(210[5] 214[10])
    defparam i19555_4_lut.LUT_INIT = 16'h3022;
    SB_LUT4 rem_4_unary_minus_2_inv_0_i17_1_lut (.I0(communication_counter[16]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n17_adj_4966));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_unary_minus_2_inv_0_i17_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i12720_4_lut (.I0(n5478), .I1(r_Clock_Count_adj_5048[6]), .I2(n315), 
            .I3(r_SM_Main_adj_5047[2]), .O(n17549));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i12720_4_lut.LUT_INIT = 16'h4450;
    SB_LUT4 i13164_3_lut (.I0(\data_out_frame[19] [6]), .I1(displacement[14]), 
            .I2(n13724), .I3(GND_net), .O(n17993));   // verilog/coms.v(126[12] 293[6])
    defparam i13164_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13384_3_lut (.I0(encoder0_position[5]), .I1(n3227), .I2(count_enable), 
            .I3(GND_net), .O(n18213));   // quad.v(35[10] 41[6])
    defparam i13384_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13165_3_lut (.I0(\data_out_frame[19] [7]), .I1(displacement[15]), 
            .I2(n13724), .I3(GND_net), .O(n17994));   // verilog/coms.v(126[12] 293[6])
    defparam i13165_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13383_3_lut (.I0(encoder0_position[4]), .I1(n3228), .I2(count_enable), 
            .I3(GND_net), .O(n18212));   // quad.v(35[10] 41[6])
    defparam i13383_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13386_3_lut (.I0(encoder0_position[7]), .I1(n3225), .I2(count_enable), 
            .I3(GND_net), .O(n18215));   // quad.v(35[10] 41[6])
    defparam i13386_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13385_3_lut (.I0(encoder0_position[6]), .I1(n3226), .I2(count_enable), 
            .I3(GND_net), .O(n18214));   // quad.v(35[10] 41[6])
    defparam i13385_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i30909_2_lut (.I0(displacement[17]), .I1(control_mode[0]), .I2(GND_net), 
            .I3(GND_net), .O(n37352));   // verilog/TinyFPGA_B.v(210[5] 214[10])
    defparam i30909_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 mux_843_Mux_17_i1_3_lut (.I0(encoder0_position[17]), .I1(encoder1_position[17]), 
            .I2(control_mode[0]), .I3(GND_net), .O(n1_adj_4944));   // verilog/TinyFPGA_B.v(210[5] 214[10])
    defparam mux_843_Mux_17_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i19556_4_lut (.I0(n1_adj_4944), .I1(n34919), .I2(n37352), 
            .I3(control_mode[1]), .O(motor_state[17]));   // verilog/TinyFPGA_B.v(210[5] 214[10])
    defparam i19556_4_lut.LUT_INIT = 16'h3022;
    SB_LUT4 i13388_3_lut (.I0(encoder0_position[9]), .I1(n3223), .I2(count_enable), 
            .I3(GND_net), .O(n18217));   // quad.v(35[10] 41[6])
    defparam i13388_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13166_3_lut (.I0(\data_out_frame[20] [0]), .I1(displacement[0]), 
            .I2(n13724), .I3(GND_net), .O(n17995));   // verilog/coms.v(126[12] 293[6])
    defparam i13166_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i2218_3_lut (.I0(n3257), .I1(n3324), .I2(n3263), .I3(GND_net), 
            .O(n3356));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i2218_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12906_3_lut (.I0(n17681), .I1(r_Bit_Index[0]), .I2(n33769), 
            .I3(GND_net), .O(n17735));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i12906_3_lut.LUT_INIT = 16'h8282;
    SB_LUT4 i12902_4_lut (.I0(n17527), .I1(byte_transmit_counter[0]), .I2(n8014), 
            .I3(n25050), .O(n17731));   // verilog/coms.v(126[12] 293[6])
    defparam i12902_4_lut.LUT_INIT = 16'h4450;
    SB_LUT4 rem_4_unary_minus_2_inv_0_i18_1_lut (.I0(communication_counter[17]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n16_adj_4965));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_unary_minus_2_inv_0_i18_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 rem_4_unary_minus_2_inv_0_i19_1_lut (.I0(communication_counter[18]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n15_adj_4964));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_unary_minus_2_inv_0_i19_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i13387_3_lut (.I0(encoder0_position[8]), .I1(n3224), .I2(count_enable), 
            .I3(GND_net), .O(n18216));   // quad.v(35[10] 41[6])
    defparam i13387_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13390_3_lut (.I0(encoder0_position[11]), .I1(n3221), .I2(count_enable), 
            .I3(GND_net), .O(n18219));   // quad.v(35[10] 41[6])
    defparam i13390_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13389_3_lut (.I0(encoder0_position[10]), .I1(n3222), .I2(count_enable), 
            .I3(GND_net), .O(n18218));   // quad.v(35[10] 41[6])
    defparam i13389_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13392_3_lut (.I0(encoder0_position[13]), .I1(n3219), .I2(count_enable), 
            .I3(GND_net), .O(n18221));   // quad.v(35[10] 41[6])
    defparam i13392_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13391_3_lut (.I0(encoder0_position[12]), .I1(n3220), .I2(count_enable), 
            .I3(GND_net), .O(n18220));   // quad.v(35[10] 41[6])
    defparam i13391_3_lut.LUT_INIT = 16'hcaca;
    SB_IO PIN_19_pad (.PACKAGE_PIN(PIN_19), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(PIN_19_c_0)) /* synthesis IO_FF_OUT=TRUE */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam PIN_19_pad.PIN_TYPE = 6'b011001;
    defparam PIN_19_pad.PULLUP = 1'b0;
    defparam PIN_19_pad.NEG_TRIGGER = 1'b0;
    defparam PIN_19_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO PIN_11_pad (.PACKAGE_PIN(PIN_11), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(PIN_11_c));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam PIN_11_pad.PIN_TYPE = 6'b011001;
    defparam PIN_11_pad.PULLUP = 1'b0;
    defparam PIN_11_pad.NEG_TRIGGER = 1'b0;
    defparam PIN_11_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO PIN_8_pad (.PACKAGE_PIN(PIN_8), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(PIN_8_c));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam PIN_8_pad.PIN_TYPE = 6'b011001;
    defparam PIN_8_pad.PULLUP = 1'b0;
    defparam PIN_8_pad.NEG_TRIGGER = 1'b0;
    defparam PIN_8_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO USBPU_pad (.PACKAGE_PIN(USBPU), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(GND_net));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam USBPU_pad.PIN_TYPE = 6'b011001;
    defparam USBPU_pad.PULLUP = 1'b0;
    defparam USBPU_pad.NEG_TRIGGER = 1'b0;
    defparam USBPU_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO LED_pad (.PACKAGE_PIN(LED), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(LED_c));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam LED_pad.PIN_TYPE = 6'b011001;
    defparam LED_pad.PULLUP = 1'b0;
    defparam LED_pad.NEG_TRIGGER = 1'b0;
    defparam LED_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO PIN_22_pad (.PACKAGE_PIN(PIN_22), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(PIN_22_c)) /* synthesis IO_FF_OUT=TRUE */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam PIN_22_pad.PIN_TYPE = 6'b011001;
    defparam PIN_22_pad.PULLUP = 1'b0;
    defparam PIN_22_pad.NEG_TRIGGER = 1'b0;
    defparam PIN_22_pad.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 rem_4_unary_minus_2_add_3_27_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n8_adj_4957), .I3(n29593), .O(n8_adj_4876)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_unary_minus_2_add_3_27_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_unary_minus_2_add_3_27 (.CI(n29593), .I0(GND_net), .I1(n8_adj_4957), 
            .CO(n29594));
    SB_LUT4 add_5647_6_lut (.I0(GND_net), .I1(n3354), .I2(GND_net), .I3(n28043), 
            .O(n10391)) /* synthesis syn_instantiated=1 */ ;
    defparam add_5647_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_unary_minus_2_add_3_26_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n9_adj_4958), .I3(n29592), .O(n9_adj_4875)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_unary_minus_2_add_3_26_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5647_6 (.CI(n28043), .I0(n3354), .I1(GND_net), .CO(n28044));
    SB_LUT4 add_582_17_lut (.I0(duty[15]), .I1(n38238), .I2(n10), .I3(n28170), 
            .O(pwm_setpoint_22__N_57[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_582_17_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 i12899_3_lut (.I0(n17534), .I1(r_Bit_Index_adj_5049[0]), .I2(n17362), 
            .I3(GND_net), .O(n17728));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i12899_3_lut.LUT_INIT = 16'h1414;
    SB_LUT4 i23_3_lut (.I0(bit_ctr[1]), .I1(n37241), .I2(n33701), .I3(GND_net), 
            .O(n31527));   // verilog/neopixel.v(35[12] 117[6])
    defparam i23_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY rem_4_unary_minus_2_add_3_26 (.CI(n29592), .I0(GND_net), .I1(n9_adj_4958), 
            .CO(n29593));
    SB_LUT4 i23_3_lut_adj_1603 (.I0(bit_ctr[2]), .I1(n37251), .I2(n33701), 
            .I3(GND_net), .O(n31529));   // verilog/neopixel.v(35[12] 117[6])
    defparam i23_3_lut_adj_1603.LUT_INIT = 16'hacac;
    SB_LUT4 rem_4_unary_minus_2_add_3_25_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n10_adj_4959), .I3(n29591), .O(n10_adj_4874)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_unary_minus_2_add_3_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_unary_minus_2_add_3_25 (.CI(n29591), .I0(GND_net), .I1(n10_adj_4959), 
            .CO(n29592));
    SB_LUT4 rem_4_unary_minus_2_add_3_24_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n11_adj_4960), .I3(n29590), .O(n11_adj_4873)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_unary_minus_2_add_3_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_unary_minus_2_inv_0_i20_1_lut (.I0(communication_counter[19]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n14_adj_4963));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_unary_minus_2_inv_0_i20_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i13167_3_lut (.I0(\data_out_frame[20] [1]), .I1(displacement[1]), 
            .I2(n13724), .I3(GND_net), .O(n17996));   // verilog/coms.v(126[12] 293[6])
    defparam i13167_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_add_1787_4_lut (.I0(n2656), .I1(n2656), .I2(n2669), 
            .I3(n27876), .O(n2755)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1787_4_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 unary_minus_28_inv_0_i2_1_lut (.I0(duty[1]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n24));   // verilog/TinyFPGA_B.v(149[23:28])
    defparam unary_minus_28_inv_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i13168_3_lut (.I0(\data_out_frame[20] [2]), .I1(displacement[2]), 
            .I2(n13724), .I3(GND_net), .O(n17997));   // verilog/coms.v(126[12] 293[6])
    defparam i13168_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 unary_minus_28_inv_0_i3_1_lut (.I0(duty[2]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n23));   // verilog/TinyFPGA_B.v(149[23:28])
    defparam unary_minus_28_inv_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i13169_3_lut (.I0(\data_out_frame[20] [3]), .I1(displacement[3]), 
            .I2(n13724), .I3(GND_net), .O(n17998));   // verilog/coms.v(126[12] 293[6])
    defparam i13169_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i22_3_lut (.I0(bit_ctr[3]), .I1(n37232), .I2(n33701), .I3(GND_net), 
            .O(n31531));   // verilog/neopixel.v(35[12] 117[6])
    defparam i22_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i22_3_lut_adj_1604 (.I0(bit_ctr[4]), .I1(n37231), .I2(n33701), 
            .I3(GND_net), .O(n31533));   // verilog/neopixel.v(35[12] 117[6])
    defparam i22_3_lut_adj_1604.LUT_INIT = 16'hacac;
    SB_CARRY rem_4_unary_minus_2_add_3_24 (.CI(n29590), .I0(GND_net), .I1(n11_adj_4960), 
            .CO(n29591));
    SB_LUT4 add_5647_5_lut (.I0(GND_net), .I1(n3355), .I2(GND_net), .I3(n28042), 
            .O(n10392)) /* synthesis syn_instantiated=1 */ ;
    defparam add_5647_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1385_18_lut (.I0(n2075), .I1(n2042), .I2(VCC_net), 
            .I3(n28247), .O(n2141)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1385_18_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i13396_3_lut (.I0(encoder0_position[17]), .I1(n3215), .I2(count_enable), 
            .I3(GND_net), .O(n18225));   // quad.v(35[10] 41[6])
    defparam i13396_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13395_3_lut (.I0(encoder0_position[16]), .I1(n3216), .I2(count_enable), 
            .I3(GND_net), .O(n18224));   // quad.v(35[10] 41[6])
    defparam i13395_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_unary_minus_2_inv_0_i21_1_lut (.I0(communication_counter[20]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n13_adj_4962));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_unary_minus_2_inv_0_i21_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i13394_3_lut (.I0(encoder0_position[15]), .I1(n3217), .I2(count_enable), 
            .I3(GND_net), .O(n18223));   // quad.v(35[10] 41[6])
    defparam i13394_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13393_3_lut (.I0(encoder0_position[14]), .I1(n3218), .I2(count_enable), 
            .I3(GND_net), .O(n18222));   // quad.v(35[10] 41[6])
    defparam i13393_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12884_4_lut (.I0(n5478), .I1(r_Clock_Count_adj_5048[7]), .I2(n314), 
            .I3(r_SM_Main_adj_5047[2]), .O(n17713));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i12884_4_lut.LUT_INIT = 16'h4450;
    SB_LUT4 rem_4_unary_minus_2_inv_0_i22_1_lut (.I0(communication_counter[21]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n12_adj_4961));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_unary_minus_2_inv_0_i22_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 rem_4_unary_minus_2_add_3_23_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n12_adj_4961), .I3(n29589), .O(n12_adj_4872)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_unary_minus_2_add_3_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_unary_minus_2_add_3_23 (.CI(n29589), .I0(GND_net), .I1(n12_adj_4961), 
            .CO(n29590));
    SB_LUT4 rem_4_add_1385_17_lut (.I0(GND_net), .I1(n2043), .I2(VCC_net), 
            .I3(n28246), .O(n2110)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1385_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_unary_minus_2_add_3_22_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n13_adj_4962), .I3(n29588), .O(n13_adj_4871)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_unary_minus_2_add_3_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i13170_3_lut (.I0(\data_out_frame[20] [4]), .I1(displacement[4]), 
            .I2(n13724), .I3(GND_net), .O(n17999));   // verilog/coms.v(126[12] 293[6])
    defparam i13170_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY rem_4_unary_minus_2_add_3_22 (.CI(n29588), .I0(GND_net), .I1(n13_adj_4962), 
            .CO(n29589));
    SB_CARRY rem_4_add_1385_17 (.CI(n28246), .I0(n2043), .I1(VCC_net), 
            .CO(n28247));
    SB_LUT4 i12879_4_lut (.I0(n5478), .I1(r_Clock_Count_adj_5048[8]), .I2(n313), 
            .I3(r_SM_Main_adj_5047[2]), .O(n17708));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i12879_4_lut.LUT_INIT = 16'h4450;
    SB_LUT4 rem_4_unary_minus_2_add_3_21_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n14_adj_4963), .I3(n29587), .O(n14_adj_4870)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_unary_minus_2_add_3_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_unary_minus_2_add_3_21 (.CI(n29587), .I0(GND_net), .I1(n14_adj_4963), 
            .CO(n29588));
    SB_CARRY add_5647_5 (.CI(n28042), .I0(n3355), .I1(GND_net), .CO(n28043));
    SB_LUT4 rem_4_unary_minus_2_add_3_20_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n15_adj_4964), .I3(n29586), .O(n15_adj_4869)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_unary_minus_2_add_3_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_unary_minus_2_add_3_20 (.CI(n29586), .I0(GND_net), .I1(n15_adj_4964), 
            .CO(n29587));
    SB_LUT4 rem_4_unary_minus_2_add_3_19_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n16_adj_4965), .I3(n29585), .O(n16_adj_4868)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_unary_minus_2_add_3_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1385_16_lut (.I0(GND_net), .I1(n2044), .I2(VCC_net), 
            .I3(n28245), .O(n2111)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1385_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_28_inv_0_i4_1_lut (.I0(duty[3]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n22));   // verilog/TinyFPGA_B.v(149[23:28])
    defparam unary_minus_28_inv_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY rem_4_unary_minus_2_add_3_19 (.CI(n29585), .I0(GND_net), .I1(n16_adj_4965), 
            .CO(n29586));
    SB_LUT4 add_5647_4_lut (.I0(GND_net), .I1(n3356), .I2(VCC_net), .I3(n28041), 
            .O(n10393)) /* synthesis syn_instantiated=1 */ ;
    defparam add_5647_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5647_4 (.CI(n28041), .I0(n3356), .I1(VCC_net), .CO(n28042));
    SB_LUT4 i12853_4_lut (.I0(n17681), .I1(r_Bit_Index[1]), .I2(r_Bit_Index[0]), 
            .I3(n33769), .O(n17682));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i12853_4_lut.LUT_INIT = 16'h8828;
    SB_LUT4 rem_4_unary_minus_2_add_3_18_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n17_adj_4966), .I3(n29584), .O(n17_adj_4867)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_unary_minus_2_add_3_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_unary_minus_2_add_3_18 (.CI(n29584), .I0(GND_net), .I1(n17_adj_4966), 
            .CO(n29585));
    SB_LUT4 i12977_3_lut (.I0(\data_in[2] [0]), .I1(\data_in[3] [0]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n17806));   // verilog/coms.v(126[12] 293[6])
    defparam i12977_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_unary_minus_2_add_3_17_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n18_adj_4967), .I3(n29583), .O(n18_adj_4866)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_unary_minus_2_add_3_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_unary_minus_2_add_3_17 (.CI(n29583), .I0(GND_net), .I1(n18_adj_4967), 
            .CO(n29584));
    SB_CARRY rem_4_add_1385_16 (.CI(n28245), .I0(n2044), .I1(VCC_net), 
            .CO(n28246));
    SB_LUT4 rem_4_unary_minus_2_add_3_16_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n19_adj_4968), .I3(n29582), .O(n19_adj_4865)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_unary_minus_2_add_3_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_unary_minus_2_add_3_16 (.CI(n29582), .I0(GND_net), .I1(n19_adj_4968), 
            .CO(n29583));
    SB_LUT4 rem_4_unary_minus_2_add_3_15_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n20_adj_4969), .I3(n29581), .O(n20_adj_4864)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_unary_minus_2_add_3_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_i2217_3_lut (.I0(n3256), .I1(n3323), .I2(n3263), .I3(GND_net), 
            .O(n3355));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i2217_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_582_17 (.CI(n28170), .I0(n38238), .I1(n10), .CO(n28171));
    SB_LUT4 i12850_4_lut (.I0(n17681), .I1(r_Bit_Index[2]), .I2(n5578), 
            .I3(n33769), .O(n17679));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i12850_4_lut.LUT_INIT = 16'h8828;
    SB_CARRY rem_4_unary_minus_2_add_3_15 (.CI(n29581), .I0(GND_net), .I1(n20_adj_4969), 
            .CO(n29582));
    SB_LUT4 i12847_2_lut (.I0(n17527), .I1(n17674), .I2(GND_net), .I3(GND_net), 
            .O(n17676));   // verilog/coms.v(126[12] 293[6])
    defparam i12847_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 rem_4_add_1385_15_lut (.I0(GND_net), .I1(n2045), .I2(VCC_net), 
            .I3(n28244), .O(n2112)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1385_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1787_4 (.CI(n27876), .I0(n2656), .I1(n2669), .CO(n27877));
    SB_LUT4 i13405_3_lut (.I0(encoder1_position[1]), .I1(n3181), .I2(count_enable_adj_4807), 
            .I3(GND_net), .O(n18234));   // quad.v(35[10] 41[6])
    defparam i13405_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13171_3_lut (.I0(\data_out_frame[20] [5]), .I1(displacement[5]), 
            .I2(n13724), .I3(GND_net), .O(n18000));   // verilog/coms.v(126[12] 293[6])
    defparam i13171_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12844_2_lut (.I0(n17527), .I1(n17671), .I2(GND_net), .I3(GND_net), 
            .O(n17673));   // verilog/coms.v(126[12] 293[6])
    defparam i12844_2_lut.LUT_INIT = 16'h4444;
    SB_CARRY rem_4_add_1385_15 (.CI(n28244), .I0(n2045), .I1(VCC_net), 
            .CO(n28245));
    SB_LUT4 i12979_3_lut (.I0(\data_in[2] [2]), .I1(\data_in[3] [2]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n17808));   // verilog/coms.v(126[12] 293[6])
    defparam i12979_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13172_3_lut (.I0(\data_out_frame[20] [6]), .I1(displacement[6]), 
            .I2(n13724), .I3(GND_net), .O(n18001));   // verilog/coms.v(126[12] 293[6])
    defparam i13172_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_582_16_lut (.I0(duty[14]), .I1(n38238), .I2(n11), .I3(n28169), 
            .O(pwm_setpoint_22__N_57[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_582_16_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 rem_4_unary_minus_2_add_3_14_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n21_adj_4970), .I3(n29580), .O(n21_adj_4863)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_unary_minus_2_add_3_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1385_14_lut (.I0(GND_net), .I1(n2046), .I2(VCC_net), 
            .I3(n28243), .O(n2113)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1385_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i30910_2_lut (.I0(displacement[18]), .I1(control_mode[0]), .I2(GND_net), 
            .I3(GND_net), .O(n37353));   // verilog/TinyFPGA_B.v(210[5] 214[10])
    defparam i30910_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i12981_3_lut (.I0(\data_in[2] [4]), .I1(\data_in[3] [4]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n17810));   // verilog/coms.v(126[12] 293[6])
    defparam i12981_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY rem_4_unary_minus_2_add_3_14 (.CI(n29580), .I0(GND_net), .I1(n21_adj_4970), 
            .CO(n29581));
    SB_LUT4 mux_843_Mux_18_i1_3_lut (.I0(encoder0_position[18]), .I1(encoder1_position[18]), 
            .I2(control_mode[0]), .I3(GND_net), .O(n1_adj_4945));   // verilog/TinyFPGA_B.v(210[5] 214[10])
    defparam mux_843_Mux_18_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_add_1787_3_lut (.I0(n2657), .I1(n2657), .I2(n2669), 
            .I3(n27875), .O(n2756)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1787_3_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i19557_4_lut (.I0(n1_adj_4945), .I1(n34919), .I2(n37353), 
            .I3(control_mode[1]), .O(motor_state[18]));   // verilog/TinyFPGA_B.v(210[5] 214[10])
    defparam i19557_4_lut.LUT_INIT = 16'h3022;
    SB_LUT4 rem_4_unary_minus_2_add_3_13_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n22_adj_4971), .I3(n29579), .O(n22_adj_4862)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_unary_minus_2_add_3_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_unary_minus_2_add_3_13 (.CI(n29579), .I0(GND_net), .I1(n22_adj_4971), 
            .CO(n29580));
    SB_CARRY add_582_16 (.CI(n28169), .I0(n38238), .I1(n11), .CO(n28170));
    SB_CARRY rem_4_add_1787_3 (.CI(n27875), .I0(n2657), .I1(n2669), .CO(n27876));
    SB_LUT4 i13173_3_lut (.I0(\data_out_frame[20] [7]), .I1(displacement[7]), 
            .I2(n13724), .I3(GND_net), .O(n18002));   // verilog/coms.v(126[12] 293[6])
    defparam i13173_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_unary_minus_2_add_3_12_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n23_adj_4972), .I3(n29578), .O(n23_adj_4861)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_unary_minus_2_add_3_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i12841_2_lut (.I0(n17527), .I1(n17668), .I2(GND_net), .I3(GND_net), 
            .O(n17670));   // verilog/coms.v(126[12] 293[6])
    defparam i12841_2_lut.LUT_INIT = 16'h4444;
    SB_CARRY rem_4_add_1385_14 (.CI(n28243), .I0(n2046), .I1(VCC_net), 
            .CO(n28244));
    SB_LUT4 add_582_15_lut (.I0(duty[13]), .I1(n38238), .I2(n12_adj_4773), 
            .I3(n28168), .O(pwm_setpoint_22__N_57[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_582_15_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 i12838_2_lut (.I0(n17527), .I1(n17665), .I2(GND_net), .I3(GND_net), 
            .O(n17667));   // verilog/coms.v(126[12] 293[6])
    defparam i12838_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i12983_3_lut (.I0(\data_in[2] [6]), .I1(\data_in[3] [6]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n17812));   // verilog/coms.v(126[12] 293[6])
    defparam i12983_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12984_3_lut (.I0(\data_in[2] [7]), .I1(\data_in[3] [7]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n17813));   // verilog/coms.v(126[12] 293[6])
    defparam i12984_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY rem_4_unary_minus_2_add_3_12 (.CI(n29578), .I0(GND_net), .I1(n23_adj_4972), 
            .CO(n29579));
    SB_LUT4 rem_4_unary_minus_2_add_3_11_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n24_adj_4973), .I3(n29577), .O(n24_adj_4860)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_unary_minus_2_add_3_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i12985_3_lut (.I0(\data_in[3] [0]), .I1(rx_data[0]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n17814));   // verilog/coms.v(126[12] 293[6])
    defparam i12985_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY rem_4_unary_minus_2_add_3_11 (.CI(n29577), .I0(GND_net), .I1(n24_adj_4973), 
            .CO(n29578));
    SB_LUT4 i12835_2_lut (.I0(n17527), .I1(n17662), .I2(GND_net), .I3(GND_net), 
            .O(n17664));   // verilog/coms.v(126[12] 293[6])
    defparam i12835_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 rem_4_add_1787_2_lut (.I0(n2658), .I1(n2658), .I2(n38232), 
            .I3(VCC_net), .O(n2757)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1787_2_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 rem_4_unary_minus_2_add_3_10_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n25_adj_4974), .I3(n29576), .O(n25_adj_4859)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_unary_minus_2_add_3_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i12987_3_lut (.I0(\data_in[3] [2]), .I1(rx_data[2]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n17816));   // verilog/coms.v(126[12] 293[6])
    defparam i12987_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_add_1385_13_lut (.I0(GND_net), .I1(n2047), .I2(VCC_net), 
            .I3(n28242), .O(n2114)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1385_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i12832_2_lut (.I0(n17527), .I1(n17659), .I2(GND_net), .I3(GND_net), 
            .O(n17661));   // verilog/coms.v(126[12] 293[6])
    defparam i12832_2_lut.LUT_INIT = 16'h4444;
    SB_CARRY rem_4_add_1787_2 (.CI(VCC_net), .I0(n2658), .I1(n38232), 
            .CO(n27875));
    SB_CARRY rem_4_unary_minus_2_add_3_10 (.CI(n29576), .I0(GND_net), .I1(n25_adj_4974), 
            .CO(n29577));
    SB_LUT4 rem_4_unary_minus_2_add_3_9_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n26_adj_4975), .I3(n29575), .O(n26_adj_4858)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_unary_minus_2_add_3_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i12989_3_lut (.I0(\data_in[3] [4]), .I1(rx_data[4]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n17818));   // verilog/coms.v(126[12] 293[6])
    defparam i12989_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF communication_counter_1522__i0 (.Q(communication_counter[0]), .C(LED_c), 
           .D(n165));   // verilog/TinyFPGA_B.v(52[28:51])
    SB_LUT4 add_5647_3_lut (.I0(GND_net), .I1(n3357), .I2(VCC_net), .I3(n28040), 
            .O(n10394)) /* synthesis syn_instantiated=1 */ ;
    defparam add_5647_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i30911_2_lut (.I0(displacement[19]), .I1(control_mode[0]), .I2(GND_net), 
            .I3(GND_net), .O(n37354));   // verilog/TinyFPGA_B.v(210[5] 214[10])
    defparam i30911_2_lut.LUT_INIT = 16'h2222;
    SB_CARRY add_582_15 (.CI(n28168), .I0(n38238), .I1(n12_adj_4773), 
            .CO(n28169));
    SB_CARRY rem_4_add_1385_13 (.CI(n28242), .I0(n2047), .I1(VCC_net), 
            .CO(n28243));
    SB_LUT4 i12991_3_lut (.I0(\data_in[3] [6]), .I1(rx_data[6]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n17820));   // verilog/coms.v(126[12] 293[6])
    defparam i12991_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_843_Mux_19_i1_3_lut (.I0(encoder0_position[19]), .I1(encoder1_position[19]), 
            .I2(control_mode[0]), .I3(GND_net), .O(n1_adj_4946));   // verilog/TinyFPGA_B.v(210[5] 214[10])
    defparam mux_843_Mux_19_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_5647_3 (.CI(n28040), .I0(n3357), .I1(VCC_net), .CO(n28041));
    SB_LUT4 add_582_14_lut (.I0(duty[12]), .I1(n38238), .I2(n13), .I3(n28167), 
            .O(pwm_setpoint_22__N_57[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_582_14_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 i19558_4_lut (.I0(n1_adj_4946), .I1(n34919), .I2(n37354), 
            .I3(control_mode[1]), .O(motor_state[19]));   // verilog/TinyFPGA_B.v(210[5] 214[10])
    defparam i19558_4_lut.LUT_INIT = 16'h3022;
    SB_CARRY rem_4_unary_minus_2_add_3_9 (.CI(n29575), .I0(GND_net), .I1(n26_adj_4975), 
            .CO(n29576));
    SB_LUT4 add_5647_2_lut (.I0(GND_net), .I1(n3358), .I2(GND_net), .I3(VCC_net), 
            .O(n10395)) /* synthesis syn_instantiated=1 */ ;
    defparam add_5647_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i12992_3_lut (.I0(\data_in[3] [7]), .I1(rx_data[7]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n17821));   // verilog/coms.v(126[12] 293[6])
    defparam i12992_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_unary_minus_2_add_3_8_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n27_adj_4976), .I3(n29574), .O(n27_adj_4857)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_unary_minus_2_add_3_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_unary_minus_2_add_3_8 (.CI(n29574), .I0(GND_net), .I1(n27_adj_4976), 
            .CO(n29575));
    SB_CARRY add_5647_2 (.CI(VCC_net), .I0(n3358), .I1(GND_net), .CO(n28040));
    SB_LUT4 i12829_2_lut (.I0(n17527), .I1(n17656), .I2(GND_net), .I3(GND_net), 
            .O(n17658));   // verilog/coms.v(126[12] 293[6])
    defparam i12829_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 unary_minus_28_inv_0_i5_1_lut (.I0(duty[4]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n21));   // verilog/TinyFPGA_B.v(149[23:28])
    defparam unary_minus_28_inv_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i12993_3_lut (.I0(Kp[1]), .I1(\data_in_frame[3] [1]), .I2(n34066), 
            .I3(GND_net), .O(n17822));   // verilog/coms.v(126[12] 293[6])
    defparam i12993_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12826_4_lut (.I0(n17534), .I1(r_Bit_Index_adj_5049[1]), .I2(r_Bit_Index_adj_5049[0]), 
            .I3(n17362), .O(n17655));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i12826_4_lut.LUT_INIT = 16'h1444;
    SB_CARRY add_582_14 (.CI(n28167), .I0(n38238), .I1(n13), .CO(n28168));
    SB_LUT4 rem_4_unary_minus_2_add_3_7_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n28_adj_4977), .I3(n29573), .O(n28_adj_4856)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_unary_minus_2_add_3_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_unary_minus_2_add_3_7 (.CI(n29573), .I0(GND_net), .I1(n28_adj_4977), 
            .CO(n29574));
    SB_LUT4 rem_4_unary_minus_2_add_3_6_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n29_adj_4978), .I3(n29572), .O(n29_adj_4855)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_unary_minus_2_add_3_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i12823_4_lut (.I0(n17534), .I1(r_Bit_Index_adj_5049[2]), .I2(n5600), 
            .I3(n17362), .O(n17652));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i12823_4_lut.LUT_INIT = 16'h1444;
    SB_LUT4 i22_3_lut_adj_1605 (.I0(bit_ctr[5]), .I1(n37230), .I2(n33701), 
            .I3(GND_net), .O(n31535));   // verilog/neopixel.v(35[12] 117[6])
    defparam i22_3_lut_adj_1605.LUT_INIT = 16'hacac;
    SB_LUT4 i22_3_lut_adj_1606 (.I0(bit_ctr[6]), .I1(n37229), .I2(n33701), 
            .I3(GND_net), .O(n31537));   // verilog/neopixel.v(35[12] 117[6])
    defparam i22_3_lut_adj_1606.LUT_INIT = 16'hacac;
    SB_CARRY rem_4_unary_minus_2_add_3_6 (.CI(n29572), .I0(GND_net), .I1(n29_adj_4978), 
            .CO(n29573));
    SB_DFF h1_67 (.Q(PIN_20_c), .C(clk32MHz), .D(hall1));   // verilog/TinyFPGA_B.v(139[10] 152[6])
    SB_LUT4 i22_3_lut_adj_1607 (.I0(bit_ctr[7]), .I1(n37228), .I2(n33701), 
            .I3(GND_net), .O(n31539));   // verilog/neopixel.v(35[12] 117[6])
    defparam i22_3_lut_adj_1607.LUT_INIT = 16'hacac;
    SB_LUT4 i30912_2_lut (.I0(displacement[20]), .I1(control_mode[0]), .I2(GND_net), 
            .I3(GND_net), .O(n37355));   // verilog/TinyFPGA_B.v(210[5] 214[10])
    defparam i30912_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 mux_843_Mux_20_i1_3_lut (.I0(encoder0_position[20]), .I1(encoder1_position[20]), 
            .I2(control_mode[0]), .I3(GND_net), .O(n1_adj_4947));   // verilog/TinyFPGA_B.v(210[5] 214[10])
    defparam mux_843_Mux_20_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i19559_4_lut (.I0(n1_adj_4947), .I1(n34919), .I2(n37355), 
            .I3(control_mode[1]), .O(motor_state[20]));   // verilog/TinyFPGA_B.v(210[5] 214[10])
    defparam i19559_4_lut.LUT_INIT = 16'h3022;
    SB_LUT4 i12994_3_lut (.I0(Kp[2]), .I1(\data_in_frame[3] [2]), .I2(n34066), 
            .I3(GND_net), .O(n17823));   // verilog/coms.v(126[12] 293[6])
    defparam i12994_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12_3_lut (.I0(bit_ctr[8]), .I1(n37227), .I2(n33701), .I3(GND_net), 
            .O(n31541));   // verilog/neopixel.v(35[12] 117[6])
    defparam i12_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 rem_4_unary_minus_2_add_3_5_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n30_adj_4979), .I3(n29571), .O(n30_adj_4854)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_unary_minus_2_add_3_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i12_3_lut_adj_1608 (.I0(bit_ctr[9]), .I1(n37226), .I2(n33701), 
            .I3(GND_net), .O(n31543));   // verilog/neopixel.v(35[12] 117[6])
    defparam i12_3_lut_adj_1608.LUT_INIT = 16'hacac;
    SB_LUT4 i12_3_lut_adj_1609 (.I0(bit_ctr[10]), .I1(n37225), .I2(n33701), 
            .I3(GND_net), .O(n31545));   // verilog/neopixel.v(35[12] 117[6])
    defparam i12_3_lut_adj_1609.LUT_INIT = 16'hacac;
    SB_LUT4 i30913_2_lut (.I0(displacement[21]), .I1(control_mode[0]), .I2(GND_net), 
            .I3(GND_net), .O(n37356));   // verilog/TinyFPGA_B.v(210[5] 214[10])
    defparam i30913_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 rem_4_add_1385_12_lut (.I0(GND_net), .I1(n2048), .I2(VCC_net), 
            .I3(n28241), .O(n2115)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1385_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mux_843_Mux_21_i1_3_lut (.I0(encoder0_position[21]), .I1(encoder1_position[21]), 
            .I2(control_mode[0]), .I3(GND_net), .O(n1_adj_4948));   // verilog/TinyFPGA_B.v(210[5] 214[10])
    defparam mux_843_Mux_21_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i19560_4_lut (.I0(n1_adj_4948), .I1(n34919), .I2(n37356), 
            .I3(control_mode[1]), .O(motor_state[21]));   // verilog/TinyFPGA_B.v(210[5] 214[10])
    defparam i19560_4_lut.LUT_INIT = 16'h3022;
    SB_LUT4 i30914_2_lut (.I0(displacement[22]), .I1(control_mode[0]), .I2(GND_net), 
            .I3(GND_net), .O(n37357));   // verilog/TinyFPGA_B.v(210[5] 214[10])
    defparam i30914_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 mux_843_Mux_22_i1_3_lut (.I0(encoder0_position[22]), .I1(encoder1_position[22]), 
            .I2(control_mode[0]), .I3(GND_net), .O(n1_adj_4949));   // verilog/TinyFPGA_B.v(210[5] 214[10])
    defparam mux_843_Mux_22_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2_4_lut (.I0(n32973), .I1(n16154), .I2(n3893), .I3(\FRAME_MATCHER.state_31__N_2566 [2]), 
            .O(n6_adj_4984));   // verilog/coms.v(126[12] 293[6])
    defparam i2_4_lut.LUT_INIT = 16'hbbba;
    SB_LUT4 i3_4_lut (.I0(\FRAME_MATCHER.state_31__N_2566 [2]), .I1(n6_adj_4984), 
            .I2(n34531), .I3(n32849), .O(n38508));   // verilog/coms.v(126[12] 293[6])
    defparam i3_4_lut.LUT_INIT = 16'hfefc;
    SB_LUT4 i13438_3_lut (.I0(\half_duty[0] [3]), .I1(half_duty_new[3]), 
            .I2(n1466), .I3(GND_net), .O(n18267));   // vhdl/pwm.vhd(59[5] 95[12])
    defparam i13438_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13436_3_lut (.I0(\half_duty[0] [1]), .I1(half_duty_new[1]), 
            .I2(n1466), .I3(GND_net), .O(n18265));   // vhdl/pwm.vhd(59[5] 95[12])
    defparam i13436_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i19561_4_lut (.I0(n1_adj_4949), .I1(n34919), .I2(n37357), 
            .I3(control_mode[1]), .O(motor_state[22]));   // verilog/TinyFPGA_B.v(210[5] 214[10])
    defparam i19561_4_lut.LUT_INIT = 16'h3022;
    SB_LUT4 i12_3_lut_adj_1610 (.I0(bit_ctr[11]), .I1(n37224), .I2(n33701), 
            .I3(GND_net), .O(n31547));   // verilog/neopixel.v(35[12] 117[6])
    defparam i12_3_lut_adj_1610.LUT_INIT = 16'hacac;
    SB_CARRY rem_4_unary_minus_2_add_3_5 (.CI(n29571), .I0(GND_net), .I1(n30_adj_4979), 
            .CO(n29572));
    SB_LUT4 i4_4_lut (.I0(control_mode[5]), .I1(control_mode[7]), .I2(control_mode[4]), 
            .I3(control_mode[6]), .O(n10_adj_4782));
    defparam i4_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i5_3_lut (.I0(control_mode[3]), .I1(n10_adj_4782), .I2(control_mode[2]), 
            .I3(GND_net), .O(n34919));
    defparam i5_3_lut.LUT_INIT = 16'hfefe;
    SB_CARRY rem_4_add_1385_12 (.CI(n28241), .I0(n2048), .I1(VCC_net), 
            .CO(n28242));
    SB_LUT4 i30915_2_lut (.I0(displacement[23]), .I1(control_mode[0]), .I2(GND_net), 
            .I3(GND_net), .O(n37358));   // verilog/TinyFPGA_B.v(210[5] 214[10])
    defparam i30915_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i12995_3_lut (.I0(Kp[3]), .I1(\data_in_frame[3] [3]), .I2(n34066), 
            .I3(GND_net), .O(n17824));   // verilog/coms.v(126[12] 293[6])
    defparam i12995_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mux_843_Mux_23_i1_3_lut (.I0(encoder0_position[23]), .I1(encoder1_position[23]), 
            .I2(control_mode[0]), .I3(GND_net), .O(n1_adj_4950));   // verilog/TinyFPGA_B.v(210[5] 214[10])
    defparam mux_843_Mux_23_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12996_3_lut (.I0(Kp[4]), .I1(\data_in_frame[3] [4]), .I2(n34066), 
            .I3(GND_net), .O(n17825));   // verilog/coms.v(126[12] 293[6])
    defparam i12996_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i19562_4_lut (.I0(n1_adj_4950), .I1(n34919), .I2(n37358), 
            .I3(control_mode[1]), .O(motor_state[23]));   // verilog/TinyFPGA_B.v(210[5] 214[10])
    defparam i19562_4_lut.LUT_INIT = 16'h3022;
    SB_LUT4 i12997_3_lut (.I0(Kp[5]), .I1(\data_in_frame[3] [5]), .I2(n34066), 
            .I3(GND_net), .O(n17826));   // verilog/coms.v(126[12] 293[6])
    defparam i12997_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12_3_lut_adj_1611 (.I0(bit_ctr[12]), .I1(n37369), .I2(n33701), 
            .I3(GND_net), .O(n31549));   // verilog/neopixel.v(35[12] 117[6])
    defparam i12_3_lut_adj_1611.LUT_INIT = 16'hacac;
    SB_LUT4 i12_3_lut_adj_1612 (.I0(bit_ctr[13]), .I1(n37368), .I2(n33701), 
            .I3(GND_net), .O(n31551));   // verilog/neopixel.v(35[12] 117[6])
    defparam i12_3_lut_adj_1612.LUT_INIT = 16'hacac;
    SB_LUT4 rem_4_add_1385_11_lut (.I0(GND_net), .I1(n2049), .I2(VCC_net), 
            .I3(n28240), .O(n2116)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1385_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i12_3_lut_adj_1613 (.I0(bit_ctr[14]), .I1(n37365), .I2(n33701), 
            .I3(GND_net), .O(n31553));   // verilog/neopixel.v(35[12] 117[6])
    defparam i12_3_lut_adj_1613.LUT_INIT = 16'hacac;
    SB_LUT4 i12998_3_lut (.I0(Kp[6]), .I1(\data_in_frame[3] [6]), .I2(n34066), 
            .I3(GND_net), .O(n17827));   // verilog/coms.v(126[12] 293[6])
    defparam i12998_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12_3_lut_adj_1614 (.I0(bit_ctr[15]), .I1(n37364), .I2(n33701), 
            .I3(GND_net), .O(n31555));   // verilog/neopixel.v(35[12] 117[6])
    defparam i12_3_lut_adj_1614.LUT_INIT = 16'hacac;
    SB_LUT4 add_582_13_lut (.I0(duty[11]), .I1(n38238), .I2(n14), .I3(n28166), 
            .O(pwm_setpoint_22__N_57[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_582_13_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_582_13 (.CI(n28166), .I0(n38238), .I1(n14), .CO(n28167));
    SB_CARRY rem_4_add_1385_11 (.CI(n28240), .I0(n2049), .I1(VCC_net), 
            .CO(n28241));
    SB_LUT4 rem_4_add_1385_10_lut (.I0(GND_net), .I1(n2050), .I2(VCC_net), 
            .I3(n28239), .O(n2117)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1385_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_582_12_lut (.I0(duty[10]), .I1(n38238), .I2(n15), .I3(n28165), 
            .O(pwm_setpoint_22__N_57[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_582_12_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY rem_4_add_1385_10 (.CI(n28239), .I0(n2050), .I1(VCC_net), 
            .CO(n28240));
    SB_LUT4 i12_3_lut_adj_1615 (.I0(bit_ctr[16]), .I1(n37363), .I2(n33701), 
            .I3(GND_net), .O(n31557));   // verilog/neopixel.v(35[12] 117[6])
    defparam i12_3_lut_adj_1615.LUT_INIT = 16'hacac;
    SB_CARRY add_582_12 (.CI(n28165), .I0(n38238), .I1(n15), .CO(n28166));
    SB_LUT4 rem_4_add_1385_9_lut (.I0(GND_net), .I1(n2051), .I2(VCC_net), 
            .I3(n28238), .O(n2118)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1385_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1385_9 (.CI(n28238), .I0(n2051), .I1(VCC_net), 
            .CO(n28239));
    SB_LUT4 add_582_11_lut (.I0(duty[9]), .I1(n38238), .I2(n16), .I3(n28164), 
            .O(pwm_setpoint_22__N_57[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_582_11_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 rem_4_add_1385_8_lut (.I0(GND_net), .I1(n2052), .I2(VCC_net), 
            .I3(n28237), .O(n2119)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1385_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i12_3_lut_adj_1616 (.I0(bit_ctr[17]), .I1(n37245), .I2(n33701), 
            .I3(GND_net), .O(n31559));   // verilog/neopixel.v(35[12] 117[6])
    defparam i12_3_lut_adj_1616.LUT_INIT = 16'hacac;
    SB_CARRY rem_4_add_1385_8 (.CI(n28237), .I0(n2052), .I1(VCC_net), 
            .CO(n28238));
    SB_LUT4 i12_3_lut_adj_1617 (.I0(bit_ctr[18]), .I1(n37362), .I2(n33701), 
            .I3(GND_net), .O(n31561));   // verilog/neopixel.v(35[12] 117[6])
    defparam i12_3_lut_adj_1617.LUT_INIT = 16'hacac;
    SB_CARRY add_582_11 (.CI(n28164), .I0(n38238), .I1(n16), .CO(n28165));
    SB_LUT4 rem_4_add_1385_7_lut (.I0(GND_net), .I1(n2053), .I2(VCC_net), 
            .I3(n28236), .O(n2120)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1385_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i12999_3_lut (.I0(Kp[7]), .I1(\data_in_frame[3] [7]), .I2(n34066), 
            .I3(GND_net), .O(n17828));   // verilog/coms.v(126[12] 293[6])
    defparam i12999_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12_3_lut_adj_1618 (.I0(bit_ctr[19]), .I1(n37361), .I2(n33701), 
            .I3(GND_net), .O(n31563));   // verilog/neopixel.v(35[12] 117[6])
    defparam i12_3_lut_adj_1618.LUT_INIT = 16'hacac;
    SB_CARRY rem_4_add_1385_7 (.CI(n28236), .I0(n2053), .I1(VCC_net), 
            .CO(n28237));
    SB_LUT4 i12_3_lut_adj_1619 (.I0(bit_ctr[20]), .I1(n37360), .I2(n33701), 
            .I3(GND_net), .O(n31565));   // verilog/neopixel.v(35[12] 117[6])
    defparam i12_3_lut_adj_1619.LUT_INIT = 16'hacac;
    SB_LUT4 add_582_10_lut (.I0(duty[8]), .I1(n38238), .I2(n17), .I3(n28163), 
            .O(pwm_setpoint_22__N_57[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_582_10_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 rem_4_add_1385_6_lut (.I0(GND_net), .I1(n2054), .I2(GND_net), 
            .I3(n28235), .O(n2121)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1385_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i13000_3_lut (.I0(Kp[8]), .I1(\data_in_frame[2] [0]), .I2(n34066), 
            .I3(GND_net), .O(n17829));   // verilog/coms.v(126[12] 293[6])
    defparam i13000_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12_3_lut_adj_1620 (.I0(bit_ctr[21]), .I1(n37359), .I2(n33701), 
            .I3(GND_net), .O(n31567));   // verilog/neopixel.v(35[12] 117[6])
    defparam i12_3_lut_adj_1620.LUT_INIT = 16'hacac;
    SB_LUT4 i12_3_lut_adj_1621 (.I0(bit_ctr[22]), .I1(n37335), .I2(n33701), 
            .I3(GND_net), .O(n31569));   // verilog/neopixel.v(35[12] 117[6])
    defparam i12_3_lut_adj_1621.LUT_INIT = 16'hacac;
    SB_LUT4 i12_3_lut_adj_1622 (.I0(bit_ctr[23]), .I1(n37330), .I2(n33701), 
            .I3(GND_net), .O(n31571));   // verilog/neopixel.v(35[12] 117[6])
    defparam i12_3_lut_adj_1622.LUT_INIT = 16'hacac;
    SB_LUT4 rem_4_unary_minus_2_add_3_4_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n31_adj_4980), .I3(n29570), .O(n31_adj_4853)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_unary_minus_2_add_3_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i12_3_lut_adj_1623 (.I0(bit_ctr[24]), .I1(n37309), .I2(n33701), 
            .I3(GND_net), .O(n31573));   // verilog/neopixel.v(35[12] 117[6])
    defparam i12_3_lut_adj_1623.LUT_INIT = 16'hacac;
    SB_CARRY rem_4_unary_minus_2_add_3_4 (.CI(n29570), .I0(GND_net), .I1(n31_adj_4980), 
            .CO(n29571));
    SB_LUT4 i12_3_lut_adj_1624 (.I0(bit_ctr[25]), .I1(n37308), .I2(n33701), 
            .I3(GND_net), .O(n31575));   // verilog/neopixel.v(35[12] 117[6])
    defparam i12_3_lut_adj_1624.LUT_INIT = 16'hacac;
    SB_LUT4 rem_4_unary_minus_2_add_3_3_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n32_adj_4981), .I3(n29569), .O(n32_adj_4852)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_unary_minus_2_add_3_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i12_3_lut_adj_1625 (.I0(bit_ctr[26]), .I1(n37304), .I2(n33701), 
            .I3(GND_net), .O(n31577));   // verilog/neopixel.v(35[12] 117[6])
    defparam i12_3_lut_adj_1625.LUT_INIT = 16'hacac;
    SB_CARRY rem_4_unary_minus_2_add_3_3 (.CI(n29569), .I0(GND_net), .I1(n32_adj_4981), 
            .CO(n29570));
    SB_LUT4 rem_4_unary_minus_2_add_3_2_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n33_adj_4982), .I3(VCC_net), .O(n33_adj_4851)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_unary_minus_2_add_3_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_unary_minus_2_add_3_2 (.CI(VCC_net), .I0(GND_net), .I1(n33_adj_4982), 
            .CO(n29569));
    SB_LUT4 i12_3_lut_adj_1626 (.I0(bit_ctr[27]), .I1(n37263), .I2(n33701), 
            .I3(GND_net), .O(n31583));   // verilog/neopixel.v(35[12] 117[6])
    defparam i12_3_lut_adj_1626.LUT_INIT = 16'hacac;
    SB_CARRY rem_4_add_1385_6 (.CI(n28235), .I0(n2054), .I1(GND_net), 
            .CO(n28236));
    SB_LUT4 rem_4_mux_3_i1_3_lut (.I0(communication_counter[0]), .I1(n33_adj_4851), 
            .I2(communication_counter[31]), .I3(GND_net), .O(n2865));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_mux_3_i1_3_lut.LUT_INIT = 16'h3535;
    SB_CARRY add_582_10 (.CI(n28163), .I0(n38238), .I1(n17), .CO(n28164));
    SB_LUT4 add_582_9_lut (.I0(duty[7]), .I1(n38238), .I2(n18), .I3(n28162), 
            .O(pwm_setpoint_22__N_57[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_582_9_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_582_9 (.CI(n28162), .I0(n38238), .I1(n18), .CO(n28163));
    SB_LUT4 i12_3_lut_adj_1627 (.I0(bit_ctr[28]), .I1(n37262), .I2(n33701), 
            .I3(GND_net), .O(n31585));   // verilog/neopixel.v(35[12] 117[6])
    defparam i12_3_lut_adj_1627.LUT_INIT = 16'hacac;
    SB_LUT4 i12_3_lut_adj_1628 (.I0(bit_ctr[29]), .I1(n37261), .I2(n33701), 
            .I3(GND_net), .O(n31587));   // verilog/neopixel.v(35[12] 117[6])
    defparam i12_3_lut_adj_1628.LUT_INIT = 16'hacac;
    SB_LUT4 i12_3_lut_adj_1629 (.I0(bit_ctr[30]), .I1(n37260), .I2(n33701), 
            .I3(GND_net), .O(n31589));   // verilog/neopixel.v(35[12] 117[6])
    defparam i12_3_lut_adj_1629.LUT_INIT = 16'hacac;
    SB_IO PIN_23_pad (.PACKAGE_PIN(PIN_23), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(PIN_23_c)) /* synthesis IO_FF_OUT=TRUE */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam PIN_23_pad.PIN_TYPE = 6'b011001;
    defparam PIN_23_pad.PULLUP = 1'b0;
    defparam PIN_23_pad.NEG_TRIGGER = 1'b0;
    defparam PIN_23_pad.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 i12_3_lut_adj_1630 (.I0(bit_ctr[0]), .I1(n37252), .I2(n33701), 
            .I3(GND_net), .O(n31591));   // verilog/neopixel.v(35[12] 117[6])
    defparam i12_3_lut_adj_1630.LUT_INIT = 16'hacac;
    SB_LUT4 add_582_8_lut (.I0(duty[6]), .I1(n38238), .I2(n19), .I3(n28161), 
            .O(pwm_setpoint_22__N_57[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_582_8_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 rem_4_add_1385_5_lut (.I0(GND_net), .I1(n2055), .I2(GND_net), 
            .I3(n28234), .O(n2122)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1385_5_lut.LUT_INIT = 16'hC33C;
    SB_DFF pwm_setpoint_i1 (.Q(pwm_setpoint[1]), .C(clk32MHz), .D(pwm_setpoint_22__N_57[1]));   // verilog/TinyFPGA_B.v(139[10] 152[6])
    SB_LUT4 encoder1_position_23__I_0_inv_0_i1_1_lut (.I0(encoder0_position[0]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n25_adj_4849));   // verilog/TinyFPGA_B.v(248[21:58])
    defparam encoder1_position_23__I_0_inv_0_i1_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder1_position_23__I_0_inv_0_i2_1_lut (.I0(encoder0_position[1]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n24_adj_4848));   // verilog/TinyFPGA_B.v(248[21:58])
    defparam encoder1_position_23__I_0_inv_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder1_position_23__I_0_inv_0_i3_1_lut (.I0(encoder0_position[2]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n23_adj_4847));   // verilog/TinyFPGA_B.v(248[21:58])
    defparam encoder1_position_23__I_0_inv_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder1_position_23__I_0_inv_0_i4_1_lut (.I0(encoder0_position[3]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n22_adj_4846));   // verilog/TinyFPGA_B.v(248[21:58])
    defparam encoder1_position_23__I_0_inv_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder1_position_23__I_0_inv_0_i5_1_lut (.I0(encoder0_position[4]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n21_adj_4845));   // verilog/TinyFPGA_B.v(248[21:58])
    defparam encoder1_position_23__I_0_inv_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder1_position_23__I_0_inv_0_i6_1_lut (.I0(encoder0_position[5]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n20_adj_4844));   // verilog/TinyFPGA_B.v(248[21:58])
    defparam encoder1_position_23__I_0_inv_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder1_position_23__I_0_inv_0_i7_1_lut (.I0(encoder0_position[6]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n19_adj_4843));   // verilog/TinyFPGA_B.v(248[21:58])
    defparam encoder1_position_23__I_0_inv_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder1_position_23__I_0_inv_0_i8_1_lut (.I0(encoder0_position[7]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n18_adj_4842));   // verilog/TinyFPGA_B.v(248[21:58])
    defparam encoder1_position_23__I_0_inv_0_i8_1_lut.LUT_INIT = 16'h5555;
    SB_IO PIN_24_pad (.PACKAGE_PIN(PIN_24), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(VCC_net));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam PIN_24_pad.PIN_TYPE = 6'b011001;
    defparam PIN_24_pad.PULLUP = 1'b0;
    defparam PIN_24_pad.NEG_TRIGGER = 1'b0;
    defparam PIN_24_pad.IO_STANDARD = "SB_LVCMOS";
    SB_GB_IO CLK_pad (.PACKAGE_PIN(CLK), .OUTPUT_ENABLE(VCC_net), .GLOBAL_BUFFER_OUTPUT(CLK_c));   // verilog/TinyFPGA_B.v(3[9:12])
    defparam CLK_pad.PIN_TYPE = 6'b000001;
    defparam CLK_pad.PULLUP = 1'b0;
    defparam CLK_pad.NEG_TRIGGER = 1'b0;
    defparam CLK_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO PIN_1_pad (.PACKAGE_PIN(PIN_1), .OUTPUT_ENABLE(VCC_net), .D_IN_0(PIN_1_c_1)) /* synthesis IO_FF_IN=TRUE */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam PIN_1_pad.PIN_TYPE = 6'b000001;
    defparam PIN_1_pad.PULLUP = 1'b0;
    defparam PIN_1_pad.NEG_TRIGGER = 1'b0;
    defparam PIN_1_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO PIN_2_pad (.PACKAGE_PIN(PIN_2), .OUTPUT_ENABLE(VCC_net), .D_IN_0(PIN_2_c_0)) /* synthesis IO_FF_IN=TRUE */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam PIN_2_pad.PIN_TYPE = 6'b000001;
    defparam PIN_2_pad.PULLUP = 1'b0;
    defparam PIN_2_pad.NEG_TRIGGER = 1'b0;
    defparam PIN_2_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO PIN_9_pad (.PACKAGE_PIN(PIN_9), .OUTPUT_ENABLE(VCC_net), .D_IN_0(PIN_9_c_1)) /* synthesis IO_FF_IN=TRUE */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam PIN_9_pad.PIN_TYPE = 6'b000001;
    defparam PIN_9_pad.PULLUP = 1'b0;
    defparam PIN_9_pad.NEG_TRIGGER = 1'b0;
    defparam PIN_9_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO PIN_10_pad (.PACKAGE_PIN(PIN_10), .OUTPUT_ENABLE(VCC_net), .D_IN_0(PIN_10_c_0)) /* synthesis IO_FF_IN=TRUE */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam PIN_10_pad.PIN_TYPE = 6'b000001;
    defparam PIN_10_pad.PULLUP = 1'b0;
    defparam PIN_10_pad.NEG_TRIGGER = 1'b0;
    defparam PIN_10_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO PIN_13_pad (.PACKAGE_PIN(PIN_13), .OUTPUT_ENABLE(VCC_net), .D_IN_0(PIN_13_c));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam PIN_13_pad.PIN_TYPE = 6'b000001;
    defparam PIN_13_pad.PULLUP = 1'b0;
    defparam PIN_13_pad.NEG_TRIGGER = 1'b0;
    defparam PIN_13_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO PIN_21_pad (.PACKAGE_PIN(PIN_21), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(PIN_21_c)) /* synthesis IO_FF_OUT=TRUE */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam PIN_21_pad.PIN_TYPE = 6'b011001;
    defparam PIN_21_pad.PULLUP = 1'b0;
    defparam PIN_21_pad.NEG_TRIGGER = 1'b0;
    defparam PIN_21_pad.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 encoder1_position_23__I_0_inv_0_i9_1_lut (.I0(encoder0_position[8]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n17_adj_4841));   // verilog/TinyFPGA_B.v(248[21:58])
    defparam encoder1_position_23__I_0_inv_0_i9_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 rem_4_add_2298_9_lut (.I0(n38197), .I1(n2_adj_4951), .I2(n3452), 
            .I3(n28714), .O(color_23__N_209[7])) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2298_9_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 rem_4_add_2298_8_lut (.I0(n38194), .I1(n2_adj_4951), .I2(n3453), 
            .I3(n28713), .O(color_23__N_209[6])) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2298_8_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY rem_4_add_2298_8 (.CI(n28713), .I0(n2_adj_4951), .I1(n3453), 
            .CO(n28714));
    SB_LUT4 rem_4_add_2298_7_lut (.I0(n38191), .I1(n2_adj_4951), .I2(n3454), 
            .I3(n28712), .O(color_23__N_209[5])) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2298_7_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY rem_4_add_2298_7 (.CI(n28712), .I0(n2_adj_4951), .I1(n3454), 
            .CO(n28713));
    SB_CARRY add_582_8 (.CI(n28161), .I0(n38238), .I1(n19), .CO(n28162));
    SB_CARRY rem_4_add_1385_5 (.CI(n28234), .I0(n2055), .I1(GND_net), 
            .CO(n28235));
    SB_LUT4 add_582_7_lut (.I0(duty[5]), .I1(n38238), .I2(n20_adj_4774), 
            .I3(n28160), .O(pwm_setpoint_22__N_57[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_582_7_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 rem_4_add_1385_4_lut (.I0(GND_net), .I1(n2056), .I2(VCC_net), 
            .I3(n28233), .O(n2123)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1385_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1385_4 (.CI(n28233), .I0(n2056), .I1(VCC_net), 
            .CO(n28234));
    SB_LUT4 rem_4_add_2298_6_lut (.I0(n38188), .I1(n2_adj_4951), .I2(n3455), 
            .I3(n28711), .O(color_23__N_209[4])) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2298_6_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY rem_4_add_2298_6 (.CI(n28711), .I0(n2_adj_4951), .I1(n3455), 
            .CO(n28712));
    SB_CARRY add_582_7 (.CI(n28160), .I0(n38238), .I1(n20_adj_4774), .CO(n28161));
    SB_LUT4 rem_4_mux_3_i2_3_lut (.I0(communication_counter[1]), .I1(n32_adj_4852), 
            .I2(communication_counter[31]), .I3(GND_net), .O(n3458));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_mux_3_i2_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 encoder1_position_23__I_0_inv_0_i10_1_lut (.I0(encoder0_position[9]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n16_adj_4840));   // verilog/TinyFPGA_B.v(248[21:58])
    defparam encoder1_position_23__I_0_inv_0_i10_1_lut.LUT_INIT = 16'h5555;
    SB_DFF pwm_setpoint_i2 (.Q(pwm_setpoint[2]), .C(clk32MHz), .D(pwm_setpoint_22__N_57[2]));   // verilog/TinyFPGA_B.v(139[10] 152[6])
    SB_LUT4 i23_3_lut_adj_1631 (.I0(bit_ctr[31]), .I1(n37244), .I2(n33701), 
            .I3(GND_net), .O(n31521));   // verilog/neopixel.v(35[12] 117[6])
    defparam i23_3_lut_adj_1631.LUT_INIT = 16'hacac;
    SB_LUT4 rem_4_i1737_3_lut (.I0(n2552), .I1(n2619), .I2(n2570), .I3(GND_net), 
            .O(n2651));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1737_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1738_3_lut (.I0(n2553), .I1(n2620), .I2(n2570), .I3(GND_net), 
            .O(n2652));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1738_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1736_3_lut (.I0(n2551), .I1(n2618), .I2(n2570), .I3(GND_net), 
            .O(n2650));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1736_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1727_3_lut (.I0(n2542), .I1(n2609), .I2(n2570), .I3(GND_net), 
            .O(n2641));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1727_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1731_3_lut (.I0(n2546), .I1(n2613), .I2(n2570), .I3(GND_net), 
            .O(n2645));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1731_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1723_3_lut (.I0(n2538), .I1(n2605), .I2(n2570), .I3(GND_net), 
            .O(n2637));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1723_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1732_3_lut (.I0(n2547), .I1(n2614), .I2(n2570), .I3(GND_net), 
            .O(n2646));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1732_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1724_3_lut (.I0(n2539), .I1(n2606), .I2(n2570), .I3(GND_net), 
            .O(n2638));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1724_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1729_3_lut (.I0(n2544), .I1(n2611), .I2(n2570), .I3(GND_net), 
            .O(n2643));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1729_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1739_3_lut (.I0(n2554), .I1(n2621), .I2(n2570), .I3(GND_net), 
            .O(n2653));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1739_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1730_3_lut (.I0(n2545), .I1(n2612), .I2(n2570), .I3(GND_net), 
            .O(n2644));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1730_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1728_3_lut (.I0(n2543), .I1(n2610), .I2(n2570), .I3(GND_net), 
            .O(n2642));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1728_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1743_3_lut (.I0(n2558), .I1(n2625), .I2(n2570), .I3(GND_net), 
            .O(n2657));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1743_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1741_3_lut (.I0(n2556), .I1(n2623), .I2(n2570), .I3(GND_net), 
            .O(n2655));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1741_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1740_3_lut (.I0(n2555), .I1(n2622), .I2(n2570), .I3(GND_net), 
            .O(n2654));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1740_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF pwm_setpoint_i3 (.Q(pwm_setpoint[3]), .C(clk32MHz), .D(pwm_setpoint_22__N_57[3]));   // verilog/TinyFPGA_B.v(139[10] 152[6])
    SB_DFF pwm_setpoint_i4 (.Q(pwm_setpoint[4]), .C(clk32MHz), .D(pwm_setpoint_22__N_57[4]));   // verilog/TinyFPGA_B.v(139[10] 152[6])
    SB_DFF pwm_setpoint_i5 (.Q(pwm_setpoint[5]), .C(clk32MHz), .D(pwm_setpoint_22__N_57[5]));   // verilog/TinyFPGA_B.v(139[10] 152[6])
    SB_DFF pwm_setpoint_i6 (.Q(pwm_setpoint[6]), .C(clk32MHz), .D(pwm_setpoint_22__N_57[6]));   // verilog/TinyFPGA_B.v(139[10] 152[6])
    SB_DFF pwm_setpoint_i7 (.Q(pwm_setpoint[7]), .C(clk32MHz), .D(pwm_setpoint_22__N_57[7]));   // verilog/TinyFPGA_B.v(139[10] 152[6])
    SB_DFF pwm_setpoint_i8 (.Q(pwm_setpoint[8]), .C(clk32MHz), .D(pwm_setpoint_22__N_57[8]));   // verilog/TinyFPGA_B.v(139[10] 152[6])
    SB_DFF pwm_setpoint_i9 (.Q(pwm_setpoint[9]), .C(clk32MHz), .D(pwm_setpoint_22__N_57[9]));   // verilog/TinyFPGA_B.v(139[10] 152[6])
    SB_DFF pwm_setpoint_i10 (.Q(pwm_setpoint[10]), .C(clk32MHz), .D(pwm_setpoint_22__N_57[10]));   // verilog/TinyFPGA_B.v(139[10] 152[6])
    SB_DFF pwm_setpoint_i11 (.Q(pwm_setpoint[11]), .C(clk32MHz), .D(pwm_setpoint_22__N_57[11]));   // verilog/TinyFPGA_B.v(139[10] 152[6])
    SB_DFF pwm_setpoint_i12 (.Q(pwm_setpoint[12]), .C(clk32MHz), .D(pwm_setpoint_22__N_57[12]));   // verilog/TinyFPGA_B.v(139[10] 152[6])
    SB_DFF pwm_setpoint_i13 (.Q(pwm_setpoint[13]), .C(clk32MHz), .D(pwm_setpoint_22__N_57[13]));   // verilog/TinyFPGA_B.v(139[10] 152[6])
    SB_DFF pwm_setpoint_i14 (.Q(pwm_setpoint[14]), .C(clk32MHz), .D(pwm_setpoint_22__N_57[14]));   // verilog/TinyFPGA_B.v(139[10] 152[6])
    SB_DFF pwm_setpoint_i15 (.Q(pwm_setpoint[15]), .C(clk32MHz), .D(pwm_setpoint_22__N_57[15]));   // verilog/TinyFPGA_B.v(139[10] 152[6])
    SB_DFF pwm_setpoint_i16 (.Q(pwm_setpoint[16]), .C(clk32MHz), .D(pwm_setpoint_22__N_57[16]));   // verilog/TinyFPGA_B.v(139[10] 152[6])
    SB_DFF pwm_setpoint_i17 (.Q(pwm_setpoint[17]), .C(clk32MHz), .D(pwm_setpoint_22__N_57[17]));   // verilog/TinyFPGA_B.v(139[10] 152[6])
    SB_DFF pwm_setpoint_i18 (.Q(pwm_setpoint[18]), .C(clk32MHz), .D(pwm_setpoint_22__N_57[18]));   // verilog/TinyFPGA_B.v(139[10] 152[6])
    SB_DFF pwm_setpoint_i19 (.Q(pwm_setpoint[19]), .C(clk32MHz), .D(pwm_setpoint_22__N_57[19]));   // verilog/TinyFPGA_B.v(139[10] 152[6])
    SB_DFF pwm_setpoint_i20 (.Q(pwm_setpoint[20]), .C(clk32MHz), .D(pwm_setpoint_22__N_57[20]));   // verilog/TinyFPGA_B.v(139[10] 152[6])
    SB_DFF pwm_setpoint_i21 (.Q(pwm_setpoint[21]), .C(clk32MHz), .D(pwm_setpoint_22__N_57[21]));   // verilog/TinyFPGA_B.v(139[10] 152[6])
    SB_DFF pwm_setpoint_i22 (.Q(pwm_setpoint[22]), .C(clk32MHz), .D(pwm_setpoint_22__N_57[22]));   // verilog/TinyFPGA_B.v(139[10] 152[6])
    SB_DFF displacement_i1 (.Q(displacement[1]), .C(clk32MHz), .D(displacement_23__N_80[1]));   // verilog/TinyFPGA_B.v(247[10] 249[6])
    SB_DFF displacement_i2 (.Q(displacement[2]), .C(clk32MHz), .D(displacement_23__N_80[2]));   // verilog/TinyFPGA_B.v(247[10] 249[6])
    SB_DFF displacement_i3 (.Q(displacement[3]), .C(clk32MHz), .D(displacement_23__N_80[3]));   // verilog/TinyFPGA_B.v(247[10] 249[6])
    SB_DFF displacement_i4 (.Q(displacement[4]), .C(clk32MHz), .D(displacement_23__N_80[4]));   // verilog/TinyFPGA_B.v(247[10] 249[6])
    SB_DFF displacement_i5 (.Q(displacement[5]), .C(clk32MHz), .D(displacement_23__N_80[5]));   // verilog/TinyFPGA_B.v(247[10] 249[6])
    SB_DFF displacement_i6 (.Q(displacement[6]), .C(clk32MHz), .D(displacement_23__N_80[6]));   // verilog/TinyFPGA_B.v(247[10] 249[6])
    SB_DFF displacement_i7 (.Q(displacement[7]), .C(clk32MHz), .D(displacement_23__N_80[7]));   // verilog/TinyFPGA_B.v(247[10] 249[6])
    SB_DFF displacement_i8 (.Q(displacement[8]), .C(clk32MHz), .D(displacement_23__N_80[8]));   // verilog/TinyFPGA_B.v(247[10] 249[6])
    SB_DFF displacement_i9 (.Q(displacement[9]), .C(clk32MHz), .D(displacement_23__N_80[9]));   // verilog/TinyFPGA_B.v(247[10] 249[6])
    SB_DFF displacement_i10 (.Q(displacement[10]), .C(clk32MHz), .D(displacement_23__N_80[10]));   // verilog/TinyFPGA_B.v(247[10] 249[6])
    SB_DFF displacement_i11 (.Q(displacement[11]), .C(clk32MHz), .D(displacement_23__N_80[11]));   // verilog/TinyFPGA_B.v(247[10] 249[6])
    SB_DFF displacement_i12 (.Q(displacement[12]), .C(clk32MHz), .D(displacement_23__N_80[12]));   // verilog/TinyFPGA_B.v(247[10] 249[6])
    SB_DFF displacement_i13 (.Q(displacement[13]), .C(clk32MHz), .D(displacement_23__N_80[13]));   // verilog/TinyFPGA_B.v(247[10] 249[6])
    SB_DFF displacement_i14 (.Q(displacement[14]), .C(clk32MHz), .D(displacement_23__N_80[14]));   // verilog/TinyFPGA_B.v(247[10] 249[6])
    SB_DFF displacement_i15 (.Q(displacement[15]), .C(clk32MHz), .D(displacement_23__N_80[15]));   // verilog/TinyFPGA_B.v(247[10] 249[6])
    SB_DFF displacement_i16 (.Q(displacement[16]), .C(clk32MHz), .D(displacement_23__N_80[16]));   // verilog/TinyFPGA_B.v(247[10] 249[6])
    SB_DFF displacement_i17 (.Q(displacement[17]), .C(clk32MHz), .D(displacement_23__N_80[17]));   // verilog/TinyFPGA_B.v(247[10] 249[6])
    SB_DFF displacement_i18 (.Q(displacement[18]), .C(clk32MHz), .D(displacement_23__N_80[18]));   // verilog/TinyFPGA_B.v(247[10] 249[6])
    SB_DFF displacement_i19 (.Q(displacement[19]), .C(clk32MHz), .D(displacement_23__N_80[19]));   // verilog/TinyFPGA_B.v(247[10] 249[6])
    SB_DFF displacement_i20 (.Q(displacement[20]), .C(clk32MHz), .D(displacement_23__N_80[20]));   // verilog/TinyFPGA_B.v(247[10] 249[6])
    SB_DFF displacement_i21 (.Q(displacement[21]), .C(clk32MHz), .D(displacement_23__N_80[21]));   // verilog/TinyFPGA_B.v(247[10] 249[6])
    SB_DFF displacement_i22 (.Q(displacement[22]), .C(clk32MHz), .D(displacement_23__N_80[22]));   // verilog/TinyFPGA_B.v(247[10] 249[6])
    SB_DFF displacement_i23 (.Q(displacement[23]), .C(clk32MHz), .D(displacement_23__N_80[23]));   // verilog/TinyFPGA_B.v(247[10] 249[6])
    SB_LUT4 rem_4_add_2298_5_lut (.I0(n38185), .I1(n2_adj_4951), .I2(n3456), 
            .I3(n28710), .O(color_23__N_209[3])) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2298_5_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY rem_4_add_2298_5 (.CI(n28710), .I0(n2_adj_4951), .I1(n3456), 
            .CO(n28711));
    SB_LUT4 rem_4_add_2298_4_lut (.I0(n38182), .I1(n2_adj_4951), .I2(n3457), 
            .I3(n28709), .O(color_23__N_209[2])) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2298_4_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY rem_4_add_2298_4 (.CI(n28709), .I0(n2_adj_4951), .I1(n3457), 
            .CO(n28710));
    SB_LUT4 rem_4_add_2298_3_lut (.I0(communication_counter[1]), .I1(n2_adj_4951), 
            .I2(n3458), .I3(n28708), .O(color_23__N_209[1])) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2298_3_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY rem_4_add_2298_3 (.CI(n28708), .I0(n2_adj_4951), .I1(n3458), 
            .CO(n28709));
    SB_LUT4 rem_4_add_2298_2_lut (.I0(communication_counter[0]), .I1(n2_adj_4951), 
            .I2(n2865), .I3(VCC_net), .O(color_23__N_209[0])) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2298_2_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 rem_4_add_1385_3_lut (.I0(GND_net), .I1(n2057), .I2(VCC_net), 
            .I3(n28232), .O(n2124)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1385_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1385_3 (.CI(n28232), .I0(n2057), .I1(VCC_net), 
            .CO(n28233));
    SB_CARRY rem_4_add_2298_2 (.CI(VCC_net), .I0(n2_adj_4951), .I1(n2865), 
            .CO(n28708));
    SB_LUT4 rem_4_add_1385_2_lut (.I0(GND_net), .I1(n2058), .I2(GND_net), 
            .I3(VCC_net), .O(n2125)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1385_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1385_2 (.CI(VCC_net), .I0(n2058), .I1(GND_net), 
            .CO(n28232));
    SB_LUT4 rem_4_add_2189_31_lut (.I0(n3263), .I1(n3230_adj_4902), .I2(VCC_net), 
            .I3(n28707), .O(n36391)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2189_31_lut.LUT_INIT = 16'h8228;
    SB_LUT4 rem_4_add_1452_19_lut (.I0(n2174), .I1(n2141), .I2(VCC_net), 
            .I3(n28231), .O(n2240)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1452_19_lut.LUT_INIT = 16'h8228;
    SB_LUT4 rem_4_add_2189_30_lut (.I0(GND_net), .I1(n3231_adj_4903), .I2(VCC_net), 
            .I3(n28706), .O(n3298)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2189_30_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i31500_1_lut (.I0(n3457), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n38182));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam i31500_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY rem_4_add_2189_30 (.CI(n28706), .I0(n3231_adj_4903), .I1(VCC_net), 
            .CO(n28707));
    SB_LUT4 rem_4_i2287_3_lut (.I0(n3358), .I1(n10395), .I2(n3362), .I3(GND_net), 
            .O(n3457));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i2287_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 rem_4_add_1452_18_lut (.I0(GND_net), .I1(n2142), .I2(VCC_net), 
            .I3(n28230), .O(n2209)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1452_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_2189_29_lut (.I0(GND_net), .I1(n3232_adj_4904), .I2(VCC_net), 
            .I3(n28705), .O(n3299)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2189_29_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_2189_29 (.CI(n28705), .I0(n3232_adj_4904), .I1(VCC_net), 
            .CO(n28706));
    SB_LUT4 rem_4_add_2189_28_lut (.I0(GND_net), .I1(n3233), .I2(VCC_net), 
            .I3(n28704), .O(n3300)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2189_28_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_2189_28 (.CI(n28704), .I0(n3233), .I1(VCC_net), 
            .CO(n28705));
    SB_LUT4 rem_4_add_2189_27_lut (.I0(GND_net), .I1(n3234), .I2(VCC_net), 
            .I3(n28703), .O(n3301)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2189_27_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_2189_27 (.CI(n28703), .I0(n3234), .I1(VCC_net), 
            .CO(n28704));
    SB_LUT4 add_582_6_lut (.I0(duty[4]), .I1(n38238), .I2(n21), .I3(n28159), 
            .O(pwm_setpoint_22__N_57[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_582_6_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 encoder1_position_23__I_0_inv_0_i11_1_lut (.I0(encoder0_position[10]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n15_adj_4839));   // verilog/TinyFPGA_B.v(248[21:58])
    defparam encoder1_position_23__I_0_inv_0_i11_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 rem_4_add_2189_26_lut (.I0(GND_net), .I1(n3235), .I2(VCC_net), 
            .I3(n28702), .O(n3302)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2189_26_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder1_position_23__I_0_inv_0_i12_1_lut (.I0(encoder0_position[11]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n14_adj_4838));   // verilog/TinyFPGA_B.v(248[21:58])
    defparam encoder1_position_23__I_0_inv_0_i12_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_582_6 (.CI(n28159), .I0(n38238), .I1(n21), .CO(n28160));
    SB_LUT4 encoder1_position_23__I_0_inv_0_i13_1_lut (.I0(encoder0_position[12]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n13_adj_4837));   // verilog/TinyFPGA_B.v(248[21:58])
    defparam encoder1_position_23__I_0_inv_0_i13_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder1_position_23__I_0_inv_0_i14_1_lut (.I0(encoder0_position[13]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n12_adj_4836));   // verilog/TinyFPGA_B.v(248[21:58])
    defparam encoder1_position_23__I_0_inv_0_i14_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY rem_4_add_1452_18 (.CI(n28230), .I0(n2142), .I1(VCC_net), 
            .CO(n28231));
    SB_CARRY rem_4_add_2189_26 (.CI(n28702), .I0(n3235), .I1(VCC_net), 
            .CO(n28703));
    SB_LUT4 add_582_5_lut (.I0(duty[3]), .I1(n38238), .I2(n22), .I3(n28158), 
            .O(pwm_setpoint_22__N_57[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_582_5_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_582_5 (.CI(n28158), .I0(n38238), .I1(n22), .CO(n28159));
    SB_LUT4 rem_4_add_2189_25_lut (.I0(GND_net), .I1(n3236), .I2(VCC_net), 
            .I3(n28701), .O(n3303)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2189_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder1_position_23__I_0_inv_0_i15_1_lut (.I0(encoder0_position[14]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n11_adj_4835));   // verilog/TinyFPGA_B.v(248[21:58])
    defparam encoder1_position_23__I_0_inv_0_i15_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_582_4_lut (.I0(duty[2]), .I1(n38238), .I2(n23), .I3(n28157), 
            .O(pwm_setpoint_22__N_57[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_582_4_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_582_4 (.CI(n28157), .I0(n38238), .I1(n23), .CO(n28158));
    SB_LUT4 add_582_3_lut (.I0(duty[1]), .I1(n38238), .I2(n24), .I3(n28156), 
            .O(pwm_setpoint_22__N_57[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_582_3_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 encoder1_position_23__I_0_inv_0_i16_1_lut (.I0(encoder0_position[15]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n10_adj_4809));   // verilog/TinyFPGA_B.v(248[21:58])
    defparam encoder1_position_23__I_0_inv_0_i16_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_582_3 (.CI(n28156), .I0(n38238), .I1(n24), .CO(n28157));
    SB_LUT4 encoder1_position_23__I_0_inv_0_i17_1_lut (.I0(encoder0_position[16]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n9_adj_4812));   // verilog/TinyFPGA_B.v(248[21:58])
    defparam encoder1_position_23__I_0_inv_0_i17_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder1_position_23__I_0_inv_0_i18_1_lut (.I0(encoder0_position[17]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n8_adj_4823));   // verilog/TinyFPGA_B.v(248[21:58])
    defparam encoder1_position_23__I_0_inv_0_i18_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder1_position_23__I_0_inv_0_i19_1_lut (.I0(encoder0_position[18]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n7_adj_4824));   // verilog/TinyFPGA_B.v(248[21:58])
    defparam encoder1_position_23__I_0_inv_0_i19_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder1_position_23__I_0_inv_0_i20_1_lut (.I0(encoder0_position[19]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n6_adj_4825));   // verilog/TinyFPGA_B.v(248[21:58])
    defparam encoder1_position_23__I_0_inv_0_i20_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i13449_4_lut (.I0(n5478), .I1(r_Clock_Count_adj_5048[0]), .I2(n321), 
            .I3(r_SM_Main_adj_5047[2]), .O(n18278));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i13449_4_lut.LUT_INIT = 16'h4450;
    SB_LUT4 encoder1_position_23__I_0_inv_0_i21_1_lut (.I0(encoder0_position[20]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n5_adj_4827));   // verilog/TinyFPGA_B.v(248[21:58])
    defparam encoder1_position_23__I_0_inv_0_i21_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder1_position_23__I_0_inv_0_i22_1_lut (.I0(encoder0_position[21]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n4_adj_4830));   // verilog/TinyFPGA_B.v(248[21:58])
    defparam encoder1_position_23__I_0_inv_0_i22_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder1_position_23__I_0_inv_0_i23_1_lut (.I0(encoder0_position[22]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n3_adj_4834));   // verilog/TinyFPGA_B.v(248[21:58])
    defparam encoder1_position_23__I_0_inv_0_i23_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder1_position_23__I_0_inv_0_i24_1_lut (.I0(encoder0_position[23]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n2));   // verilog/TinyFPGA_B.v(248[21:58])
    defparam encoder1_position_23__I_0_inv_0_i24_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i12854_4_lut (.I0(r_Rx_Data), .I1(rx_data[7]), .I2(n24193), 
            .I3(n16148), .O(n17683));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i12854_4_lut.LUT_INIT = 16'hccac;
    SB_LUT4 rem_4_mux_3_i10_3_lut (.I0(communication_counter[9]), .I1(n24_adj_4860), 
            .I2(communication_counter[31]), .I3(GND_net), .O(n2658));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_mux_3_i10_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1742_3_lut (.I0(n2557), .I1(n2624), .I2(n2570), .I3(GND_net), 
            .O(n2656));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1742_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i31025_3_lut (.I0(n2353), .I1(n2420), .I2(n2372), .I3(GND_net), 
            .O(n2452));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam i31025_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i31026_3_lut (.I0(n2452), .I1(n2519), .I2(n2471), .I3(GND_net), 
            .O(n2551));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam i31026_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i31027_3_lut (.I0(n2352), .I1(n2419), .I2(n2372), .I3(GND_net), 
            .O(n2451));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam i31027_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i31028_3_lut (.I0(n2451), .I1(n2518), .I2(n2471), .I3(GND_net), 
            .O(n2550));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam i31028_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1660_3_lut (.I0(n2443), .I1(n2510), .I2(n2471), .I3(GND_net), 
            .O(n2542));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1660_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12855_4_lut (.I0(r_Rx_Data), .I1(rx_data[6]), .I2(n24193), 
            .I3(n16143), .O(n17684));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i12855_4_lut.LUT_INIT = 16'hccac;
    SB_LUT4 i12856_4_lut (.I0(r_Rx_Data), .I1(rx_data[5]), .I2(n4_adj_4808), 
            .I3(n16148), .O(n17685));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i12856_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 rem_4_i1658_3_lut (.I0(n2441), .I1(n2508), .I2(n2471), .I3(GND_net), 
            .O(n2540));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1658_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1656_3_lut (.I0(n2439), .I1(n2506), .I2(n2471), .I3(GND_net), 
            .O(n2538));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1656_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1659_3_lut (.I0(n2442), .I1(n2509), .I2(n2471), .I3(GND_net), 
            .O(n2541));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1659_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1657_3_lut (.I0(n2440), .I1(n2507), .I2(n2471), .I3(GND_net), 
            .O(n2539));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1657_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1662_3_lut (.I0(n2445), .I1(n2512), .I2(n2471), .I3(GND_net), 
            .O(n2544));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1662_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1671_3_lut (.I0(n2454), .I1(n2521), .I2(n2471), .I3(GND_net), 
            .O(n2553));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1671_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1663_3_lut (.I0(n2446), .I1(n2513), .I2(n2471), .I3(GND_net), 
            .O(n2545));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1663_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i31009_3_lut (.I0(n2372), .I1(n2273), .I2(n2174), .I3(GND_net), 
            .O(n36654));
    defparam i31009_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i12857_4_lut (.I0(r_Rx_Data), .I1(rx_data[4]), .I2(n4_adj_4808), 
            .I3(n16143), .O(n17686));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i12857_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i31503_1_lut (.I0(n3456), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n38185));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam i31503_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i13174_4_lut (.I0(\data_out_frame[23] [6]), .I1(n4_adj_4909), 
            .I2(n17308), .I3(n33228), .O(n18003));   // verilog/coms.v(126[12] 293[6])
    defparam i13174_4_lut.LUT_INIT = 16'h3aca;
    SB_LUT4 rem_4_i2286_3_lut (.I0(n3357), .I1(n10394), .I2(n3362), .I3(GND_net), 
            .O(n3456));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i2286_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 i12858_4_lut (.I0(r_Rx_Data), .I1(rx_data[3]), .I2(n4_adj_4798), 
            .I3(n16148), .O(n17687));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i12858_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i13001_3_lut (.I0(Kp[9]), .I1(\data_in_frame[2] [1]), .I2(n34066), 
            .I3(GND_net), .O(n17830));   // verilog/coms.v(126[12] 293[6])
    defparam i13001_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13175_3_lut (.I0(control_mode[1]), .I1(\data_in_frame[1] [1]), 
            .I2(n5439), .I3(GND_net), .O(n18004));   // verilog/coms.v(126[12] 293[6])
    defparam i13175_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12859_4_lut (.I0(r_Rx_Data), .I1(rx_data[2]), .I2(n4_adj_4798), 
            .I3(n16143), .O(n17688));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i12859_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i12860_4_lut (.I0(r_Rx_Data), .I1(rx_data[1]), .I2(n4_adj_4822), 
            .I3(n16148), .O(n17689));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i12860_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 rem_4_unary_minus_2_inv_0_i23_1_lut (.I0(communication_counter[22]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n11_adj_4960));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_unary_minus_2_inv_0_i23_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 rem_4_unary_minus_2_inv_0_i24_1_lut (.I0(communication_counter[23]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n10_adj_4959));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_unary_minus_2_inv_0_i24_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i12861_3_lut (.I0(\data_in[0] [0]), .I1(\data_in[1] [0]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n17690));   // verilog/coms.v(126[12] 293[6])
    defparam i12861_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12862_3_lut (.I0(Kp[0]), .I1(\data_in_frame[3] [0]), .I2(n34066), 
            .I3(GND_net), .O(n17691));   // verilog/coms.v(126[12] 293[6])
    defparam i12862_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 rem_4_i1673_3_lut (.I0(n2456), .I1(n2523), .I2(n2471), .I3(GND_net), 
            .O(n2555));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1673_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1661_3_lut (.I0(n2444), .I1(n2511), .I2(n2471), .I3(GND_net), 
            .O(n2543));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1661_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1672_3_lut (.I0(n2455), .I1(n2522), .I2(n2471), .I3(GND_net), 
            .O(n2554));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1672_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i31040_3_lut (.I0(n2249), .I1(n2316), .I2(n2273), .I3(GND_net), 
            .O(n2348));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam i31040_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i31036_3_lut (.I0(n2252), .I1(n2319), .I2(n2273), .I3(GND_net), 
            .O(n2351));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam i31036_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1593_3_lut (.I0(n2344), .I1(n2411), .I2(n2372), .I3(GND_net), 
            .O(n2443));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1593_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1591_3_lut (.I0(n2342), .I1(n2409), .I2(n2372), .I3(GND_net), 
            .O(n2441));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1591_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12863_3_lut (.I0(Ki[0]), .I1(\data_in_frame[5] [0]), .I2(n34066), 
            .I3(GND_net), .O(n17692));   // verilog/coms.v(126[12] 293[6])
    defparam i12863_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_1632 (.I0(\FRAME_MATCHER.state_31__N_2566 [1]), .I1(n32849), 
            .I2(n33657), .I3(n16159), .O(n12));   // verilog/coms.v(126[12] 293[6])
    defparam i1_4_lut_adj_1632.LUT_INIT = 16'h8aaa;
    SB_LUT4 i12864_3_lut (.I0(setpoint[0]), .I1(n4996), .I2(n35492), .I3(GND_net), 
            .O(n17693));   // verilog/coms.v(126[12] 293[6])
    defparam i12864_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12865_3_lut (.I0(control_mode[0]), .I1(\data_in_frame[1] [0]), 
            .I2(n5439), .I3(GND_net), .O(n17694));   // verilog/coms.v(126[12] 293[6])
    defparam i12865_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12867_3_lut (.I0(PWMLimit[0]), .I1(\data_in_frame[10] [0]), 
            .I2(n5439), .I3(GND_net), .O(n17696));   // verilog/coms.v(126[12] 293[6])
    defparam i12867_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12868_3_lut (.I0(encoder0_position[0]), .I1(n3232), .I2(count_enable), 
            .I3(GND_net), .O(n17697));   // quad.v(35[10] 41[6])
    defparam i12868_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2_4_lut_adj_1633 (.I0(n12), .I1(n16159), .I2(n32973), .I3(n737), 
            .O(n34206));   // verilog/coms.v(126[12] 293[6])
    defparam i2_4_lut_adj_1633.LUT_INIT = 16'hfbfa;
    SB_LUT4 rem_4_i1592_3_lut (.I0(n2343), .I1(n2410), .I2(n2372), .I3(GND_net), 
            .O(n2442));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1592_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1590_3_lut (.I0(n2341), .I1(n2408), .I2(n2372), .I3(GND_net), 
            .O(n2440));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1590_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i31234_3_lut (.I0(n2351), .I1(n2418), .I2(n2372), .I3(GND_net), 
            .O(n2450));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam i31234_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1603_3_lut (.I0(n2354), .I1(n2421), .I2(n2372), .I3(GND_net), 
            .O(n2453));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1603_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1607_3_lut (.I0(n2358), .I1(n2425), .I2(n2372), .I3(GND_net), 
            .O(n2457));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1607_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1605_3_lut (.I0(n2356), .I1(n2423), .I2(n2372), .I3(GND_net), 
            .O(n2455));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1605_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1604_3_lut (.I0(n2355), .I1(n2422), .I2(n2372), .I3(GND_net), 
            .O(n2454));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1604_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12870_3_lut (.I0(encoder1_position[0]), .I1(n3182), .I2(count_enable_adj_4807), 
            .I3(GND_net), .O(n17699));   // quad.v(35[10] 41[6])
    defparam i12870_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13402_3_lut (.I0(encoder0_position[23]), .I1(n3209), .I2(count_enable), 
            .I3(GND_net), .O(n18231));   // quad.v(35[10] 41[6])
    defparam i13402_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12871_3_lut (.I0(quadB_debounced), .I1(reg_B[0]), .I2(n34970), 
            .I3(GND_net), .O(n17700));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(186[9] 190[16])
    defparam i12871_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 unary_minus_28_inv_0_i16_1_lut (.I0(duty[15]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n10));   // verilog/TinyFPGA_B.v(149[23:28])
    defparam unary_minus_28_inv_0_i16_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i12872_4_lut (.I0(r_SM_Main[2]), .I1(n1_adj_4923), .I2(n25070), 
            .I3(r_SM_Main[1]), .O(n17701));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i12872_4_lut.LUT_INIT = 16'h0544;
    SB_LUT4 rem_4_mux_3_i12_3_lut (.I0(communication_counter[11]), .I1(n22_adj_4862), 
            .I2(communication_counter[31]), .I3(GND_net), .O(n2458));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_mux_3_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1606_3_lut (.I0(n2357), .I1(n2424), .I2(n2372), .I3(GND_net), 
            .O(n2456));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1606_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i31318_3_lut (.I0(n2251), .I1(n2318), .I2(n2273), .I3(GND_net), 
            .O(n2350));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam i31318_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i31236_3_lut (.I0(n2350), .I1(n2417), .I2(n2372), .I3(GND_net), 
            .O(n2449));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam i31236_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i31238_3_lut (.I0(n2349), .I1(n2416), .I2(n2372), .I3(GND_net), 
            .O(n2448));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam i31238_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1528_3_lut (.I0(n2247), .I1(n2314), .I2(n2273), .I3(GND_net), 
            .O(n2346));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1528_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1596_3_lut (.I0(n2347), .I1(n2414), .I2(n2372), .I3(GND_net), 
            .O(n2446));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1596_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1595_3_lut (.I0(n2346), .I1(n2413), .I2(n2372), .I3(GND_net), 
            .O(n2445));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1595_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13401_3_lut (.I0(encoder0_position[22]), .I1(n3210), .I2(count_enable), 
            .I3(GND_net), .O(n18230));   // quad.v(35[10] 41[6])
    defparam i13401_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13400_3_lut (.I0(encoder0_position[21]), .I1(n3211), .I2(count_enable), 
            .I3(GND_net), .O(n18229));   // quad.v(35[10] 41[6])
    defparam i13400_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13399_3_lut (.I0(encoder0_position[20]), .I1(n3212), .I2(count_enable), 
            .I3(GND_net), .O(n18228));   // quad.v(35[10] 41[6])
    defparam i13399_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13398_3_lut (.I0(encoder0_position[19]), .I1(n3213), .I2(count_enable), 
            .I3(GND_net), .O(n18227));   // quad.v(35[10] 41[6])
    defparam i13398_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12876_3_lut (.I0(quadB_debounced_adj_4806), .I1(reg_B_adj_5056[0]), 
            .I2(n34971), .I3(GND_net), .O(n17705));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(186[9] 190[16])
    defparam i12876_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 rem_4_i1594_3_lut (.I0(n2345), .I1(n2412), .I2(n2372), .I3(GND_net), 
            .O(n2444));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1594_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1589_3_lut (.I0(n2340), .I1(n2407), .I2(n2372), .I3(GND_net), 
            .O(n2439));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1589_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_adj_1634 (.I0(n2439), .I1(n2438), .I2(GND_net), .I3(GND_net), 
            .O(n18_adj_4785));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam i1_2_lut_adj_1634.LUT_INIT = 16'heeee;
    SB_LUT4 i1_2_lut_adj_1635 (.I0(n2456), .I1(n2458), .I2(GND_net), .I3(GND_net), 
            .O(n36297));
    defparam i1_2_lut_adj_1635.LUT_INIT = 16'heeee;
    SB_LUT4 i1_4_lut_adj_1636 (.I0(n2454), .I1(n36297), .I2(n2455), .I3(n2457), 
            .O(n34007));
    defparam i1_4_lut_adj_1636.LUT_INIT = 16'ha080;
    SB_LUT4 i13_4_lut (.I0(n2452), .I1(n2453), .I2(n2450), .I3(n18_adj_4785), 
            .O(n30));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam i13_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i11_4_lut (.I0(n2444), .I1(n2445), .I2(n34007), .I3(n2446), 
            .O(n28_adj_4783));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam i11_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i12_4_lut (.I0(n2448), .I1(n2447), .I2(n2449), .I3(n2451), 
            .O(n29));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam i12_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i10_4_lut (.I0(n2440), .I1(n2442), .I2(n2441), .I3(n2443), 
            .O(n27_adj_4784));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam i10_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i16_4_lut (.I0(n27_adj_4784), .I1(n29), .I2(n28_adj_4783), 
            .I3(n30), .O(n2471));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam i16_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i13397_3_lut (.I0(encoder0_position[18]), .I1(n3214), .I2(count_enable), 
            .I3(GND_net), .O(n18226));   // quad.v(35[10] 41[6])
    defparam i13397_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13409_3_lut (.I0(encoder1_position[5]), .I1(n3177), .I2(count_enable_adj_4807), 
            .I3(GND_net), .O(n18238));   // quad.v(35[10] 41[6])
    defparam i13409_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13408_3_lut (.I0(encoder1_position[4]), .I1(n3178), .I2(count_enable_adj_4807), 
            .I3(GND_net), .O(n18237));   // quad.v(35[10] 41[6])
    defparam i13408_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12881_3_lut (.I0(\half_duty[0] [0]), .I1(half_duty_new[0]), 
            .I2(n1466), .I3(GND_net), .O(n17710));   // vhdl/pwm.vhd(59[5] 95[12])
    defparam i12881_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i31240_3_lut (.I0(n2348), .I1(n2415), .I2(n2372), .I3(GND_net), 
            .O(n2447));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam i31240_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1526_3_lut (.I0(n2245), .I1(n2312), .I2(n2273), .I3(GND_net), 
            .O(n2344));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1526_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1527_3_lut (.I0(n2246), .I1(n2313), .I2(n2273), .I3(GND_net), 
            .O(n2345));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1527_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1525_3_lut (.I0(n2244), .I1(n2311), .I2(n2273), .I3(GND_net), 
            .O(n2343));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1525_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1534_rep_48_3_lut (.I0(n2253), .I1(n2320), .I2(n2273), 
            .I3(GND_net), .O(n2352));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1534_rep_48_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1535_3_lut (.I0(n2254), .I1(n2321), .I2(n2273), .I3(GND_net), 
            .O(n2353));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1535_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1524_3_lut (.I0(n2243), .I1(n2310), .I2(n2273), .I3(GND_net), 
            .O(n2342));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1524_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1523_3_lut (.I0(n2242), .I1(n2309), .I2(n2273), .I3(GND_net), 
            .O(n2341));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1523_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1522_3_lut (.I0(n2241), .I1(n2308), .I2(n2273), .I3(GND_net), 
            .O(n2340));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1522_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1539_3_lut (.I0(n2258), .I1(n2325), .I2(n2273), .I3(GND_net), 
            .O(n2357));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1539_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13407_3_lut (.I0(encoder1_position[3]), .I1(n3179), .I2(count_enable_adj_4807), 
            .I3(GND_net), .O(n18236));   // quad.v(35[10] 41[6])
    defparam i13407_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1537_3_lut (.I0(n2256), .I1(n2323), .I2(n2273), .I3(GND_net), 
            .O(n2355));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1537_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1536_3_lut (.I0(n2255), .I1(n2322), .I2(n2273), .I3(GND_net), 
            .O(n2354));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1536_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_mux_3_i13_3_lut (.I0(communication_counter[12]), .I1(n21_adj_4863), 
            .I2(communication_counter[31]), .I3(GND_net), .O(n2358));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_mux_3_i13_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1538_3_lut (.I0(n2257), .I1(n2324), .I2(n2273), .I3(GND_net), 
            .O(n2356));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1538_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_adj_1637 (.I0(n2356), .I1(n2358), .I2(GND_net), .I3(GND_net), 
            .O(n36067));
    defparam i1_2_lut_adj_1637.LUT_INIT = 16'heeee;
    SB_LUT4 i1_4_lut_adj_1638 (.I0(n2354), .I1(n36067), .I2(n2355), .I3(n2357), 
            .O(n33944));
    defparam i1_4_lut_adj_1638.LUT_INIT = 16'ha080;
    SB_LUT4 i12_4_lut_adj_1639 (.I0(n2353), .I1(n2349), .I2(n2350), .I3(n2352), 
            .O(n28_adj_4905));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam i12_4_lut_adj_1639.LUT_INIT = 16'hfffe;
    SB_LUT4 i10_4_lut_adj_1640 (.I0(n2343), .I1(n2345), .I2(n2344), .I3(n33944), 
            .O(n26_adj_4907));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam i10_4_lut_adj_1640.LUT_INIT = 16'hfffe;
    SB_LUT4 i11_4_lut_adj_1641 (.I0(n2346), .I1(n2351), .I2(n2347), .I3(n2348), 
            .O(n27_adj_4906));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam i11_4_lut_adj_1641.LUT_INIT = 16'hfffe;
    SB_LUT4 i9_4_lut (.I0(n2340), .I1(n2341), .I2(n2339), .I3(n2342), 
            .O(n25_adj_4908));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam i9_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i15_4_lut (.I0(n25_adj_4908), .I1(n27_adj_4906), .I2(n26_adj_4907), 
            .I3(n28_adj_4905), .O(n2372));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam i15_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i31313_3_lut (.I0(n2250), .I1(n2317), .I2(n2273), .I3(GND_net), 
            .O(n2349));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam i31313_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i31232_3_lut (.I0(n2448), .I1(n2515), .I2(n2471), .I3(GND_net), 
            .O(n2547));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam i31232_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_unary_minus_2_inv_0_i25_1_lut (.I0(communication_counter[24]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n9_adj_4958));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_unary_minus_2_inv_0_i25_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 rem_4_i1664_3_lut (.I0(n2447), .I1(n2514), .I2(n2471), .I3(GND_net), 
            .O(n2546));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1664_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1670_3_lut (.I0(n2453), .I1(n2520), .I2(n2471), .I3(GND_net), 
            .O(n2552));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1670_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1466_rep_55_3_lut (.I0(n2220), .I1(n2319), .I2(n2273), 
            .I3(GND_net), .O(n36489));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1466_rep_55_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1533_rep_47_3_lut (.I0(n36489), .I1(n2418), .I2(n2372), 
            .I3(GND_net), .O(n36481));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1533_rep_47_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i31029_3_lut (.I0(n36481), .I1(n2153), .I2(n36654), .I3(GND_net), 
            .O(n37711));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam i31029_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i31030_3_lut (.I0(n37711), .I1(n2517), .I2(n2471), .I3(GND_net), 
            .O(n2549));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam i31030_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_mux_3_i11_3_lut (.I0(communication_counter[10]), .I1(n23_adj_4861), 
            .I2(communication_counter[31]), .I3(GND_net), .O(n2558));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_mux_3_i11_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1675_3_lut (.I0(n2458), .I1(n2525), .I2(n2471), .I3(GND_net), 
            .O(n2557));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1675_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1674_3_lut (.I0(n2457), .I1(n2524), .I2(n2471), .I3(GND_net), 
            .O(n2556));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1674_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_3_lut_adj_1642 (.I0(n2556), .I1(n2557), .I2(n2558), .I3(GND_net), 
            .O(n33949));
    defparam i1_3_lut_adj_1642.LUT_INIT = 16'hfefe;
    SB_LUT4 i10_4_lut_adj_1643 (.I0(n2538), .I1(n2540), .I2(n2537), .I3(n2542), 
            .O(n28_adj_4921));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam i10_4_lut_adj_1643.LUT_INIT = 16'hfffe;
    SB_LUT4 i13_4_lut_adj_1644 (.I0(n2549), .I1(n2552), .I2(n2546), .I3(n2547), 
            .O(n31_adj_4919));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam i13_4_lut_adj_1644.LUT_INIT = 16'hfffe;
    SB_LUT4 i4_4_lut_adj_1645 (.I0(n2554), .I1(n2543), .I2(n33949), .I3(n2555), 
            .O(n22_adj_4922));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam i4_4_lut_adj_1645.LUT_INIT = 16'heccc;
    SB_LUT4 i12_4_lut_adj_1646 (.I0(n2545), .I1(n2553), .I2(n2544), .I3(n2548), 
            .O(n30_adj_4920));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam i12_4_lut_adj_1646.LUT_INIT = 16'hfffe;
    SB_LUT4 i16_4_lut_adj_1647 (.I0(n31_adj_4919), .I1(n2550), .I2(n28_adj_4921), 
            .I3(n2551), .O(n34_adj_4918));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam i16_4_lut_adj_1647.LUT_INIT = 16'hfffe;
    SB_LUT4 rem_4_i1058_3_lut (.I0(n1553), .I1(n1620), .I2(n1580), .I3(GND_net), 
            .O(n1652));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1058_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13406_3_lut (.I0(encoder1_position[2]), .I1(n3180), .I2(count_enable_adj_4807), 
            .I3(GND_net), .O(n18235));   // quad.v(35[10] 41[6])
    defparam i13406_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13411_3_lut (.I0(encoder1_position[7]), .I1(n3175), .I2(count_enable_adj_4807), 
            .I3(GND_net), .O(n18240));   // quad.v(35[10] 41[6])
    defparam i13411_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13410_3_lut (.I0(encoder1_position[6]), .I1(n3176), .I2(count_enable_adj_4807), 
            .I3(GND_net), .O(n18239));   // quad.v(35[10] 41[6])
    defparam i13410_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1057_3_lut (.I0(n1552), .I1(n1619), .I2(n1580), .I3(GND_net), 
            .O(n1651));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1057_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13414_3_lut (.I0(encoder1_position[10]), .I1(n3172), .I2(count_enable_adj_4807), 
            .I3(GND_net), .O(n18243));   // quad.v(35[10] 41[6])
    defparam i13414_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13317_3_lut (.I0(\data_in_frame[17] [0]), .I1(rx_data[0]), 
            .I2(n32957), .I3(GND_net), .O(n18146));   // verilog/coms.v(126[12] 293[6])
    defparam i13317_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13413_3_lut (.I0(encoder1_position[9]), .I1(n3173), .I2(count_enable_adj_4807), 
            .I3(GND_net), .O(n18242));   // quad.v(35[10] 41[6])
    defparam i13413_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3_2_lut_adj_1648 (.I0(n2539), .I1(n2541), .I2(GND_net), .I3(GND_net), 
            .O(n21_adj_4924));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam i3_2_lut_adj_1648.LUT_INIT = 16'heeee;
    SB_LUT4 i17_4_lut (.I0(n21_adj_4924), .I1(n34_adj_4918), .I2(n30_adj_4920), 
            .I3(n22_adj_4922), .O(n2570));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam i17_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 rem_4_i1465_rep_60_3_lut (.I0(n2219), .I1(n2318), .I2(n2273), 
            .I3(GND_net), .O(n36494));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1465_rep_60_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1532_rep_51_3_lut (.I0(n36494), .I1(n2417), .I2(n2372), 
            .I3(GND_net), .O(n36485));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1532_rep_51_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i31031_3_lut (.I0(n36485), .I1(n2152), .I2(n36654), .I3(GND_net), 
            .O(n37713));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam i31031_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i31032_3_lut (.I0(n37713), .I1(n2516), .I2(n2471), .I3(GND_net), 
            .O(n2548));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam i31032_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1733_3_lut (.I0(n2548), .I1(n2615), .I2(n2570), .I3(GND_net), 
            .O(n2647));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1733_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1734_3_lut (.I0(n2549), .I1(n2616), .I2(n2570), .I3(GND_net), 
            .O(n2648));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1734_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1725_3_lut (.I0(n2540), .I1(n2607), .I2(n2570), .I3(GND_net), 
            .O(n2639));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1725_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1726_3_lut (.I0(n2541), .I1(n2608), .I2(n2570), .I3(GND_net), 
            .O(n2640));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1726_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11_4_lut_adj_1649 (.I0(n2640), .I1(n2639), .I2(n2648), .I3(n2647), 
            .O(n30_adj_4833));
    defparam i11_4_lut_adj_1649.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_adj_1650 (.I0(n2656), .I1(n2658), .I2(GND_net), .I3(GND_net), 
            .O(n36301));
    defparam i1_2_lut_adj_1650.LUT_INIT = 16'heeee;
    SB_LUT4 i1_4_lut_adj_1651 (.I0(n2654), .I1(n36301), .I2(n2655), .I3(n2657), 
            .O(n34021));
    defparam i1_4_lut_adj_1651.LUT_INIT = 16'ha080;
    SB_LUT4 i15_4_lut_adj_1652 (.I0(n2638), .I1(n30_adj_4833), .I2(n2649), 
            .I3(n2646), .O(n34_adj_4828));
    defparam i15_4_lut_adj_1652.LUT_INIT = 16'hfffe;
    SB_LUT4 i13_4_lut_adj_1653 (.I0(n2642), .I1(n2644), .I2(n2653), .I3(n2643), 
            .O(n32_adj_4831));
    defparam i13_4_lut_adj_1653.LUT_INIT = 16'hfffe;
    SB_LUT4 rem_4_add_1452_17_lut (.I0(GND_net), .I1(n2143), .I2(VCC_net), 
            .I3(n28229), .O(n2210)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1452_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_i2216_3_lut (.I0(n3255), .I1(n3322), .I2(n3263), .I3(GND_net), 
            .O(n3354));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i2216_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_unary_minus_2_inv_0_i26_1_lut (.I0(communication_counter[25]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n8_adj_4957));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_unary_minus_2_inv_0_i26_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i13412_3_lut (.I0(encoder1_position[8]), .I1(n3174), .I2(count_enable_adj_4807), 
            .I3(GND_net), .O(n18241));   // quad.v(35[10] 41[6])
    defparam i13412_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14_4_lut (.I0(n2637), .I1(n2645), .I2(n2636), .I3(n2641), 
            .O(n33_adj_4829));
    defparam i14_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i12_4_lut_adj_1654 (.I0(n2650), .I1(n2652), .I2(n34021), .I3(n2651), 
            .O(n31_adj_4832));
    defparam i12_4_lut_adj_1654.LUT_INIT = 16'hfffe;
    SB_LUT4 i18_4_lut_adj_1655 (.I0(n31_adj_4832), .I1(n33_adj_4829), .I2(n32_adj_4831), 
            .I3(n34_adj_4828), .O(n2669));
    defparam i18_4_lut_adj_1655.LUT_INIT = 16'hfffe;
    SB_LUT4 rem_4_i1735_3_lut (.I0(n2550), .I1(n2617), .I2(n2570), .I3(GND_net), 
            .O(n2649));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1735_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1463_3_lut (.I0(n2150), .I1(n2217), .I2(n2174), .I3(GND_net), 
            .O(n2249));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1463_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1459_3_lut (.I0(n2146), .I1(n2213), .I2(n2174), .I3(GND_net), 
            .O(n2245));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1459_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1457_3_lut (.I0(n2144), .I1(n2211), .I2(n2174), .I3(GND_net), 
            .O(n2243));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1457_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1458_3_lut (.I0(n2145), .I1(n2212), .I2(n2174), .I3(GND_net), 
            .O(n2244));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1458_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1456_3_lut (.I0(n2143), .I1(n2210), .I2(n2174), .I3(GND_net), 
            .O(n2242));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1456_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1455_3_lut (.I0(n2142), .I1(n2209), .I2(n2174), .I3(GND_net), 
            .O(n2241));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1455_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1465_3_lut (.I0(n2152), .I1(n2219), .I2(n2174), .I3(GND_net), 
            .O(n2251));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1465_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1461_3_lut (.I0(n2148), .I1(n2215), .I2(n2174), .I3(GND_net), 
            .O(n2247));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1461_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1469_3_lut (.I0(n2156), .I1(n2223), .I2(n2174), .I3(GND_net), 
            .O(n2255));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1469_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1460_3_lut (.I0(n2147), .I1(n2214), .I2(n2174), .I3(GND_net), 
            .O(n2246));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1460_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1468_3_lut (.I0(n2155), .I1(n2222), .I2(n2174), .I3(GND_net), 
            .O(n2254));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1468_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1467_3_lut (.I0(n2154), .I1(n2221), .I2(n2174), .I3(GND_net), 
            .O(n2253));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1467_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1464_3_lut (.I0(n2151), .I1(n2218), .I2(n2174), .I3(GND_net), 
            .O(n2250));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1464_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1466_3_lut (.I0(n2153), .I1(n2220), .I2(n2174), .I3(GND_net), 
            .O(n2252));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1466_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1390_3_lut (.I0(n2045), .I1(n2112), .I2(n2075), .I3(GND_net), 
            .O(n2144));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1390_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1389_3_lut (.I0(n2044), .I1(n2111), .I2(n2075), .I3(GND_net), 
            .O(n2143));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1389_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1388_3_lut (.I0(n2043), .I1(n2110), .I2(n2075), .I3(GND_net), 
            .O(n2142));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1388_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1395_3_lut (.I0(n2050), .I1(n2117), .I2(n2075), .I3(GND_net), 
            .O(n2149));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1395_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1396_3_lut (.I0(n2051), .I1(n2118), .I2(n2075), .I3(GND_net), 
            .O(n2150));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1396_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1397_3_lut (.I0(n2052), .I1(n2119), .I2(n2075), .I3(GND_net), 
            .O(n2151));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1397_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1399_3_lut (.I0(n2054), .I1(n2121), .I2(n2075), .I3(GND_net), 
            .O(n2153));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1399_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1398_3_lut (.I0(n2053), .I1(n2120), .I2(n2075), .I3(GND_net), 
            .O(n2152));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1398_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1394_3_lut (.I0(n2049), .I1(n2116), .I2(n2075), .I3(GND_net), 
            .O(n2148));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1394_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1401_3_lut (.I0(n2056), .I1(n2123), .I2(n2075), .I3(GND_net), 
            .O(n2155));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1401_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1393_3_lut (.I0(n2048), .I1(n2115), .I2(n2075), .I3(GND_net), 
            .O(n2147));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1393_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1400_3_lut (.I0(n2055), .I1(n2122), .I2(n2075), .I3(GND_net), 
            .O(n2154));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1400_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1392_3_lut (.I0(n2047), .I1(n2114), .I2(n2075), .I3(GND_net), 
            .O(n2146));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1392_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1391_3_lut (.I0(n2046), .I1(n2113), .I2(n2075), .I3(GND_net), 
            .O(n2145));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1391_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13176_3_lut (.I0(control_mode[2]), .I1(\data_in_frame[1] [2]), 
            .I2(n5439), .I3(GND_net), .O(n18005));   // verilog/coms.v(126[12] 293[6])
    defparam i13176_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_582_2_lut (.I0(duty[0]), .I1(n38238), .I2(n25_adj_4775), 
            .I3(VCC_net), .O(pwm_setpoint_22__N_57[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_582_2_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 rem_4_i1323_3_lut (.I0(n1946), .I1(n2013), .I2(n1976), .I3(GND_net), 
            .O(n2045));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1323_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1322_3_lut (.I0(n1945), .I1(n2012), .I2(n1976), .I3(GND_net), 
            .O(n2044));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1322_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1321_3_lut (.I0(n1944), .I1(n2011), .I2(n1976), .I3(GND_net), 
            .O(n2043));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1321_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1331_3_lut (.I0(n1954), .I1(n2021), .I2(n1976), .I3(GND_net), 
            .O(n2053));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1331_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1329_3_lut (.I0(n1952), .I1(n2019), .I2(n1976), .I3(GND_net), 
            .O(n2051));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1329_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1326_3_lut (.I0(n1949), .I1(n2016), .I2(n1976), .I3(GND_net), 
            .O(n2048));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1326_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1330_3_lut (.I0(n1953), .I1(n2020), .I2(n1976), .I3(GND_net), 
            .O(n2052));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1330_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1325_3_lut (.I0(n1948), .I1(n2015), .I2(n1976), .I3(GND_net), 
            .O(n2047));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1325_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1333_3_lut (.I0(n1956), .I1(n2023), .I2(n1976), .I3(GND_net), 
            .O(n2055));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1333_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1332_3_lut (.I0(n1955), .I1(n2022), .I2(n1976), .I3(GND_net), 
            .O(n2054));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1332_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1324_3_lut (.I0(n1947), .I1(n2014), .I2(n1976), .I3(GND_net), 
            .O(n2046));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1324_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1328_3_lut (.I0(n1951), .I1(n2018), .I2(n1976), .I3(GND_net), 
            .O(n2050));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1328_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1327_3_lut (.I0(n1950), .I1(n2017), .I2(n1976), .I3(GND_net), 
            .O(n2049));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1327_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1261_3_lut (.I0(n1852), .I1(n1919), .I2(n1877), .I3(GND_net), 
            .O(n1951));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1261_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1259_3_lut (.I0(n1850), .I1(n1917), .I2(n1877), .I3(GND_net), 
            .O(n1949));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1259_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1263_3_lut (.I0(n1854), .I1(n1921), .I2(n1877), .I3(GND_net), 
            .O(n1953));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1263_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1262_3_lut (.I0(n1853), .I1(n1920), .I2(n1877), .I3(GND_net), 
            .O(n1952));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1262_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1260_3_lut (.I0(n1851), .I1(n1918), .I2(n1877), .I3(GND_net), 
            .O(n1950));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1260_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1258_3_lut (.I0(n1849), .I1(n1916), .I2(n1877), .I3(GND_net), 
            .O(n1948));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1258_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_582_2 (.CI(VCC_net), .I0(n38238), .I1(n25_adj_4775), 
            .CO(n28156));
    SB_LUT4 rem_4_i1256_3_lut (.I0(n1847), .I1(n1914), .I2(n1877), .I3(GND_net), 
            .O(n1946));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1256_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1255_3_lut (.I0(n1846), .I1(n1913), .I2(n1877), .I3(GND_net), 
            .O(n1945));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1255_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1254_3_lut (.I0(n1845), .I1(n1912), .I2(n1877), .I3(GND_net), 
            .O(n1944));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1254_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1265_3_lut (.I0(n1856), .I1(n1923), .I2(n1877), .I3(GND_net), 
            .O(n1955));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1265_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1264_3_lut (.I0(n1855), .I1(n1922), .I2(n1877), .I3(GND_net), 
            .O(n1954));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1264_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1257_3_lut (.I0(n1848), .I1(n1915), .I2(n1877), .I3(GND_net), 
            .O(n1947));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1257_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_mux_3_i20_3_lut (.I0(communication_counter[19]), .I1(n14_adj_4870), 
            .I2(communication_counter[31]), .I3(GND_net), .O(n1658));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_mux_3_i20_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1131_3_lut (.I0(n1658), .I1(n1725), .I2(n1679), .I3(GND_net), 
            .O(n1757));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1131_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i785_3_lut (.I0(n1152), .I1(n1219), .I2(n1184), .I3(GND_net), 
            .O(n1251));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i785_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i852_3_lut (.I0(n1251), .I1(n1318), .I2(n1283), .I3(GND_net), 
            .O(n1350));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i852_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i919_3_lut (.I0(n1350), .I1(n1417), .I2(n1382), .I3(GND_net), 
            .O(n1449));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i919_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i986_3_lut (.I0(n1449), .I1(n1516), .I2(n1481), .I3(GND_net), 
            .O(n1548));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i986_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1053_3_lut (.I0(n1548), .I1(n1615), .I2(n1580), .I3(GND_net), 
            .O(n1647));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1053_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1120_3_lut (.I0(n1647), .I1(n1714), .I2(n1679), .I3(GND_net), 
            .O(n1746));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1120_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1187_3_lut (.I0(n1746), .I1(n1813), .I2(n1778), .I3(GND_net), 
            .O(n1845));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1187_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1193_3_lut (.I0(n1752), .I1(n1819), .I2(n1778), .I3(GND_net), 
            .O(n1851));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1193_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1194_3_lut (.I0(n1753), .I1(n1820), .I2(n1778), .I3(GND_net), 
            .O(n1852));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1194_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1195_3_lut (.I0(n1754), .I1(n1821), .I2(n1778), .I3(GND_net), 
            .O(n1853));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1195_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_mux_3_i21_3_lut (.I0(communication_counter[20]), .I1(n13_adj_4871), 
            .I2(communication_counter[31]), .I3(GND_net), .O(n1558));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_mux_3_i21_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1063_3_lut (.I0(n1558), .I1(n1625), .I2(n1580), .I3(GND_net), 
            .O(n1657));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1063_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i991_3_lut (.I0(n1454), .I1(n1521), .I2(n1481), .I3(GND_net), 
            .O(n1553));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i991_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13177_3_lut (.I0(control_mode[3]), .I1(\data_in_frame[1] [3]), 
            .I2(n5439), .I3(GND_net), .O(n18006));   // verilog/coms.v(126[12] 293[6])
    defparam i13177_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i990_3_lut (.I0(n1453), .I1(n1520), .I2(n1481), .I3(GND_net), 
            .O(n1552));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i990_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_mux_3_i19_3_lut (.I0(communication_counter[18]), .I1(n15_adj_4869), 
            .I2(communication_counter[31]), .I3(GND_net), .O(n1758));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_mux_3_i19_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1130_3_lut (.I0(n1657), .I1(n1724), .I2(n1679), .I3(GND_net), 
            .O(n1756));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1130_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1199_3_lut (.I0(n1758), .I1(n1825), .I2(n1778), .I3(GND_net), 
            .O(n1857));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1199_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1197_3_lut (.I0(n1756), .I1(n1823), .I2(n1778), .I3(GND_net), 
            .O(n1855));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1197_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1196_3_lut (.I0(n1755), .I1(n1822), .I2(n1778), .I3(GND_net), 
            .O(n1854));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1196_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1192_3_lut (.I0(n1751), .I1(n1818), .I2(n1778), .I3(GND_net), 
            .O(n1850));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1192_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1191_3_lut (.I0(n1750), .I1(n1817), .I2(n1778), .I3(GND_net), 
            .O(n1849));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1191_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_mux_3_i29_3_lut (.I0(communication_counter[28]), .I1(n5_adj_4879), 
            .I2(communication_counter[31]), .I3(GND_net), .O(n749));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_mux_3_i29_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i653_3_lut (.I0(n956), .I1(n1023), .I2(n986), .I3(GND_net), 
            .O(n1055));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i653_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i720_3_lut (.I0(n1055), .I1(n1122), .I2(n1085), .I3(GND_net), 
            .O(n1154));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i720_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i787_3_lut (.I0(n1154), .I1(n1221), .I2(n1184), .I3(GND_net), 
            .O(n1253));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i787_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i854_3_lut (.I0(n1253), .I1(n1320), .I2(n1283), .I3(GND_net), 
            .O(n1352));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i854_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i921_3_lut (.I0(n1352), .I1(n1419), .I2(n1382), .I3(GND_net), 
            .O(n1451));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i921_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i988_3_lut (.I0(n1451), .I1(n1518), .I2(n1481), .I3(GND_net), 
            .O(n1550));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i988_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1055_3_lut (.I0(n1550), .I1(n1617), .I2(n1580), .I3(GND_net), 
            .O(n1649));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1055_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i786_3_lut (.I0(n1153), .I1(n1220), .I2(n1184), .I3(GND_net), 
            .O(n1252));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i786_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i853_3_lut (.I0(n1252), .I1(n1319), .I2(n1283), .I3(GND_net), 
            .O(n1351));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i853_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i920_3_lut (.I0(n1351), .I1(n1418), .I2(n1382), .I3(GND_net), 
            .O(n1450));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i920_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i987_3_lut (.I0(n1450), .I1(n1517), .I2(n1481), .I3(GND_net), 
            .O(n1549));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i987_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1054_3_lut (.I0(n1549), .I1(n1616), .I2(n1580), .I3(GND_net), 
            .O(n1648));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1054_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i31506_1_lut (.I0(n3455), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n38188));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam i31506_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 rem_4_i2285_3_lut (.I0(n3356), .I1(n10393), .I2(n3362), .I3(GND_net), 
            .O(n3455));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i2285_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 i13178_3_lut (.I0(control_mode[4]), .I1(\data_in_frame[1] [4]), 
            .I2(n5439), .I3(GND_net), .O(n18007));   // verilog/coms.v(126[12] 293[6])
    defparam i13178_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY rem_4_add_1452_17 (.CI(n28229), .I0(n2143), .I1(VCC_net), 
            .CO(n28230));
    SB_LUT4 unary_minus_28_inv_0_i6_1_lut (.I0(duty[5]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n20_adj_4774));   // verilog/TinyFPGA_B.v(149[23:28])
    defparam unary_minus_28_inv_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i13179_3_lut (.I0(control_mode[5]), .I1(\data_in_frame[1] [5]), 
            .I2(n5439), .I3(GND_net), .O(n18008));   // verilog/coms.v(126[12] 293[6])
    defparam i13179_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_unary_minus_2_inv_0_i27_1_lut (.I0(communication_counter[26]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n7_adj_4956));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_unary_minus_2_inv_0_i27_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i13180_3_lut (.I0(control_mode[6]), .I1(\data_in_frame[1] [6]), 
            .I2(n5439), .I3(GND_net), .O(n18009));   // verilog/coms.v(126[12] 293[6])
    defparam i13180_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_unary_minus_2_inv_0_i28_1_lut (.I0(communication_counter[27]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n6_adj_4955));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_unary_minus_2_inv_0_i28_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 rem_4_i1121_3_lut (.I0(n1648), .I1(n1715), .I2(n1679), .I3(GND_net), 
            .O(n1747));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1121_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_mux_3_i28_3_lut (.I0(communication_counter[27]), .I1(n6_adj_4878), 
            .I2(communication_counter[31]), .I3(GND_net), .O(n855));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_mux_3_i28_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i654_3_lut (.I0(n957), .I1(n1024), .I2(n986), .I3(GND_net), 
            .O(n1056));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i654_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i721_3_lut (.I0(n1056), .I1(n1123), .I2(n1085), .I3(GND_net), 
            .O(n1155));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i721_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i788_3_lut (.I0(n1155), .I1(n1222), .I2(n1184), .I3(GND_net), 
            .O(n1254));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i788_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i855_3_lut (.I0(n1254), .I1(n1321), .I2(n1283), .I3(GND_net), 
            .O(n1353));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i855_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i922_3_lut (.I0(n1353), .I1(n1420), .I2(n1382), .I3(GND_net), 
            .O(n1452));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i922_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i989_3_lut (.I0(n1452), .I1(n1519), .I2(n1481), .I3(GND_net), 
            .O(n1551));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i989_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_mux_3_i23_3_lut (.I0(communication_counter[22]), .I1(n11_adj_4873), 
            .I2(communication_counter[31]), .I3(GND_net), .O(n1358));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_mux_3_i23_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i927_3_lut (.I0(n1358), .I1(n1425), .I2(n1382), .I3(GND_net), 
            .O(n1457));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i927_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i994_3_lut (.I0(n1457), .I1(n1524), .I2(n1481), .I3(GND_net), 
            .O(n1556));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i994_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1061_3_lut (.I0(n1556), .I1(n1623), .I2(n1580), .I3(GND_net), 
            .O(n1655));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1061_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_mux_3_i22_3_lut (.I0(communication_counter[21]), .I1(n12_adj_4872), 
            .I2(communication_counter[31]), .I3(GND_net), .O(n1458));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_mux_3_i22_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i995_3_lut (.I0(n1458), .I1(n1525), .I2(n1481), .I3(GND_net), 
            .O(n1557));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i995_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1062_3_lut (.I0(n1557), .I1(n1624), .I2(n1580), .I3(GND_net), 
            .O(n1656));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1062_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1056_3_lut (.I0(n1551), .I1(n1618), .I2(n1580), .I3(GND_net), 
            .O(n1650));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1056_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1129_3_lut (.I0(n1656), .I1(n1723), .I2(n1679), .I3(GND_net), 
            .O(n1755));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1129_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1123_3_lut (.I0(n1650), .I1(n1717), .I2(n1679), .I3(GND_net), 
            .O(n1749));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1123_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1128_3_lut (.I0(n1655), .I1(n1722), .I2(n1679), .I3(GND_net), 
            .O(n1754));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1128_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i31509_1_lut (.I0(n3454), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n38191));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam i31509_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 rem_4_i2284_3_lut (.I0(n3355), .I1(n10392), .I2(n3362), .I3(GND_net), 
            .O(n3454));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i2284_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 i13416_3_lut (.I0(encoder1_position[12]), .I1(n3170), .I2(count_enable_adj_4807), 
            .I3(GND_net), .O(n18245));   // quad.v(35[10] 41[6])
    defparam i13416_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13415_3_lut (.I0(encoder1_position[11]), .I1(n3171), .I2(count_enable_adj_4807), 
            .I3(GND_net), .O(n18244));   // quad.v(35[10] 41[6])
    defparam i13415_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13418_3_lut (.I0(encoder1_position[14]), .I1(n3168), .I2(count_enable_adj_4807), 
            .I3(GND_net), .O(n18247));   // quad.v(35[10] 41[6])
    defparam i13418_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13417_3_lut (.I0(encoder1_position[13]), .I1(n3169), .I2(count_enable_adj_4807), 
            .I3(GND_net), .O(n18246));   // quad.v(35[10] 41[6])
    defparam i13417_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_mux_3_i31_3_lut (.I0(communication_counter[30]), .I1(n3_adj_4881), 
            .I2(communication_counter[31]), .I3(GND_net), .O(n852));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_mux_3_i31_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_3_lut_adj_1656 (.I0(n957), .I1(n956), .I2(n958), .I3(GND_net), 
            .O(n33879));
    defparam i1_3_lut_adj_1656.LUT_INIT = 16'hfefe;
    SB_LUT4 i20066_4_lut (.I0(n954), .I1(n953), .I2(n33879), .I3(n955), 
            .O(n986));
    defparam i20066_4_lut.LUT_INIT = 16'heccc;
    SB_LUT4 i1_3_lut_adj_1657 (.I0(n1056), .I1(n1057), .I2(n1058), .I3(GND_net), 
            .O(n33877));
    defparam i1_3_lut_adj_1657.LUT_INIT = 16'hfefe;
    SB_LUT4 i1_2_lut_adj_1658 (.I0(n1054), .I1(n1055), .I2(GND_net), .I3(GND_net), 
            .O(n35913));
    defparam i1_2_lut_adj_1658.LUT_INIT = 16'h8888;
    SB_LUT4 i1_4_lut_adj_1659 (.I0(n1052), .I1(n35913), .I2(n1053), .I3(n33877), 
            .O(n1085));
    defparam i1_4_lut_adj_1659.LUT_INIT = 16'hfefa;
    SB_LUT4 rem_4_i651_3_lut (.I0(n954), .I1(n1021), .I2(n986), .I3(GND_net), 
            .O(n1053));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i651_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i719_3_lut (.I0(n1054), .I1(n1121), .I2(n1085), .I3(GND_net), 
            .O(n1153));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i719_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i718_3_lut (.I0(n1053), .I1(n1120), .I2(n1085), .I3(GND_net), 
            .O(n1152));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i718_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_adj_1660 (.I0(n1156), .I1(n1158), .I2(GND_net), .I3(GND_net), 
            .O(n35917));
    defparam i1_2_lut_adj_1660.LUT_INIT = 16'heeee;
    SB_LUT4 i1_4_lut_adj_1661 (.I0(n1154), .I1(n35917), .I2(n1155), .I3(n1157), 
            .O(n33873));
    defparam i1_4_lut_adj_1661.LUT_INIT = 16'ha080;
    SB_LUT4 i3_4_lut_adj_1662 (.I0(n33873), .I1(n1152), .I2(n1151), .I3(n1153), 
            .O(n1184));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam i3_4_lut_adj_1662.LUT_INIT = 16'hfffe;
    SB_LUT4 rem_4_mux_3_i25_3_lut (.I0(communication_counter[24]), .I1(n9_adj_4875), 
            .I2(communication_counter[31]), .I3(GND_net), .O(n1158));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_mux_3_i25_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i791_3_lut (.I0(n1158), .I1(n1225), .I2(n1184), .I3(GND_net), 
            .O(n1257));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i791_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i858_3_lut (.I0(n1257), .I1(n1324), .I2(n1283), .I3(GND_net), 
            .O(n1356));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i858_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i925_3_lut (.I0(n1356), .I1(n1423), .I2(n1382), .I3(GND_net), 
            .O(n1455));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i925_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i992_3_lut (.I0(n1455), .I1(n1522), .I2(n1481), .I3(GND_net), 
            .O(n1554));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i992_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1059_3_lut (.I0(n1554), .I1(n1621), .I2(n1580), .I3(GND_net), 
            .O(n1653));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1059_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_3_lut_adj_1663 (.I0(n1256), .I1(n1257), .I2(n1258), .I3(GND_net), 
            .O(n33871));
    defparam i1_3_lut_adj_1663.LUT_INIT = 16'hfefe;
    SB_LUT4 i1_4_lut_adj_1664 (.I0(n1254), .I1(n1250), .I2(n33871), .I3(n1255), 
            .O(n6_adj_4987));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam i1_4_lut_adj_1664.LUT_INIT = 16'heccc;
    SB_LUT4 i4_4_lut_adj_1665 (.I0(n1251), .I1(n1253), .I2(n1252), .I3(n6_adj_4987), 
            .O(n1283));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam i4_4_lut_adj_1665.LUT_INIT = 16'hfffe;
    SB_LUT4 rem_4_mux_3_i24_3_lut (.I0(communication_counter[23]), .I1(n10_adj_4874), 
            .I2(communication_counter[31]), .I3(GND_net), .O(n1258));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_mux_3_i24_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_add_1452_16_lut (.I0(GND_net), .I1(n2144), .I2(VCC_net), 
            .I3(n28228), .O(n2211)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1452_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i13420_3_lut (.I0(encoder1_position[16]), .I1(n3166), .I2(count_enable_adj_4807), 
            .I3(GND_net), .O(n18249));   // quad.v(35[10] 41[6])
    defparam i13420_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i31512_1_lut (.I0(n3453), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n38194));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam i31512_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 rem_4_i2283_3_lut (.I0(n3354), .I1(n10391), .I2(n3362), .I3(GND_net), 
            .O(n3453));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i2283_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 rem_4_unary_minus_2_inv_0_i29_1_lut (.I0(communication_counter[28]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n5_adj_4954));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_unary_minus_2_inv_0_i29_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1_3_lut_adj_1666 (.I0(n1356), .I1(n1357), .I2(n1358), .I3(GND_net), 
            .O(n33867));
    defparam i1_3_lut_adj_1666.LUT_INIT = 16'hfefe;
    SB_LUT4 i2_4_lut_adj_1667 (.I0(n1351), .I1(n1354), .I2(n33867), .I3(n1355), 
            .O(n8_adj_4985));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam i2_4_lut_adj_1667.LUT_INIT = 16'heaaa;
    SB_LUT4 i1_2_lut_adj_1668 (.I0(n1350), .I1(n1349), .I2(GND_net), .I3(GND_net), 
            .O(n7_adj_4986));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam i1_2_lut_adj_1668.LUT_INIT = 16'heeee;
    SB_LUT4 i5_4_lut (.I0(n1352), .I1(n7_adj_4986), .I2(n1353), .I3(n8_adj_4985), 
            .O(n1382));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam i5_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 rem_4_i859_3_lut (.I0(n1258), .I1(n1325), .I2(n1283), .I3(GND_net), 
            .O(n1357));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i859_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_adj_1669 (.I0(n1456), .I1(n1458), .I2(GND_net), .I3(GND_net), 
            .O(n36011));
    defparam i1_2_lut_adj_1669.LUT_INIT = 16'heeee;
    SB_LUT4 i1_4_lut_adj_1670 (.I0(n1454), .I1(n36011), .I2(n1455), .I3(n1457), 
            .O(n33901));
    defparam i1_4_lut_adj_1670.LUT_INIT = 16'ha080;
    SB_LUT4 i5_4_lut_adj_1671 (.I0(n33901), .I1(n1451), .I2(n1450), .I3(n1452), 
            .O(n12_adj_4983));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam i5_4_lut_adj_1671.LUT_INIT = 16'hfffe;
    SB_LUT4 i6_4_lut (.I0(n1453), .I1(n12_adj_4983), .I2(n1449), .I3(n1448), 
            .O(n1481));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam i6_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 rem_4_i926_3_lut (.I0(n1357), .I1(n1424), .I2(n1382), .I3(GND_net), 
            .O(n1456));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i926_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_3_lut_adj_1672 (.I0(n1556), .I1(n1557), .I2(n1558), .I3(GND_net), 
            .O(n33898));
    defparam i1_3_lut_adj_1672.LUT_INIT = 16'hfefe;
    SB_LUT4 i3_4_lut_adj_1673 (.I0(n1554), .I1(n1551), .I2(n33898), .I3(n1555), 
            .O(n11_adj_4796));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam i3_4_lut_adj_1673.LUT_INIT = 16'heccc;
    SB_LUT4 i5_4_lut_adj_1674 (.I0(n1548), .I1(n1549), .I2(n1547), .I3(n1550), 
            .O(n13_adj_4795));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam i5_4_lut_adj_1674.LUT_INIT = 16'hfffe;
    SB_LUT4 i7_4_lut (.I0(n13_adj_4795), .I1(n11_adj_4796), .I2(n1553), 
            .I3(n1552), .O(n1580));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam i7_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 rem_4_i993_3_lut (.I0(n1456), .I1(n1523), .I2(n1481), .I3(GND_net), 
            .O(n1555));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i993_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_adj_1675 (.I0(n1647), .I1(n1646), .I2(GND_net), .I3(GND_net), 
            .O(n10_adj_5003));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam i1_2_lut_adj_1675.LUT_INIT = 16'heeee;
    SB_LUT4 i1_3_lut_adj_1676 (.I0(n1656), .I1(n1657), .I2(n1658), .I3(GND_net), 
            .O(n33917));
    defparam i1_3_lut_adj_1676.LUT_INIT = 16'hfefe;
    SB_LUT4 i7_4_lut_adj_1677 (.I0(n1653), .I1(n1652), .I2(n1651), .I3(n10_adj_5003), 
            .O(n16_adj_5001));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam i7_4_lut_adj_1677.LUT_INIT = 16'hfffe;
    SB_LUT4 i2_4_lut_adj_1678 (.I0(n1648), .I1(n1654), .I2(n33917), .I3(n1655), 
            .O(n11_adj_5002));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam i2_4_lut_adj_1678.LUT_INIT = 16'heaaa;
    SB_LUT4 i8_4_lut (.I0(n11_adj_5002), .I1(n16_adj_5001), .I2(n1649), 
            .I3(n1650), .O(n1679));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam i8_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 rem_4_i1060_3_lut (.I0(n1555), .I1(n1622), .I2(n1580), .I3(GND_net), 
            .O(n1654));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1060_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1125_3_lut (.I0(n1652), .I1(n1719), .I2(n1679), .I3(GND_net), 
            .O(n1751));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1125_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1127_3_lut (.I0(n1654), .I1(n1721), .I2(n1679), .I3(GND_net), 
            .O(n1753));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1127_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1124_3_lut (.I0(n1651), .I1(n1718), .I2(n1679), .I3(GND_net), 
            .O(n1750));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1124_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13181_3_lut (.I0(control_mode[7]), .I1(\data_in_frame[1] [7]), 
            .I2(n5439), .I3(GND_net), .O(n18010));   // verilog/coms.v(126[12] 293[6])
    defparam i13181_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY rem_4_add_2189_25 (.CI(n28701), .I0(n3236), .I1(VCC_net), 
            .CO(n28702));
    SB_LUT4 i13419_3_lut (.I0(encoder1_position[15]), .I1(n3167), .I2(count_enable_adj_4807), 
            .I3(GND_net), .O(n18248));   // quad.v(35[10] 41[6])
    defparam i13419_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i2208_3_lut (.I0(n3247), .I1(n3314), .I2(n3263), .I3(GND_net), 
            .O(n3346));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i2208_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i2207_3_lut (.I0(n3246), .I1(n3313), .I2(n3263), .I3(GND_net), 
            .O(n3345));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i2207_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1126_3_lut (.I0(n1653), .I1(n1720), .I2(n1679), .I3(GND_net), 
            .O(n1752));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1126_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i6_4_lut_adj_1679 (.I0(n1746), .I1(n1747), .I2(n1745), .I3(n1748), 
            .O(n16_adj_4998));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam i6_4_lut_adj_1679.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_3_lut_adj_1680 (.I0(n1756), .I1(n1757), .I2(n1758), .I3(GND_net), 
            .O(n33909));
    defparam i1_3_lut_adj_1680.LUT_INIT = 16'hfefe;
    SB_LUT4 i8_3_lut (.I0(n1753), .I1(n16_adj_4998), .I2(n1751), .I3(GND_net), 
            .O(n18_adj_4997));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam i8_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i3_4_lut_adj_1681 (.I0(n1754), .I1(n1749), .I2(n33909), .I3(n1755), 
            .O(n13_adj_4999));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam i3_4_lut_adj_1681.LUT_INIT = 16'heccc;
    SB_LUT4 i9_4_lut_adj_1682 (.I0(n13_adj_4999), .I1(n18_adj_4997), .I2(n1752), 
            .I3(n1750), .O(n1778));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam i9_4_lut_adj_1682.LUT_INIT = 16'hfffe;
    SB_LUT4 rem_4_i1122_3_lut (.I0(n1649), .I1(n1716), .I2(n1679), .I3(GND_net), 
            .O(n1748));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1122_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1190_3_lut (.I0(n1749), .I1(n1816), .I2(n1778), .I3(GND_net), 
            .O(n1848));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1190_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1189_3_lut (.I0(n1748), .I1(n1815), .I2(n1778), .I3(GND_net), 
            .O(n1847));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1189_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1188_3_lut (.I0(n1747), .I1(n1814), .I2(n1778), .I3(GND_net), 
            .O(n1846));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1188_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1198_3_lut (.I0(n1757), .I1(n1824), .I2(n1778), .I3(GND_net), 
            .O(n1856));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1198_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_adj_1683 (.I0(n1856), .I1(n1858), .I2(GND_net), .I3(GND_net), 
            .O(n36177));
    defparam i1_2_lut_adj_1683.LUT_INIT = 16'heeee;
    SB_LUT4 i1_4_lut_adj_1684 (.I0(n1854), .I1(n36177), .I2(n1855), .I3(n1857), 
            .O(n33942));
    defparam i1_4_lut_adj_1684.LUT_INIT = 16'ha080;
    SB_LUT4 i7_4_lut_adj_1685 (.I0(n1846), .I1(n33942), .I2(n1847), .I3(n1848), 
            .O(n18_adj_4994));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam i7_4_lut_adj_1685.LUT_INIT = 16'hfffe;
    SB_LUT4 i5_2_lut (.I0(n1853), .I1(n1852), .I2(GND_net), .I3(GND_net), 
            .O(n16_adj_4995));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam i5_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i9_4_lut_adj_1686 (.I0(n1851), .I1(n18_adj_4994), .I2(n1845), 
            .I3(n1844), .O(n20_adj_4991));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam i9_4_lut_adj_1686.LUT_INIT = 16'hfffe;
    SB_LUT4 i10_4_lut_adj_1687 (.I0(n1849), .I1(n20_adj_4991), .I2(n16_adj_4995), 
            .I3(n1850), .O(n1877));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam i10_4_lut_adj_1687.LUT_INIT = 16'hfffe;
    SB_LUT4 rem_4_mux_3_i18_3_lut (.I0(communication_counter[17]), .I1(n16_adj_4868), 
            .I2(communication_counter[31]), .I3(GND_net), .O(n1858));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_mux_3_i18_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1267_3_lut (.I0(n1858), .I1(n1925), .I2(n1877), .I3(GND_net), 
            .O(n1957));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1267_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1266_3_lut (.I0(n1857), .I1(n1924), .I2(n1877), .I3(GND_net), 
            .O(n1956));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1266_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_3_lut_adj_1688 (.I0(n1956), .I1(n1957), .I2(n1958), .I3(GND_net), 
            .O(n33925));
    defparam i1_3_lut_adj_1688.LUT_INIT = 16'hfefe;
    SB_LUT4 i3_4_lut_adj_1689 (.I0(n1947), .I1(n1954), .I2(n33925), .I3(n1955), 
            .O(n15_adj_4917));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam i3_4_lut_adj_1689.LUT_INIT = 16'heaaa;
    SB_LUT4 i7_4_lut_adj_1690 (.I0(n1944), .I1(n1945), .I2(n1943), .I3(n1946), 
            .O(n19_adj_4915));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam i7_4_lut_adj_1690.LUT_INIT = 16'hfffe;
    SB_LUT4 i6_2_lut (.I0(n1952), .I1(n1953), .I2(GND_net), .I3(GND_net), 
            .O(n18_adj_4916));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam i6_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i10_4_lut_adj_1691 (.I0(n19_adj_4915), .I1(n15_adj_4917), .I2(n1948), 
            .I3(n1950), .O(n22_adj_4914));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam i10_4_lut_adj_1691.LUT_INIT = 16'hfffe;
    SB_LUT4 rem_4_i2204_3_lut (.I0(n3243), .I1(n3310), .I2(n3263), .I3(GND_net), 
            .O(n3342));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i2204_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_1692 (.I0(n3251), .I1(n3345), .I2(n3318), .I3(n3263), 
            .O(n35831));
    defparam i1_4_lut_adj_1692.LUT_INIT = 16'hfcee;
    SB_LUT4 i11_4_lut_adj_1693 (.I0(n1949), .I1(n22_adj_4914), .I2(n18_adj_4916), 
            .I3(n1951), .O(n1976));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam i11_4_lut_adj_1693.LUT_INIT = 16'hfffe;
    SB_LUT4 rem_4_mux_3_i17_3_lut (.I0(communication_counter[16]), .I1(n17_adj_4867), 
            .I2(communication_counter[31]), .I3(GND_net), .O(n1958));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_mux_3_i17_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1335_3_lut (.I0(n1958), .I1(n2025), .I2(n1976), .I3(GND_net), 
            .O(n2057));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1335_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1334_3_lut (.I0(n1957), .I1(n2024), .I2(n1976), .I3(GND_net), 
            .O(n2056));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1334_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_3_lut_adj_1694 (.I0(n2056), .I1(n2057), .I2(n2058), .I3(GND_net), 
            .O(n33970));
    defparam i1_3_lut_adj_1694.LUT_INIT = 16'hfefe;
    SB_LUT4 i3_4_lut_adj_1695 (.I0(n2046), .I1(n2054), .I2(n33970), .I3(n2055), 
            .O(n16_adj_4913));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam i3_4_lut_adj_1695.LUT_INIT = 16'heaaa;
    SB_LUT4 i9_4_lut_adj_1696 (.I0(n2047), .I1(n2052), .I2(n2048), .I3(n2051), 
            .O(n22_adj_4911));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam i9_4_lut_adj_1696.LUT_INIT = 16'hfffe;
    SB_LUT4 i7_3_lut (.I0(n2053), .I1(n2043), .I2(n2042), .I3(GND_net), 
            .O(n20_adj_4912));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam i7_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i11_4_lut_adj_1697 (.I0(n2044), .I1(n22_adj_4911), .I2(n16_adj_4913), 
            .I3(n2045), .O(n24_adj_4910));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam i11_4_lut_adj_1697.LUT_INIT = 16'hfffe;
    SB_LUT4 i12_4_lut_adj_1698 (.I0(n2049), .I1(n24_adj_4910), .I2(n20_adj_4912), 
            .I3(n2050), .O(n2075));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam i12_4_lut_adj_1698.LUT_INIT = 16'hfffe;
    SB_LUT4 rem_4_mux_3_i16_3_lut (.I0(communication_counter[15]), .I1(n18_adj_4866), 
            .I2(communication_counter[31]), .I3(GND_net), .O(n2058));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_mux_3_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1403_3_lut (.I0(n2058), .I1(n2125), .I2(n2075), .I3(GND_net), 
            .O(n2157));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1403_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1402_3_lut (.I0(n2057), .I1(n2124), .I2(n2075), .I3(GND_net), 
            .O(n2156));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1402_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_3_lut_adj_1699 (.I0(n2156), .I1(n2157), .I2(n2158), .I3(GND_net), 
            .O(n33930));
    defparam i1_3_lut_adj_1699.LUT_INIT = 16'hfefe;
    SB_LUT4 i4_4_lut_adj_1700 (.I0(n2154), .I1(n2147), .I2(n33930), .I3(n2155), 
            .O(n18_adj_4804));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam i4_4_lut_adj_1700.LUT_INIT = 16'heccc;
    SB_LUT4 i10_4_lut_adj_1701 (.I0(n2148), .I1(n2152), .I2(n2153), .I3(n2151), 
            .O(n24_adj_4801));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam i10_4_lut_adj_1701.LUT_INIT = 16'hfffe;
    SB_LUT4 i8_4_lut_adj_1702 (.I0(n2142), .I1(n2143), .I2(n2141), .I3(n2144), 
            .O(n22_adj_4802));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam i8_4_lut_adj_1702.LUT_INIT = 16'hfffe;
    SB_LUT4 i12_4_lut_adj_1703 (.I0(n2145), .I1(n24_adj_4801), .I2(n18_adj_4804), 
            .I3(n2146), .O(n26_adj_4800));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam i12_4_lut_adj_1703.LUT_INIT = 16'hfffe;
    SB_LUT4 i13_4_lut_adj_1704 (.I0(n2150), .I1(n26_adj_4800), .I2(n22_adj_4802), 
            .I3(n2149), .O(n2174));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam i13_4_lut_adj_1704.LUT_INIT = 16'hfffe;
    SB_LUT4 rem_4_mux_3_i15_3_lut (.I0(communication_counter[14]), .I1(n19_adj_4865), 
            .I2(communication_counter[31]), .I3(GND_net), .O(n2158));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_mux_3_i15_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_mux_3_i14_3_lut (.I0(communication_counter[13]), .I1(n20_adj_4864), 
            .I2(communication_counter[31]), .I3(GND_net), .O(n2258));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_mux_3_i14_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1471_3_lut (.I0(n2158), .I1(n2225), .I2(n2174), .I3(GND_net), 
            .O(n2257));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1471_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1470_3_lut (.I0(n2157), .I1(n2224), .I2(n2174), .I3(GND_net), 
            .O(n2256));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1470_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_3_lut_adj_1705 (.I0(n2256), .I1(n2257), .I2(n2258), .I3(GND_net), 
            .O(n34002));
    defparam i1_3_lut_adj_1705.LUT_INIT = 16'hfefe;
    SB_LUT4 i11_4_lut_adj_1706 (.I0(n2248), .I1(n2252), .I2(n2250), .I3(n2253), 
            .O(n26_adj_4989));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam i11_4_lut_adj_1706.LUT_INIT = 16'hfffe;
    SB_LUT4 i4_4_lut_adj_1707 (.I0(n2254), .I1(n2246), .I2(n34002), .I3(n2255), 
            .O(n19_adj_4992));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam i4_4_lut_adj_1707.LUT_INIT = 16'heccc;
    SB_LUT4 i1_4_lut_adj_1708 (.I0(n3353), .I1(n3248), .I2(n3315), .I3(n3263), 
            .O(n35837));
    defparam i1_4_lut_adj_1708.LUT_INIT = 16'hfaee;
    SB_LUT4 rem_4_i2205_3_lut (.I0(n3244), .I1(n3311), .I2(n3263), .I3(GND_net), 
            .O(n3343));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i2205_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_adj_1709 (.I0(n2241), .I1(n2240), .I2(GND_net), .I3(GND_net), 
            .O(n16_adj_4993));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam i1_2_lut_adj_1709.LUT_INIT = 16'heeee;
    SB_LUT4 i9_4_lut_adj_1710 (.I0(n2242), .I1(n2244), .I2(n2243), .I3(n2245), 
            .O(n24_adj_4990));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam i9_4_lut_adj_1710.LUT_INIT = 16'hfffe;
    SB_LUT4 i13_4_lut_adj_1711 (.I0(n19_adj_4992), .I1(n26_adj_4989), .I2(n2247), 
            .I3(n2251), .O(n28_adj_4988));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam i13_4_lut_adj_1711.LUT_INIT = 16'hfffe;
    SB_LUT4 rem_4_i2210_3_lut (.I0(n3249), .I1(n3316), .I2(n3263), .I3(GND_net), 
            .O(n3348));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i2210_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_1712 (.I0(n3253), .I1(n3348), .I2(n3320), .I3(n3263), 
            .O(n35835));
    defparam i1_4_lut_adj_1712.LUT_INIT = 16'hfcee;
    SB_LUT4 rem_4_i2206_3_lut (.I0(n3245), .I1(n3312), .I2(n3263), .I3(GND_net), 
            .O(n3344));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i2206_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_1713 (.I0(n3250), .I1(n3346), .I2(n3317), .I3(n3263), 
            .O(n35833));
    defparam i1_4_lut_adj_1713.LUT_INIT = 16'hfcee;
    SB_LUT4 i1_4_lut_adj_1714 (.I0(n3252), .I1(n3344), .I2(n3319), .I3(n3263), 
            .O(n35829));
    defparam i1_4_lut_adj_1714.LUT_INIT = 16'hfcee;
    SB_LUT4 i1_4_lut_adj_1715 (.I0(n3343), .I1(n35837), .I2(n35831), .I3(n3342), 
            .O(n35845));
    defparam i1_4_lut_adj_1715.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1716 (.I0(n3242), .I1(n35835), .I2(n3309), .I3(n3263), 
            .O(n35843));
    defparam i1_4_lut_adj_1716.LUT_INIT = 16'hfcee;
    SB_LUT4 rem_4_add_2189_24_lut (.I0(GND_net), .I1(n3237), .I2(VCC_net), 
            .I3(n28700), .O(n3304)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2189_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i13422_3_lut (.I0(encoder1_position[18]), .I1(n3164), .I2(count_enable_adj_4807), 
            .I3(GND_net), .O(n18251));   // quad.v(35[10] 41[6])
    defparam i13422_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY rem_4_add_2189_24 (.CI(n28700), .I0(n3237), .I1(VCC_net), 
            .CO(n28701));
    SB_LUT4 rem_4_add_2189_23_lut (.I0(GND_net), .I1(n3238), .I2(VCC_net), 
            .I3(n28699), .O(n3305)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2189_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_2189_23 (.CI(n28699), .I0(n3238), .I1(VCC_net), 
            .CO(n28700));
    SB_LUT4 rem_4_add_2189_22_lut (.I0(GND_net), .I1(n3239), .I2(VCC_net), 
            .I3(n28698), .O(n3306)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2189_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_2189_22 (.CI(n28698), .I0(n3239), .I1(VCC_net), 
            .CO(n28699));
    SB_CARRY rem_4_add_1452_16 (.CI(n28228), .I0(n2144), .I1(VCC_net), 
            .CO(n28229));
    SB_LUT4 i13421_3_lut (.I0(encoder1_position[17]), .I1(n3165), .I2(count_enable_adj_4807), 
            .I3(GND_net), .O(n18250));   // quad.v(35[10] 41[6])
    defparam i13421_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_add_2189_21_lut (.I0(GND_net), .I1(n3240), .I2(VCC_net), 
            .I3(n28697), .O(n3307)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2189_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_2189_21 (.CI(n28697), .I0(n3240), .I1(VCC_net), 
            .CO(n28698));
    SB_LUT4 rem_4_add_2189_20_lut (.I0(GND_net), .I1(n3241), .I2(VCC_net), 
            .I3(n28696), .O(n3308)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2189_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_2189_20 (.CI(n28696), .I0(n3241), .I1(VCC_net), 
            .CO(n28697));
    SB_LUT4 rem_4_add_2189_19_lut (.I0(GND_net), .I1(n3242), .I2(VCC_net), 
            .I3(n28695), .O(n3309)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2189_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_2189_19 (.CI(n28695), .I0(n3242), .I1(VCC_net), 
            .CO(n28696));
    SB_LUT4 rem_4_add_2189_18_lut (.I0(GND_net), .I1(n3243), .I2(VCC_net), 
            .I3(n28694), .O(n3310)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2189_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_2189_18 (.CI(n28694), .I0(n3243), .I1(VCC_net), 
            .CO(n28695));
    SB_LUT4 rem_4_add_2189_17_lut (.I0(GND_net), .I1(n3244), .I2(VCC_net), 
            .I3(n28693), .O(n3311)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2189_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_2189_17 (.CI(n28693), .I0(n3244), .I1(VCC_net), 
            .CO(n28694));
    SB_LUT4 rem_4_add_2189_16_lut (.I0(GND_net), .I1(n3245), .I2(VCC_net), 
            .I3(n28692), .O(n3312)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2189_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_2189_16 (.CI(n28692), .I0(n3245), .I1(VCC_net), 
            .CO(n28693));
    SB_LUT4 rem_4_add_2189_15_lut (.I0(GND_net), .I1(n3246), .I2(VCC_net), 
            .I3(n28691), .O(n3313)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2189_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_2189_15 (.CI(n28691), .I0(n3246), .I1(VCC_net), 
            .CO(n28692));
    SB_LUT4 rem_4_add_2189_14_lut (.I0(GND_net), .I1(n3247), .I2(VCC_net), 
            .I3(n28690), .O(n3314)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2189_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_2189_14 (.CI(n28690), .I0(n3247), .I1(VCC_net), 
            .CO(n28691));
    SB_LUT4 rem_4_add_2189_13_lut (.I0(GND_net), .I1(n3248), .I2(VCC_net), 
            .I3(n28689), .O(n3315)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2189_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_2189_13 (.CI(n28689), .I0(n3248), .I1(VCC_net), 
            .CO(n28690));
    SB_LUT4 rem_4_add_2189_12_lut (.I0(GND_net), .I1(n3249), .I2(VCC_net), 
            .I3(n28688), .O(n3316)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2189_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_2189_12 (.CI(n28688), .I0(n3249), .I1(VCC_net), 
            .CO(n28689));
    SB_LUT4 rem_4_add_2189_11_lut (.I0(GND_net), .I1(n3250), .I2(VCC_net), 
            .I3(n28687), .O(n3317)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2189_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_2189_11 (.CI(n28687), .I0(n3250), .I1(VCC_net), 
            .CO(n28688));
    SB_LUT4 rem_4_add_2189_10_lut (.I0(GND_net), .I1(n3251), .I2(VCC_net), 
            .I3(n28686), .O(n3318)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2189_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_2189_10 (.CI(n28686), .I0(n3251), .I1(VCC_net), 
            .CO(n28687));
    SB_LUT4 rem_4_add_2189_9_lut (.I0(GND_net), .I1(n3252), .I2(VCC_net), 
            .I3(n28685), .O(n3319)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2189_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_2189_9 (.CI(n28685), .I0(n3252), .I1(VCC_net), 
            .CO(n28686));
    SB_LUT4 rem_4_add_2189_8_lut (.I0(GND_net), .I1(n3253), .I2(VCC_net), 
            .I3(n28684), .O(n3320)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2189_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_2189_8 (.CI(n28684), .I0(n3253), .I1(VCC_net), 
            .CO(n28685));
    SB_LUT4 rem_4_add_2189_7_lut (.I0(GND_net), .I1(n3254), .I2(GND_net), 
            .I3(n28683), .O(n3321)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2189_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_2189_7 (.CI(n28683), .I0(n3254), .I1(GND_net), 
            .CO(n28684));
    SB_LUT4 rem_4_add_2189_6_lut (.I0(GND_net), .I1(n3255), .I2(GND_net), 
            .I3(n28682), .O(n3322)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2189_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_2189_6 (.CI(n28682), .I0(n3255), .I1(GND_net), 
            .CO(n28683));
    SB_LUT4 rem_4_add_2189_5_lut (.I0(GND_net), .I1(n3256), .I2(VCC_net), 
            .I3(n28681), .O(n3323)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2189_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_2189_5 (.CI(n28681), .I0(n3256), .I1(VCC_net), 
            .CO(n28682));
    SB_LUT4 rem_4_add_2189_4_lut (.I0(GND_net), .I1(n3257), .I2(VCC_net), 
            .I3(n28680), .O(n3324)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2189_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i13424_3_lut (.I0(encoder1_position[20]), .I1(n3162), .I2(count_enable_adj_4807), 
            .I3(GND_net), .O(n18253));   // quad.v(35[10] 41[6])
    defparam i13424_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_add_1452_15_lut (.I0(GND_net), .I1(n2145), .I2(VCC_net), 
            .I3(n28227), .O(n2212)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1452_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i13423_3_lut (.I0(encoder1_position[19]), .I1(n3163), .I2(count_enable_adj_4807), 
            .I3(GND_net), .O(n18252));   // quad.v(35[10] 41[6])
    defparam i13423_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13370_3_lut (.I0(PWMLimit[14]), .I1(\data_in_frame[9] [6]), 
            .I2(n5439), .I3(GND_net), .O(n18199));   // verilog/coms.v(126[12] 293[6])
    defparam i13370_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i586_3_lut_4_lut (.I0(n36410), .I1(n746), .I2(n855), 
            .I3(n749), .O(n956));
    defparam rem_4_i586_3_lut_4_lut.LUT_INIT = 16'hf708;
    SB_LUT4 i13373_3_lut (.I0(PWMLimit[17]), .I1(\data_in_frame[8] [1]), 
            .I2(n5439), .I3(GND_net), .O(n18202));   // verilog/coms.v(126[12] 293[6])
    defparam i13373_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13369_3_lut (.I0(PWMLimit[13]), .I1(\data_in_frame[9] [5]), 
            .I2(n5439), .I3(GND_net), .O(n18198));   // verilog/coms.v(126[12] 293[6])
    defparam i13369_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_1717 (.I0(n35843), .I1(n35845), .I2(n35829), 
            .I3(n35833), .O(n35849));
    defparam i1_4_lut_adj_1717.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_3_lut_adj_1718 (.I0(n3356), .I1(n3357), .I2(n3358), .I3(GND_net), 
            .O(n33989));
    defparam i1_3_lut_adj_1718.LUT_INIT = 16'hfefe;
    SB_LUT4 i1_4_lut_adj_1719 (.I0(n3241), .I1(n35849), .I2(n3308), .I3(n3263), 
            .O(n35851));
    defparam i1_4_lut_adj_1719.LUT_INIT = 16'hfcee;
    SB_LUT4 i1_4_lut_adj_1720 (.I0(n3354), .I1(n35851), .I2(n33989), .I3(n3355), 
            .O(n35853));
    defparam i1_4_lut_adj_1720.LUT_INIT = 16'heccc;
    SB_LUT4 rem_4_unary_minus_2_inv_0_i30_1_lut (.I0(communication_counter[29]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n4_adj_4953));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_unary_minus_2_inv_0_i30_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i13368_3_lut (.I0(PWMLimit[12]), .I1(\data_in_frame[9] [4]), 
            .I2(n5439), .I3(GND_net), .O(n18197));   // verilog/coms.v(126[12] 293[6])
    defparam i13368_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i23020_2_lut_3_lut (.I0(n36410), .I1(n746), .I2(n855), .I3(GND_net), 
            .O(n957));
    defparam i23020_2_lut_3_lut.LUT_INIT = 16'h7878;
    SB_LUT4 rem_4_i585_3_lut_4_lut (.I0(n36410), .I1(n746), .I2(n4_adj_4781), 
            .I3(n748), .O(n955));
    defparam rem_4_i585_3_lut_4_lut.LUT_INIT = 16'hf708;
    SB_LUT4 rem_4_i584_3_lut_4_lut (.I0(n36410), .I1(n746), .I2(n6_adj_5000), 
            .I3(n852), .O(n954));
    defparam rem_4_i584_3_lut_4_lut.LUT_INIT = 16'h7f08;
    SB_CARRY rem_4_add_2189_4 (.CI(n28680), .I0(n3257), .I1(VCC_net), 
            .CO(n28681));
    SB_LUT4 rem_4_add_2189_3_lut (.I0(GND_net), .I1(n3258), .I2(GND_net), 
            .I3(n28679), .O(n3325)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2189_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_4_lut_adj_1721 (.I0(n3240), .I1(n35853), .I2(n3307), .I3(n3263), 
            .O(n35855));
    defparam i1_4_lut_adj_1721.LUT_INIT = 16'hfcee;
    SB_LUT4 i1_4_lut_adj_1722 (.I0(n3239), .I1(n35855), .I2(n3306), .I3(n3263), 
            .O(n35857));
    defparam i1_4_lut_adj_1722.LUT_INIT = 16'hfcee;
    SB_LUT4 rem_4_unary_minus_2_inv_0_i31_1_lut (.I0(communication_counter[30]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n3_adj_4952));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_unary_minus_2_inv_0_i31_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY rem_4_add_1452_15 (.CI(n28227), .I0(n2145), .I1(VCC_net), 
            .CO(n28228));
    SB_LUT4 rem_4_add_1452_14_lut (.I0(GND_net), .I1(n2146), .I2(VCC_net), 
            .I3(n28226), .O(n2213)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1452_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_2189_3 (.CI(n28679), .I0(n3258), .I1(GND_net), 
            .CO(n28680));
    SB_CARRY rem_4_add_1452_14 (.CI(n28226), .I0(n2146), .I1(VCC_net), 
            .CO(n28227));
    SB_LUT4 rem_4_add_1452_13_lut (.I0(GND_net), .I1(n2147), .I2(VCC_net), 
            .I3(n28225), .O(n2214)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1452_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1452_13 (.CI(n28225), .I0(n2147), .I1(VCC_net), 
            .CO(n28226));
    SB_CARRY rem_4_add_2189_2 (.CI(VCC_net), .I0(n3358), .I1(VCC_net), 
            .CO(n28679));
    SB_LUT4 rem_4_add_2122_30_lut (.I0(n3164_adj_4884), .I1(n3131), .I2(VCC_net), 
            .I3(n28678), .O(n3230_adj_4902)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2122_30_lut.LUT_INIT = 16'h8228;
    SB_LUT4 rem_4_add_1452_12_lut (.I0(GND_net), .I1(n2148), .I2(VCC_net), 
            .I3(n28224), .O(n2215)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1452_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_2122_29_lut (.I0(GND_net), .I1(n3132), .I2(VCC_net), 
            .I3(n28677), .O(n3199)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2122_29_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_4_lut_adj_1723 (.I0(n3238), .I1(n35857), .I2(n3305), .I3(n3263), 
            .O(n35859));
    defparam i1_4_lut_adj_1723.LUT_INIT = 16'hfcee;
    SB_CARRY rem_4_add_2122_29 (.CI(n28677), .I0(n3132), .I1(VCC_net), 
            .CO(n28678));
    SB_CARRY rem_4_add_1452_12 (.CI(n28224), .I0(n2148), .I1(VCC_net), 
            .CO(n28225));
    SB_LUT4 rem_4_add_2122_28_lut (.I0(GND_net), .I1(n3133), .I2(VCC_net), 
            .I3(n28676), .O(n3200)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2122_28_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_2122_28 (.CI(n28676), .I0(n3133), .I1(VCC_net), 
            .CO(n28677));
    SB_LUT4 rem_4_add_2122_27_lut (.I0(GND_net), .I1(n3134), .I2(VCC_net), 
            .I3(n28675), .O(n3201)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2122_27_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1452_11_lut (.I0(GND_net), .I1(n2149), .I2(VCC_net), 
            .I3(n28223), .O(n2216)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1452_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_2122_27 (.CI(n28675), .I0(n3134), .I1(VCC_net), 
            .CO(n28676));
    SB_LUT4 rem_4_add_2122_26_lut (.I0(GND_net), .I1(n3135), .I2(VCC_net), 
            .I3(n28674), .O(n3202)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2122_26_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i13367_3_lut (.I0(PWMLimit[11]), .I1(\data_in_frame[9] [3]), 
            .I2(n5439), .I3(GND_net), .O(n18196));   // verilog/coms.v(126[12] 293[6])
    defparam i13367_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13366_3_lut (.I0(PWMLimit[10]), .I1(\data_in_frame[9] [2]), 
            .I2(n5439), .I3(GND_net), .O(n18195));   // verilog/coms.v(126[12] 293[6])
    defparam i13366_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_1724 (.I0(n3237), .I1(n35859), .I2(n3304), .I3(n3263), 
            .O(n35861));
    defparam i1_4_lut_adj_1724.LUT_INIT = 16'hfcee;
    SB_LUT4 i13365_3_lut (.I0(PWMLimit[9]), .I1(\data_in_frame[9] [1]), 
            .I2(n5439), .I3(GND_net), .O(n18194));   // verilog/coms.v(126[12] 293[6])
    defparam i13365_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_unary_minus_2_inv_0_i32_1_lut (.I0(communication_counter[31]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n2_adj_4951));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_unary_minus_2_inv_0_i32_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i13379_3_lut (.I0(PWMLimit[23]), .I1(\data_in_frame[8] [7]), 
            .I2(n5439), .I3(GND_net), .O(n18208));   // verilog/coms.v(126[12] 293[6])
    defparam i13379_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13378_3_lut (.I0(PWMLimit[22]), .I1(\data_in_frame[8] [6]), 
            .I2(n5439), .I3(GND_net), .O(n18207));   // verilog/coms.v(126[12] 293[6])
    defparam i13378_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13377_3_lut (.I0(PWMLimit[21]), .I1(\data_in_frame[8] [5]), 
            .I2(n5439), .I3(GND_net), .O(n18206));   // verilog/coms.v(126[12] 293[6])
    defparam i13377_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13376_3_lut (.I0(PWMLimit[20]), .I1(\data_in_frame[8] [4]), 
            .I2(n5439), .I3(GND_net), .O(n18205));   // verilog/coms.v(126[12] 293[6])
    defparam i13376_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12730_4_lut (.I0(n5478), .I1(r_Clock_Count_adj_5048[3]), .I2(n318), 
            .I3(r_SM_Main_adj_5047[2]), .O(n17559));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i12730_4_lut.LUT_INIT = 16'h4450;
    SB_LUT4 i13375_3_lut (.I0(PWMLimit[19]), .I1(\data_in_frame[8] [3]), 
            .I2(n5439), .I3(GND_net), .O(n18204));   // verilog/coms.v(126[12] 293[6])
    defparam i13375_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13374_3_lut (.I0(PWMLimit[18]), .I1(\data_in_frame[8] [2]), 
            .I2(n5439), .I3(GND_net), .O(n18203));   // verilog/coms.v(126[12] 293[6])
    defparam i13374_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_1725 (.I0(n3236), .I1(n35861), .I2(n3303), .I3(n3263), 
            .O(n35863));
    defparam i1_4_lut_adj_1725.LUT_INIT = 16'hfcee;
    SB_LUT4 i1_4_lut_adj_1726 (.I0(n3235), .I1(n35863), .I2(n3302), .I3(n3263), 
            .O(n35865));
    defparam i1_4_lut_adj_1726.LUT_INIT = 16'hfcee;
    SB_LUT4 unary_minus_28_inv_0_i17_1_lut (.I0(duty[16]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n9));   // verilog/TinyFPGA_B.v(149[23:28])
    defparam unary_minus_28_inv_0_i17_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i12908_3_lut (.I0(\neo_pixel_transmitter.t0 [1]), .I1(timer[1]), 
            .I2(n20), .I3(GND_net), .O(n17737));   // verilog/neopixel.v(35[12] 117[6])
    defparam i12908_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_1727 (.I0(n3234), .I1(n35865), .I2(n3301), .I3(n3263), 
            .O(n35867));
    defparam i1_4_lut_adj_1727.LUT_INIT = 16'hfcee;
    SB_LUT4 i1_4_lut_adj_1728 (.I0(n3233), .I1(n35867), .I2(n3300), .I3(n3263), 
            .O(n35869));
    defparam i1_4_lut_adj_1728.LUT_INIT = 16'hfcee;
    SB_LUT4 i12909_3_lut (.I0(\neo_pixel_transmitter.t0 [2]), .I1(timer[2]), 
            .I2(n20), .I3(GND_net), .O(n17738));   // verilog/neopixel.v(35[12] 117[6])
    defparam i12909_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 unary_minus_28_inv_0_i18_1_lut (.I0(duty[17]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n8));   // verilog/TinyFPGA_B.v(149[23:28])
    defparam unary_minus_28_inv_0_i18_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_28_inv_0_i19_1_lut (.I0(duty[18]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n7));   // verilog/TinyFPGA_B.v(149[23:28])
    defparam unary_minus_28_inv_0_i19_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i12910_3_lut (.I0(\neo_pixel_transmitter.t0 [3]), .I1(timer[3]), 
            .I2(n20), .I3(GND_net), .O(n17739));   // verilog/neopixel.v(35[12] 117[6])
    defparam i12910_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 rem_4_i2193_3_lut (.I0(n3232_adj_4904), .I1(n3299), .I2(n3263), 
            .I3(GND_net), .O(n3331));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i2193_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i2192_3_lut (.I0(n3231_adj_4903), .I1(n3298), .I2(n3263), 
            .I3(GND_net), .O(n3330));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i2192_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i31552_1_lut (.I0(n2669), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n38232));
    defparam i31552_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i12911_3_lut (.I0(\neo_pixel_transmitter.t0 [4]), .I1(timer[4]), 
            .I2(n20), .I3(GND_net), .O(n17740));   // verilog/neopixel.v(35[12] 117[6])
    defparam i12911_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY rem_4_add_1452_11 (.CI(n28223), .I0(n2149), .I1(VCC_net), 
            .CO(n28224));
    SB_LUT4 unary_minus_28_inv_0_i20_1_lut (.I0(duty[19]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n6));   // verilog/TinyFPGA_B.v(149[23:28])
    defparam unary_minus_28_inv_0_i20_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1_4_lut_adj_1729 (.I0(n3330), .I1(n36391), .I2(n3331), .I3(n35869), 
            .O(n3362));
    defparam i1_4_lut_adj_1729.LUT_INIT = 16'hfffe;
    SB_LUT4 i12912_3_lut (.I0(\neo_pixel_transmitter.t0 [5]), .I1(timer[5]), 
            .I2(n20), .I3(GND_net), .O(n17741));   // verilog/neopixel.v(35[12] 117[6])
    defparam i12912_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12913_3_lut (.I0(\neo_pixel_transmitter.t0 [6]), .I1(timer[6]), 
            .I2(n20), .I3(GND_net), .O(n17742));   // verilog/neopixel.v(35[12] 117[6])
    defparam i12913_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12914_3_lut (.I0(\neo_pixel_transmitter.t0 [7]), .I1(timer[7]), 
            .I2(n20), .I3(GND_net), .O(n17743));   // verilog/neopixel.v(35[12] 117[6])
    defparam i12914_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 rem_4_i2282_3_lut (.I0(n3353), .I1(n10390), .I2(n3362), .I3(GND_net), 
            .O(n3452));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i2282_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 i13427_3_lut (.I0(encoder1_position[23]), .I1(n3159), .I2(count_enable_adj_4807), 
            .I3(GND_net), .O(n18256));   // quad.v(35[10] 41[6])
    defparam i13427_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12915_3_lut (.I0(\neo_pixel_transmitter.t0 [8]), .I1(timer[8]), 
            .I2(n20), .I3(GND_net), .O(n17744));   // verilog/neopixel.v(35[12] 117[6])
    defparam i12915_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12916_3_lut (.I0(\neo_pixel_transmitter.t0 [9]), .I1(timer[9]), 
            .I2(n20), .I3(GND_net), .O(n17745));   // verilog/neopixel.v(35[12] 117[6])
    defparam i12916_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12917_3_lut (.I0(\neo_pixel_transmitter.t0 [10]), .I1(timer[10]), 
            .I2(n20), .I3(GND_net), .O(n17746));   // verilog/neopixel.v(35[12] 117[6])
    defparam i12917_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13189_3_lut (.I0(\data_in_frame[1] [0]), .I1(rx_data[0]), .I2(n32962), 
            .I3(GND_net), .O(n18018));   // verilog/coms.v(126[12] 293[6])
    defparam i13189_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12918_3_lut (.I0(\neo_pixel_transmitter.t0 [11]), .I1(timer[11]), 
            .I2(n20), .I3(GND_net), .O(n17747));   // verilog/neopixel.v(35[12] 117[6])
    defparam i12918_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 unary_minus_28_inv_0_i21_1_lut (.I0(duty[20]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n5));   // verilog/TinyFPGA_B.v(149[23:28])
    defparam unary_minus_28_inv_0_i21_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 rem_4_i2129_3_lut (.I0(n3136), .I1(n3203), .I2(n3164_adj_4884), 
            .I3(GND_net), .O(n3235));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i2129_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12919_3_lut (.I0(\neo_pixel_transmitter.t0 [12]), .I1(timer[12]), 
            .I2(n20), .I3(GND_net), .O(n17748));   // verilog/neopixel.v(35[12] 117[6])
    defparam i12919_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12920_3_lut (.I0(\neo_pixel_transmitter.t0 [13]), .I1(timer[13]), 
            .I2(n20), .I3(GND_net), .O(n17749));   // verilog/neopixel.v(35[12] 117[6])
    defparam i12920_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 rem_4_i2127_3_lut (.I0(n3134), .I1(n3201), .I2(n3164_adj_4884), 
            .I3(GND_net), .O(n3233));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i2127_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY rem_4_add_2122_26 (.CI(n28674), .I0(n3135), .I1(VCC_net), 
            .CO(n28675));
    SB_LUT4 rem_4_add_2122_25_lut (.I0(GND_net), .I1(n3136), .I2(VCC_net), 
            .I3(n28673), .O(n3203)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2122_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i12921_3_lut (.I0(\neo_pixel_transmitter.t0 [14]), .I1(timer[14]), 
            .I2(n20), .I3(GND_net), .O(n17750));   // verilog/neopixel.v(35[12] 117[6])
    defparam i12921_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 rem_4_add_1452_10_lut (.I0(GND_net), .I1(n2150), .I2(VCC_net), 
            .I3(n28222), .O(n2217)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1452_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1452_10 (.CI(n28222), .I0(n2150), .I1(VCC_net), 
            .CO(n28223));
    SB_CARRY rem_4_add_2122_25 (.CI(n28673), .I0(n3136), .I1(VCC_net), 
            .CO(n28674));
    SB_LUT4 rem_4_add_1452_9_lut (.I0(GND_net), .I1(n2151), .I2(VCC_net), 
            .I3(n28221), .O(n2218)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1452_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i12922_3_lut (.I0(\neo_pixel_transmitter.t0 [15]), .I1(timer[15]), 
            .I2(n20), .I3(GND_net), .O(n17751));   // verilog/neopixel.v(35[12] 117[6])
    defparam i12922_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 rem_4_i2128_3_lut (.I0(n3135), .I1(n3202), .I2(n3164_adj_4884), 
            .I3(GND_net), .O(n3234));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i2128_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12923_3_lut (.I0(\neo_pixel_transmitter.t0 [16]), .I1(timer[16]), 
            .I2(n20), .I3(GND_net), .O(n17752));   // verilog/neopixel.v(35[12] 117[6])
    defparam i12923_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 rem_4_i2126_3_lut (.I0(n3133), .I1(n3200), .I2(n3164_adj_4884), 
            .I3(GND_net), .O(n3232_adj_4904));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i2126_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12924_3_lut (.I0(\neo_pixel_transmitter.t0 [17]), .I1(timer[17]), 
            .I2(n20), .I3(GND_net), .O(n17753));   // verilog/neopixel.v(35[12] 117[6])
    defparam i12924_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12925_3_lut (.I0(\neo_pixel_transmitter.t0 [18]), .I1(timer[18]), 
            .I2(n20), .I3(GND_net), .O(n17754));   // verilog/neopixel.v(35[12] 117[6])
    defparam i12925_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12926_3_lut (.I0(\neo_pixel_transmitter.t0 [19]), .I1(timer[19]), 
            .I2(n20), .I3(GND_net), .O(n17755));   // verilog/neopixel.v(35[12] 117[6])
    defparam i12926_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 rem_4_i2135_3_lut (.I0(n3142), .I1(n3209_adj_4885), .I2(n3164_adj_4884), 
            .I3(GND_net), .O(n3241));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i2135_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12927_3_lut (.I0(\neo_pixel_transmitter.t0 [20]), .I1(timer[20]), 
            .I2(n20), .I3(GND_net), .O(n17756));   // verilog/neopixel.v(35[12] 117[6])
    defparam i12927_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12928_3_lut (.I0(\neo_pixel_transmitter.t0 [21]), .I1(timer[21]), 
            .I2(n20), .I3(GND_net), .O(n17757));   // verilog/neopixel.v(35[12] 117[6])
    defparam i12928_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12929_3_lut (.I0(\neo_pixel_transmitter.t0 [22]), .I1(timer[22]), 
            .I2(n20), .I3(GND_net), .O(n17758));   // verilog/neopixel.v(35[12] 117[6])
    defparam i12929_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12930_3_lut (.I0(\neo_pixel_transmitter.t0 [23]), .I1(timer[23]), 
            .I2(n20), .I3(GND_net), .O(n17759));   // verilog/neopixel.v(35[12] 117[6])
    defparam i12930_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12931_3_lut (.I0(\neo_pixel_transmitter.t0 [24]), .I1(timer[24]), 
            .I2(n20), .I3(GND_net), .O(n17760));   // verilog/neopixel.v(35[12] 117[6])
    defparam i12931_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 rem_4_i2134_3_lut (.I0(n3141), .I1(n3208), .I2(n3164_adj_4884), 
            .I3(GND_net), .O(n3240));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i2134_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i2145_3_lut (.I0(n3152), .I1(n3219_adj_4895), .I2(n3164_adj_4884), 
            .I3(GND_net), .O(n3251));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i2145_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i2141_3_lut (.I0(n3148), .I1(n3215_adj_4891), .I2(n3164_adj_4884), 
            .I3(GND_net), .O(n3247));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i2141_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i2133_3_lut (.I0(n3140), .I1(n3207), .I2(n3164_adj_4884), 
            .I3(GND_net), .O(n3239));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i2133_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12932_3_lut (.I0(\neo_pixel_transmitter.t0 [25]), .I1(timer[25]), 
            .I2(n20), .I3(GND_net), .O(n17761));   // verilog/neopixel.v(35[12] 117[6])
    defparam i12932_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12933_3_lut (.I0(\neo_pixel_transmitter.t0 [26]), .I1(timer[26]), 
            .I2(n20), .I3(GND_net), .O(n17762));   // verilog/neopixel.v(35[12] 117[6])
    defparam i12933_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12934_3_lut (.I0(\neo_pixel_transmitter.t0 [27]), .I1(timer[27]), 
            .I2(n20), .I3(GND_net), .O(n17763));   // verilog/neopixel.v(35[12] 117[6])
    defparam i12934_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 rem_4_i2131_3_lut (.I0(n3138), .I1(n3205), .I2(n3164_adj_4884), 
            .I3(GND_net), .O(n3237));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i2131_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i2132_3_lut (.I0(n3139), .I1(n3206), .I2(n3164_adj_4884), 
            .I3(GND_net), .O(n3238));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i2132_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12935_3_lut (.I0(\neo_pixel_transmitter.t0 [28]), .I1(timer[28]), 
            .I2(n20), .I3(GND_net), .O(n17764));   // verilog/neopixel.v(35[12] 117[6])
    defparam i12935_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12936_3_lut (.I0(\neo_pixel_transmitter.t0 [29]), .I1(timer[29]), 
            .I2(n20), .I3(GND_net), .O(n17765));   // verilog/neopixel.v(35[12] 117[6])
    defparam i12936_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 rem_4_i2130_3_lut (.I0(n3137), .I1(n3204), .I2(n3164_adj_4884), 
            .I3(GND_net), .O(n3236));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i2130_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_add_2122_24_lut (.I0(GND_net), .I1(n3137), .I2(VCC_net), 
            .I3(n28672), .O(n3204)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2122_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i12937_3_lut (.I0(\neo_pixel_transmitter.t0 [30]), .I1(timer[30]), 
            .I2(n20), .I3(GND_net), .O(n17766));   // verilog/neopixel.v(35[12] 117[6])
    defparam i12937_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12938_3_lut (.I0(\neo_pixel_transmitter.t0 [31]), .I1(timer[31]), 
            .I2(n20), .I3(GND_net), .O(n17767));   // verilog/neopixel.v(35[12] 117[6])
    defparam i12938_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY rem_4_add_2122_24 (.CI(n28672), .I0(n3137), .I1(VCC_net), 
            .CO(n28673));
    SB_LUT4 rem_4_add_2122_23_lut (.I0(GND_net), .I1(n3138), .I2(VCC_net), 
            .I3(n28671), .O(n3205)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2122_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i12939_3_lut (.I0(IntegralLimit[1]), .I1(\data_in_frame[13] [1]), 
            .I2(n5439), .I3(GND_net), .O(n17768));   // verilog/coms.v(126[12] 293[6])
    defparam i12939_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12940_3_lut (.I0(IntegralLimit[2]), .I1(\data_in_frame[13] [2]), 
            .I2(n5439), .I3(GND_net), .O(n17769));   // verilog/coms.v(126[12] 293[6])
    defparam i12940_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12941_3_lut (.I0(IntegralLimit[3]), .I1(\data_in_frame[13] [3]), 
            .I2(n5439), .I3(GND_net), .O(n17770));   // verilog/coms.v(126[12] 293[6])
    defparam i12941_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12942_3_lut (.I0(IntegralLimit[4]), .I1(\data_in_frame[13] [4]), 
            .I2(n5439), .I3(GND_net), .O(n17771));   // verilog/coms.v(126[12] 293[6])
    defparam i12942_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12943_3_lut (.I0(IntegralLimit[5]), .I1(\data_in_frame[13] [5]), 
            .I2(n5439), .I3(GND_net), .O(n17772));   // verilog/coms.v(126[12] 293[6])
    defparam i12943_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12944_3_lut (.I0(IntegralLimit[6]), .I1(\data_in_frame[13] [6]), 
            .I2(n5439), .I3(GND_net), .O(n17773));   // verilog/coms.v(126[12] 293[6])
    defparam i12944_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY rem_4_add_2122_23 (.CI(n28671), .I0(n3138), .I1(VCC_net), 
            .CO(n28672));
    SB_LUT4 rem_4_add_2122_22_lut (.I0(GND_net), .I1(n3139), .I2(VCC_net), 
            .I3(n28670), .O(n3206)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2122_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1452_9 (.CI(n28221), .I0(n2151), .I1(VCC_net), 
            .CO(n28222));
    SB_LUT4 rem_4_add_1452_8_lut (.I0(GND_net), .I1(n2152), .I2(VCC_net), 
            .I3(n28220), .O(n2219)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1452_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1452_8 (.CI(n28220), .I0(n2152), .I1(VCC_net), 
            .CO(n28221));
    SB_CARRY rem_4_add_2122_22 (.CI(n28670), .I0(n3139), .I1(VCC_net), 
            .CO(n28671));
    SB_LUT4 rem_4_add_2122_21_lut (.I0(GND_net), .I1(n3140), .I2(VCC_net), 
            .I3(n28669), .O(n3207)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2122_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i12717_3_lut (.I0(\neo_pixel_transmitter.t0 [0]), .I1(timer[0]), 
            .I2(n20), .I3(GND_net), .O(n17546));   // verilog/neopixel.v(35[12] 117[6])
    defparam i12717_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12721_3_lut (.I0(IntegralLimit[0]), .I1(\data_in_frame[13] [0]), 
            .I2(n5439), .I3(GND_net), .O(n17550));   // verilog/coms.v(126[12] 293[6])
    defparam i12721_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY rem_4_add_2122_21 (.CI(n28669), .I0(n3140), .I1(VCC_net), 
            .CO(n28670));
    SB_LUT4 i13318_3_lut (.I0(\data_in_frame[17] [1]), .I1(rx_data[1]), 
            .I2(n32957), .I3(GND_net), .O(n18147));   // verilog/coms.v(126[12] 293[6])
    defparam i13318_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13319_3_lut (.I0(\data_in_frame[17] [2]), .I1(rx_data[2]), 
            .I2(n32957), .I3(GND_net), .O(n18148));   // verilog/coms.v(126[12] 293[6])
    defparam i13319_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 rem_4_i924_3_lut (.I0(n1355), .I1(n1422), .I2(n1382), .I3(GND_net), 
            .O(n1454));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i924_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i923_3_lut (.I0(n1354), .I1(n1421), .I2(n1382), .I3(GND_net), 
            .O(n1453));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i923_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 unary_minus_28_inv_0_i7_1_lut (.I0(duty[6]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n19));   // verilog/TinyFPGA_B.v(149[23:28])
    defparam unary_minus_28_inv_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i13253_3_lut (.I0(\data_in_frame[9] [0]), .I1(rx_data[0]), .I2(n32941), 
            .I3(GND_net), .O(n18082));   // verilog/coms.v(126[12] 293[6])
    defparam i13253_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 rem_4_i2138_3_lut (.I0(n3145), .I1(n3212_adj_4888), .I2(n3164_adj_4884), 
            .I3(GND_net), .O(n3244));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i2138_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13254_3_lut (.I0(\data_in_frame[9] [1]), .I1(rx_data[1]), .I2(n32941), 
            .I3(GND_net), .O(n18083));   // verilog/coms.v(126[12] 293[6])
    defparam i13254_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13255_3_lut (.I0(\data_in_frame[9] [2]), .I1(rx_data[2]), .I2(n32941), 
            .I3(GND_net), .O(n18084));   // verilog/coms.v(126[12] 293[6])
    defparam i13255_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 rem_4_i857_3_lut (.I0(n1256), .I1(n1323), .I2(n1283), .I3(GND_net), 
            .O(n1355));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i857_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13002_3_lut (.I0(Kp[10]), .I1(\data_in_frame[2] [2]), .I2(n34066), 
            .I3(GND_net), .O(n17831));   // verilog/coms.v(126[12] 293[6])
    defparam i13002_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 rem_4_i856_3_lut (.I0(n1255), .I1(n1322), .I2(n1283), .I3(GND_net), 
            .O(n1354));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i856_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13256_3_lut (.I0(\data_in_frame[9] [3]), .I1(rx_data[3]), .I2(n32941), 
            .I3(GND_net), .O(n18085));   // verilog/coms.v(126[12] 293[6])
    defparam i13256_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13257_3_lut (.I0(\data_in_frame[9] [4]), .I1(rx_data[4]), .I2(n32941), 
            .I3(GND_net), .O(n18086));   // verilog/coms.v(126[12] 293[6])
    defparam i13257_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 rem_4_i2144_3_lut (.I0(n3151), .I1(n3218_adj_4894), .I2(n3164_adj_4884), 
            .I3(GND_net), .O(n3250));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i2144_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i2147_3_lut (.I0(n3154), .I1(n3221_adj_4897), .I2(n3164_adj_4884), 
            .I3(GND_net), .O(n3253));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i2147_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i2143_3_lut (.I0(n3150), .I1(n3217_adj_4893), .I2(n3164_adj_4884), 
            .I3(GND_net), .O(n3249));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i2143_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i2125_3_lut (.I0(n3132), .I1(n3199), .I2(n3164_adj_4884), 
            .I3(GND_net), .O(n3231_adj_4903));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i2125_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY rem_4_add_1787_14 (.CI(n27886), .I0(n2646), .I1(n2669), .CO(n27887));
    SB_LUT4 i13426_3_lut (.I0(encoder1_position[22]), .I1(n3160), .I2(count_enable_adj_4807), 
            .I3(GND_net), .O(n18255));   // quad.v(35[10] 41[6])
    defparam i13426_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13258_3_lut (.I0(\data_in_frame[9] [5]), .I1(rx_data[5]), .I2(n32941), 
            .I3(GND_net), .O(n18087));   // verilog/coms.v(126[12] 293[6])
    defparam i13258_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 rem_4_i790_3_lut (.I0(n1157), .I1(n1224), .I2(n1184), .I3(GND_net), 
            .O(n1256));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i790_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13003_3_lut (.I0(Kp[11]), .I1(\data_in_frame[2] [3]), .I2(n34066), 
            .I3(GND_net), .O(n17832));   // verilog/coms.v(126[12] 293[6])
    defparam i13003_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 rem_4_i789_3_lut (.I0(n1156), .I1(n1223), .I2(n1184), .I3(GND_net), 
            .O(n1255));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i789_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i2139_3_lut (.I0(n3146), .I1(n3213_adj_4889), .I2(n3164_adj_4884), 
            .I3(GND_net), .O(n3245));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i2139_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i723_3_lut (.I0(n1058), .I1(n1125), .I2(n1085), .I3(GND_net), 
            .O(n1157));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i723_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i722_3_lut (.I0(n1057), .I1(n1124), .I2(n1085), .I3(GND_net), 
            .O(n1156));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i722_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_mux_3_i26_3_lut (.I0(communication_counter[25]), .I1(n8_adj_4876), 
            .I2(communication_counter[31]), .I3(GND_net), .O(n1058));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_mux_3_i26_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_add_2122_20_lut (.I0(GND_net), .I1(n3141), .I2(VCC_net), 
            .I3(n28668), .O(n3208)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2122_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_i2146_3_lut (.I0(n3153), .I1(n3220_adj_4896), .I2(n3164_adj_4884), 
            .I3(GND_net), .O(n3252));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i2146_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i655_3_lut (.I0(n958), .I1(n1025), .I2(n986), .I3(GND_net), 
            .O(n1057));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i655_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i652_3_lut (.I0(n955), .I1(n1022), .I2(n986), .I3(GND_net), 
            .O(n1054));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i652_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i2140_3_lut (.I0(n3147), .I1(n3214_adj_4890), .I2(n3164_adj_4884), 
            .I3(GND_net), .O(n3246));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i2140_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_mux_3_i27_3_lut (.I0(communication_counter[26]), .I1(n7_adj_4877), 
            .I2(communication_counter[31]), .I3(GND_net), .O(n958));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_mux_3_i27_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_mux_3_i30_3_lut (.I0(communication_counter[29]), .I1(n4_adj_4880), 
            .I2(communication_counter[31]), .I3(GND_net), .O(n748));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_mux_3_i30_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i27066_2_lut (.I0(n36410), .I1(n746), .I2(GND_net), .I3(GND_net), 
            .O(n953));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam i27066_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 rem_4_add_1452_7_lut (.I0(GND_net), .I1(n2153), .I2(VCC_net), 
            .I3(n28219), .O(n2220)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1452_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_2122_20 (.CI(n28668), .I0(n3141), .I1(VCC_net), 
            .CO(n28669));
    SB_LUT4 rem_4_add_2122_19_lut (.I0(GND_net), .I1(n3142), .I2(VCC_net), 
            .I3(n28667), .O(n3209_adj_4885)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2122_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i13425_3_lut (.I0(encoder1_position[21]), .I1(n3161), .I2(count_enable_adj_4807), 
            .I3(GND_net), .O(n18254));   // quad.v(35[10] 41[6])
    defparam i13425_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY rem_4_add_2122_19 (.CI(n28667), .I0(n3142), .I1(VCC_net), 
            .CO(n28668));
    SB_LUT4 rem_4_add_2122_18_lut (.I0(GND_net), .I1(n3143), .I2(VCC_net), 
            .I3(n28666), .O(n3210_adj_4886)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2122_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i13432_3_lut (.I0(quadA_debounced), .I1(reg_B[1]), .I2(n34970), 
            .I3(GND_net), .O(n18261));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(186[9] 190[16])
    defparam i13432_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13435_3_lut (.I0(quadA_debounced_adj_4805), .I1(reg_B_adj_5056[1]), 
            .I2(n34971), .I3(GND_net), .O(n18264));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(186[9] 190[16])
    defparam i13435_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY rem_4_add_1452_7 (.CI(n28219), .I0(n2153), .I1(VCC_net), 
            .CO(n28220));
    SB_CARRY rem_4_add_2122_18 (.CI(n28666), .I0(n3143), .I1(VCC_net), 
            .CO(n28667));
    SB_LUT4 rem_4_add_2122_17_lut (.I0(GND_net), .I1(n3144), .I2(VCC_net), 
            .I3(n28665), .O(n3211_adj_4887)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2122_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_2122_17 (.CI(n28665), .I0(n3144), .I1(VCC_net), 
            .CO(n28666));
    SB_LUT4 rem_4_add_2122_16_lut (.I0(GND_net), .I1(n3145), .I2(VCC_net), 
            .I3(n28664), .O(n3212_adj_4888)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2122_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_2122_16 (.CI(n28664), .I0(n3145), .I1(VCC_net), 
            .CO(n28665));
    SB_LUT4 rem_4_add_2122_15_lut (.I0(GND_net), .I1(n3146), .I2(VCC_net), 
            .I3(n28663), .O(n3213_adj_4889)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2122_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_2122_15 (.CI(n28663), .I0(n3146), .I1(VCC_net), 
            .CO(n28664));
    SB_LUT4 rem_4_add_2122_14_lut (.I0(GND_net), .I1(n3147), .I2(VCC_net), 
            .I3(n28662), .O(n3214_adj_4890)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2122_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_2122_14 (.CI(n28662), .I0(n3147), .I1(VCC_net), 
            .CO(n28663));
    SB_LUT4 rem_4_add_2122_13_lut (.I0(GND_net), .I1(n3148), .I2(VCC_net), 
            .I3(n28661), .O(n3215_adj_4891)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2122_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_i2142_3_lut (.I0(n3149), .I1(n3216_adj_4892), .I2(n3164_adj_4884), 
            .I3(GND_net), .O(n3248));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i2142_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i2137_3_lut (.I0(n3144), .I1(n3211_adj_4887), .I2(n3164_adj_4884), 
            .I3(GND_net), .O(n3243));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i2137_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13004_3_lut (.I0(Kp[12]), .I1(\data_in_frame[2] [4]), .I2(n34066), 
            .I3(GND_net), .O(n17833));   // verilog/coms.v(126[12] 293[6])
    defparam i13004_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 rem_4_mux_3_i4_3_lut (.I0(communication_counter[3]), .I1(n30_adj_4854), 
            .I2(communication_counter[31]), .I3(GND_net), .O(n3258));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_mux_3_i4_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i2151_3_lut (.I0(n3158), .I1(n3225_adj_4901), .I2(n3164_adj_4884), 
            .I3(GND_net), .O(n3257));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i2151_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i2150_3_lut (.I0(n3157), .I1(n3224_adj_4900), .I2(n3164_adj_4884), 
            .I3(GND_net), .O(n3256));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i2150_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i2058_3_lut (.I0(n3033), .I1(n3100), .I2(n3065), .I3(GND_net), 
            .O(n3132));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i2058_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i2079_3_lut (.I0(n3054), .I1(n3121), .I2(n3065), .I3(GND_net), 
            .O(n3153));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i2079_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_add_1452_6_lut (.I0(GND_net), .I1(n2154), .I2(GND_net), 
            .I3(n28218), .O(n2221)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1452_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i13005_3_lut (.I0(Kp[13]), .I1(\data_in_frame[2] [5]), .I2(n34066), 
            .I3(GND_net), .O(n17834));   // verilog/coms.v(126[12] 293[6])
    defparam i13005_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13006_3_lut (.I0(Kp[14]), .I1(\data_in_frame[2] [6]), .I2(n34066), 
            .I3(GND_net), .O(n17835));   // verilog/coms.v(126[12] 293[6])
    defparam i13006_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13007_3_lut (.I0(Kp[15]), .I1(\data_in_frame[2] [7]), .I2(n34066), 
            .I3(GND_net), .O(n17836));   // verilog/coms.v(126[12] 293[6])
    defparam i13007_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13008_3_lut (.I0(Ki[1]), .I1(\data_in_frame[5] [1]), .I2(n34066), 
            .I3(GND_net), .O(n17837));   // verilog/coms.v(126[12] 293[6])
    defparam i13008_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 rem_4_i2072_3_lut (.I0(n3047), .I1(n3114), .I2(n3065), .I3(GND_net), 
            .O(n3146));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i2072_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i2069_3_lut (.I0(n3044), .I1(n3111), .I2(n3065), .I3(GND_net), 
            .O(n3143));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i2069_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i2071_3_lut (.I0(n3046), .I1(n3113), .I2(n3065), .I3(GND_net), 
            .O(n3145));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i2071_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i2074_3_lut (.I0(n3049), .I1(n3116), .I2(n3065), .I3(GND_net), 
            .O(n3148));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i2074_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY rem_4_add_2122_13 (.CI(n28661), .I0(n3148), .I1(VCC_net), 
            .CO(n28662));
    SB_LUT4 rem_4_i2073_3_lut (.I0(n3048), .I1(n3115), .I2(n3065), .I3(GND_net), 
            .O(n3147));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i2073_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i2075_3_lut (.I0(n3050), .I1(n3117), .I2(n3065), .I3(GND_net), 
            .O(n3149));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i2075_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i2078_3_lut (.I0(n3053), .I1(n3120), .I2(n3065), .I3(GND_net), 
            .O(n3152));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i2078_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i2064_3_lut (.I0(n3039), .I1(n3106), .I2(n3065), .I3(GND_net), 
            .O(n3138));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i2064_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13259_3_lut (.I0(\data_in_frame[9] [6]), .I1(rx_data[6]), .I2(n32941), 
            .I3(GND_net), .O(n18088));   // verilog/coms.v(126[12] 293[6])
    defparam i13259_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 rem_4_add_2122_12_lut (.I0(GND_net), .I1(n3149), .I2(VCC_net), 
            .I3(n28660), .O(n3216_adj_4892)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2122_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_2122_12 (.CI(n28660), .I0(n3149), .I1(VCC_net), 
            .CO(n28661));
    SB_LUT4 rem_4_add_2122_11_lut (.I0(GND_net), .I1(n3150), .I2(VCC_net), 
            .I3(n28659), .O(n3217_adj_4893)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2122_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_2122_11 (.CI(n28659), .I0(n3150), .I1(VCC_net), 
            .CO(n28660));
    SB_LUT4 rem_4_add_2122_10_lut (.I0(GND_net), .I1(n3151), .I2(VCC_net), 
            .I3(n28658), .O(n3218_adj_4894)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2122_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_2122_10 (.CI(n28658), .I0(n3151), .I1(VCC_net), 
            .CO(n28659));
    SB_LUT4 i12945_3_lut (.I0(IntegralLimit[7]), .I1(\data_in_frame[13] [7]), 
            .I2(n5439), .I3(GND_net), .O(n17774));   // verilog/coms.v(126[12] 293[6])
    defparam i12945_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13009_3_lut (.I0(Ki[2]), .I1(\data_in_frame[5] [2]), .I2(n34066), 
            .I3(GND_net), .O(n17838));   // verilog/coms.v(126[12] 293[6])
    defparam i13009_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12946_3_lut (.I0(IntegralLimit[8]), .I1(\data_in_frame[12] [0]), 
            .I2(n5439), .I3(GND_net), .O(n17775));   // verilog/coms.v(126[12] 293[6])
    defparam i12946_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i2062_3_lut (.I0(n3037), .I1(n3104), .I2(n3065), .I3(GND_net), 
            .O(n3136));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i2062_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_add_2122_9_lut (.I0(GND_net), .I1(n3152), .I2(VCC_net), 
            .I3(n28657), .O(n3219_adj_4895)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2122_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_2122_9 (.CI(n28657), .I0(n3152), .I1(VCC_net), 
            .CO(n28658));
    SB_LUT4 rem_4_add_2122_8_lut (.I0(GND_net), .I1(n3153), .I2(VCC_net), 
            .I3(n28656), .O(n3220_adj_4896)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2122_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_2122_8 (.CI(n28656), .I0(n3153), .I1(VCC_net), 
            .CO(n28657));
    SB_LUT4 rem_4_add_2122_7_lut (.I0(GND_net), .I1(n3154), .I2(GND_net), 
            .I3(n28655), .O(n3221_adj_4897)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2122_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_2122_7 (.CI(n28655), .I0(n3154), .I1(GND_net), 
            .CO(n28656));
    SB_LUT4 rem_4_add_2122_6_lut (.I0(GND_net), .I1(n3155), .I2(GND_net), 
            .I3(n28654), .O(n3222_adj_4898)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2122_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_2122_6 (.CI(n28654), .I0(n3155), .I1(GND_net), 
            .CO(n28655));
    SB_LUT4 rem_4_add_2122_5_lut (.I0(GND_net), .I1(n3156), .I2(VCC_net), 
            .I3(n28653), .O(n3223_adj_4899)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2122_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_2122_5 (.CI(n28653), .I0(n3156), .I1(VCC_net), 
            .CO(n28654));
    SB_LUT4 rem_4_add_2122_4_lut (.I0(GND_net), .I1(n3157), .I2(VCC_net), 
            .I3(n28652), .O(n3224_adj_4900)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2122_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_2122_4 (.CI(n28652), .I0(n3157), .I1(VCC_net), 
            .CO(n28653));
    SB_LUT4 rem_4_add_1787_24_lut (.I0(n2636), .I1(n2636), .I2(n2669), 
            .I3(n27896), .O(n2735)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1787_24_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 rem_4_add_2122_3_lut (.I0(GND_net), .I1(n3158), .I2(GND_net), 
            .I3(n28651), .O(n3225_adj_4901)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2122_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_i2063_3_lut (.I0(n3038), .I1(n3105), .I2(n3065), .I3(GND_net), 
            .O(n3137));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i2063_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13260_3_lut (.I0(\data_in_frame[9] [7]), .I1(rx_data[7]), .I2(n32941), 
            .I3(GND_net), .O(n18089));   // verilog/coms.v(126[12] 293[6])
    defparam i13260_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 rem_4_i2061_3_lut (.I0(n3036), .I1(n3103), .I2(n3065), .I3(GND_net), 
            .O(n3135));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i2061_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i2066_3_lut (.I0(n3041), .I1(n3108), .I2(n3065), .I3(GND_net), 
            .O(n3140));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i2066_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY rem_4_add_2122_3 (.CI(n28651), .I0(n3158), .I1(GND_net), 
            .CO(n28652));
    SB_CARRY rem_4_add_2122_2 (.CI(VCC_net), .I0(n3258), .I1(VCC_net), 
            .CO(n28651));
    SB_LUT4 rem_4_add_2055_29_lut (.I0(n3065), .I1(n3032), .I2(VCC_net), 
            .I3(n28650), .O(n3131)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2055_29_lut.LUT_INIT = 16'h8228;
    SB_LUT4 rem_4_add_1787_23_lut (.I0(n2637), .I1(n2637), .I2(n2669), 
            .I3(n27895), .O(n2736)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1787_23_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 rem_4_add_2055_28_lut (.I0(GND_net), .I1(n3033), .I2(VCC_net), 
            .I3(n28649), .O(n3100)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2055_28_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_2055_28 (.CI(n28649), .I0(n3033), .I1(VCC_net), 
            .CO(n28650));
    SB_LUT4 rem_4_add_2055_27_lut (.I0(GND_net), .I1(n3034), .I2(VCC_net), 
            .I3(n28648), .O(n3101)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2055_27_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_2055_27 (.CI(n28648), .I0(n3034), .I1(VCC_net), 
            .CO(n28649));
    SB_LUT4 rem_4_add_2055_26_lut (.I0(GND_net), .I1(n3035), .I2(VCC_net), 
            .I3(n28647), .O(n3102)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2055_26_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_2055_26 (.CI(n28647), .I0(n3035), .I1(VCC_net), 
            .CO(n28648));
    SB_LUT4 rem_4_add_2055_25_lut (.I0(GND_net), .I1(n3036), .I2(VCC_net), 
            .I3(n28646), .O(n3103)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2055_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_2055_25 (.CI(n28646), .I0(n3036), .I1(VCC_net), 
            .CO(n28647));
    SB_LUT4 rem_4_i2065_3_lut (.I0(n3040), .I1(n3107), .I2(n3065), .I3(GND_net), 
            .O(n3139));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i2065_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF communication_counter_1522__i1 (.Q(communication_counter[1]), .C(LED_c), 
           .D(n164));   // verilog/TinyFPGA_B.v(52[28:51])
    SB_LUT4 rem_4_i2060_3_lut (.I0(n3035), .I1(n3102), .I2(n3065), .I3(GND_net), 
            .O(n3134));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i2060_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i2059_3_lut (.I0(n3034), .I1(n3101), .I2(n3065), .I3(GND_net), 
            .O(n3133));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i2059_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i2081_3_lut (.I0(n3056), .I1(n3123), .I2(n3065), .I3(GND_net), 
            .O(n3155));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i2081_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i2067_3_lut (.I0(n3042), .I1(n3109), .I2(n3065), .I3(GND_net), 
            .O(n3141));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i2067_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i2080_3_lut (.I0(n3055), .I1(n3122), .I2(n3065), .I3(GND_net), 
            .O(n3154));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i2080_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i2007_3_lut (.I0(n2950), .I1(n3017), .I2(n2966), .I3(GND_net), 
            .O(n3049));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i2007_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_add_2055_24_lut (.I0(GND_net), .I1(n3037), .I2(VCC_net), 
            .I3(n28645), .O(n3104)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2055_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i13320_3_lut (.I0(\data_in_frame[17] [3]), .I1(rx_data[3]), 
            .I2(n32957), .I3(GND_net), .O(n18149));   // verilog/coms.v(126[12] 293[6])
    defparam i13320_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13321_3_lut (.I0(\data_in_frame[17] [4]), .I1(rx_data[4]), 
            .I2(n32957), .I3(GND_net), .O(n18150));   // verilog/coms.v(126[12] 293[6])
    defparam i13321_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY rem_4_add_2055_24 (.CI(n28645), .I0(n3037), .I1(VCC_net), 
            .CO(n28646));
    SB_LUT4 rem_4_add_2055_23_lut (.I0(GND_net), .I1(n3038), .I2(VCC_net), 
            .I3(n28644), .O(n3105)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2055_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i13322_3_lut (.I0(\data_in_frame[17] [5]), .I1(rx_data[5]), 
            .I2(n32957), .I3(GND_net), .O(n18151));   // verilog/coms.v(126[12] 293[6])
    defparam i13322_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY rem_4_add_1787_23 (.CI(n27895), .I0(n2637), .I1(n2669), .CO(n27896));
    SB_LUT4 i13323_3_lut (.I0(\data_in_frame[17] [6]), .I1(rx_data[6]), 
            .I2(n32957), .I3(GND_net), .O(n18152));   // verilog/coms.v(126[12] 293[6])
    defparam i13323_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 rem_4_i2010_3_lut (.I0(n2953), .I1(n3020), .I2(n2966), .I3(GND_net), 
            .O(n3052));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i2010_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13324_3_lut (.I0(\data_in_frame[17] [7]), .I1(rx_data[7]), 
            .I2(n32957), .I3(GND_net), .O(n18153));   // verilog/coms.v(126[12] 293[6])
    defparam i13324_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 rem_4_i2003_3_lut (.I0(n2946), .I1(n3013), .I2(n2966), .I3(GND_net), 
            .O(n3045));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i2003_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY rem_4_add_2055_23 (.CI(n28644), .I0(n3038), .I1(VCC_net), 
            .CO(n28645));
    SB_LUT4 rem_4_add_1787_22_lut (.I0(n2638), .I1(n2638), .I2(n2669), 
            .I3(n27894), .O(n2737)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1787_22_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 rem_4_add_2055_22_lut (.I0(GND_net), .I1(n3039), .I2(VCC_net), 
            .I3(n28643), .O(n3106)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2055_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_2055_22 (.CI(n28643), .I0(n3039), .I1(VCC_net), 
            .CO(n28644));
    SB_CARRY rem_4_add_1787_22 (.CI(n27894), .I0(n2638), .I1(n2669), .CO(n27895));
    SB_LUT4 rem_4_add_2055_21_lut (.I0(GND_net), .I1(n3040), .I2(VCC_net), 
            .I3(n28642), .O(n3107)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2055_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1452_6 (.CI(n28218), .I0(n2154), .I1(GND_net), 
            .CO(n28219));
    SB_CARRY rem_4_add_2055_21 (.CI(n28642), .I0(n3040), .I1(VCC_net), 
            .CO(n28643));
    SB_LUT4 rem_4_add_2055_20_lut (.I0(GND_net), .I1(n3041), .I2(VCC_net), 
            .I3(n28641), .O(n3108)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2055_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_i2004_3_lut (.I0(n2947), .I1(n3014), .I2(n2966), .I3(GND_net), 
            .O(n3046));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i2004_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_add_1787_21_lut (.I0(n2639), .I1(n2639), .I2(n2669), 
            .I3(n27893), .O(n2738)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1787_21_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 rem_4_add_1653_22_lut (.I0(n2471), .I1(n2438), .I2(VCC_net), 
            .I3(n28085), .O(n2537)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1653_22_lut.LUT_INIT = 16'h8228;
    SB_CARRY rem_4_add_2055_20 (.CI(n28641), .I0(n3041), .I1(VCC_net), 
            .CO(n28642));
    SB_LUT4 rem_4_add_2055_19_lut (.I0(GND_net), .I1(n3042), .I2(VCC_net), 
            .I3(n28640), .O(n3109)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2055_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_2055_19 (.CI(n28640), .I0(n3042), .I1(VCC_net), 
            .CO(n28641));
    SB_LUT4 rem_4_add_1653_21_lut (.I0(GND_net), .I1(n2439), .I2(VCC_net), 
            .I3(n28084), .O(n2506)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1653_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_2055_18_lut (.I0(GND_net), .I1(n3043), .I2(VCC_net), 
            .I3(n28639), .O(n3110)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2055_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_2055_18 (.CI(n28639), .I0(n3043), .I1(VCC_net), 
            .CO(n28640));
    SB_LUT4 rem_4_add_2055_17_lut (.I0(GND_net), .I1(n3044), .I2(VCC_net), 
            .I3(n28638), .O(n3111)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2055_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_2055_17 (.CI(n28638), .I0(n3044), .I1(VCC_net), 
            .CO(n28639));
    SB_LUT4 rem_4_add_2055_16_lut (.I0(GND_net), .I1(n3045), .I2(VCC_net), 
            .I3(n28637), .O(n3112)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2055_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_2055_16 (.CI(n28637), .I0(n3045), .I1(VCC_net), 
            .CO(n28638));
    SB_LUT4 rem_4_add_2055_15_lut (.I0(GND_net), .I1(n3046), .I2(VCC_net), 
            .I3(n28636), .O(n3113)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2055_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_2055_15 (.CI(n28636), .I0(n3046), .I1(VCC_net), 
            .CO(n28637));
    SB_LUT4 rem_4_add_2055_14_lut (.I0(GND_net), .I1(n3047), .I2(VCC_net), 
            .I3(n28635), .O(n3114)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2055_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_2055_14 (.CI(n28635), .I0(n3047), .I1(VCC_net), 
            .CO(n28636));
    SB_LUT4 rem_4_add_2055_13_lut (.I0(GND_net), .I1(n3048), .I2(VCC_net), 
            .I3(n28634), .O(n3115)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2055_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_2055_13 (.CI(n28634), .I0(n3048), .I1(VCC_net), 
            .CO(n28635));
    SB_LUT4 rem_4_add_2055_12_lut (.I0(GND_net), .I1(n3049), .I2(VCC_net), 
            .I3(n28633), .O(n3116)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2055_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_2055_12 (.CI(n28633), .I0(n3049), .I1(VCC_net), 
            .CO(n28634));
    SB_LUT4 rem_4_add_2055_11_lut (.I0(GND_net), .I1(n3050), .I2(VCC_net), 
            .I3(n28632), .O(n3117)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2055_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_2055_11 (.CI(n28632), .I0(n3050), .I1(VCC_net), 
            .CO(n28633));
    SB_LUT4 rem_4_add_2055_10_lut (.I0(GND_net), .I1(n3051), .I2(VCC_net), 
            .I3(n28631), .O(n3118)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2055_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_2055_10 (.CI(n28631), .I0(n3051), .I1(VCC_net), 
            .CO(n28632));
    SB_LUT4 rem_4_add_2055_9_lut (.I0(GND_net), .I1(n3052), .I2(VCC_net), 
            .I3(n28630), .O(n3119)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2055_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_2055_9 (.CI(n28630), .I0(n3052), .I1(VCC_net), 
            .CO(n28631));
    SB_LUT4 rem_4_add_2055_8_lut (.I0(GND_net), .I1(n3053), .I2(VCC_net), 
            .I3(n28629), .O(n3120)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2055_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_2055_8 (.CI(n28629), .I0(n3053), .I1(VCC_net), 
            .CO(n28630));
    SB_LUT4 rem_4_add_2055_7_lut (.I0(GND_net), .I1(n3054), .I2(GND_net), 
            .I3(n28628), .O(n3121)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2055_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_2055_7 (.CI(n28628), .I0(n3054), .I1(GND_net), 
            .CO(n28629));
    SB_LUT4 rem_4_add_2055_6_lut (.I0(GND_net), .I1(n3055), .I2(GND_net), 
            .I3(n28627), .O(n3122)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2055_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_2055_6 (.CI(n28627), .I0(n3055), .I1(GND_net), 
            .CO(n28628));
    SB_LUT4 rem_4_add_2055_5_lut (.I0(GND_net), .I1(n3056), .I2(VCC_net), 
            .I3(n28626), .O(n3123)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2055_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_2055_5 (.CI(n28626), .I0(n3056), .I1(VCC_net), 
            .CO(n28627));
    SB_LUT4 rem_4_add_2055_4_lut (.I0(GND_net), .I1(n3057), .I2(VCC_net), 
            .I3(n28625), .O(n3124)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2055_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_2055_4 (.CI(n28625), .I0(n3057), .I1(VCC_net), 
            .CO(n28626));
    SB_LUT4 rem_4_add_2055_3_lut (.I0(GND_net), .I1(n3058), .I2(GND_net), 
            .I3(n28624), .O(n3125)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2055_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_2055_3 (.CI(n28624), .I0(n3058), .I1(GND_net), 
            .CO(n28625));
    SB_CARRY rem_4_add_2055_2 (.CI(VCC_net), .I0(n3158), .I1(VCC_net), 
            .CO(n28624));
    SB_LUT4 rem_4_add_1988_28_lut (.I0(n2966), .I1(n2933), .I2(VCC_net), 
            .I3(n28623), .O(n3032)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1988_28_lut.LUT_INIT = 16'h8228;
    SB_LUT4 rem_4_add_1988_27_lut (.I0(GND_net), .I1(n2934), .I2(VCC_net), 
            .I3(n28622), .O(n3001)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1988_27_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1988_27 (.CI(n28622), .I0(n2934), .I1(VCC_net), 
            .CO(n28623));
    SB_LUT4 rem_4_add_1988_26_lut (.I0(GND_net), .I1(n2935), .I2(VCC_net), 
            .I3(n28621), .O(n3002)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1988_26_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1988_26 (.CI(n28621), .I0(n2935), .I1(VCC_net), 
            .CO(n28622));
    SB_LUT4 rem_4_add_1988_25_lut (.I0(GND_net), .I1(n2936), .I2(VCC_net), 
            .I3(n28620), .O(n3003)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1988_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_i2011_3_lut (.I0(n2954), .I1(n3021), .I2(n2966), .I3(GND_net), 
            .O(n3053));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i2011_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i2005_3_lut (.I0(n2948), .I1(n3015), .I2(n2966), .I3(GND_net), 
            .O(n3047));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i2005_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY rem_4_add_1988_25 (.CI(n28620), .I0(n2936), .I1(VCC_net), 
            .CO(n28621));
    SB_LUT4 rem_4_add_1988_24_lut (.I0(GND_net), .I1(n2937), .I2(VCC_net), 
            .I3(n28619), .O(n3004)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1988_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1787_21 (.CI(n27893), .I0(n2639), .I1(n2669), .CO(n27894));
    SB_CARRY rem_4_add_1988_24 (.CI(n28619), .I0(n2937), .I1(VCC_net), 
            .CO(n28620));
    SB_LUT4 rem_4_add_1787_20_lut (.I0(n2640), .I1(n2640), .I2(n2669), 
            .I3(n27892), .O(n2739)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1787_20_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 rem_4_i2008_3_lut (.I0(n2951), .I1(n3018), .I2(n2966), .I3(GND_net), 
            .O(n3050));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i2008_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_add_1988_23_lut (.I0(GND_net), .I1(n2938), .I2(VCC_net), 
            .I3(n28618), .O(n3005)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1988_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1988_23 (.CI(n28618), .I0(n2938), .I1(VCC_net), 
            .CO(n28619));
    SB_LUT4 rem_4_i2001_3_lut (.I0(n2944), .I1(n3011), .I2(n2966), .I3(GND_net), 
            .O(n3043));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i2001_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_add_1988_22_lut (.I0(GND_net), .I1(n2939), .I2(VCC_net), 
            .I3(n28617), .O(n3006)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1988_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1988_22 (.CI(n28617), .I0(n2939), .I1(VCC_net), 
            .CO(n28618));
    SB_LUT4 rem_4_add_1988_21_lut (.I0(GND_net), .I1(n2940), .I2(VCC_net), 
            .I3(n28616), .O(n3007_adj_4883)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1988_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i29807_2_lut_4_lut (.I0(communication_counter[30]), .I1(n3_adj_4881), 
            .I2(communication_counter[31]), .I3(n6_adj_5000), .O(n36410));
    defparam i29807_2_lut_4_lut.LUT_INIT = 16'hca00;
    SB_LUT4 i22873_2_lut_4_lut (.I0(communication_counter[28]), .I1(n5_adj_4879), 
            .I2(communication_counter[31]), .I3(n855), .O(n4_adj_4781));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam i22873_2_lut_4_lut.LUT_INIT = 16'hffca;
    SB_LUT4 rem_4_i2000_3_lut (.I0(n2943), .I1(n3010), .I2(n2966), .I3(GND_net), 
            .O(n3042));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i2000_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1991_3_lut (.I0(n2934), .I1(n3001), .I2(n2966), .I3(GND_net), 
            .O(n3033));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1991_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i2006_3_lut (.I0(n2949), .I1(n3016), .I2(n2966), .I3(GND_net), 
            .O(n3048));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i2006_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1995_3_lut (.I0(n2938), .I1(n3005), .I2(n2966), .I3(GND_net), 
            .O(n3037));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1995_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY rem_4_add_1988_21 (.CI(n28616), .I0(n2940), .I1(VCC_net), 
            .CO(n28617));
    SB_LUT4 rem_4_add_1988_20_lut (.I0(GND_net), .I1(n2941), .I2(VCC_net), 
            .I3(n28615), .O(n3008)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1988_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1988_20 (.CI(n28615), .I0(n2941), .I1(VCC_net), 
            .CO(n28616));
    SB_LUT4 rem_4_add_1988_19_lut (.I0(GND_net), .I1(n2942), .I2(VCC_net), 
            .I3(n28614), .O(n3009)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1988_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1452_5_lut (.I0(GND_net), .I1(n2155), .I2(GND_net), 
            .I3(n28217), .O(n2222)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1452_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1653_21 (.CI(n28084), .I0(n2439), .I1(VCC_net), 
            .CO(n28085));
    SB_LUT4 rem_4_i1993_3_lut (.I0(n2936), .I1(n3003), .I2(n2966), .I3(GND_net), 
            .O(n3035));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1993_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1994_3_lut (.I0(n2937), .I1(n3004), .I2(n2966), .I3(GND_net), 
            .O(n3036));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1994_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1992_3_lut (.I0(n2935), .I1(n3002), .I2(n2966), .I3(GND_net), 
            .O(n3034));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1992_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1999_3_lut (.I0(n2942), .I1(n3009), .I2(n2966), .I3(GND_net), 
            .O(n3041));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1999_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i31515_1_lut_3_lut (.I0(n3353), .I1(n10390), .I2(n3362), .I3(GND_net), 
            .O(n38197));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam i31515_1_lut_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1997_3_lut (.I0(n2940), .I1(n3007_adj_4883), .I2(n2966), 
            .I3(GND_net), .O(n3039));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1997_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1998_3_lut (.I0(n2941), .I1(n3008), .I2(n2966), .I3(GND_net), 
            .O(n3040));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1998_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1996_3_lut (.I0(n2939), .I1(n3006), .I2(n2966), .I3(GND_net), 
            .O(n3038));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1996_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i2013_3_lut (.I0(n2956), .I1(n3023), .I2(n2966), .I3(GND_net), 
            .O(n3055));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i2013_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i2002_3_lut (.I0(n2945), .I1(n3012), .I2(n2966), .I3(GND_net), 
            .O(n3044));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i2002_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i2012_3_lut (.I0(n2955), .I1(n3022), .I2(n2966), .I3(GND_net), 
            .O(n3054));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i2012_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i31089_3_lut (.I0(n2750), .I1(n2817), .I2(n2768), .I3(GND_net), 
            .O(n2849));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam i31089_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i31090_3_lut (.I0(n2849), .I1(n2916), .I2(n2867), .I3(GND_net), 
            .O(n2948));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam i31090_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1943_3_lut (.I0(n2854), .I1(n2921), .I2(n2867), .I3(GND_net), 
            .O(n2953));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1943_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1934_3_lut (.I0(n2845), .I1(n2912), .I2(n2867), .I3(GND_net), 
            .O(n2944));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1934_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i31093_3_lut (.I0(n2753), .I1(n2820), .I2(n2768), .I3(GND_net), 
            .O(n2852));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam i31093_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i31094_3_lut (.I0(n2852), .I1(n2919), .I2(n2867), .I3(GND_net), 
            .O(n2951));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam i31094_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY rem_4_add_1988_19 (.CI(n28614), .I0(n2942), .I1(VCC_net), 
            .CO(n28615));
    SB_LUT4 rem_4_add_1988_18_lut (.I0(GND_net), .I1(n2943), .I2(VCC_net), 
            .I3(n28613), .O(n3010)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1988_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1988_18 (.CI(n28613), .I0(n2943), .I1(VCC_net), 
            .CO(n28614));
    SB_LUT4 rem_4_add_1988_17_lut (.I0(GND_net), .I1(n2944), .I2(VCC_net), 
            .I3(n28612), .O(n3011)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1988_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1988_17 (.CI(n28612), .I0(n2944), .I1(VCC_net), 
            .CO(n28613));
    SB_LUT4 rem_4_add_1988_16_lut (.I0(GND_net), .I1(n2945), .I2(VCC_net), 
            .I3(n28611), .O(n3012)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1988_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1988_16 (.CI(n28611), .I0(n2945), .I1(VCC_net), 
            .CO(n28612));
    SB_LUT4 rem_4_add_1988_15_lut (.I0(GND_net), .I1(n2946), .I2(VCC_net), 
            .I3(n28610), .O(n3013)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1988_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1988_15 (.CI(n28610), .I0(n2946), .I1(VCC_net), 
            .CO(n28611));
    SB_LUT4 rem_4_add_1988_14_lut (.I0(GND_net), .I1(n2947), .I2(VCC_net), 
            .I3(n28609), .O(n3014)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1988_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1988_14 (.CI(n28609), .I0(n2947), .I1(VCC_net), 
            .CO(n28610));
    SB_LUT4 rem_4_add_1988_13_lut (.I0(GND_net), .I1(n2948), .I2(VCC_net), 
            .I3(n28608), .O(n3015)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1988_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1988_13 (.CI(n28608), .I0(n2948), .I1(VCC_net), 
            .CO(n28609));
    SB_LUT4 rem_4_add_1988_12_lut (.I0(GND_net), .I1(n2949), .I2(VCC_net), 
            .I3(n28607), .O(n3016)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1988_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1988_12 (.CI(n28607), .I0(n2949), .I1(VCC_net), 
            .CO(n28608));
    SB_LUT4 rem_4_add_1988_11_lut (.I0(GND_net), .I1(n2950), .I2(VCC_net), 
            .I3(n28606), .O(n3017)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1988_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1988_11 (.CI(n28606), .I0(n2950), .I1(VCC_net), 
            .CO(n28607));
    SB_LUT4 rem_4_add_1988_10_lut (.I0(GND_net), .I1(n2951), .I2(VCC_net), 
            .I3(n28605), .O(n3018)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1988_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1988_10 (.CI(n28605), .I0(n2951), .I1(VCC_net), 
            .CO(n28606));
    SB_LUT4 rem_4_add_1988_9_lut (.I0(GND_net), .I1(n2952), .I2(VCC_net), 
            .I3(n28604), .O(n3019)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1988_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1988_9 (.CI(n28604), .I0(n2952), .I1(VCC_net), 
            .CO(n28605));
    SB_LUT4 rem_4_add_1988_8_lut (.I0(GND_net), .I1(n2953), .I2(VCC_net), 
            .I3(n28603), .O(n3020)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1988_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1988_8 (.CI(n28603), .I0(n2953), .I1(VCC_net), 
            .CO(n28604));
    SB_LUT4 rem_4_add_1988_7_lut (.I0(GND_net), .I1(n2954), .I2(GND_net), 
            .I3(n28602), .O(n3021)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1988_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1988_7 (.CI(n28602), .I0(n2954), .I1(GND_net), 
            .CO(n28603));
    SB_LUT4 rem_4_add_1988_6_lut (.I0(GND_net), .I1(n2955), .I2(GND_net), 
            .I3(n28601), .O(n3022)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1988_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1988_6 (.CI(n28601), .I0(n2955), .I1(GND_net), 
            .CO(n28602));
    SB_LUT4 rem_4_add_1988_5_lut (.I0(GND_net), .I1(n2956), .I2(VCC_net), 
            .I3(n28600), .O(n3023)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1988_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1988_5 (.CI(n28600), .I0(n2956), .I1(VCC_net), 
            .CO(n28601));
    SB_LUT4 rem_4_add_1988_4_lut (.I0(GND_net), .I1(n2957), .I2(VCC_net), 
            .I3(n28599), .O(n3024)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1988_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1988_4 (.CI(n28599), .I0(n2957), .I1(VCC_net), 
            .CO(n28600));
    SB_LUT4 rem_4_add_1988_3_lut (.I0(GND_net), .I1(n2958_adj_4882), .I2(GND_net), 
            .I3(n28598), .O(n3025)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1988_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1988_3 (.CI(n28598), .I0(n2958_adj_4882), .I1(GND_net), 
            .CO(n28599));
    SB_CARRY rem_4_add_1988_2 (.CI(VCC_net), .I0(n3058), .I1(VCC_net), 
            .CO(n28598));
    SB_LUT4 rem_4_add_1921_27_lut (.I0(n2867), .I1(n2834), .I2(VCC_net), 
            .I3(n28597), .O(n2933)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1921_27_lut.LUT_INIT = 16'h8228;
    SB_LUT4 rem_4_add_1921_26_lut (.I0(GND_net), .I1(n2835), .I2(VCC_net), 
            .I3(n28596), .O(n2902)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1921_26_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1921_26 (.CI(n28596), .I0(n2835), .I1(VCC_net), 
            .CO(n28597));
    SB_LUT4 rem_4_add_1921_25_lut (.I0(GND_net), .I1(n2836), .I2(VCC_net), 
            .I3(n28595), .O(n2903)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1921_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1921_25 (.CI(n28595), .I0(n2836), .I1(VCC_net), 
            .CO(n28596));
    SB_LUT4 rem_4_add_1921_24_lut (.I0(GND_net), .I1(n2837), .I2(VCC_net), 
            .I3(n28594), .O(n2904)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1921_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1921_24 (.CI(n28594), .I0(n2837), .I1(VCC_net), 
            .CO(n28595));
    SB_LUT4 rem_4_add_1921_23_lut (.I0(GND_net), .I1(n2838), .I2(VCC_net), 
            .I3(n28593), .O(n2905)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1921_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1921_23 (.CI(n28593), .I0(n2838), .I1(VCC_net), 
            .CO(n28594));
    SB_LUT4 rem_4_add_1921_22_lut (.I0(GND_net), .I1(n2839), .I2(VCC_net), 
            .I3(n28592), .O(n2906)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1921_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1921_22 (.CI(n28592), .I0(n2839), .I1(VCC_net), 
            .CO(n28593));
    SB_LUT4 rem_4_add_1921_21_lut (.I0(GND_net), .I1(n2840), .I2(VCC_net), 
            .I3(n28591), .O(n2907)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1921_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1921_21 (.CI(n28591), .I0(n2840), .I1(VCC_net), 
            .CO(n28592));
    SB_LUT4 rem_4_add_1921_20_lut (.I0(GND_net), .I1(n2841), .I2(VCC_net), 
            .I3(n28590), .O(n2908)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1921_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1921_20 (.CI(n28590), .I0(n2841), .I1(VCC_net), 
            .CO(n28591));
    SB_LUT4 rem_4_add_1921_19_lut (.I0(GND_net), .I1(n2842), .I2(VCC_net), 
            .I3(n28589), .O(n2909)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1921_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1921_19 (.CI(n28589), .I0(n2842), .I1(VCC_net), 
            .CO(n28590));
    SB_LUT4 rem_4_add_1921_18_lut (.I0(GND_net), .I1(n2843), .I2(VCC_net), 
            .I3(n28588), .O(n2910)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1921_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1921_18 (.CI(n28588), .I0(n2843), .I1(VCC_net), 
            .CO(n28589));
    SB_LUT4 rem_4_add_1921_17_lut (.I0(GND_net), .I1(n2844), .I2(VCC_net), 
            .I3(n28587), .O(n2911)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1921_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1921_17 (.CI(n28587), .I0(n2844), .I1(VCC_net), 
            .CO(n28588));
    SB_LUT4 rem_4_add_1921_16_lut (.I0(GND_net), .I1(n2845), .I2(VCC_net), 
            .I3(n28586), .O(n2912)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1921_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1921_16 (.CI(n28586), .I0(n2845), .I1(VCC_net), 
            .CO(n28587));
    SB_LUT4 rem_4_add_1921_15_lut (.I0(GND_net), .I1(n2846), .I2(VCC_net), 
            .I3(n28585), .O(n2913)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1921_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1921_15 (.CI(n28585), .I0(n2846), .I1(VCC_net), 
            .CO(n28586));
    SB_LUT4 rem_4_add_1921_14_lut (.I0(GND_net), .I1(n2847), .I2(VCC_net), 
            .I3(n28584), .O(n2914)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1921_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1921_14 (.CI(n28584), .I0(n2847), .I1(VCC_net), 
            .CO(n28585));
    SB_LUT4 rem_4_add_1921_13_lut (.I0(GND_net), .I1(n2848), .I2(VCC_net), 
            .I3(n28583), .O(n2915)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1921_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1921_13 (.CI(n28583), .I0(n2848), .I1(VCC_net), 
            .CO(n28584));
    SB_LUT4 rem_4_add_1921_12_lut (.I0(GND_net), .I1(n2849), .I2(VCC_net), 
            .I3(n28582), .O(n2916)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1921_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1921_12 (.CI(n28582), .I0(n2849), .I1(VCC_net), 
            .CO(n28583));
    SB_LUT4 rem_4_add_1921_11_lut (.I0(GND_net), .I1(n2850), .I2(VCC_net), 
            .I3(n28581), .O(n2917)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1921_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1921_11 (.CI(n28581), .I0(n2850), .I1(VCC_net), 
            .CO(n28582));
    SB_LUT4 rem_4_add_1921_10_lut (.I0(GND_net), .I1(n2851), .I2(VCC_net), 
            .I3(n28580), .O(n2918)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1921_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1921_10 (.CI(n28580), .I0(n2851), .I1(VCC_net), 
            .CO(n28581));
    SB_LUT4 rem_4_add_1921_9_lut (.I0(GND_net), .I1(n2852), .I2(VCC_net), 
            .I3(n28579), .O(n2919)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1921_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1921_9 (.CI(n28579), .I0(n2852), .I1(VCC_net), 
            .CO(n28580));
    SB_LUT4 rem_4_add_1921_8_lut (.I0(GND_net), .I1(n2853), .I2(VCC_net), 
            .I3(n28578), .O(n2920)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1921_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1921_8 (.CI(n28578), .I0(n2853), .I1(VCC_net), 
            .CO(n28579));
    SB_LUT4 rem_4_add_1921_7_lut (.I0(GND_net), .I1(n2854), .I2(GND_net), 
            .I3(n28577), .O(n2921)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1921_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1921_7 (.CI(n28577), .I0(n2854), .I1(GND_net), 
            .CO(n28578));
    SB_LUT4 rem_4_add_1921_6_lut (.I0(GND_net), .I1(n2855), .I2(GND_net), 
            .I3(n28576), .O(n2922)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1921_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1921_6 (.CI(n28576), .I0(n2855), .I1(GND_net), 
            .CO(n28577));
    SB_LUT4 rem_4_add_1921_5_lut (.I0(GND_net), .I1(n2856), .I2(VCC_net), 
            .I3(n28575), .O(n2923)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1921_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1921_5 (.CI(n28575), .I0(n2856), .I1(VCC_net), 
            .CO(n28576));
    SB_LUT4 rem_4_add_1921_4_lut (.I0(GND_net), .I1(n2857), .I2(VCC_net), 
            .I3(n28574), .O(n2924)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1921_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1921_4 (.CI(n28574), .I0(n2857), .I1(VCC_net), 
            .CO(n28575));
    SB_LUT4 rem_4_add_1921_3_lut (.I0(GND_net), .I1(n2759), .I2(GND_net), 
            .I3(n28573), .O(n2925)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1921_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1921_3 (.CI(n28573), .I0(n2759), .I1(GND_net), 
            .CO(n28574));
    SB_CARRY rem_4_add_1921_2 (.CI(VCC_net), .I0(n2958_adj_4882), .I1(VCC_net), 
            .CO(n28573));
    SB_LUT4 rem_4_add_1854_26_lut (.I0(n2768), .I1(n2735), .I2(VCC_net), 
            .I3(n28572), .O(n2834)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1854_26_lut.LUT_INIT = 16'h8228;
    SB_LUT4 rem_4_add_1854_25_lut (.I0(GND_net), .I1(n2736), .I2(VCC_net), 
            .I3(n28571), .O(n2803)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1854_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1854_25 (.CI(n28571), .I0(n2736), .I1(VCC_net), 
            .CO(n28572));
    SB_LUT4 rem_4_add_1854_24_lut (.I0(GND_net), .I1(n2737), .I2(VCC_net), 
            .I3(n28570), .O(n2804)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1854_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1854_24 (.CI(n28570), .I0(n2737), .I1(VCC_net), 
            .CO(n28571));
    SB_LUT4 rem_4_add_1854_23_lut (.I0(GND_net), .I1(n2738), .I2(VCC_net), 
            .I3(n28569), .O(n2805)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1854_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1854_23 (.CI(n28569), .I0(n2738), .I1(VCC_net), 
            .CO(n28570));
    SB_LUT4 rem_4_add_1854_22_lut (.I0(GND_net), .I1(n2739), .I2(VCC_net), 
            .I3(n28568), .O(n2806)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1854_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1854_22 (.CI(n28568), .I0(n2739), .I1(VCC_net), 
            .CO(n28569));
    SB_LUT4 rem_4_i1933_3_lut (.I0(n2844), .I1(n2911), .I2(n2867), .I3(GND_net), 
            .O(n2943));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1933_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i31085_3_lut (.I0(n2748), .I1(n2815), .I2(n2768), .I3(GND_net), 
            .O(n2847));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam i31085_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i31086_3_lut (.I0(n2847), .I1(n2914), .I2(n2867), .I3(GND_net), 
            .O(n2946));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam i31086_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_add_1854_21_lut (.I0(GND_net), .I1(n2740), .I2(VCC_net), 
            .I3(n28567), .O(n2807)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1854_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1854_21 (.CI(n28567), .I0(n2740), .I1(VCC_net), 
            .CO(n28568));
    SB_CARRY rem_4_add_1452_5 (.CI(n28217), .I0(n2155), .I1(GND_net), 
            .CO(n28218));
    SB_LUT4 rem_4_i1932_3_lut (.I0(n2843), .I1(n2910), .I2(n2867), .I3(GND_net), 
            .O(n2942));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1932_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_add_1854_20_lut (.I0(GND_net), .I1(n2741), .I2(VCC_net), 
            .I3(n28566), .O(n2808)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1854_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1653_20_lut (.I0(GND_net), .I1(n2440), .I2(VCC_net), 
            .I3(n28083), .O(n2507)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1653_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1854_20 (.CI(n28566), .I0(n2741), .I1(VCC_net), 
            .CO(n28567));
    SB_CARRY rem_4_add_1653_20 (.CI(n28083), .I0(n2440), .I1(VCC_net), 
            .CO(n28084));
    SB_LUT4 rem_4_add_1854_19_lut (.I0(GND_net), .I1(n2742), .I2(VCC_net), 
            .I3(n28565), .O(n2809)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1854_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1653_19_lut (.I0(GND_net), .I1(n2441), .I2(VCC_net), 
            .I3(n28082), .O(n2508)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1653_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1653_19 (.CI(n28082), .I0(n2441), .I1(VCC_net), 
            .CO(n28083));
    SB_CARRY rem_4_add_1854_19 (.CI(n28565), .I0(n2742), .I1(VCC_net), 
            .CO(n28566));
    SB_LUT4 rem_4_i1931_3_lut (.I0(n2842), .I1(n2909), .I2(n2867), .I3(GND_net), 
            .O(n2941));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1931_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i31083_3_lut (.I0(n2747), .I1(n2814), .I2(n2768), .I3(GND_net), 
            .O(n2846));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam i31083_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_add_1854_18_lut (.I0(GND_net), .I1(n2743), .I2(VCC_net), 
            .I3(n28564), .O(n2810)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1854_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1452_4_lut (.I0(GND_net), .I1(n2156), .I2(VCC_net), 
            .I3(n28216), .O(n2223)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1452_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1452_4 (.CI(n28216), .I0(n2156), .I1(VCC_net), 
            .CO(n28217));
    SB_LUT4 rem_4_add_1452_3_lut (.I0(GND_net), .I1(n2157), .I2(VCC_net), 
            .I3(n28215), .O(n2224)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1452_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1854_18 (.CI(n28564), .I0(n2743), .I1(VCC_net), 
            .CO(n28565));
    SB_LUT4 rem_4_add_1854_17_lut (.I0(GND_net), .I1(n2744), .I2(VCC_net), 
            .I3(n28563), .O(n2811)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1854_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1854_17 (.CI(n28563), .I0(n2744), .I1(VCC_net), 
            .CO(n28564));
    SB_CARRY rem_4_add_1452_3 (.CI(n28215), .I0(n2157), .I1(VCC_net), 
            .CO(n28216));
    SB_LUT4 rem_4_add_1854_16_lut (.I0(GND_net), .I1(n2745), .I2(VCC_net), 
            .I3(n28562), .O(n2812)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1854_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1854_16 (.CI(n28562), .I0(n2745), .I1(VCC_net), 
            .CO(n28563));
    SB_LUT4 rem_4_add_1452_2_lut (.I0(GND_net), .I1(n2158), .I2(GND_net), 
            .I3(VCC_net), .O(n2225)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1452_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i13010_3_lut (.I0(Ki[3]), .I1(\data_in_frame[5] [3]), .I2(n34066), 
            .I3(GND_net), .O(n17839));   // verilog/coms.v(126[12] 293[6])
    defparam i13010_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 rem_4_add_1854_15_lut (.I0(GND_net), .I1(n2746), .I2(VCC_net), 
            .I3(n28561), .O(n2813)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1854_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i31084_3_lut (.I0(n2846), .I1(n2913), .I2(n2867), .I3(GND_net), 
            .O(n2945));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam i31084_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY rem_4_add_1854_15 (.CI(n28561), .I0(n2746), .I1(VCC_net), 
            .CO(n28562));
    SB_LUT4 rem_4_add_1854_14_lut (.I0(GND_net), .I1(n2747), .I2(VCC_net), 
            .I3(n28560), .O(n2814)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1854_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1854_14 (.CI(n28560), .I0(n2747), .I1(VCC_net), 
            .CO(n28561));
    SB_LUT4 rem_4_add_1854_13_lut (.I0(GND_net), .I1(n2748), .I2(VCC_net), 
            .I3(n28559), .O(n2815)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1854_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1854_13 (.CI(n28559), .I0(n2748), .I1(VCC_net), 
            .CO(n28560));
    SB_LUT4 rem_4_i1940_3_lut (.I0(n2851), .I1(n2918), .I2(n2867), .I3(GND_net), 
            .O(n2950));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1940_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_add_1854_12_lut (.I0(GND_net), .I1(n2749), .I2(VCC_net), 
            .I3(n28558), .O(n2816)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1854_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_i1942_3_lut (.I0(n2853), .I1(n2920), .I2(n2867), .I3(GND_net), 
            .O(n2952));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1942_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i31091_3_lut (.I0(n2751), .I1(n2818), .I2(n2768), .I3(GND_net), 
            .O(n2850));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam i31091_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY rem_4_add_1854_12 (.CI(n28558), .I0(n2749), .I1(VCC_net), 
            .CO(n28559));
    SB_LUT4 rem_4_add_1854_11_lut (.I0(GND_net), .I1(n2750), .I2(VCC_net), 
            .I3(n28557), .O(n2817)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1854_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1854_11 (.CI(n28557), .I0(n2750), .I1(VCC_net), 
            .CO(n28558));
    SB_LUT4 rem_4_add_1854_10_lut (.I0(GND_net), .I1(n2751), .I2(VCC_net), 
            .I3(n28556), .O(n2818)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1854_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1787_20 (.CI(n27892), .I0(n2640), .I1(n2669), .CO(n27893));
    SB_CARRY rem_4_add_1452_2 (.CI(VCC_net), .I0(n2158), .I1(GND_net), 
            .CO(n28215));
    SB_LUT4 rem_4_add_1519_20_lut (.I0(n2273), .I1(n2240), .I2(VCC_net), 
            .I3(n28214), .O(n2339)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1519_20_lut.LUT_INIT = 16'h8228;
    SB_CARRY rem_4_add_1854_10 (.CI(n28556), .I0(n2751), .I1(VCC_net), 
            .CO(n28557));
    SB_LUT4 rem_4_add_1653_18_lut (.I0(GND_net), .I1(n2442), .I2(VCC_net), 
            .I3(n28081), .O(n2509)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1653_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1653_18 (.CI(n28081), .I0(n2442), .I1(VCC_net), 
            .CO(n28082));
    SB_LUT4 i31092_3_lut (.I0(n2850), .I1(n2917), .I2(n2867), .I3(GND_net), 
            .O(n2949));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam i31092_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1930_3_lut (.I0(n2841), .I1(n2908), .I2(n2867), .I3(GND_net), 
            .O(n2940));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1930_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_add_1854_9_lut (.I0(GND_net), .I1(n2752), .I2(VCC_net), 
            .I3(n28555), .O(n2819)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1854_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1854_9 (.CI(n28555), .I0(n2752), .I1(VCC_net), 
            .CO(n28556));
    SB_LUT4 rem_4_add_1653_17_lut (.I0(GND_net), .I1(n2443), .I2(VCC_net), 
            .I3(n28080), .O(n2510)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1653_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1653_17 (.CI(n28080), .I0(n2443), .I1(VCC_net), 
            .CO(n28081));
    SB_LUT4 rem_4_add_1854_8_lut (.I0(GND_net), .I1(n2753), .I2(VCC_net), 
            .I3(n28554), .O(n2820)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1854_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1854_8 (.CI(n28554), .I0(n2753), .I1(VCC_net), 
            .CO(n28555));
    SB_LUT4 rem_4_add_1854_7_lut (.I0(GND_net), .I1(n2754), .I2(GND_net), 
            .I3(n28553), .O(n2821)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1854_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1854_7 (.CI(n28553), .I0(n2754), .I1(GND_net), 
            .CO(n28554));
    SB_LUT4 rem_4_add_1854_6_lut (.I0(GND_net), .I1(n2755), .I2(GND_net), 
            .I3(n28552), .O(n2822)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1854_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1854_6 (.CI(n28552), .I0(n2755), .I1(GND_net), 
            .CO(n28553));
    SB_LUT4 rem_4_add_1854_5_lut (.I0(GND_net), .I1(n2756), .I2(VCC_net), 
            .I3(n28551), .O(n2823)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1854_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1854_5 (.CI(n28551), .I0(n2756), .I1(VCC_net), 
            .CO(n28552));
    SB_LUT4 rem_4_add_1854_4_lut (.I0(GND_net), .I1(n2757), .I2(VCC_net), 
            .I3(n28550), .O(n2824)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1854_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1854_4 (.CI(n28550), .I0(n2757), .I1(VCC_net), 
            .CO(n28551));
    SB_LUT4 rem_4_add_1854_3_lut (.I0(GND_net), .I1(n2758), .I2(GND_net), 
            .I3(n28549), .O(n2825)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1854_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1854_3 (.CI(n28549), .I0(n2758), .I1(GND_net), 
            .CO(n28550));
    SB_CARRY rem_4_add_1854_2 (.CI(VCC_net), .I0(n2759), .I1(VCC_net), 
            .CO(n28549));
    SB_LUT4 rem_4_add_648_7_lut (.I0(n986), .I1(n953), .I2(VCC_net), .I3(n28548), 
            .O(n1052)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_648_7_lut.LUT_INIT = 16'h8228;
    SB_LUT4 rem_4_add_648_6_lut (.I0(GND_net), .I1(n954), .I2(GND_net), 
            .I3(n28547), .O(n1021)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_648_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_648_6 (.CI(n28547), .I0(n954), .I1(GND_net), .CO(n28548));
    SB_LUT4 rem_4_add_648_5_lut (.I0(GND_net), .I1(n955), .I2(GND_net), 
            .I3(n28546), .O(n1022)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_648_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_648_5 (.CI(n28546), .I0(n955), .I1(GND_net), .CO(n28547));
    SB_LUT4 rem_4_add_648_4_lut (.I0(GND_net), .I1(n956), .I2(VCC_net), 
            .I3(n28545), .O(n1023)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_648_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_648_4 (.CI(n28545), .I0(n956), .I1(VCC_net), .CO(n28546));
    SB_LUT4 rem_4_add_648_3_lut (.I0(GND_net), .I1(n957), .I2(VCC_net), 
            .I3(n28544), .O(n1024)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_648_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_648_3 (.CI(n28544), .I0(n957), .I1(VCC_net), .CO(n28545));
    SB_LUT4 rem_4_add_648_2_lut (.I0(GND_net), .I1(n958), .I2(GND_net), 
            .I3(VCC_net), .O(n1025)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_648_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_648_2 (.CI(VCC_net), .I0(n958), .I1(GND_net), .CO(n28544));
    SB_LUT4 rem_4_add_715_9_lut (.I0(n1085), .I1(n1052), .I2(VCC_net), 
            .I3(n28543), .O(n1151)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_715_9_lut.LUT_INIT = 16'h8228;
    SB_LUT4 rem_4_add_715_8_lut (.I0(GND_net), .I1(n1053), .I2(VCC_net), 
            .I3(n28542), .O(n1120)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_715_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_715_8 (.CI(n28542), .I0(n1053), .I1(VCC_net), .CO(n28543));
    SB_LUT4 rem_4_add_715_7_lut (.I0(GND_net), .I1(n1054), .I2(GND_net), 
            .I3(n28541), .O(n1121)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_715_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_715_7 (.CI(n28541), .I0(n1054), .I1(GND_net), .CO(n28542));
    SB_LUT4 rem_4_add_715_6_lut (.I0(GND_net), .I1(n1055), .I2(GND_net), 
            .I3(n28540), .O(n1122)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_715_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_715_6 (.CI(n28540), .I0(n1055), .I1(GND_net), .CO(n28541));
    SB_LUT4 rem_4_add_715_5_lut (.I0(GND_net), .I1(n1056), .I2(VCC_net), 
            .I3(n28539), .O(n1123)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_715_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_715_5 (.CI(n28539), .I0(n1056), .I1(VCC_net), .CO(n28540));
    SB_LUT4 rem_4_add_715_4_lut (.I0(GND_net), .I1(n1057), .I2(VCC_net), 
            .I3(n28538), .O(n1124)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_715_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_715_4 (.CI(n28538), .I0(n1057), .I1(VCC_net), .CO(n28539));
    SB_LUT4 i22881_2_lut_4_lut (.I0(communication_counter[29]), .I1(n4_adj_4880), 
            .I2(communication_counter[31]), .I3(n4_adj_4781), .O(n6_adj_5000));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam i22881_2_lut_4_lut.LUT_INIT = 16'hffca;
    SB_LUT4 rem_4_add_715_3_lut (.I0(GND_net), .I1(n1058), .I2(GND_net), 
            .I3(n28537), .O(n1125)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_715_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_715_3 (.CI(n28537), .I0(n1058), .I1(GND_net), .CO(n28538));
    SB_CARRY rem_4_add_715_2 (.CI(VCC_net), .I0(n1158), .I1(VCC_net), 
            .CO(n28537));
    SB_LUT4 rem_4_add_782_10_lut (.I0(n1184), .I1(n1151), .I2(VCC_net), 
            .I3(n28536), .O(n1250)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_782_10_lut.LUT_INIT = 16'h8228;
    SB_LUT4 rem_4_add_782_9_lut (.I0(GND_net), .I1(n1152), .I2(VCC_net), 
            .I3(n28535), .O(n1219)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_782_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_782_9 (.CI(n28535), .I0(n1152), .I1(VCC_net), .CO(n28536));
    SB_LUT4 rem_4_add_782_8_lut (.I0(GND_net), .I1(n1153), .I2(VCC_net), 
            .I3(n28534), .O(n1220)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_782_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_782_8 (.CI(n28534), .I0(n1153), .I1(VCC_net), .CO(n28535));
    SB_LUT4 rem_4_add_782_7_lut (.I0(GND_net), .I1(n1154), .I2(GND_net), 
            .I3(n28533), .O(n1221)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_782_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_782_7 (.CI(n28533), .I0(n1154), .I1(GND_net), .CO(n28534));
    SB_LUT4 rem_4_add_782_6_lut (.I0(GND_net), .I1(n1155), .I2(GND_net), 
            .I3(n28532), .O(n1222)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_782_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_782_6 (.CI(n28532), .I0(n1155), .I1(GND_net), .CO(n28533));
    SB_LUT4 rem_4_add_782_5_lut (.I0(GND_net), .I1(n1156), .I2(VCC_net), 
            .I3(n28531), .O(n1223)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_782_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_782_5 (.CI(n28531), .I0(n1156), .I1(VCC_net), .CO(n28532));
    SB_LUT4 rem_4_add_782_4_lut (.I0(GND_net), .I1(n1157), .I2(VCC_net), 
            .I3(n28530), .O(n1224)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_782_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_782_4 (.CI(n28530), .I0(n1157), .I1(VCC_net), .CO(n28531));
    SB_LUT4 rem_4_add_782_3_lut (.I0(GND_net), .I1(n1158), .I2(GND_net), 
            .I3(n28529), .O(n1225)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_782_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_782_3 (.CI(n28529), .I0(n1158), .I1(GND_net), .CO(n28530));
    SB_CARRY rem_4_add_782_2 (.CI(VCC_net), .I0(n1258), .I1(VCC_net), 
            .CO(n28529));
    SB_LUT4 rem_4_add_849_11_lut (.I0(n1283), .I1(n1250), .I2(VCC_net), 
            .I3(n28528), .O(n1349)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_849_11_lut.LUT_INIT = 16'h8228;
    SB_LUT4 rem_4_add_849_10_lut (.I0(GND_net), .I1(n1251), .I2(VCC_net), 
            .I3(n28527), .O(n1318)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_849_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_849_10 (.CI(n28527), .I0(n1251), .I1(VCC_net), 
            .CO(n28528));
    SB_LUT4 rem_4_add_849_9_lut (.I0(GND_net), .I1(n1252), .I2(VCC_net), 
            .I3(n28526), .O(n1319)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_849_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_849_9 (.CI(n28526), .I0(n1252), .I1(VCC_net), .CO(n28527));
    SB_LUT4 rem_4_add_849_8_lut (.I0(GND_net), .I1(n1253), .I2(VCC_net), 
            .I3(n28525), .O(n1320)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_849_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_849_8 (.CI(n28525), .I0(n1253), .I1(VCC_net), .CO(n28526));
    SB_LUT4 rem_4_add_849_7_lut (.I0(GND_net), .I1(n1254), .I2(GND_net), 
            .I3(n28524), .O(n1321)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_849_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_849_7 (.CI(n28524), .I0(n1254), .I1(GND_net), .CO(n28525));
    SB_LUT4 rem_4_add_849_6_lut (.I0(GND_net), .I1(n1255), .I2(GND_net), 
            .I3(n28523), .O(n1322)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_849_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_849_6 (.CI(n28523), .I0(n1255), .I1(GND_net), .CO(n28524));
    SB_LUT4 rem_4_add_849_5_lut (.I0(GND_net), .I1(n1256), .I2(VCC_net), 
            .I3(n28522), .O(n1323)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_849_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_849_5 (.CI(n28522), .I0(n1256), .I1(VCC_net), .CO(n28523));
    SB_LUT4 rem_4_add_849_4_lut (.I0(GND_net), .I1(n1257), .I2(VCC_net), 
            .I3(n28521), .O(n1324)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_849_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_849_4 (.CI(n28521), .I0(n1257), .I1(VCC_net), .CO(n28522));
    SB_LUT4 rem_4_add_849_3_lut (.I0(GND_net), .I1(n1258), .I2(GND_net), 
            .I3(n28520), .O(n1325)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_849_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_849_3 (.CI(n28520), .I0(n1258), .I1(GND_net), .CO(n28521));
    SB_CARRY rem_4_add_849_2 (.CI(VCC_net), .I0(n1358), .I1(VCC_net), 
            .CO(n28520));
    SB_LUT4 rem_4_add_916_12_lut (.I0(n1382), .I1(n1349), .I2(VCC_net), 
            .I3(n28519), .O(n1448)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_916_12_lut.LUT_INIT = 16'h8228;
    SB_LUT4 rem_4_add_916_11_lut (.I0(GND_net), .I1(n1350), .I2(VCC_net), 
            .I3(n28518), .O(n1417)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_916_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_916_11 (.CI(n28518), .I0(n1350), .I1(VCC_net), 
            .CO(n28519));
    SB_LUT4 rem_4_add_916_10_lut (.I0(GND_net), .I1(n1351), .I2(VCC_net), 
            .I3(n28517), .O(n1418)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_916_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_916_10 (.CI(n28517), .I0(n1351), .I1(VCC_net), 
            .CO(n28518));
    SB_LUT4 i13011_3_lut (.I0(Ki[4]), .I1(\data_in_frame[5] [4]), .I2(n34066), 
            .I3(GND_net), .O(n17840));   // verilog/coms.v(126[12] 293[6])
    defparam i13011_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 rem_4_i1928_3_lut (.I0(n2839), .I1(n2906), .I2(n2867), .I3(GND_net), 
            .O(n2938));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1928_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13012_3_lut (.I0(Ki[5]), .I1(\data_in_frame[5] [5]), .I2(n34066), 
            .I3(GND_net), .O(n17841));   // verilog/coms.v(126[12] 293[6])
    defparam i13012_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 rem_4_i1929_3_lut (.I0(n2840), .I1(n2907), .I2(n2867), .I3(GND_net), 
            .O(n2939));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1929_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1927_3_lut (.I0(n2838), .I1(n2905), .I2(n2867), .I3(GND_net), 
            .O(n2937));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1927_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1926_3_lut (.I0(n2837), .I1(n2904), .I2(n2867), .I3(GND_net), 
            .O(n2936));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1926_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1925_3_lut (.I0(n2836), .I1(n2903), .I2(n2867), .I3(GND_net), 
            .O(n2935));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1925_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1924_3_lut (.I0(n2835), .I1(n2902), .I2(n2867), .I3(GND_net), 
            .O(n2934));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1924_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13013_3_lut (.I0(Ki[6]), .I1(\data_in_frame[5] [6]), .I2(n34066), 
            .I3(GND_net), .O(n17842));   // verilog/coms.v(126[12] 293[6])
    defparam i13013_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 rem_4_i1947_3_lut (.I0(n2759), .I1(n2925), .I2(n2867), .I3(GND_net), 
            .O(n2957));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1947_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1946_3_lut (.I0(n2857), .I1(n2924), .I2(n2867), .I3(GND_net), 
            .O(n2956));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1946_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1865_3_lut (.I0(n2744), .I1(n2811), .I2(n2768), .I3(GND_net), 
            .O(n2843));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1865_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_3_lut_4_lut (.I0(n63), .I1(n24786), .I2(n16158), .I3(n3007), 
            .O(n32973));   // verilog/coms.v(126[12] 293[6])
    defparam i1_3_lut_4_lut.LUT_INIT = 16'h5d55;
    SB_LUT4 rem_4_i1863_3_lut (.I0(n2742), .I1(n2809), .I2(n2768), .I3(GND_net), 
            .O(n2841));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1863_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1864_3_lut (.I0(n2743), .I1(n2810), .I2(n2768), .I3(GND_net), 
            .O(n2842));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1864_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_add_916_9_lut (.I0(GND_net), .I1(n1352), .I2(VCC_net), 
            .I3(n28516), .O(n1419)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_916_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_916_9 (.CI(n28516), .I0(n1352), .I1(VCC_net), .CO(n28517));
    SB_LUT4 rem_4_i1862_3_lut (.I0(n2741), .I1(n2808), .I2(n2768), .I3(GND_net), 
            .O(n2840));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1862_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_add_916_8_lut (.I0(GND_net), .I1(n1353), .I2(VCC_net), 
            .I3(n28515), .O(n1420)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_916_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_916_8 (.CI(n28515), .I0(n1353), .I1(VCC_net), .CO(n28516));
    SB_LUT4 rem_4_i1867_3_lut (.I0(n2746), .I1(n2813), .I2(n2768), .I3(GND_net), 
            .O(n2845));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1867_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_add_916_7_lut (.I0(GND_net), .I1(n1354), .I2(GND_net), 
            .I3(n28514), .O(n1421)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_916_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_i1875_3_lut (.I0(n2754), .I1(n2821), .I2(n2768), .I3(GND_net), 
            .O(n2853));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1875_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13014_3_lut (.I0(Ki[7]), .I1(\data_in_frame[5] [7]), .I2(n34066), 
            .I3(GND_net), .O(n17843));   // verilog/coms.v(126[12] 293[6])
    defparam i13014_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 rem_4_i1873_3_lut (.I0(n2752), .I1(n2819), .I2(n2768), .I3(GND_net), 
            .O(n2851));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1873_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1861_3_lut (.I0(n2740), .I1(n2807), .I2(n2768), .I3(GND_net), 
            .O(n2839));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1861_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1859_3_lut (.I0(n2738), .I1(n2805), .I2(n2768), .I3(GND_net), 
            .O(n2837));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1859_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_add_1519_19_lut (.I0(GND_net), .I1(n2241), .I2(VCC_net), 
            .I3(n28213), .O(n2308)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1519_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i13015_3_lut (.I0(Ki[8]), .I1(\data_in_frame[4] [0]), .I2(n34066), 
            .I3(GND_net), .O(n17844));   // verilog/coms.v(126[12] 293[6])
    defparam i13015_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 rem_4_i1860_3_lut (.I0(n2739), .I1(n2806), .I2(n2768), .I3(GND_net), 
            .O(n2838));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1860_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY rem_4_add_916_7 (.CI(n28514), .I0(n1354), .I1(GND_net), .CO(n28515));
    SB_LUT4 rem_4_add_916_6_lut (.I0(GND_net), .I1(n1355), .I2(GND_net), 
            .I3(n28513), .O(n1422)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_916_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1787_19_lut (.I0(n2641), .I1(n2641), .I2(n2669), 
            .I3(n27891), .O(n2740)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1787_19_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 rem_4_add_1653_16_lut (.I0(GND_net), .I1(n2444), .I2(VCC_net), 
            .I3(n28079), .O(n2511)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1653_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_916_6 (.CI(n28513), .I0(n1355), .I1(GND_net), .CO(n28514));
    SB_LUT4 rem_4_add_916_5_lut (.I0(GND_net), .I1(n1356), .I2(VCC_net), 
            .I3(n28512), .O(n1423)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_916_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1787_19 (.CI(n27891), .I0(n2641), .I1(n2669), .CO(n27892));
    SB_CARRY rem_4_add_916_5 (.CI(n28512), .I0(n1356), .I1(VCC_net), .CO(n28513));
    SB_LUT4 rem_4_add_916_4_lut (.I0(GND_net), .I1(n1357), .I2(VCC_net), 
            .I3(n28511), .O(n1424)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_916_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1653_16 (.CI(n28079), .I0(n2444), .I1(VCC_net), 
            .CO(n28080));
    SB_LUT4 rem_4_add_1653_15_lut (.I0(GND_net), .I1(n2445), .I2(VCC_net), 
            .I3(n28078), .O(n2512)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1653_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_916_4 (.CI(n28511), .I0(n1357), .I1(VCC_net), .CO(n28512));
    SB_LUT4 rem_4_add_916_3_lut (.I0(GND_net), .I1(n1358), .I2(GND_net), 
            .I3(n28510), .O(n1425)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_916_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_916_3 (.CI(n28510), .I0(n1358), .I1(GND_net), .CO(n28511));
    SB_LUT4 rem_4_i1858_3_lut (.I0(n2737), .I1(n2804), .I2(n2768), .I3(GND_net), 
            .O(n2836));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1858_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY rem_4_add_916_2 (.CI(VCC_net), .I0(n1458), .I1(VCC_net), 
            .CO(n28510));
    SB_LUT4 rem_4_add_983_13_lut (.I0(n1481), .I1(n1448), .I2(VCC_net), 
            .I3(n28509), .O(n1547)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_983_13_lut.LUT_INIT = 16'h8228;
    SB_LUT4 rem_4_add_983_12_lut (.I0(GND_net), .I1(n1449), .I2(VCC_net), 
            .I3(n28508), .O(n1516)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_983_12_lut.LUT_INIT = 16'hC33C;
    SB_DFF communication_counter_1522__i2 (.Q(communication_counter[2]), .C(LED_c), 
           .D(n163));   // verilog/TinyFPGA_B.v(52[28:51])
    SB_CARRY rem_4_add_983_12 (.CI(n28508), .I0(n1449), .I1(VCC_net), 
            .CO(n28509));
    SB_LUT4 rem_4_i1870_3_lut (.I0(n2749), .I1(n2816), .I2(n2768), .I3(GND_net), 
            .O(n2848));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1870_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_add_1787_18_lut (.I0(n2642), .I1(n2642), .I2(n2669), 
            .I3(n27890), .O(n2741)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1787_18_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY rem_4_add_1519_19 (.CI(n28213), .I0(n2241), .I1(VCC_net), 
            .CO(n28214));
    SB_CARRY rem_4_add_1653_15 (.CI(n28078), .I0(n2445), .I1(VCC_net), 
            .CO(n28079));
    SB_LUT4 rem_4_add_1653_14_lut (.I0(GND_net), .I1(n2446), .I2(VCC_net), 
            .I3(n28077), .O(n2513)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1653_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_i1877_3_lut (.I0(n2756), .I1(n2823), .I2(n2768), .I3(GND_net), 
            .O(n2855));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1877_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1876_3_lut (.I0(n2755), .I1(n2822), .I2(n2768), .I3(GND_net), 
            .O(n2854));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1876_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_add_983_11_lut (.I0(GND_net), .I1(n1450), .I2(VCC_net), 
            .I3(n28507), .O(n1517)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_983_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_i1866_3_lut (.I0(n2745), .I1(n2812), .I2(n2768), .I3(GND_net), 
            .O(n2844));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1866_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_3_lut_adj_1730 (.I0(n2756), .I1(n2757), .I2(n2758), .I3(GND_net), 
            .O(n33960));
    defparam i1_3_lut_adj_1730.LUT_INIT = 16'hfefe;
    SB_LUT4 i14_4_lut_adj_1731 (.I0(n2751), .I1(n2748), .I2(n2752), .I3(n2746), 
            .O(n34));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam i14_4_lut_adj_1731.LUT_INIT = 16'hfffe;
    SB_LUT4 i5_4_lut_adj_1732 (.I0(n2754), .I1(n2743), .I2(n33960), .I3(n2755), 
            .O(n25));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam i5_4_lut_adj_1732.LUT_INIT = 16'heccc;
    SB_LUT4 i12_4_lut_adj_1733 (.I0(n2739), .I1(n2741), .I2(n2740), .I3(n2742), 
            .O(n32));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam i12_4_lut_adj_1733.LUT_INIT = 16'hfffe;
    SB_LUT4 i11_4_lut_adj_1734 (.I0(n2736), .I1(n2737), .I2(n2735), .I3(n2738), 
            .O(n31));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam i11_4_lut_adj_1734.LUT_INIT = 16'hfffe;
    SB_LUT4 i15_4_lut_adj_1735 (.I0(n2750), .I1(n2745), .I2(n2753), .I3(n2749), 
            .O(n35));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam i15_4_lut_adj_1735.LUT_INIT = 16'hfffe;
    SB_LUT4 i17_4_lut_adj_1736 (.I0(n25), .I1(n34), .I2(n2747), .I3(n2744), 
            .O(n37));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam i17_4_lut_adj_1736.LUT_INIT = 16'hfffe;
    SB_LUT4 i19_4_lut (.I0(n37), .I1(n35), .I2(n31), .I3(n32), .O(n2768));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam i19_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 rem_4_mux_3_i9_3_lut (.I0(communication_counter[8]), .I1(n25_adj_4859), 
            .I2(communication_counter[31]), .I3(GND_net), .O(n2758));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_mux_3_i9_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_mux_3_i8_3_lut (.I0(communication_counter[7]), .I1(n26_adj_4858), 
            .I2(communication_counter[31]), .I3(GND_net), .O(n2759));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_mux_3_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1879_3_lut (.I0(n2758), .I1(n2825), .I2(n2768), .I3(GND_net), 
            .O(n2857));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1879_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1857_3_lut (.I0(n2736), .I1(n2803), .I2(n2768), .I3(GND_net), 
            .O(n2835));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1857_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY rem_4_add_983_11 (.CI(n28507), .I0(n1450), .I1(VCC_net), 
            .CO(n28508));
    SB_LUT4 i1_2_lut_adj_1737 (.I0(n2835), .I1(n2834), .I2(GND_net), .I3(GND_net), 
            .O(n22_adj_4776));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam i1_2_lut_adj_1737.LUT_INIT = 16'heeee;
    SB_LUT4 i1_3_lut_adj_1738 (.I0(n2856), .I1(n2857), .I2(n2759), .I3(GND_net), 
            .O(n34029));
    defparam i1_3_lut_adj_1738.LUT_INIT = 16'hfefe;
    SB_LUT4 i15_4_lut_adj_1739 (.I0(n2849), .I1(n2848), .I2(n2852), .I3(n2847), 
            .O(n36));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam i15_4_lut_adj_1739.LUT_INIT = 16'hfffe;
    SB_LUT4 i6_4_lut_adj_1740 (.I0(n2844), .I1(n2854), .I2(n34029), .I3(n2855), 
            .O(n27));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam i6_4_lut_adj_1740.LUT_INIT = 16'heaaa;
    SB_LUT4 i13_4_lut_adj_1741 (.I0(n2840), .I1(n2842), .I2(n2841), .I3(n2843), 
            .O(n34_adj_4771));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam i13_4_lut_adj_1741.LUT_INIT = 16'hfffe;
    SB_LUT4 i12_4_lut_adj_1742 (.I0(n2836), .I1(n2838), .I2(n2837), .I3(n2839), 
            .O(n33));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam i12_4_lut_adj_1742.LUT_INIT = 16'hfffe;
    SB_LUT4 i16_4_lut_adj_1743 (.I0(n2851), .I1(n2853), .I2(n2846), .I3(n22_adj_4776), 
            .O(n37_adj_4770));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam i16_4_lut_adj_1743.LUT_INIT = 16'hfffe;
    SB_LUT4 i18_4_lut_adj_1744 (.I0(n27), .I1(n36), .I2(n2850), .I3(n2845), 
            .O(n39));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam i18_4_lut_adj_1744.LUT_INIT = 16'hfffe;
    SB_LUT4 i20_4_lut (.I0(n39), .I1(n37_adj_4770), .I2(n33), .I3(n34_adj_4771), 
            .O(n2867));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam i20_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 rem_4_i1878_3_lut (.I0(n2757), .I1(n2824), .I2(n2768), .I3(GND_net), 
            .O(n2856));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1878_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1945_3_lut (.I0(n2856), .I1(n2923), .I2(n2867), .I3(GND_net), 
            .O(n2955));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1945_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_add_983_10_lut (.I0(GND_net), .I1(n1451), .I2(VCC_net), 
            .I3(n28506), .O(n1518)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_983_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_983_10 (.CI(n28506), .I0(n1451), .I1(VCC_net), 
            .CO(n28507));
    SB_LUT4 rem_4_add_983_9_lut (.I0(GND_net), .I1(n1452), .I2(VCC_net), 
            .I3(n28505), .O(n1519)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_983_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1653_14 (.CI(n28077), .I0(n2446), .I1(VCC_net), 
            .CO(n28078));
    SB_CARRY rem_4_add_1787_18 (.CI(n27890), .I0(n2642), .I1(n2669), .CO(n27891));
    SB_CARRY rem_4_add_983_9 (.CI(n28505), .I0(n1452), .I1(VCC_net), .CO(n28506));
    SB_LUT4 rem_4_add_983_8_lut (.I0(GND_net), .I1(n1453), .I2(VCC_net), 
            .I3(n28504), .O(n1520)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_983_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_983_8 (.CI(n28504), .I0(n1453), .I1(VCC_net), .CO(n28505));
    SB_LUT4 rem_4_add_983_7_lut (.I0(GND_net), .I1(n1454), .I2(GND_net), 
            .I3(n28503), .O(n1521)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_983_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1787_17_lut (.I0(n2643), .I1(n2643), .I2(n2669), 
            .I3(n27889), .O(n2742)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1787_17_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY rem_4_add_983_7 (.CI(n28503), .I0(n1454), .I1(GND_net), .CO(n28504));
    SB_LUT4 i14_4_lut_adj_1745 (.I0(n2249), .I1(n28_adj_4988), .I2(n24_adj_4990), 
            .I3(n16_adj_4993), .O(n2273));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam i14_4_lut_adj_1745.LUT_INIT = 16'hfffe;
    SB_LUT4 rem_4_add_983_6_lut (.I0(GND_net), .I1(n1455), .I2(GND_net), 
            .I3(n28502), .O(n1522)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_983_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_983_6 (.CI(n28502), .I0(n1455), .I1(GND_net), .CO(n28503));
    SB_LUT4 rem_4_add_983_5_lut (.I0(GND_net), .I1(n1456), .I2(VCC_net), 
            .I3(n28501), .O(n1523)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_983_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_983_5 (.CI(n28501), .I0(n1456), .I1(VCC_net), .CO(n28502));
    SB_CARRY rem_4_add_1787_17 (.CI(n27889), .I0(n2643), .I1(n2669), .CO(n27890));
    SB_LUT4 rem_4_add_1653_13_lut (.I0(GND_net), .I1(n2447), .I2(VCC_net), 
            .I3(n28076), .O(n2514)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1653_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1653_13 (.CI(n28076), .I0(n2447), .I1(VCC_net), 
            .CO(n28077));
    SB_LUT4 rem_4_i1944_3_lut (.I0(n2855), .I1(n2922), .I2(n2867), .I3(GND_net), 
            .O(n2954));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1944_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i31088_3_lut (.I0(n2848), .I1(n2915), .I2(n2867), .I3(GND_net), 
            .O(n2947));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam i31088_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_3_lut_adj_1746 (.I0(n2956), .I1(n2957), .I2(n2958_adj_4882), 
            .I3(GND_net), .O(n33975));
    defparam i1_3_lut_adj_1746.LUT_INIT = 16'hfefe;
    SB_LUT4 rem_4_add_983_4_lut (.I0(GND_net), .I1(n1457), .I2(VCC_net), 
            .I3(n28500), .O(n1524)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_983_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i6_4_lut_adj_1747 (.I0(n2947), .I1(n2954), .I2(n33975), .I3(n2955), 
            .O(n28));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam i6_4_lut_adj_1747.LUT_INIT = 16'heaaa;
    SB_CARRY rem_4_add_983_4 (.CI(n28500), .I0(n1457), .I1(VCC_net), .CO(n28501));
    SB_LUT4 rem_4_add_1653_12_lut (.I0(GND_net), .I1(n2448), .I2(VCC_net), 
            .I3(n28075), .O(n2515)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1653_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i13_4_lut_adj_1748 (.I0(n2937), .I1(n2939), .I2(n2938), .I3(n2940), 
            .O(n35_adj_4779));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam i13_4_lut_adj_1748.LUT_INIT = 16'hfffe;
    SB_LUT4 i13437_3_lut (.I0(\half_duty[0] [2]), .I1(half_duty_new[2]), 
            .I2(n1466), .I3(GND_net), .O(n18266));   // vhdl/pwm.vhd(59[5] 95[12])
    defparam i13437_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF communication_counter_1522__i3 (.Q(communication_counter[3]), .C(LED_c), 
           .D(n162));   // verilog/TinyFPGA_B.v(52[28:51])
    SB_DFF communication_counter_1522__i4 (.Q(communication_counter[4]), .C(LED_c), 
           .D(n161));   // verilog/TinyFPGA_B.v(52[28:51])
    SB_DFF communication_counter_1522__i5 (.Q(communication_counter[5]), .C(LED_c), 
           .D(n160));   // verilog/TinyFPGA_B.v(52[28:51])
    SB_DFF communication_counter_1522__i6 (.Q(communication_counter[6]), .C(LED_c), 
           .D(n159));   // verilog/TinyFPGA_B.v(52[28:51])
    SB_DFF communication_counter_1522__i7 (.Q(communication_counter[7]), .C(LED_c), 
           .D(n158));   // verilog/TinyFPGA_B.v(52[28:51])
    SB_DFF communication_counter_1522__i8 (.Q(communication_counter[8]), .C(LED_c), 
           .D(n157));   // verilog/TinyFPGA_B.v(52[28:51])
    SB_DFF communication_counter_1522__i9 (.Q(communication_counter[9]), .C(LED_c), 
           .D(n156));   // verilog/TinyFPGA_B.v(52[28:51])
    SB_DFF communication_counter_1522__i10 (.Q(communication_counter[10]), 
           .C(LED_c), .D(n155));   // verilog/TinyFPGA_B.v(52[28:51])
    SB_DFF communication_counter_1522__i11 (.Q(communication_counter[11]), 
           .C(LED_c), .D(n154));   // verilog/TinyFPGA_B.v(52[28:51])
    SB_DFF communication_counter_1522__i12 (.Q(communication_counter[12]), 
           .C(LED_c), .D(n153));   // verilog/TinyFPGA_B.v(52[28:51])
    SB_DFF communication_counter_1522__i13 (.Q(communication_counter[13]), 
           .C(LED_c), .D(n152));   // verilog/TinyFPGA_B.v(52[28:51])
    SB_DFF communication_counter_1522__i14 (.Q(communication_counter[14]), 
           .C(LED_c), .D(n151));   // verilog/TinyFPGA_B.v(52[28:51])
    SB_DFF communication_counter_1522__i15 (.Q(communication_counter[15]), 
           .C(LED_c), .D(n150));   // verilog/TinyFPGA_B.v(52[28:51])
    SB_DFF communication_counter_1522__i16 (.Q(communication_counter[16]), 
           .C(LED_c), .D(n149));   // verilog/TinyFPGA_B.v(52[28:51])
    SB_DFF communication_counter_1522__i17 (.Q(communication_counter[17]), 
           .C(LED_c), .D(n148));   // verilog/TinyFPGA_B.v(52[28:51])
    SB_DFF communication_counter_1522__i18 (.Q(communication_counter[18]), 
           .C(LED_c), .D(n147));   // verilog/TinyFPGA_B.v(52[28:51])
    SB_DFF communication_counter_1522__i19 (.Q(communication_counter[19]), 
           .C(LED_c), .D(n146));   // verilog/TinyFPGA_B.v(52[28:51])
    SB_DFF communication_counter_1522__i20 (.Q(communication_counter[20]), 
           .C(LED_c), .D(n145));   // verilog/TinyFPGA_B.v(52[28:51])
    SB_DFF communication_counter_1522__i21 (.Q(communication_counter[21]), 
           .C(LED_c), .D(n144));   // verilog/TinyFPGA_B.v(52[28:51])
    SB_DFF communication_counter_1522__i22 (.Q(communication_counter[22]), 
           .C(LED_c), .D(n143));   // verilog/TinyFPGA_B.v(52[28:51])
    SB_DFF communication_counter_1522__i23 (.Q(communication_counter[23]), 
           .C(LED_c), .D(n142));   // verilog/TinyFPGA_B.v(52[28:51])
    SB_DFF communication_counter_1522__i24 (.Q(communication_counter[24]), 
           .C(LED_c), .D(n141));   // verilog/TinyFPGA_B.v(52[28:51])
    SB_DFF communication_counter_1522__i25 (.Q(communication_counter[25]), 
           .C(LED_c), .D(n140));   // verilog/TinyFPGA_B.v(52[28:51])
    SB_DFF communication_counter_1522__i26 (.Q(communication_counter[26]), 
           .C(LED_c), .D(n139));   // verilog/TinyFPGA_B.v(52[28:51])
    SB_DFF communication_counter_1522__i27 (.Q(communication_counter[27]), 
           .C(LED_c), .D(n138));   // verilog/TinyFPGA_B.v(52[28:51])
    SB_DFF communication_counter_1522__i28 (.Q(communication_counter[28]), 
           .C(LED_c), .D(n137));   // verilog/TinyFPGA_B.v(52[28:51])
    SB_DFF communication_counter_1522__i29 (.Q(communication_counter[29]), 
           .C(LED_c), .D(n136));   // verilog/TinyFPGA_B.v(52[28:51])
    SB_DFF communication_counter_1522__i30 (.Q(communication_counter[30]), 
           .C(LED_c), .D(n135));   // verilog/TinyFPGA_B.v(52[28:51])
    SB_DFF communication_counter_1522__i31 (.Q(communication_counter[31]), 
           .C(LED_c), .D(n134));   // verilog/TinyFPGA_B.v(52[28:51])
    SB_LUT4 rem_4_add_983_3_lut (.I0(GND_net), .I1(n1458), .I2(GND_net), 
            .I3(n28499), .O(n1525)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_983_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_983_3 (.CI(n28499), .I0(n1458), .I1(GND_net), .CO(n28500));
    SB_LUT4 rem_4_add_1787_16_lut (.I0(n2644), .I1(n2644), .I2(n2669), 
            .I3(n27888), .O(n2743)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1787_16_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY rem_4_add_1653_12 (.CI(n28075), .I0(n2448), .I1(VCC_net), 
            .CO(n28076));
    SB_CARRY rem_4_add_983_2 (.CI(VCC_net), .I0(n1558), .I1(VCC_net), 
            .CO(n28499));
    SB_LUT4 rem_4_add_1519_18_lut (.I0(GND_net), .I1(n2242), .I2(VCC_net), 
            .I3(n28212), .O(n2309)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1519_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i12_4_lut_adj_1749 (.I0(n2934), .I1(n2935), .I2(n2933), .I3(n2936), 
            .O(n34_adj_4780));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam i12_4_lut_adj_1749.LUT_INIT = 16'hfffe;
    SB_LUT4 i18_4_lut_adj_1750 (.I0(n35_adj_4779), .I1(n2941), .I2(n28), 
            .I3(n2942), .O(n40));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam i18_4_lut_adj_1750.LUT_INIT = 16'hfffe;
    SB_LUT4 i16_4_lut_adj_1751 (.I0(n2949), .I1(n2952), .I2(n2950), .I3(n2945), 
            .O(n38));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam i16_4_lut_adj_1751.LUT_INIT = 16'hfffe;
    SB_LUT4 i17_3_lut (.I0(n2953), .I1(n34_adj_4780), .I2(n2948), .I3(GND_net), 
            .O(n39_adj_4777));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam i17_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i15_4_lut_adj_1752 (.I0(n2946), .I1(n2943), .I2(n2951), .I3(n2944), 
            .O(n37_adj_4778));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam i15_4_lut_adj_1752.LUT_INIT = 16'hfffe;
    SB_LUT4 i21_4_lut (.I0(n37_adj_4778), .I1(n39_adj_4777), .I2(n38), 
            .I3(n40), .O(n2966));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam i21_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 rem_4_mux_3_i7_3_lut (.I0(communication_counter[6]), .I1(n27_adj_4857), 
            .I2(communication_counter[31]), .I3(GND_net), .O(n2958_adj_4882));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_mux_3_i7_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_mux_3_i6_3_lut (.I0(communication_counter[5]), .I1(n28_adj_4856), 
            .I2(communication_counter[31]), .I3(GND_net), .O(n3058));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_mux_3_i6_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i2015_3_lut (.I0(n2958_adj_4882), .I1(n3025), .I2(n2966), 
            .I3(GND_net), .O(n3057));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i2015_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i2014_3_lut (.I0(n2957), .I1(n3024), .I2(n2966), .I3(GND_net), 
            .O(n3056));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i2014_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_3_lut_adj_1753 (.I0(n3056), .I1(n3057), .I2(n3058), .I3(GND_net), 
            .O(n34037));
    defparam i1_3_lut_adj_1753.LUT_INIT = 16'hfefe;
    SB_LUT4 i7_4_lut_adj_1754 (.I0(n3054), .I1(n3044), .I2(n34037), .I3(n3055), 
            .O(n30_adj_4791));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam i7_4_lut_adj_1754.LUT_INIT = 16'heccc;
    SB_LUT4 i14_4_lut_adj_1755 (.I0(n3038), .I1(n3040), .I2(n3039), .I3(n3041), 
            .O(n37_adj_4789));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam i14_4_lut_adj_1755.LUT_INIT = 16'hfffe;
    SB_LUT4 i13_4_lut_adj_1756 (.I0(n3034), .I1(n3036), .I2(n3035), .I3(n3037), 
            .O(n36_adj_4790));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam i13_4_lut_adj_1756.LUT_INIT = 16'hfffe;
    SB_CARRY rem_4_add_1519_18 (.CI(n28212), .I0(n2242), .I1(VCC_net), 
            .CO(n28213));
    SB_LUT4 i19_4_lut_adj_1757 (.I0(n37_adj_4789), .I1(n3042), .I2(n30_adj_4791), 
            .I3(n3043), .O(n42));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam i19_4_lut_adj_1757.LUT_INIT = 16'hfffe;
    SB_LUT4 i17_4_lut_adj_1758 (.I0(n3050), .I1(n3047), .I2(n3053), .I3(n3046), 
            .O(n40_adj_4787));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam i17_4_lut_adj_1758.LUT_INIT = 16'hfffe;
    SB_LUT4 i18_4_lut_adj_1759 (.I0(n3048), .I1(n36_adj_4790), .I2(n3033), 
            .I3(n3032), .O(n41));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam i18_4_lut_adj_1759.LUT_INIT = 16'hfffe;
    SB_LUT4 i16_4_lut_adj_1760 (.I0(n3051), .I1(n3045), .I2(n3052), .I3(n3049), 
            .O(n39_adj_4788));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam i16_4_lut_adj_1760.LUT_INIT = 16'hfffe;
    SB_LUT4 i22_4_lut (.I0(n39_adj_4788), .I1(n41), .I2(n40_adj_4787), 
            .I3(n42), .O(n3065));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam i22_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 rem_4_add_1653_11_lut (.I0(GND_net), .I1(n2449), .I2(VCC_net), 
            .I3(n28074), .O(n2516)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1653_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_i2009_3_lut (.I0(n2952), .I1(n3019), .I2(n2966), .I3(GND_net), 
            .O(n3051));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i2009_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i2076_3_lut (.I0(n3051), .I1(n3118), .I2(n3065), .I3(GND_net), 
            .O(n3150));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i2076_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i2077_3_lut (.I0(n3052), .I1(n3119), .I2(n3065), .I3(GND_net), 
            .O(n3151));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i2077_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_add_1519_17_lut (.I0(GND_net), .I1(n2243), .I2(VCC_net), 
            .I3(n28211), .O(n2310)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1519_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1787_16 (.CI(n27888), .I0(n2644), .I1(n2669), .CO(n27889));
    SB_LUT4 rem_4_add_1787_15_lut (.I0(n2645), .I1(n2645), .I2(n2669), 
            .I3(n27887), .O(n2744)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1787_15_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY rem_4_add_1519_17 (.CI(n28211), .I0(n2243), .I1(VCC_net), 
            .CO(n28212));
    SB_LUT4 i13441_3_lut (.I0(\half_duty[0] [6]), .I1(half_duty_new[6]), 
            .I2(n1466), .I3(GND_net), .O(n18270));   // vhdl/pwm.vhd(59[5] 95[12])
    defparam i13441_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_add_1519_16_lut (.I0(GND_net), .I1(n2244), .I2(VCC_net), 
            .I3(n28210), .O(n2311)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1519_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_i2068_3_lut (.I0(n3043), .I1(n3110), .I2(n3065), .I3(GND_net), 
            .O(n3142));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i2068_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY rem_4_add_1519_16 (.CI(n28210), .I0(n2244), .I1(VCC_net), 
            .CO(n28211));
    SB_CARRY rem_4_add_1653_11 (.CI(n28074), .I0(n2449), .I1(VCC_net), 
            .CO(n28075));
    SB_LUT4 rem_4_i2070_3_lut (.I0(n3045), .I1(n3112), .I2(n3065), .I3(GND_net), 
            .O(n3144));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i2070_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_mux_3_i5_3_lut (.I0(communication_counter[4]), .I1(n29_adj_4855), 
            .I2(communication_counter[31]), .I3(GND_net), .O(n3158));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_mux_3_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_add_1653_10_lut (.I0(GND_net), .I1(n2450), .I2(VCC_net), 
            .I3(n28073), .O(n2517)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1653_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_i2083_3_lut (.I0(n3058), .I1(n3125), .I2(n3065), .I3(GND_net), 
            .O(n3157));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i2083_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY rem_4_add_1787_15 (.CI(n27887), .I0(n2645), .I1(n2669), .CO(n27888));
    SB_LUT4 rem_4_add_1519_15_lut (.I0(GND_net), .I1(n2245), .I2(VCC_net), 
            .I3(n28209), .O(n2312)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1519_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_3_lut_adj_1761 (.I0(n3156), .I1(n3157), .I2(n3158), .I3(GND_net), 
            .O(n33985));
    defparam i1_3_lut_adj_1761.LUT_INIT = 16'hfefe;
    SB_CARRY rem_4_add_1519_15 (.CI(n28209), .I0(n2245), .I1(VCC_net), 
            .CO(n28210));
    SB_CARRY rem_4_add_1653_10 (.CI(n28073), .I0(n2450), .I1(VCC_net), 
            .CO(n28074));
    SB_LUT4 i6_4_lut_adj_1762 (.I0(n3154), .I1(n3141), .I2(n33985), .I3(n3155), 
            .O(n30_adj_4799));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam i6_4_lut_adj_1762.LUT_INIT = 16'heccc;
    SB_LUT4 i16_4_lut_adj_1763 (.I0(n3144), .I1(n3142), .I2(n3151), .I3(n3150), 
            .O(n40_adj_4794));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam i16_4_lut_adj_1763.LUT_INIT = 16'hfffe;
    SB_LUT4 rem_4_add_1519_14_lut (.I0(GND_net), .I1(n2246), .I2(VCC_net), 
            .I3(n28208), .O(n2313)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1519_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i2_2_lut (.I0(n3133), .I1(n3134), .I2(GND_net), .I3(GND_net), 
            .O(n26));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam i2_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 rem_4_add_1787_14_lut (.I0(n2646), .I1(n2646), .I2(n2669), 
            .I3(n27886), .O(n2745)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1787_14_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY rem_4_add_1519_14 (.CI(n28208), .I0(n2246), .I1(VCC_net), 
            .CO(n28209));
    SB_LUT4 rem_4_add_1519_13_lut (.I0(GND_net), .I1(n2247), .I2(VCC_net), 
            .I3(n28207), .O(n2314)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1519_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i14_4_lut_adj_1764 (.I0(n3135), .I1(n3137), .I2(n3136), .I3(n3138), 
            .O(n38_adj_4797));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam i14_4_lut_adj_1764.LUT_INIT = 16'hfffe;
    SB_LUT4 i2_3_lut_4_lut (.I0(n24786), .I1(n16158), .I2(n5_adj_4786), 
            .I3(n2958), .O(n32849));   // verilog/coms.v(126[12] 293[6])
    defparam i2_3_lut_4_lut.LUT_INIT = 16'hfff2;
    SB_CARRY rem_4_add_1787_12 (.CI(n27884), .I0(n2648), .I1(n2669), .CO(n27885));
    SB_LUT4 i20_4_lut_adj_1765 (.I0(n3139), .I1(n40_adj_4794), .I2(n30_adj_4799), 
            .I3(n3140), .O(n44));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam i20_4_lut_adj_1765.LUT_INIT = 16'hfffe;
    SB_LUT4 i18_4_lut_adj_1766 (.I0(n3152), .I1(n3149), .I2(n3147), .I3(n3148), 
            .O(n42_adj_4792));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam i18_4_lut_adj_1766.LUT_INIT = 16'hfffe;
    SB_CARRY rem_4_add_1519_13 (.CI(n28207), .I0(n2247), .I1(VCC_net), 
            .CO(n28208));
    SB_LUT4 i19_4_lut_adj_1767 (.I0(n3132), .I1(n38_adj_4797), .I2(n26), 
            .I3(n3131), .O(n43));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam i19_4_lut_adj_1767.LUT_INIT = 16'hfffe;
    SB_LUT4 rem_4_add_1653_9_lut (.I0(GND_net), .I1(n2451), .I2(VCC_net), 
            .I3(n28072), .O(n2518)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1653_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i17_4_lut_adj_1768 (.I0(n3145), .I1(n3143), .I2(n3146), .I3(n3153), 
            .O(n41_adj_4793));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam i17_4_lut_adj_1768.LUT_INIT = 16'hfffe;
    SB_CARRY rem_4_add_1653_9 (.CI(n28072), .I0(n2451), .I1(VCC_net), 
            .CO(n28073));
    SB_LUT4 i23_4_lut (.I0(n41_adj_4793), .I1(n43), .I2(n42_adj_4792), 
            .I3(n44), .O(n3164_adj_4884));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam i23_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 rem_4_i2082_3_lut (.I0(n3057), .I1(n3124), .I2(n3065), .I3(GND_net), 
            .O(n3156));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i2082_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_add_1653_8_lut (.I0(GND_net), .I1(n2452), .I2(VCC_net), 
            .I3(n28071), .O(n2519)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1653_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1519_12_lut (.I0(GND_net), .I1(n2248), .I2(VCC_net), 
            .I3(n28206), .O(n2315)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1519_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_i2149_3_lut (.I0(n3156), .I1(n3223_adj_4899), .I2(n3164_adj_4884), 
            .I3(GND_net), .O(n3255));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i2149_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY rem_4_add_1653_8 (.CI(n28071), .I0(n2452), .I1(VCC_net), 
            .CO(n28072));
    SB_LUT4 rem_4_i2136_3_lut (.I0(n3143), .I1(n3210_adj_4886), .I2(n3164_adj_4884), 
            .I3(GND_net), .O(n3242));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i2136_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_3_lut_adj_1769 (.I0(n3256), .I1(n3257), .I2(n3258), .I3(GND_net), 
            .O(n34042));
    defparam i1_3_lut_adj_1769.LUT_INIT = 16'hfefe;
    SB_LUT4 rem_4_add_1787_13_lut (.I0(n2647), .I1(n2647), .I2(n2669), 
            .I3(n27885), .O(n2746)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1787_13_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i7_4_lut_adj_1770 (.I0(n3242), .I1(n3254), .I2(n34042), .I3(n3255), 
            .O(n32_adj_4826));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam i7_4_lut_adj_1770.LUT_INIT = 16'heaaa;
    SB_LUT4 i17_4_lut_adj_1771 (.I0(n3243), .I1(n3248), .I2(n3246), .I3(n3252), 
            .O(n42_adj_4811));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam i17_4_lut_adj_1771.LUT_INIT = 16'hfffe;
    SB_CARRY rem_4_add_1519_12 (.CI(n28206), .I0(n2248), .I1(VCC_net), 
            .CO(n28207));
    SB_LUT4 i1_2_lut_4_lut (.I0(tx_active), .I1(r_SM_Main_2__N_3458[0]), 
            .I2(tx_transmit_N_3355), .I3(n16157), .O(n5_adj_4786));   // verilog/coms.v(126[12] 293[6])
    defparam i1_2_lut_4_lut.LUT_INIT = 16'h00fe;
    SB_LUT4 rem_4_add_1519_11_lut (.I0(GND_net), .I1(n2249), .I2(VCC_net), 
            .I3(n28205), .O(n2316)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1519_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1050_14_lut (.I0(n1580), .I1(n1547), .I2(VCC_net), 
            .I3(n28434), .O(n1646)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1050_14_lut.LUT_INIT = 16'h8228;
    SB_LUT4 rem_4_add_1050_13_lut (.I0(GND_net), .I1(n1548), .I2(VCC_net), 
            .I3(n28433), .O(n1615)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1050_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i13_3_lut (.I0(n3245), .I1(n3231_adj_4903), .I2(n3230_adj_4902), 
            .I3(GND_net), .O(n38_adj_4819));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam i13_3_lut.LUT_INIT = 16'hfefe;
    SB_CARRY rem_4_add_1050_13 (.CI(n28433), .I0(n1548), .I1(VCC_net), 
            .CO(n28434));
    SB_LUT4 i18_4_lut_adj_1772 (.I0(n3249), .I1(n3253), .I2(n3250), .I3(n3244), 
            .O(n43_adj_4810));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam i18_4_lut_adj_1772.LUT_INIT = 16'hfffe;
    SB_LUT4 rem_4_add_1050_12_lut (.I0(GND_net), .I1(n1549), .I2(VCC_net), 
            .I3(n28432), .O(n1616)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1050_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1050_12 (.CI(n28432), .I0(n1549), .I1(VCC_net), 
            .CO(n28433));
    SB_LUT4 rem_4_add_1653_7_lut (.I0(GND_net), .I1(n2453), .I2(VCC_net), 
            .I3(n28070), .O(n2520)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1653_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i15_4_lut_adj_1773 (.I0(n3236), .I1(n3238), .I2(n3237), .I3(n3239), 
            .O(n40_adj_4813));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam i15_4_lut_adj_1773.LUT_INIT = 16'hfffe;
    SB_LUT4 rem_4_add_1050_11_lut (.I0(GND_net), .I1(n1550), .I2(VCC_net), 
            .I3(n28431), .O(n1617)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1050_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1050_11 (.CI(n28431), .I0(n1550), .I1(VCC_net), 
            .CO(n28432));
    SB_LUT4 rem_4_add_1050_10_lut (.I0(GND_net), .I1(n1551), .I2(VCC_net), 
            .I3(n28430), .O(n1618)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1050_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1050_10 (.CI(n28430), .I0(n1551), .I1(VCC_net), 
            .CO(n28431));
    SB_LUT4 rem_4_add_1050_9_lut (.I0(GND_net), .I1(n1552), .I2(VCC_net), 
            .I3(n28429), .O(n1619)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1050_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i21_4_lut_adj_1774 (.I0(n3240), .I1(n42_adj_4811), .I2(n32_adj_4826), 
            .I3(n3241), .O(n46));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam i21_4_lut_adj_1774.LUT_INIT = 16'hfffe;
    SB_LUT4 i14_4_lut_adj_1775 (.I0(n3232_adj_4904), .I1(n3234), .I2(n3233), 
            .I3(n3235), .O(n39_adj_4814));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam i14_4_lut_adj_1775.LUT_INIT = 16'hfffe;
    SB_CARRY rem_4_add_1050_9 (.CI(n28429), .I0(n1552), .I1(VCC_net), 
            .CO(n28430));
    SB_LUT4 i22_4_lut_adj_1776 (.I0(n43_adj_4810), .I1(n3247), .I2(n38_adj_4819), 
            .I3(n3251), .O(n47));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam i22_4_lut_adj_1776.LUT_INIT = 16'hfffe;
    SB_LUT4 i24_4_lut (.I0(n47), .I1(n39_adj_4814), .I2(n46), .I3(n40_adj_4813), 
            .O(n3263));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam i24_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 rem_4_i2148_3_lut (.I0(n3155), .I1(n3222_adj_4898), .I2(n3164_adj_4884), 
            .I3(GND_net), .O(n3254));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i2148_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i2215_3_lut (.I0(n3254), .I1(n3321), .I2(n3263), .I3(GND_net), 
            .O(n3353));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i2215_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_add_1050_8_lut (.I0(GND_net), .I1(n1553), .I2(VCC_net), 
            .I3(n28428), .O(n1620)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1050_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1050_8 (.CI(n28428), .I0(n1553), .I1(VCC_net), 
            .CO(n28429));
    SB_LUT4 rem_4_add_1050_7_lut (.I0(GND_net), .I1(n1554), .I2(GND_net), 
            .I3(n28427), .O(n1621)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1050_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1050_7 (.CI(n28427), .I0(n1554), .I1(GND_net), 
            .CO(n28428));
    SB_LUT4 rem_4_add_1050_6_lut (.I0(GND_net), .I1(n1555), .I2(GND_net), 
            .I3(n28426), .O(n1622)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1050_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1050_6 (.CI(n28426), .I0(n1555), .I1(GND_net), 
            .CO(n28427));
    SB_LUT4 rem_4_add_1050_5_lut (.I0(GND_net), .I1(n1556), .I2(VCC_net), 
            .I3(n28425), .O(n1623)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1050_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1050_5 (.CI(n28425), .I0(n1556), .I1(VCC_net), 
            .CO(n28426));
    SB_LUT4 rem_4_add_1050_4_lut (.I0(GND_net), .I1(n1557), .I2(VCC_net), 
            .I3(n28424), .O(n1624)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1050_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i13190_3_lut (.I0(\data_in_frame[1] [1]), .I1(rx_data[1]), .I2(n32962), 
            .I3(GND_net), .O(n18019));   // verilog/coms.v(126[12] 293[6])
    defparam i13190_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY rem_4_add_1050_4 (.CI(n28424), .I0(n1557), .I1(VCC_net), 
            .CO(n28425));
    SB_LUT4 rem_4_add_1050_3_lut (.I0(GND_net), .I1(n1558), .I2(GND_net), 
            .I3(n28423), .O(n1625)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1050_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1050_3 (.CI(n28423), .I0(n1558), .I1(GND_net), 
            .CO(n28424));
    SB_CARRY rem_4_add_1050_2 (.CI(VCC_net), .I0(n1658), .I1(VCC_net), 
            .CO(n28423));
    SB_LUT4 communication_counter_1522_add_4_33_lut (.I0(GND_net), .I1(GND_net), 
            .I2(communication_counter[31]), .I3(n28422), .O(n134)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_1522_add_4_33_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 communication_counter_1522_add_4_32_lut (.I0(GND_net), .I1(GND_net), 
            .I2(communication_counter[30]), .I3(n28421), .O(n135)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_1522_add_4_32_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_1522_add_4_32 (.CI(n28421), .I0(GND_net), 
            .I1(communication_counter[30]), .CO(n28422));
    SB_LUT4 communication_counter_1522_add_4_31_lut (.I0(GND_net), .I1(GND_net), 
            .I2(communication_counter[29]), .I3(n28420), .O(n136)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_1522_add_4_31_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_1522_add_4_31 (.CI(n28420), .I0(GND_net), 
            .I1(communication_counter[29]), .CO(n28421));
    SB_LUT4 communication_counter_1522_add_4_30_lut (.I0(GND_net), .I1(GND_net), 
            .I2(communication_counter[28]), .I3(n28419), .O(n137)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_1522_add_4_30_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_1522_add_4_30 (.CI(n28419), .I0(GND_net), 
            .I1(communication_counter[28]), .CO(n28420));
    SB_LUT4 communication_counter_1522_add_4_29_lut (.I0(GND_net), .I1(GND_net), 
            .I2(communication_counter[27]), .I3(n28418), .O(n138)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_1522_add_4_29_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_1522_add_4_29 (.CI(n28418), .I0(GND_net), 
            .I1(communication_counter[27]), .CO(n28419));
    SB_LUT4 communication_counter_1522_add_4_28_lut (.I0(GND_net), .I1(GND_net), 
            .I2(communication_counter[26]), .I3(n28417), .O(n139)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_1522_add_4_28_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_1522_add_4_28 (.CI(n28417), .I0(GND_net), 
            .I1(communication_counter[26]), .CO(n28418));
    SB_LUT4 communication_counter_1522_add_4_27_lut (.I0(GND_net), .I1(GND_net), 
            .I2(communication_counter[25]), .I3(n28416), .O(n140)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_1522_add_4_27_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_1522_add_4_27 (.CI(n28416), .I0(GND_net), 
            .I1(communication_counter[25]), .CO(n28417));
    SB_LUT4 communication_counter_1522_add_4_26_lut (.I0(GND_net), .I1(GND_net), 
            .I2(communication_counter[24]), .I3(n28415), .O(n141)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_1522_add_4_26_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_1522_add_4_26 (.CI(n28415), .I0(GND_net), 
            .I1(communication_counter[24]), .CO(n28416));
    SB_LUT4 communication_counter_1522_add_4_25_lut (.I0(GND_net), .I1(GND_net), 
            .I2(communication_counter[23]), .I3(n28414), .O(n142)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_1522_add_4_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_1522_add_4_25 (.CI(n28414), .I0(GND_net), 
            .I1(communication_counter[23]), .CO(n28415));
    SB_LUT4 PIN_13_I_0_1_lut (.I0(PIN_13_c), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(PIN_13_N_105));   // verilog/TinyFPGA_B.v(189[10:15])
    defparam PIN_13_I_0_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 communication_counter_1522_add_4_24_lut (.I0(GND_net), .I1(GND_net), 
            .I2(communication_counter[22]), .I3(n28413), .O(n143)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_1522_add_4_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_1522_add_4_24 (.CI(n28413), .I0(GND_net), 
            .I1(communication_counter[22]), .CO(n28414));
    SB_LUT4 communication_counter_1522_add_4_23_lut (.I0(GND_net), .I1(GND_net), 
            .I2(communication_counter[21]), .I3(n28412), .O(n144)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_1522_add_4_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_1522_add_4_23 (.CI(n28412), .I0(GND_net), 
            .I1(communication_counter[21]), .CO(n28413));
    SB_LUT4 communication_counter_1522_add_4_22_lut (.I0(GND_net), .I1(GND_net), 
            .I2(communication_counter[20]), .I3(n28411), .O(n145)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_1522_add_4_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_1522_add_4_22 (.CI(n28411), .I0(GND_net), 
            .I1(communication_counter[20]), .CO(n28412));
    SB_LUT4 communication_counter_1522_add_4_21_lut (.I0(GND_net), .I1(GND_net), 
            .I2(communication_counter[19]), .I3(n28410), .O(n146)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_1522_add_4_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_1522_add_4_21 (.CI(n28410), .I0(GND_net), 
            .I1(communication_counter[19]), .CO(n28411));
    SB_LUT4 communication_counter_1522_add_4_20_lut (.I0(GND_net), .I1(GND_net), 
            .I2(communication_counter[18]), .I3(n28409), .O(n147)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_1522_add_4_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_1522_add_4_20 (.CI(n28409), .I0(GND_net), 
            .I1(communication_counter[18]), .CO(n28410));
    SB_LUT4 communication_counter_1522_add_4_19_lut (.I0(GND_net), .I1(GND_net), 
            .I2(communication_counter[17]), .I3(n28408), .O(n148)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_1522_add_4_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_1522_add_4_19 (.CI(n28408), .I0(GND_net), 
            .I1(communication_counter[17]), .CO(n28409));
    SB_LUT4 communication_counter_1522_add_4_18_lut (.I0(GND_net), .I1(GND_net), 
            .I2(communication_counter[16]), .I3(n28407), .O(n149)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_1522_add_4_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_1522_add_4_18 (.CI(n28407), .I0(GND_net), 
            .I1(communication_counter[16]), .CO(n28408));
    SB_LUT4 communication_counter_1522_add_4_17_lut (.I0(GND_net), .I1(GND_net), 
            .I2(communication_counter[15]), .I3(n28406), .O(n150)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_1522_add_4_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_1522_add_4_17 (.CI(n28406), .I0(GND_net), 
            .I1(communication_counter[15]), .CO(n28407));
    SB_LUT4 communication_counter_1522_add_4_16_lut (.I0(GND_net), .I1(GND_net), 
            .I2(communication_counter[14]), .I3(n28405), .O(n151)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_1522_add_4_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_1522_add_4_16 (.CI(n28405), .I0(GND_net), 
            .I1(communication_counter[14]), .CO(n28406));
    SB_LUT4 communication_counter_1522_add_4_15_lut (.I0(GND_net), .I1(GND_net), 
            .I2(communication_counter[13]), .I3(n28404), .O(n152)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_1522_add_4_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_1522_add_4_15 (.CI(n28404), .I0(GND_net), 
            .I1(communication_counter[13]), .CO(n28405));
    SB_LUT4 communication_counter_1522_add_4_14_lut (.I0(GND_net), .I1(GND_net), 
            .I2(communication_counter[12]), .I3(n28403), .O(n153)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_1522_add_4_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_1522_add_4_14 (.CI(n28403), .I0(GND_net), 
            .I1(communication_counter[12]), .CO(n28404));
    SB_LUT4 communication_counter_1522_add_4_13_lut (.I0(GND_net), .I1(GND_net), 
            .I2(communication_counter[11]), .I3(n28402), .O(n154)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_1522_add_4_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1519_11 (.CI(n28205), .I0(n2249), .I1(VCC_net), 
            .CO(n28206));
    SB_CARRY communication_counter_1522_add_4_13 (.CI(n28402), .I0(GND_net), 
            .I1(communication_counter[11]), .CO(n28403));
    SB_LUT4 communication_counter_1522_add_4_12_lut (.I0(GND_net), .I1(GND_net), 
            .I2(communication_counter[10]), .I3(n28401), .O(n155)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_1522_add_4_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_1522_add_4_12 (.CI(n28401), .I0(GND_net), 
            .I1(communication_counter[10]), .CO(n28402));
    SB_CARRY rem_4_add_1787_13 (.CI(n27885), .I0(n2647), .I1(n2669), .CO(n27886));
    SB_LUT4 communication_counter_1522_add_4_11_lut (.I0(GND_net), .I1(GND_net), 
            .I2(communication_counter[9]), .I3(n28400), .O(n156)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_1522_add_4_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_1522_add_4_11 (.CI(n28400), .I0(GND_net), 
            .I1(communication_counter[9]), .CO(n28401));
    SB_LUT4 communication_counter_1522_add_4_10_lut (.I0(GND_net), .I1(GND_net), 
            .I2(communication_counter[8]), .I3(n28399), .O(n157)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_1522_add_4_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_1522_add_4_10 (.CI(n28399), .I0(GND_net), 
            .I1(communication_counter[8]), .CO(n28400));
    SB_LUT4 communication_counter_1522_add_4_9_lut (.I0(GND_net), .I1(GND_net), 
            .I2(communication_counter[7]), .I3(n28398), .O(n158)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_1522_add_4_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_1522_add_4_9 (.CI(n28398), .I0(GND_net), 
            .I1(communication_counter[7]), .CO(n28399));
    SB_LUT4 communication_counter_1522_add_4_8_lut (.I0(GND_net), .I1(GND_net), 
            .I2(communication_counter[6]), .I3(n28397), .O(n159)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_1522_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_1522_add_4_8 (.CI(n28397), .I0(GND_net), 
            .I1(communication_counter[6]), .CO(n28398));
    SB_LUT4 rem_4_add_1519_10_lut (.I0(GND_net), .I1(n2250), .I2(VCC_net), 
            .I3(n28204), .O(n2317)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1519_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 communication_counter_1522_add_4_7_lut (.I0(GND_net), .I1(GND_net), 
            .I2(communication_counter[5]), .I3(n28396), .O(n160)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_1522_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_1522_add_4_7 (.CI(n28396), .I0(GND_net), 
            .I1(communication_counter[5]), .CO(n28397));
    SB_LUT4 communication_counter_1522_add_4_6_lut (.I0(GND_net), .I1(GND_net), 
            .I2(communication_counter[4]), .I3(n28395), .O(n161)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_1522_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_1522_add_4_6 (.CI(n28395), .I0(GND_net), 
            .I1(communication_counter[4]), .CO(n28396));
    SB_LUT4 communication_counter_1522_add_4_5_lut (.I0(GND_net), .I1(GND_net), 
            .I2(communication_counter[3]), .I3(n28394), .O(n162)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_1522_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_1522_add_4_5 (.CI(n28394), .I0(GND_net), 
            .I1(communication_counter[3]), .CO(n28395));
    SB_LUT4 communication_counter_1522_add_4_4_lut (.I0(GND_net), .I1(GND_net), 
            .I2(communication_counter[2]), .I3(n28393), .O(n163)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_1522_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_1522_add_4_4 (.CI(n28393), .I0(GND_net), 
            .I1(communication_counter[2]), .CO(n28394));
    SB_LUT4 communication_counter_1522_add_4_3_lut (.I0(GND_net), .I1(GND_net), 
            .I2(communication_counter[1]), .I3(n28392), .O(n164)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_1522_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_1522_add_4_3 (.CI(n28392), .I0(GND_net), 
            .I1(communication_counter[1]), .CO(n28393));
    SB_LUT4 communication_counter_1522_add_4_2_lut (.I0(GND_net), .I1(GND_net), 
            .I2(communication_counter[0]), .I3(VCC_net), .O(n165)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_1522_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_1522_add_4_2 (.CI(VCC_net), .I0(GND_net), 
            .I1(communication_counter[0]), .CO(n28392));
    SB_LUT4 rem_4_add_1117_15_lut (.I0(n1679), .I1(n1646), .I2(VCC_net), 
            .I3(n28391), .O(n1745)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1117_15_lut.LUT_INIT = 16'h8228;
    SB_LUT4 rem_4_add_1117_14_lut (.I0(GND_net), .I1(n1647), .I2(VCC_net), 
            .I3(n28390), .O(n1714)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1117_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1117_14 (.CI(n28390), .I0(n1647), .I1(VCC_net), 
            .CO(n28391));
    SB_LUT4 rem_4_add_1117_13_lut (.I0(GND_net), .I1(n1648), .I2(VCC_net), 
            .I3(n28389), .O(n1715)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1117_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1519_10 (.CI(n28204), .I0(n2250), .I1(VCC_net), 
            .CO(n28205));
    SB_CARRY rem_4_add_1653_7 (.CI(n28070), .I0(n2453), .I1(VCC_net), 
            .CO(n28071));
    SB_CARRY rem_4_add_1117_13 (.CI(n28389), .I0(n1648), .I1(VCC_net), 
            .CO(n28390));
    SB_LUT4 rem_4_add_1117_12_lut (.I0(GND_net), .I1(n1649), .I2(VCC_net), 
            .I3(n28388), .O(n1716)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1117_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1117_12 (.CI(n28388), .I0(n1649), .I1(VCC_net), 
            .CO(n28389));
    SB_LUT4 rem_4_add_1117_11_lut (.I0(GND_net), .I1(n1650), .I2(VCC_net), 
            .I3(n28387), .O(n1717)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1117_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1117_11 (.CI(n28387), .I0(n1650), .I1(VCC_net), 
            .CO(n28388));
    SB_LUT4 rem_4_add_1117_10_lut (.I0(GND_net), .I1(n1651), .I2(VCC_net), 
            .I3(n28386), .O(n1718)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1117_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1117_10 (.CI(n28386), .I0(n1651), .I1(VCC_net), 
            .CO(n28387));
    SB_LUT4 rem_4_add_1117_9_lut (.I0(GND_net), .I1(n1652), .I2(VCC_net), 
            .I3(n28385), .O(n1719)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1117_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1653_6_lut (.I0(GND_net), .I1(n2454), .I2(GND_net), 
            .I3(n28069), .O(n2521)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1653_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1117_9 (.CI(n28385), .I0(n1652), .I1(VCC_net), 
            .CO(n28386));
    SB_LUT4 rem_4_add_1117_8_lut (.I0(GND_net), .I1(n1653), .I2(VCC_net), 
            .I3(n28384), .O(n1720)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1117_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1117_8 (.CI(n28384), .I0(n1653), .I1(VCC_net), 
            .CO(n28385));
    SB_LUT4 rem_4_add_1117_7_lut (.I0(GND_net), .I1(n1654), .I2(GND_net), 
            .I3(n28383), .O(n1721)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1117_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1117_7 (.CI(n28383), .I0(n1654), .I1(GND_net), 
            .CO(n28384));
    SB_LUT4 rem_4_add_1117_6_lut (.I0(GND_net), .I1(n1655), .I2(GND_net), 
            .I3(n28382), .O(n1722)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1117_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1117_6 (.CI(n28382), .I0(n1655), .I1(GND_net), 
            .CO(n28383));
    SB_LUT4 rem_4_add_1117_5_lut (.I0(GND_net), .I1(n1656), .I2(VCC_net), 
            .I3(n28381), .O(n1723)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1117_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1519_9_lut (.I0(GND_net), .I1(n2251), .I2(VCC_net), 
            .I3(n28203), .O(n2318)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1519_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1117_5 (.CI(n28381), .I0(n1656), .I1(VCC_net), 
            .CO(n28382));
    SB_CARRY rem_4_add_1653_6 (.CI(n28069), .I0(n2454), .I1(GND_net), 
            .CO(n28070));
    SB_LUT4 rem_4_add_1117_4_lut (.I0(GND_net), .I1(n1657), .I2(VCC_net), 
            .I3(n28380), .O(n1724)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1117_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1117_4 (.CI(n28380), .I0(n1657), .I1(VCC_net), 
            .CO(n28381));
    SB_LUT4 rem_4_add_1117_3_lut (.I0(GND_net), .I1(n1658), .I2(GND_net), 
            .I3(n28379), .O(n1725)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1117_3_lut.LUT_INIT = 16'hC33C;
    GND i1 (.Y(GND_net));
    SB_CARRY rem_4_add_1117_3 (.CI(n28379), .I0(n1658), .I1(GND_net), 
            .CO(n28380));
    SB_CARRY rem_4_add_1117_2 (.CI(VCC_net), .I0(n1758), .I1(VCC_net), 
            .CO(n28379));
    SB_LUT4 rem_4_add_1184_15_lut (.I0(n1778), .I1(n1745), .I2(VCC_net), 
            .I3(n28378), .O(n1844)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1184_15_lut.LUT_INIT = 16'h8228;
    SB_LUT4 rem_4_add_1184_14_lut (.I0(GND_net), .I1(n1746), .I2(VCC_net), 
            .I3(n28377), .O(n1813)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1184_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1184_14 (.CI(n28377), .I0(n1746), .I1(VCC_net), 
            .CO(n28378));
    SB_LUT4 rem_4_add_1184_13_lut (.I0(GND_net), .I1(n1747), .I2(VCC_net), 
            .I3(n28376), .O(n1814)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1184_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1184_13 (.CI(n28376), .I0(n1747), .I1(VCC_net), 
            .CO(n28377));
    SB_LUT4 rem_4_add_1184_12_lut (.I0(GND_net), .I1(n1748), .I2(VCC_net), 
            .I3(n28375), .O(n1815)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1184_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1184_12 (.CI(n28375), .I0(n1748), .I1(VCC_net), 
            .CO(n28376));
    SB_LUT4 rem_4_add_1184_11_lut (.I0(GND_net), .I1(n1749), .I2(VCC_net), 
            .I3(n28374), .O(n1816)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1184_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1184_11 (.CI(n28374), .I0(n1749), .I1(VCC_net), 
            .CO(n28375));
    SB_LUT4 rem_4_add_1184_10_lut (.I0(GND_net), .I1(n1750), .I2(VCC_net), 
            .I3(n28373), .O(n1817)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1184_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1184_10 (.CI(n28373), .I0(n1750), .I1(VCC_net), 
            .CO(n28374));
    SB_LUT4 rem_4_add_1184_9_lut (.I0(GND_net), .I1(n1751), .I2(VCC_net), 
            .I3(n28372), .O(n1818)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1184_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1184_9 (.CI(n28372), .I0(n1751), .I1(VCC_net), 
            .CO(n28373));
    SB_LUT4 rem_4_add_1653_5_lut (.I0(GND_net), .I1(n2455), .I2(GND_net), 
            .I3(n28068), .O(n2522)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1653_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1184_8_lut (.I0(GND_net), .I1(n1752), .I2(VCC_net), 
            .I3(n28371), .O(n1819)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1184_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1184_8 (.CI(n28371), .I0(n1752), .I1(VCC_net), 
            .CO(n28372));
    SB_LUT4 rem_4_add_1184_7_lut (.I0(GND_net), .I1(n1753), .I2(VCC_net), 
            .I3(n28370), .O(n1820)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1184_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1184_7 (.CI(n28370), .I0(n1753), .I1(VCC_net), 
            .CO(n28371));
    SB_LUT4 rem_4_add_1184_6_lut (.I0(GND_net), .I1(n1754), .I2(GND_net), 
            .I3(n28369), .O(n1821)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1184_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1184_6 (.CI(n28369), .I0(n1754), .I1(GND_net), 
            .CO(n28370));
    SB_LUT4 rem_4_add_1184_5_lut (.I0(GND_net), .I1(n1755), .I2(GND_net), 
            .I3(n28368), .O(n1822)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1184_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1184_5 (.CI(n28368), .I0(n1755), .I1(GND_net), 
            .CO(n28369));
    SB_LUT4 rem_4_add_1184_4_lut (.I0(GND_net), .I1(n1756), .I2(VCC_net), 
            .I3(n28367), .O(n1823)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1184_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1184_4 (.CI(n28367), .I0(n1756), .I1(VCC_net), 
            .CO(n28368));
    SB_LUT4 rem_4_add_1184_3_lut (.I0(GND_net), .I1(n1757), .I2(VCC_net), 
            .I3(n28366), .O(n1824)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1184_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1184_3 (.CI(n28366), .I0(n1757), .I1(VCC_net), 
            .CO(n28367));
    SB_LUT4 rem_4_add_1184_2_lut (.I0(GND_net), .I1(n1758), .I2(GND_net), 
            .I3(VCC_net), .O(n1825)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1184_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1184_2 (.CI(VCC_net), .I0(n1758), .I1(GND_net), 
            .CO(n28366));
    SB_LUT4 rem_4_add_1251_16_lut (.I0(n1877), .I1(n1844), .I2(VCC_net), 
            .I3(n28365), .O(n1943)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1251_16_lut.LUT_INIT = 16'h8228;
    SB_LUT4 rem_4_add_1787_12_lut (.I0(n2648), .I1(n2648), .I2(n2669), 
            .I3(n27884), .O(n2747)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1787_12_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 rem_4_add_1251_15_lut (.I0(GND_net), .I1(n1845), .I2(VCC_net), 
            .I3(n28364), .O(n1912)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1251_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1251_15 (.CI(n28364), .I0(n1845), .I1(VCC_net), 
            .CO(n28365));
    SB_LUT4 rem_4_add_1251_14_lut (.I0(GND_net), .I1(n1846), .I2(VCC_net), 
            .I3(n28363), .O(n1913)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1251_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1251_14 (.CI(n28363), .I0(n1846), .I1(VCC_net), 
            .CO(n28364));
    SB_LUT4 rem_4_add_1251_13_lut (.I0(GND_net), .I1(n1847), .I2(VCC_net), 
            .I3(n28362), .O(n1914)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1251_13_lut.LUT_INIT = 16'hC33C;
    pll32MHz pll32MHz_inst (.GND_net(GND_net), .CLK_c(CLK_c), .VCC_net(VCC_net), 
            .clk32MHz(clk32MHz)) /* synthesis lattice_noprune=1, syn_preserve=0, syn_module_defined=1, syn_noprune=0 */ ;   // verilog/TinyFPGA_B.v(35[10] 38[2])
    SB_CARRY rem_4_add_1251_13 (.CI(n28362), .I0(n1847), .I1(VCC_net), 
            .CO(n28363));
    coms setpoint_23__I_0 (.\data_in_frame[10] ({\data_in_frame[10] }), .clk32MHz(clk32MHz), 
         .\data_out_frame[11] ({\data_out_frame[11] }), .\data_out_frame[9] ({\data_out_frame[9] }), 
         .GND_net(GND_net), .\data_in_frame[8] ({\data_in_frame[8] }), .\data_out_frame[6] ({\data_out_frame[6] }), 
         .rx_data({rx_data}), .\data_in_frame[5] ({\data_in_frame[5] }), 
         .\data_out_frame[8] ({\data_out_frame[8] }), .\data_out_frame[12] ({\data_out_frame[12] }), 
         .\data_out_frame[7] ({\data_out_frame[7] }), .n18202(n18202), .PWMLimit({PWMLimit}), 
         .n18203(n18203), .n18204(n18204), .n18205(n18205), .n18206(n18206), 
         .n18207(n18207), .n18208(n18208), .n18194(n18194), .n18195(n18195), 
         .n18196(n18196), .n18197(n18197), .n18198(n18198), .n18199(n18199), 
         .n34206(n34206), .n38508(n38508), .n18200(n18200), .n18201(n18201), 
         .n18186(n18186), .n18187(n18187), .n18188(n18188), .n18189(n18189), 
         .n18190(n18190), .n18191(n18191), .n18192(n18192), .n18193(n18193), 
         .\data_in_frame[13] ({\data_in_frame[13] }), .\data_out_frame[5] ({\data_out_frame[5] }), 
         .\data_in_frame[12] ({\data_in_frame[12] }), .\data_in_frame[4] ({\data_in_frame[4] }), 
         .n34066(n34066), .\data_in_frame[3] ({\data_in_frame[3] }), .n4997(n4997), 
         .n4998(n4998), .n4999(n4999), .\data_out_frame[13] ({\data_out_frame[13] }), 
         .n5000(n5000), .n5001(n5001), .\data_out_frame[10] ({\data_out_frame[10] }), 
         .n5002(n5002), .n5003(n5003), .\data_in_frame[2] ({\data_in_frame[2] }), 
         .n5004(n5004), .n5005(n5005), .n5006(n5006), .\data_out_frame[16] ({\data_out_frame[16] }), 
         .n5007(n5007), .n5008(n5008), .\data_out_frame[18] ({\data_out_frame[18] }), 
         .n5009(n5009), .n24786(n24786), .\data_out_frame[15] ({\data_out_frame[15] }), 
         .n5010(n5010), .\data_out_frame[20] ({\data_out_frame[20] }), .n5011(n5011), 
         .\data_in_frame[17] ({\data_in_frame[17] }), .\data_in_frame[1] ({\data_in_frame[1] }), 
         .n5012(n5012), .n5013(n5013), .n5014(n5014), .n5015(n5015), 
         .n5016(n5016), .n5017(n5017), .n5018(n5018), .n35492(n35492), 
         .n5019(n5019), .n18025(n18025), .n18024(n18024), .n18023(n18023), 
         .n18022(n18022), .n18021(n18021), .n18020(n18020), .\data_in[1] ({\data_in[1] }), 
         .rx_data_ready(rx_data_ready), .byte_transmit_counter({Open_0, 
         Open_1, Open_2, Open_3, Open_4, Open_5, Open_6, byte_transmit_counter[0]}), 
         .\data_out_frame[17] ({\data_out_frame[17] }), .\data_out_frame[19] ({\data_out_frame[19] }), 
         .\r_SM_Main_2__N_3458[0] (r_SM_Main_2__N_3458[0]), .n18019(n18019), 
         .n18018(n18018), .\data_in_frame[11] ({\data_in_frame[11] }), .n18010(n18010), 
         .control_mode({control_mode}), .n18009(n18009), .n18008(n18008), 
         .n18007(n18007), .n18006(n18006), .n18005(n18005), .n18004(n18004), 
         .n18003(n18003), .\data_out_frame[23][6] (\data_out_frame[23] [6]), 
         .n18002(n18002), .n18001(n18001), .n18000(n18000), .n17999(n17999), 
         .n17998(n17998), .n17997(n17997), .n17996(n17996), .n17995(n17995), 
         .n17994(n17994), .n17993(n17993), .\data_in[2] ({\data_in[2] }), 
         .n17992(n17992), .n17991(n17991), .n17990(n17990), .n13724(n13724), 
         .n17989(n17989), .n16158(n16158), .n16154(n16154), .n3893(n3893), 
         .n3007(n3007), .\data_out_frame[14] ({\data_out_frame[14] }), .n17988(n17988), 
         .n17987(n17987), .n17986(n17986), .n17985(n17985), .n17984(n17984), 
         .n17983(n17983), .\data_in_frame[9] ({\data_in_frame[9] }), .n17982(n17982), 
         .n17981(n17981), .n17980(n17980), .n17979(n17979), .n17978(n17978), 
         .n17977(n17977), .n17976(n17976), .n17975(n17975), .n17974(n17974), 
         .n17973(n17973), .n17972(n17972), .n17971(n17971), .\data_in[0][6] (\data_in[0] [6]), 
         .n17970(n17970), .n17969(n17969), .n17968(n17968), .n17967(n17967), 
         .n17966(n17966), .n17965(n17965), .n17964(n17964), .n17963(n17963), 
         .n17962(n17962), .n17961(n17961), .n17960(n17960), .n17959(n17959), 
         .n17958(n17958), .n17957(n17957), .n17956(n17956), .n33657(n33657), 
         .\data_in[3][0] (\data_in[3] [0]), .\data_in[0][3] (\data_in[0] [3]), 
         .\data_in[0][1] (\data_in[0] [1]), .\data_in[0][5] (\data_in[0] [5]), 
         .\data_in[3][2] (\data_in[3] [2]), .\data_in[3][7] (\data_in[3] [7]), 
         .n17955(n17955), .n17954(n17954), .n17953(n17953), .n17952(n17952), 
         .n17951(n17951), .n17950(n17950), .n17949(n17949), .n17948(n17948), 
         .n17947(n17947), .n17946(n17946), .n17945(n17945), .n17944(n17944), 
         .n17943(n17943), .n17942(n17942), .n17941(n17941), .n17940(n17940), 
         .n17939(n17939), .n17938(n17938), .n17937(n17937), .n17936(n17936), 
         .n17935(n17935), .n17934(n17934), .n17933(n17933), .n17932(n17932), 
         .n17931(n17931), .n17930(n17930), .n17929(n17929), .n17928(n17928), 
         .n17927(n17927), .n17926(n17926), .n17925(n17925), .n17924(n17924), 
         .n17923(n17923), .n17922(n17922), .n17921(n17921), .n17920(n17920), 
         .n17919(n17919), .n17918(n17918), .n17917(n17917), .n17916(n17916), 
         .n17915(n17915), .n17914(n17914), .n17913(n17913), .n17912(n17912), 
         .n17911(n17911), .n17910(n17910), .n17909(n17909), .n17908(n17908), 
         .n17907(n17907), .n17906(n17906), .n17905(n17905), .n17904(n17904), 
         .n17903(n17903), .n17902(n17902), .n17901(n17901), .n17900(n17900), 
         .n17899(n17899), .n17898(n17898), .n17897(n17897), .n17896(n17896), 
         .n17895(n17895), .n17894(n17894), .n17893(n17893), .n17892(n17892), 
         .n17891(n17891), .n17890(n17890), .\data_in[3][6] (\data_in[3] [6]), 
         .n17889(n17889), .n17888(n17888), .\data_in[0][7] (\data_in[0] [7]), 
         .n17887(n17887), .n17886(n17886), .n17885(n17885), .n17884(n17884), 
         .n17883(n17883), .n17882(n17882), .n17881(n17881), .n17880(n17880), 
         .n17879(n17879), .n17878(n17878), .n17877(n17877), .n17876(n17876), 
         .n17875(n17875), .n17874(n17874), .setpoint({setpoint}), .n17873(n17873), 
         .n17872(n17872), .n17871(n17871), .n17870(n17870), .n17869(n17869), 
         .n17868(n17868), .n17867(n17867), .n17866(n17866), .n17865(n17865), 
         .n17864(n17864), .n17863(n17863), .n17862(n17862), .n17861(n17861), 
         .n17860(n17860), .n17859(n17859), .n17858(n17858), .n17857(n17857), 
         .n17856(n17856), .n17855(n17855), .n17854(n17854), .n17853(n17853), 
         .n17852(n17852), .n17851(n17851), .\Ki[15] (Ki[15]), .n17850(n17850), 
         .\Ki[14] (Ki[14]), .n17849(n17849), .\Ki[13] (Ki[13]), .n17848(n17848), 
         .\Ki[12] (Ki[12]), .n17847(n17847), .\Ki[11] (Ki[11]), .n17846(n17846), 
         .\Ki[10] (Ki[10]), .n17845(n17845), .\Ki[9] (Ki[9]), .n17844(n17844), 
         .\Ki[8] (Ki[8]), .n17843(n17843), .\Ki[7] (Ki[7]), .n17842(n17842), 
         .\Ki[6] (Ki[6]), .n17841(n17841), .\Ki[5] (Ki[5]), .n17840(n17840), 
         .\Ki[4] (Ki[4]), .n17839(n17839), .\Ki[3] (Ki[3]), .n63(n63), 
         .n17838(n17838), .\Ki[2] (Ki[2]), .n17837(n17837), .\Ki[1] (Ki[1]), 
         .n17836(n17836), .\Kp[15] (Kp[15]), .n17835(n17835), .\Kp[14] (Kp[14]), 
         .n17834(n17834), .\Kp[13] (Kp[13]), .n17833(n17833), .\Kp[12] (Kp[12]), 
         .n17832(n17832), .\Kp[11] (Kp[11]), .n17831(n17831), .\Kp[10] (Kp[10]), 
         .\data_in[0][0] (\data_in[0] [0]), .\data_in[0][4] (\data_in[0] [4]), 
         .\data_in[3][4] (\data_in[3] [4]), .n17830(n17830), .\Kp[9] (Kp[9]), 
         .n17829(n17829), .\Kp[8] (Kp[8]), .n17828(n17828), .\Kp[7] (Kp[7]), 
         .n17827(n17827), .\Kp[6] (Kp[6]), .n17826(n17826), .\Kp[5] (Kp[5]), 
         .n17825(n17825), .\Kp[4] (Kp[4]), .n17824(n17824), .\Kp[3] (Kp[3]), 
         .n17823(n17823), .\Kp[2] (Kp[2]), .n17822(n17822), .\Kp[1] (Kp[1]), 
         .n17821(n17821), .n17820(n17820), .n17818(n17818), .n17816(n17816), 
         .n17814(n17814), .n17813(n17813), .n17812(n17812), .n17810(n17810), 
         .n17808(n17808), .n17806(n17806), .n33228(n33228), .n737(n737), 
         .\FRAME_MATCHER.state_31__N_2566[1] (\FRAME_MATCHER.state_31__N_2566 [1]), 
         .n4996(n4996), .n5(n5_adj_4786), .n16159(n16159), .n2958(n2958), 
         .n32962(n32962), .n32941(n32941), .n32957(n32957), .n5439(n5439), 
         .n17308(n17308), .PIN_11_c(PIN_11_c), .n17805(n17805), .n4(n4_adj_4909), 
         .n17804(n17804), .n17803(n17803), .n17802(n17802), .n17801(n17801), 
         .n17800(n17800), .n17799(n17799), .n17798(n17798), .n17797(n17797), 
         .n17796(n17796), .n17795(n17795), .n17794(n17794), .n17793(n17793), 
         .n17791(n17791), .n17790(n17790), .IntegralLimit({IntegralLimit}), 
         .n17789(n17789), .n17788(n17788), .n17787(n17787), .n17786(n17786), 
         .n17785(n17785), .n17784(n17784), .n17783(n17783), .n17782(n17782), 
         .n17781(n17781), .n17780(n17780), .n17779(n17779), .n17778(n17778), 
         .LED_c(LED_c), .n17777(n17777), .n17776(n17776), .n17527(n17527), 
         .n18153(n18153), .n18152(n18152), .n18151(n18151), .n18150(n18150), 
         .n18149(n18149), .n18089(n18089), .n17775(n17775), .n17774(n17774), 
         .n18088(n18088), .n17656(n17656), .n25050(n25050), .n17659(n17659), 
         .n18087(n18087), .n18086(n18086), .n18085(n18085), .n17662(n17662), 
         .n17665(n17665), .n18084(n18084), .n18083(n18083), .n18082(n18082), 
         .n17668(n17668), .n18148(n18148), .n18147(n18147), .n17550(n17550), 
         .n17773(n17773), .n17772(n17772), .n17771(n17771), .n17770(n17770), 
         .n17769(n17769), .n17768(n17768), .n17671(n17671), .n17674(n17674), 
         .n8014(n8014), .tx_transmit_N_3355(tx_transmit_N_3355), .n16157(n16157), 
         .n34531(n34531), .n18146(n18146), .\FRAME_MATCHER.state_31__N_2566[2] (\FRAME_MATCHER.state_31__N_2566 [2]), 
         .n17696(n17696), .n17694(n17694), .n17693(n17693), .n17692(n17692), 
         .\Ki[0] (Ki[0]), .n17691(n17691), .\Kp[0] (Kp[0]), .n17690(n17690), 
         .n17658(n17658), .n17661(n17661), .n17664(n17664), .n17667(n17667), 
         .n17670(n17670), .n17673(n17673), .n17676(n17676), .n17731(n17731), 
         .\r_SM_Main[2] (r_SM_Main_adj_5047[2]), .r_Bit_Index({r_Bit_Index_adj_5049}), 
         .n17362(n17362), .n17534(n17534), .n5600(n5600), .\r_Clock_Count[6] (r_Clock_Count_adj_5048[6]), 
         .\r_Clock_Count[7] (r_Clock_Count_adj_5048[7]), .\r_Clock_Count[8] (r_Clock_Count_adj_5048[8]), 
         .\r_Clock_Count[0] (r_Clock_Count_adj_5048[0]), .\r_Clock_Count[3] (r_Clock_Count_adj_5048[3]), 
         .n313(n313), .n314(n314), .n315(n315), .n316(n316), .\r_Clock_Count[5] (r_Clock_Count_adj_5048[5]), 
         .tx_active(tx_active), .n5478(n5478), .n318(n318), .n321(n321), 
         .VCC_net(VCC_net), .tx_o(tx_o), .tx_enable(tx_enable), .n17559(n17559), 
         .n18278(n18278), .n17652(n17652), .n17655(n17655), .n17708(n17708), 
         .n17713(n17713), .n17728(n17728), .n17549(n17549), .n17553(n17553), 
         .n25112(n25112), .\r_SM_Main[1] (r_SM_Main[1]), .n18260(n18260), 
         .r_Rx_Data(r_Rx_Data), .n37332(n37332), .PIN_13_N_105(PIN_13_N_105), 
         .\r_SM_Main[2]_adj_3 (r_SM_Main[2]), .n33769(n33769), .n17681(n17681), 
         .r_Bit_Index_adj_10({r_Bit_Index}), .n5578(n5578), .n24193(n24193), 
         .n4_adj_7(n4_adj_4808), .n4_adj_8(n4_adj_4798), .n16148(n16148), 
         .n25070(n25070), .n1(n1_adj_4923), .n37333(n37333), .n17701(n17701), 
         .n17689(n17689), .n17688(n17688), .n17687(n17687), .n17686(n17686), 
         .n17685(n17685), .n17684(n17684), .n17683(n17683), .n16143(n16143), 
         .n17679(n17679), .n17682(n17682), .n17735(n17735), .n4_adj_9(n4_adj_4822)) /* synthesis lattice_noprune=1, syn_preserve=0, syn_module_defined=1, syn_noprune=0 */ ;   // verilog/TinyFPGA_B.v(183[8] 205[4])
    SB_LUT4 rem_4_add_1251_12_lut (.I0(GND_net), .I1(n1848), .I2(VCC_net), 
            .I3(n28361), .O(n1915)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1251_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1519_9 (.CI(n28203), .I0(n2251), .I1(VCC_net), 
            .CO(n28204));
    SB_CARRY rem_4_add_1653_5 (.CI(n28068), .I0(n2455), .I1(GND_net), 
            .CO(n28069));
    SB_CARRY rem_4_add_1251_12 (.CI(n28361), .I0(n1848), .I1(VCC_net), 
            .CO(n28362));
    SB_LUT4 rem_4_add_1251_11_lut (.I0(GND_net), .I1(n1849), .I2(VCC_net), 
            .I3(n28360), .O(n1916)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1251_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1251_11 (.CI(n28360), .I0(n1849), .I1(VCC_net), 
            .CO(n28361));
    SB_LUT4 rem_4_add_1251_10_lut (.I0(GND_net), .I1(n1850), .I2(VCC_net), 
            .I3(n28359), .O(n1917)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1251_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1251_10 (.CI(n28359), .I0(n1850), .I1(VCC_net), 
            .CO(n28360));
    SB_LUT4 rem_4_add_1251_9_lut (.I0(GND_net), .I1(n1851), .I2(VCC_net), 
            .I3(n28358), .O(n1918)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1251_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1251_9 (.CI(n28358), .I0(n1851), .I1(VCC_net), 
            .CO(n28359));
    SB_LUT4 rem_4_add_1251_8_lut (.I0(GND_net), .I1(n1852), .I2(VCC_net), 
            .I3(n28357), .O(n1919)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1251_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1519_8_lut (.I0(GND_net), .I1(n2252), .I2(VCC_net), 
            .I3(n28202), .O(n2319)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1519_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1251_8 (.CI(n28357), .I0(n1852), .I1(VCC_net), 
            .CO(n28358));
    SB_LUT4 rem_4_add_1251_7_lut (.I0(GND_net), .I1(n1853), .I2(VCC_net), 
            .I3(n28356), .O(n1920)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1251_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1251_7 (.CI(n28356), .I0(n1853), .I1(VCC_net), 
            .CO(n28357));
    SB_LUT4 rem_4_add_1251_6_lut (.I0(GND_net), .I1(n1854), .I2(GND_net), 
            .I3(n28355), .O(n1921)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1251_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1251_6 (.CI(n28355), .I0(n1854), .I1(GND_net), 
            .CO(n28356));
    SB_LUT4 rem_4_add_1251_5_lut (.I0(GND_net), .I1(n1855), .I2(GND_net), 
            .I3(n28354), .O(n1922)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1251_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1251_5 (.CI(n28354), .I0(n1855), .I1(GND_net), 
            .CO(n28355));
    SB_LUT4 rem_4_add_1251_4_lut (.I0(GND_net), .I1(n1856), .I2(VCC_net), 
            .I3(n28353), .O(n1923)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1251_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1251_4 (.CI(n28353), .I0(n1856), .I1(VCC_net), 
            .CO(n28354));
    SB_LUT4 rem_4_add_1251_3_lut (.I0(GND_net), .I1(n1857), .I2(VCC_net), 
            .I3(n28352), .O(n1924)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1251_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1251_3 (.CI(n28352), .I0(n1857), .I1(VCC_net), 
            .CO(n28353));
    SB_CARRY rem_4_add_1519_8 (.CI(n28202), .I0(n2252), .I1(VCC_net), 
            .CO(n28203));
    SB_LUT4 rem_4_add_1251_2_lut (.I0(GND_net), .I1(n1858), .I2(GND_net), 
            .I3(VCC_net), .O(n1925)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1251_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1251_2 (.CI(VCC_net), .I0(n1858), .I1(GND_net), 
            .CO(n28352));
    SB_LUT4 encoder1_position_23__I_0_add_2_25_lut (.I0(GND_net), .I1(encoder1_position[23]), 
            .I2(n2), .I3(n28351), .O(displacement_23__N_80[23])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder1_position_23__I_0_add_2_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder1_position_23__I_0_add_2_24_lut (.I0(GND_net), .I1(encoder1_position[22]), 
            .I2(n3_adj_4834), .I3(n28350), .O(displacement_23__N_80[22])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder1_position_23__I_0_add_2_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder1_position_23__I_0_add_2_24 (.CI(n28350), .I0(encoder1_position[22]), 
            .I1(n3_adj_4834), .CO(n28351));
    SB_LUT4 encoder1_position_23__I_0_add_2_23_lut (.I0(GND_net), .I1(encoder1_position[21]), 
            .I2(n4_adj_4830), .I3(n28349), .O(displacement_23__N_80[21])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder1_position_23__I_0_add_2_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1653_4_lut (.I0(GND_net), .I1(n2456), .I2(VCC_net), 
            .I3(n28067), .O(n2523)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1653_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder1_position_23__I_0_add_2_23 (.CI(n28349), .I0(encoder1_position[21]), 
            .I1(n4_adj_4830), .CO(n28350));
    SB_LUT4 encoder1_position_23__I_0_add_2_22_lut (.I0(GND_net), .I1(encoder1_position[20]), 
            .I2(n5_adj_4827), .I3(n28348), .O(displacement_23__N_80[20])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder1_position_23__I_0_add_2_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder1_position_23__I_0_add_2_22 (.CI(n28348), .I0(encoder1_position[20]), 
            .I1(n5_adj_4827), .CO(n28349));
    SB_CARRY rem_4_add_1653_4 (.CI(n28067), .I0(n2456), .I1(VCC_net), 
            .CO(n28068));
    SB_LUT4 encoder1_position_23__I_0_add_2_21_lut (.I0(GND_net), .I1(encoder1_position[19]), 
            .I2(n6_adj_4825), .I3(n28347), .O(displacement_23__N_80[19])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder1_position_23__I_0_add_2_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder1_position_23__I_0_add_2_21 (.CI(n28347), .I0(encoder1_position[19]), 
            .I1(n6_adj_4825), .CO(n28348));
    SB_LUT4 encoder1_position_23__I_0_add_2_20_lut (.I0(GND_net), .I1(encoder1_position[18]), 
            .I2(n7_adj_4824), .I3(n28346), .O(displacement_23__N_80[18])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder1_position_23__I_0_add_2_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder1_position_23__I_0_add_2_20 (.CI(n28346), .I0(encoder1_position[18]), 
            .I1(n7_adj_4824), .CO(n28347));
    SB_LUT4 encoder1_position_23__I_0_add_2_19_lut (.I0(GND_net), .I1(encoder1_position[17]), 
            .I2(n8_adj_4823), .I3(n28345), .O(displacement_23__N_80[17])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder1_position_23__I_0_add_2_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder1_position_23__I_0_add_2_19 (.CI(n28345), .I0(encoder1_position[17]), 
            .I1(n8_adj_4823), .CO(n28346));
    SB_LUT4 encoder1_position_23__I_0_add_2_18_lut (.I0(GND_net), .I1(encoder1_position[16]), 
            .I2(n9_adj_4812), .I3(n28344), .O(displacement_23__N_80[16])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder1_position_23__I_0_add_2_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder1_position_23__I_0_add_2_18 (.CI(n28344), .I0(encoder1_position[16]), 
            .I1(n9_adj_4812), .CO(n28345));
    SB_LUT4 encoder1_position_23__I_0_add_2_17_lut (.I0(GND_net), .I1(encoder1_position[15]), 
            .I2(n10_adj_4809), .I3(n28343), .O(displacement_23__N_80[15])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder1_position_23__I_0_add_2_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder1_position_23__I_0_add_2_17 (.CI(n28343), .I0(encoder1_position[15]), 
            .I1(n10_adj_4809), .CO(n28344));
    SB_LUT4 encoder1_position_23__I_0_add_2_16_lut (.I0(GND_net), .I1(encoder1_position[14]), 
            .I2(n11_adj_4835), .I3(n28342), .O(displacement_23__N_80[14])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder1_position_23__I_0_add_2_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1519_7_lut (.I0(GND_net), .I1(n2253), .I2(VCC_net), 
            .I3(n28201), .O(n2320)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1519_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder1_position_23__I_0_add_2_16 (.CI(n28342), .I0(encoder1_position[14]), 
            .I1(n11_adj_4835), .CO(n28343));
    SB_LUT4 encoder1_position_23__I_0_add_2_15_lut (.I0(GND_net), .I1(encoder1_position[13]), 
            .I2(n12_adj_4836), .I3(n28341), .O(displacement_23__N_80[13])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder1_position_23__I_0_add_2_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1653_3_lut (.I0(GND_net), .I1(n2457), .I2(VCC_net), 
            .I3(n28066), .O(n2524)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1653_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder1_position_23__I_0_add_2_15 (.CI(n28341), .I0(encoder1_position[13]), 
            .I1(n12_adj_4836), .CO(n28342));
    SB_CARRY rem_4_add_1653_3 (.CI(n28066), .I0(n2457), .I1(VCC_net), 
            .CO(n28067));
    SB_LUT4 encoder1_position_23__I_0_add_2_14_lut (.I0(GND_net), .I1(encoder1_position[12]), 
            .I2(n13_adj_4837), .I3(n28340), .O(displacement_23__N_80[12])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder1_position_23__I_0_add_2_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder1_position_23__I_0_add_2_14 (.CI(n28340), .I0(encoder1_position[12]), 
            .I1(n13_adj_4837), .CO(n28341));
    SB_LUT4 encoder1_position_23__I_0_add_2_13_lut (.I0(GND_net), .I1(encoder1_position[11]), 
            .I2(n14_adj_4838), .I3(n28339), .O(displacement_23__N_80[11])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder1_position_23__I_0_add_2_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1519_7 (.CI(n28201), .I0(n2253), .I1(VCC_net), 
            .CO(n28202));
    SB_CARRY encoder1_position_23__I_0_add_2_13 (.CI(n28339), .I0(encoder1_position[11]), 
            .I1(n14_adj_4838), .CO(n28340));
    SB_LUT4 encoder1_position_23__I_0_add_2_12_lut (.I0(GND_net), .I1(encoder1_position[10]), 
            .I2(n15_adj_4839), .I3(n28338), .O(displacement_23__N_80[10])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder1_position_23__I_0_add_2_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder1_position_23__I_0_add_2_12 (.CI(n28338), .I0(encoder1_position[10]), 
            .I1(n15_adj_4839), .CO(n28339));
    SB_LUT4 encoder1_position_23__I_0_add_2_11_lut (.I0(GND_net), .I1(encoder1_position[9]), 
            .I2(n16_adj_4840), .I3(n28337), .O(displacement_23__N_80[9])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder1_position_23__I_0_add_2_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1519_6_lut (.I0(GND_net), .I1(n2254), .I2(GND_net), 
            .I3(n28200), .O(n2321)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1519_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder1_position_23__I_0_add_2_11 (.CI(n28337), .I0(encoder1_position[9]), 
            .I1(n16_adj_4840), .CO(n28338));
    SB_LUT4 encoder1_position_23__I_0_add_2_10_lut (.I0(GND_net), .I1(encoder1_position[8]), 
            .I2(n17_adj_4841), .I3(n28336), .O(displacement_23__N_80[8])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder1_position_23__I_0_add_2_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i13442_3_lut (.I0(\half_duty[0] [7]), .I1(half_duty_new[7]), 
            .I2(n1466), .I3(GND_net), .O(n18271));   // vhdl/pwm.vhd(59[5] 95[12])
    defparam i13442_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder1_position_23__I_0_add_2_10 (.CI(n28336), .I0(encoder1_position[8]), 
            .I1(n17_adj_4841), .CO(n28337));
    SB_LUT4 encoder1_position_23__I_0_add_2_9_lut (.I0(GND_net), .I1(encoder1_position[7]), 
            .I2(n18_adj_4842), .I3(n28335), .O(displacement_23__N_80[7])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder1_position_23__I_0_add_2_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder1_position_23__I_0_add_2_9 (.CI(n28335), .I0(encoder1_position[7]), 
            .I1(n18_adj_4842), .CO(n28336));
    SB_LUT4 rem_4_add_1653_2_lut (.I0(GND_net), .I1(n2458), .I2(GND_net), 
            .I3(VCC_net), .O(n2525)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1653_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder1_position_23__I_0_add_2_8_lut (.I0(GND_net), .I1(encoder1_position[6]), 
            .I2(n19_adj_4843), .I3(n28334), .O(displacement_23__N_80[6])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder1_position_23__I_0_add_2_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder1_position_23__I_0_add_2_8 (.CI(n28334), .I0(encoder1_position[6]), 
            .I1(n19_adj_4843), .CO(n28335));
    SB_CARRY rem_4_add_1653_2 (.CI(VCC_net), .I0(n2458), .I1(GND_net), 
            .CO(n28066));
    SB_LUT4 encoder1_position_23__I_0_add_2_7_lut (.I0(GND_net), .I1(encoder1_position[5]), 
            .I2(n20_adj_4844), .I3(n28333), .O(displacement_23__N_80[5])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder1_position_23__I_0_add_2_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1720_23_lut (.I0(n2570), .I1(n2537), .I2(VCC_net), 
            .I3(n28065), .O(n2636)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1720_23_lut.LUT_INIT = 16'h8228;
    SB_CARRY encoder1_position_23__I_0_add_2_7 (.CI(n28333), .I0(encoder1_position[5]), 
            .I1(n20_adj_4844), .CO(n28334));
    SB_LUT4 encoder1_position_23__I_0_add_2_6_lut (.I0(GND_net), .I1(encoder1_position[4]), 
            .I2(n21_adj_4845), .I3(n28332), .O(displacement_23__N_80[4])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder1_position_23__I_0_add_2_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder1_position_23__I_0_add_2_6 (.CI(n28332), .I0(encoder1_position[4]), 
            .I1(n21_adj_4845), .CO(n28333));
    SB_LUT4 encoder1_position_23__I_0_add_2_5_lut (.I0(GND_net), .I1(encoder1_position[3]), 
            .I2(n22_adj_4846), .I3(n28331), .O(displacement_23__N_80[3])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder1_position_23__I_0_add_2_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder1_position_23__I_0_add_2_5 (.CI(n28331), .I0(encoder1_position[3]), 
            .I1(n22_adj_4846), .CO(n28332));
    SB_LUT4 encoder1_position_23__I_0_add_2_4_lut (.I0(GND_net), .I1(encoder1_position[2]), 
            .I2(n23_adj_4847), .I3(n28330), .O(displacement_23__N_80[2])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder1_position_23__I_0_add_2_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder1_position_23__I_0_add_2_4 (.CI(n28330), .I0(encoder1_position[2]), 
            .I1(n23_adj_4847), .CO(n28331));
    SB_LUT4 encoder1_position_23__I_0_add_2_3_lut (.I0(GND_net), .I1(encoder1_position[1]), 
            .I2(n24_adj_4848), .I3(n28329), .O(displacement_23__N_80[1])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder1_position_23__I_0_add_2_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder1_position_23__I_0_add_2_3 (.CI(n28329), .I0(encoder1_position[1]), 
            .I1(n24_adj_4848), .CO(n28330));
    SB_LUT4 rem_4_add_1720_22_lut (.I0(GND_net), .I1(n2538), .I2(VCC_net), 
            .I3(n28064), .O(n2605)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1720_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1720_22 (.CI(n28064), .I0(n2538), .I1(VCC_net), 
            .CO(n28065));
    SB_LUT4 encoder1_position_23__I_0_add_2_2_lut (.I0(GND_net), .I1(encoder1_position[0]), 
            .I2(n25_adj_4849), .I3(VCC_net), .O(displacement_23__N_80[0])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder1_position_23__I_0_add_2_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder1_position_23__I_0_add_2_2 (.CI(VCC_net), .I0(encoder1_position[0]), 
            .I1(n25_adj_4849), .CO(n28329));
    SB_LUT4 rem_4_add_1318_17_lut (.I0(n1976), .I1(n1943), .I2(VCC_net), 
            .I3(n28328), .O(n2042)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1318_17_lut.LUT_INIT = 16'h8228;
    SB_LUT4 rem_4_add_1318_16_lut (.I0(GND_net), .I1(n1944), .I2(VCC_net), 
            .I3(n28327), .O(n2011)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1318_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1720_21_lut (.I0(GND_net), .I1(n2539), .I2(VCC_net), 
            .I3(n28063), .O(n2606)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1720_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1318_16 (.CI(n28327), .I0(n1944), .I1(VCC_net), 
            .CO(n28328));
    SB_CARRY rem_4_add_1720_21 (.CI(n28063), .I0(n2539), .I1(VCC_net), 
            .CO(n28064));
    SB_LUT4 rem_4_add_1318_15_lut (.I0(GND_net), .I1(n1945), .I2(VCC_net), 
            .I3(n28326), .O(n2012)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1318_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1318_15 (.CI(n28326), .I0(n1945), .I1(VCC_net), 
            .CO(n28327));
    SB_LUT4 rem_4_add_1318_14_lut (.I0(GND_net), .I1(n1946), .I2(VCC_net), 
            .I3(n28325), .O(n2013)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1318_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1519_6 (.CI(n28200), .I0(n2254), .I1(GND_net), 
            .CO(n28201));
    SB_LUT4 rem_4_add_1720_20_lut (.I0(GND_net), .I1(n2540), .I2(VCC_net), 
            .I3(n28062), .O(n2607)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1720_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1318_14 (.CI(n28325), .I0(n1946), .I1(VCC_net), 
            .CO(n28326));
    SB_LUT4 rem_4_add_1318_13_lut (.I0(GND_net), .I1(n1947), .I2(VCC_net), 
            .I3(n28324), .O(n2014)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1318_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1720_20 (.CI(n28062), .I0(n2540), .I1(VCC_net), 
            .CO(n28063));
    SB_LUT4 rem_4_add_1519_5_lut (.I0(GND_net), .I1(n2255), .I2(GND_net), 
            .I3(n28199), .O(n2322)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1519_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1318_13 (.CI(n28324), .I0(n1947), .I1(VCC_net), 
            .CO(n28325));
    SB_CARRY rem_4_add_1519_5 (.CI(n28199), .I0(n2255), .I1(GND_net), 
            .CO(n28200));
    SB_LUT4 rem_4_add_1318_12_lut (.I0(GND_net), .I1(n1948), .I2(VCC_net), 
            .I3(n28323), .O(n2015)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1318_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1318_12 (.CI(n28323), .I0(n1948), .I1(VCC_net), 
            .CO(n28324));
    SB_LUT4 rem_4_add_1318_11_lut (.I0(GND_net), .I1(n1949), .I2(VCC_net), 
            .I3(n28322), .O(n2016)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1318_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1318_11 (.CI(n28322), .I0(n1949), .I1(VCC_net), 
            .CO(n28323));
    SB_LUT4 rem_4_add_1318_10_lut (.I0(GND_net), .I1(n1950), .I2(VCC_net), 
            .I3(n28321), .O(n2017)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1318_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1318_10 (.CI(n28321), .I0(n1950), .I1(VCC_net), 
            .CO(n28322));
    SB_LUT4 rem_4_add_1519_4_lut (.I0(GND_net), .I1(n2256), .I2(VCC_net), 
            .I3(n28198), .O(n2323)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1519_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1519_4 (.CI(n28198), .I0(n2256), .I1(VCC_net), 
            .CO(n28199));
    SB_LUT4 rem_4_add_1519_3_lut (.I0(GND_net), .I1(n2257), .I2(VCC_net), 
            .I3(n28197), .O(n2324)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1519_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1318_9_lut (.I0(GND_net), .I1(n1951), .I2(VCC_net), 
            .I3(n28320), .O(n2018)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1318_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1519_3 (.CI(n28197), .I0(n2257), .I1(VCC_net), 
            .CO(n28198));
    SB_LUT4 rem_4_add_1720_19_lut (.I0(GND_net), .I1(n2541), .I2(VCC_net), 
            .I3(n28061), .O(n2608)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1720_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1318_9 (.CI(n28320), .I0(n1951), .I1(VCC_net), 
            .CO(n28321));
    SB_CARRY rem_4_add_1720_19 (.CI(n28061), .I0(n2541), .I1(VCC_net), 
            .CO(n28062));
    SB_LUT4 rem_4_add_1318_8_lut (.I0(GND_net), .I1(n1952), .I2(VCC_net), 
            .I3(n28319), .O(n2019)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1318_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1318_8 (.CI(n28319), .I0(n1952), .I1(VCC_net), 
            .CO(n28320));
    SB_LUT4 rem_4_add_1318_7_lut (.I0(GND_net), .I1(n1953), .I2(VCC_net), 
            .I3(n28318), .O(n2020)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1318_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1318_7 (.CI(n28318), .I0(n1953), .I1(VCC_net), 
            .CO(n28319));
    SB_LUT4 rem_4_add_1519_2_lut (.I0(GND_net), .I1(n2258), .I2(GND_net), 
            .I3(VCC_net), .O(n2325)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1519_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1318_6_lut (.I0(GND_net), .I1(n1954), .I2(GND_net), 
            .I3(n28317), .O(n2021)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1318_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1318_6 (.CI(n28317), .I0(n1954), .I1(GND_net), 
            .CO(n28318));
    SB_LUT4 rem_4_add_1318_5_lut (.I0(GND_net), .I1(n1955), .I2(GND_net), 
            .I3(n28316), .O(n2022)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1318_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1318_5 (.CI(n28316), .I0(n1955), .I1(GND_net), 
            .CO(n28317));
    SB_LUT4 rem_4_add_1318_4_lut (.I0(GND_net), .I1(n1956), .I2(VCC_net), 
            .I3(n28315), .O(n2023)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1318_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1318_4 (.CI(n28315), .I0(n1956), .I1(VCC_net), 
            .CO(n28316));
    SB_LUT4 rem_4_add_1318_3_lut (.I0(GND_net), .I1(n1957), .I2(VCC_net), 
            .I3(n28314), .O(n2024)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1318_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1318_3 (.CI(n28314), .I0(n1957), .I1(VCC_net), 
            .CO(n28315));
    SB_LUT4 rem_4_add_1318_2_lut (.I0(GND_net), .I1(n1958), .I2(GND_net), 
            .I3(VCC_net), .O(n2025)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1318_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1318_2 (.CI(VCC_net), .I0(n1958), .I1(GND_net), 
            .CO(n28314));
    SB_CARRY rem_4_add_1519_2 (.CI(VCC_net), .I0(n2258), .I1(GND_net), 
            .CO(n28197));
    SB_LUT4 rem_4_add_1586_21_lut (.I0(n2372), .I1(n2339), .I2(VCC_net), 
            .I3(n28196), .O(n2438)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1586_21_lut.LUT_INIT = 16'h8228;
    \quad(DEBOUNCE_TICKS=100)  quad_counter1 (.n18254(n18254), .encoder1_position({encoder1_position}), 
            .clk32MHz(clk32MHz), .n18255(n18255), .n18256(n18256), .n18252(n18252), 
            .n18253(n18253), .n18250(n18250), .n18251(n18251), .n18248(n18248), 
            .n18249(n18249), .n18246(n18246), .n18247(n18247), .n18244(n18244), 
            .n18245(n18245), .n18241(n18241), .n18242(n18242), .n18243(n18243), 
            .n18239(n18239), .n18240(n18240), .n18235(n18235), .n18236(n18236), 
            .n18237(n18237), .n18238(n18238), .n18234(n18234), .data_o({quadA_debounced_adj_4805, 
            quadB_debounced_adj_4806}), .GND_net(GND_net), .n3158({n3159, 
            n3160, n3161, n3162, n3163, n3164, n3165, n3166, n3167, 
            n3168, n3169, n3170, n3171, n3172, n3173, n3174, n3175, 
            n3176, n3177, n3178, n3179, n3180, n3181, n3182}), 
            .count_enable(count_enable_adj_4807), .n17699(n17699), .PIN_9_c_1(PIN_9_c_1), 
            .n18264(n18264), .reg_B({reg_B_adj_5056}), .n34971(n34971), 
            .PIN_10_c_0(PIN_10_c_0), .n17705(n17705)) /* synthesis lattice_noprune=1, syn_preserve=0, syn_module_defined=1, syn_noprune=0 */ ;   // verilog/TinyFPGA_B.v(240[15] 245[4])
    SB_LUT4 rem_4_add_1720_18_lut (.I0(GND_net), .I1(n2542), .I2(VCC_net), 
            .I3(n28060), .O(n2609)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1720_18_lut.LUT_INIT = 16'hC33C;
    SB_DFF color__i12 (.Q(color[12]), .C(LED_c), .D(n18275));   // verilog/TinyFPGA_B.v(51[8] 74[4])
    SB_DFF blink_65 (.Q(blink), .C(LED_c), .D(blink_N_354));   // verilog/TinyFPGA_B.v(51[8] 74[4])
    SB_CARRY rem_4_add_1720_18 (.CI(n28060), .I0(n2542), .I1(VCC_net), 
            .CO(n28061));
    SB_DFF color__i11 (.Q(color[11]), .C(LED_c), .D(n18274));   // verilog/TinyFPGA_B.v(51[8] 74[4])
    SB_DFF color__i10 (.Q(color[10]), .C(LED_c), .D(n18273));   // verilog/TinyFPGA_B.v(51[8] 74[4])
    SB_LUT4 rem_4_add_1720_17_lut (.I0(GND_net), .I1(n2543), .I2(VCC_net), 
            .I3(n28059), .O(n2610)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1720_17_lut.LUT_INIT = 16'hC33C;
    SB_DFF color__i9 (.Q(color[9]), .C(LED_c), .D(n18272));   // verilog/TinyFPGA_B.v(51[8] 74[4])
    SB_LUT4 rem_4_add_1586_20_lut (.I0(GND_net), .I1(n2340), .I2(VCC_net), 
            .I3(n28195), .O(n2407)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1586_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1720_17 (.CI(n28059), .I0(n2543), .I1(VCC_net), 
            .CO(n28060));
    SB_LUT4 rem_4_add_1720_16_lut (.I0(GND_net), .I1(n2544), .I2(VCC_net), 
            .I3(n28058), .O(n2611)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1720_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1720_16 (.CI(n28058), .I0(n2544), .I1(VCC_net), 
            .CO(n28059));
    SB_CARRY rem_4_add_1586_20 (.CI(n28195), .I0(n2340), .I1(VCC_net), 
            .CO(n28196));
    SB_LUT4 rem_4_add_1720_15_lut (.I0(GND_net), .I1(n2545), .I2(VCC_net), 
            .I3(n28057), .O(n2612)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1720_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1586_19_lut (.I0(GND_net), .I1(n2341), .I2(VCC_net), 
            .I3(n28194), .O(n2408)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1586_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1720_15 (.CI(n28057), .I0(n2545), .I1(VCC_net), 
            .CO(n28058));
    SB_LUT4 rem_4_add_1720_14_lut (.I0(GND_net), .I1(n2546), .I2(VCC_net), 
            .I3(n28056), .O(n2613)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1720_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1586_19 (.CI(n28194), .I0(n2341), .I1(VCC_net), 
            .CO(n28195));
    SB_LUT4 rem_4_add_1586_18_lut (.I0(GND_net), .I1(n2342), .I2(VCC_net), 
            .I3(n28193), .O(n2409)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1586_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1586_18 (.CI(n28193), .I0(n2342), .I1(VCC_net), 
            .CO(n28194));
    SB_LUT4 rem_4_add_1787_11_lut (.I0(n2649), .I1(n2649), .I2(n2669), 
            .I3(n27883), .O(n2748)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1787_11_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY rem_4_add_1720_14 (.CI(n28056), .I0(n2546), .I1(VCC_net), 
            .CO(n28057));
    SB_LUT4 rem_4_add_1586_17_lut (.I0(GND_net), .I1(n2343), .I2(VCC_net), 
            .I3(n28192), .O(n2410)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1586_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1720_13_lut (.I0(GND_net), .I1(n2547), .I2(VCC_net), 
            .I3(n28055), .O(n2614)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1720_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1720_13 (.CI(n28055), .I0(n2547), .I1(VCC_net), 
            .CO(n28056));
    SB_CARRY rem_4_add_1586_17 (.CI(n28192), .I0(n2343), .I1(VCC_net), 
            .CO(n28193));
    SB_LUT4 rem_4_add_1720_12_lut (.I0(GND_net), .I1(n2548), .I2(VCC_net), 
            .I3(n28054), .O(n2615)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1720_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1720_12 (.CI(n28054), .I0(n2548), .I1(VCC_net), 
            .CO(n28055));
    SB_LUT4 rem_4_add_1586_16_lut (.I0(GND_net), .I1(n2344), .I2(VCC_net), 
            .I3(n28191), .O(n2411)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1586_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1586_16 (.CI(n28191), .I0(n2344), .I1(VCC_net), 
            .CO(n28192));
    SB_LUT4 rem_4_add_1720_11_lut (.I0(GND_net), .I1(n2549), .I2(VCC_net), 
            .I3(n28053), .O(n2616)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1720_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_28_inv_0_i22_1_lut (.I0(duty[21]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n4_adj_4772));   // verilog/TinyFPGA_B.v(149[23:28])
    defparam unary_minus_28_inv_0_i22_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 rem_4_add_1586_15_lut (.I0(GND_net), .I1(n2345), .I2(VCC_net), 
            .I3(n28190), .O(n2412)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1586_15_lut.LUT_INIT = 16'hC33C;
    \quad(DEBOUNCE_TICKS=100)_U1  quad_counter0 (.n3208({n3209, n3210, n3211, 
            n3212, n3213, n3214, n3215, n3216, n3217, n3218, n3219, 
            n3220, n3221, n3222, n3223, n3224, n3225, n3226, n3227, 
            n3228, n3229, n3230, n3231, n3232}), .encoder0_position({encoder0_position}), 
            .GND_net(GND_net), .n18226(n18226), .clk32MHz(clk32MHz), .n18227(n18227), 
            .n18228(n18228), .n18229(n18229), .n18230(n18230), .n18231(n18231), 
            .n18222(n18222), .n18223(n18223), .n18224(n18224), .n18225(n18225), 
            .n18220(n18220), .n18221(n18221), .n18218(n18218), .n18219(n18219), 
            .n18216(n18216), .n18217(n18217), .n18214(n18214), .n18215(n18215), 
            .n18212(n18212), .n18213(n18213), .n18209(n18209), .n18210(n18210), 
            .n18211(n18211), .data_o({quadA_debounced, quadB_debounced}), 
            .count_enable(count_enable), .n17697(n17697), .n18261(n18261), 
            .reg_B({reg_B}), .n34970(n34970), .PIN_2_c_0(PIN_2_c_0), .PIN_1_c_1(PIN_1_c_1), 
            .n17700(n17700)) /* synthesis lattice_noprune=1, syn_preserve=0, syn_module_defined=1, syn_noprune=0 */ ;   // verilog/TinyFPGA_B.v(232[15] 237[4])
    SB_CARRY rem_4_add_1586_15 (.CI(n28190), .I0(n2345), .I1(VCC_net), 
            .CO(n28191));
    SB_LUT4 rem_4_add_1586_14_lut (.I0(GND_net), .I1(n2346), .I2(VCC_net), 
            .I3(n28189), .O(n2413)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1586_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1586_14 (.CI(n28189), .I0(n2346), .I1(VCC_net), 
            .CO(n28190));
    SB_CARRY rem_4_add_1720_11 (.CI(n28053), .I0(n2549), .I1(VCC_net), 
            .CO(n28054));
    SB_LUT4 i13431_4_lut (.I0(r_Rx_Data), .I1(rx_data[0]), .I2(n4_adj_4822), 
            .I3(n16143), .O(n18260));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i13431_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i31532_4_lut (.I0(r_SM_Main[2]), .I1(n37332), .I2(n37333), 
            .I3(r_SM_Main[1]), .O(n25112));
    defparam i31532_4_lut.LUT_INIT = 16'h0511;
    SB_LUT4 rem_4_add_1720_10_lut (.I0(GND_net), .I1(n2550), .I2(VCC_net), 
            .I3(n28052), .O(n2617)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1720_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1720_10 (.CI(n28052), .I0(n2550), .I1(VCC_net), 
            .CO(n28053));
    \pwm(32000000,20000,32000000,23,1)  PWM (.pwm_setpoint({pwm_setpoint}), 
            .GND_net(GND_net), .\half_duty_new[0] (half_duty_new[0]), .CLK_c(CLK_c), 
            .n1466(n1466), .n18268(n18268), .\half_duty[0][4] (\half_duty[0] [4]), 
            .n18270(n18270), .\half_duty[0][6] (\half_duty[0] [6]), .n18271(n18271), 
            .\half_duty[0][7] (\half_duty[0] [7]), .n18267(n18267), .\half_duty[0][3] (\half_duty[0] [3]), 
            .n18265(n18265), .\half_duty[0][1] (\half_duty[0] [1]), .n18266(n18266), 
            .\half_duty[0][2] (\half_duty[0] [2]), .\half_duty[0][0] (\half_duty[0] [0]), 
            .PIN_19_c_0(PIN_19_c_0), .VCC_net(VCC_net), .\half_duty_new[1] (half_duty_new[1]), 
            .\half_duty_new[2] (half_duty_new[2]), .\half_duty_new[3] (half_duty_new[3]), 
            .\half_duty_new[4] (half_duty_new[4]), .\half_duty_new[6] (half_duty_new[6]), 
            .\half_duty_new[7] (half_duty_new[7]), .n17710(n17710)) /* synthesis lattice_noprune=1, syn_preserve=0, syn_noprune=0 */ ;   // verilog/TinyFPGA_B.v(131[43] 137[3])
    motorControl control (.PWMLimit({PWMLimit}), .duty({duty}), .GND_net(GND_net), 
            .\Ki[11] (Ki[11]), .\Kp[15] (Kp[15]), .\Kp[9] (Kp[9]), .\Ki[6] (Ki[6]), 
            .\Ki[13] (Ki[13]), .\Ki[14] (Ki[14]), .\Ki[1] (Ki[1]), .\Ki[0] (Ki[0]), 
            .\Ki[15] (Ki[15]), .\Ki[2] (Ki[2]), .\Ki[3] (Ki[3]), .\Ki[4] (Ki[4]), 
            .IntegralLimit({IntegralLimit}), .\Ki[5] (Ki[5]), .\Kp[10] (Kp[10]), 
            .\Ki[7] (Ki[7]), .\Kp[2] (Kp[2]), .\Kp[1] (Kp[1]), .\Ki[12] (Ki[12]), 
            .\Kp[11] (Kp[11]), .\Kp[0] (Kp[0]), .n38238(n38238), .\Kp[3] (Kp[3]), 
            .\Ki[8] (Ki[8]), .\Kp[5] (Kp[5]), .\Kp[6] (Kp[6]), .\Kp[7] (Kp[7]), 
            .\Kp[8] (Kp[8]), .\Ki[9] (Ki[9]), .\Kp[4] (Kp[4]), .\Kp[12] (Kp[12]), 
            .\Kp[13] (Kp[13]), .setpoint({setpoint}), .\Kp[14] (Kp[14]), 
            .\Ki[10] (Ki[10]), .VCC_net(VCC_net), .n25(n25_adj_4775), 
            .clk32MHz(clk32MHz), .motor_state({motor_state})) /* synthesis lattice_noprune=1, syn_preserve=0, syn_module_defined=1, syn_noprune=0 */ ;   // verilog/TinyFPGA_B.v(216[16] 229[4])
    
endmodule
//
// Verilog Description of module neopixel
//

module neopixel (\neo_pixel_transmitter.done , clk32MHz, n31521, VCC_net, 
            bit_ctr, \neo_pixel_transmitter.t0 , GND_net, timer, n37232, 
            n1, n37224, \state[0] , n7, n4, \state[1] , n17229, 
            n35088, n17500, n17567, n37244, n37260, start, \state_3__N_462[1] , 
            n5, n1460, n33701, n37261, n37225, n37262, n20, n37226, 
            n37263, n37304, \color[10] , \color[11] , \color[12] , 
            \color[9] , n37308, n37309, n37330, PIN_8_c, n37251, 
            n17546, n17767, n17766, n17765, n17764, n17763, n17762, 
            n17761, n17760, n17759, n17758, n17757, n17756, n17755, 
            n17754, n17753, n17752, n17751, n17750, n17749, n17748, 
            n17747, n17746, n17745, n17744, n17743, n17742, n17741, 
            n17740, n17739, n17738, n17737, n37335, n37227, n37359, 
            n37360, n37241, n37228, n37361, n37362, n37229, n37230, 
            n37245, n37363, n37364, n31591, n31589, n31587, n31585, 
            n37252, n31583, n31577, n37365, n31575, n31573, n31571, 
            n31569, n31567, n31565, n31563, n31561, n31559, n31557, 
            n37368, n31555, n31553, n31551, n31549, n31547, n31545, 
            n31543, n31541, n31539, n31537, n31535, n31533, n31531, 
            n31529, n31527, n31599, n37231, n37369) /* synthesis lattice_noprune=1, syn_preserve=0, syn_module_defined=1, syn_noprune=0 */ ;
    output \neo_pixel_transmitter.done ;
    input clk32MHz;
    input n31521;
    input VCC_net;
    output [31:0]bit_ctr;
    output [31:0]\neo_pixel_transmitter.t0 ;
    input GND_net;
    output [31:0]timer;
    output n37232;
    input n1;
    output n37224;
    output \state[0] ;
    output n7;
    input n4;
    output \state[1] ;
    output n17229;
    output n35088;
    output n17500;
    input n17567;
    output n37244;
    output n37260;
    output start;
    output \state_3__N_462[1] ;
    output n5;
    output n1460;
    output n33701;
    output n37261;
    output n37225;
    output n37262;
    output n20;
    output n37226;
    output n37263;
    output n37304;
    input \color[10] ;
    input \color[11] ;
    input \color[12] ;
    input \color[9] ;
    output n37308;
    output n37309;
    output n37330;
    output PIN_8_c;
    output n37251;
    input n17546;
    input n17767;
    input n17766;
    input n17765;
    input n17764;
    input n17763;
    input n17762;
    input n17761;
    input n17760;
    input n17759;
    input n17758;
    input n17757;
    input n17756;
    input n17755;
    input n17754;
    input n17753;
    input n17752;
    input n17751;
    input n17750;
    input n17749;
    input n17748;
    input n17747;
    input n17746;
    input n17745;
    input n17744;
    input n17743;
    input n17742;
    input n17741;
    input n17740;
    input n17739;
    input n17738;
    input n17737;
    output n37335;
    output n37227;
    output n37359;
    output n37360;
    output n37241;
    output n37228;
    output n37361;
    output n37362;
    output n37229;
    output n37230;
    output n37245;
    output n37363;
    output n37364;
    input n31591;
    input n31589;
    input n31587;
    input n31585;
    output n37252;
    input n31583;
    input n31577;
    output n37365;
    input n31575;
    input n31573;
    input n31571;
    input n31569;
    input n31567;
    input n31565;
    input n31563;
    input n31561;
    input n31559;
    input n31557;
    output n37368;
    input n31555;
    input n31553;
    input n31551;
    input n31549;
    input n31547;
    input n31545;
    input n31543;
    input n31541;
    input n31539;
    input n31537;
    input n31535;
    input n31533;
    input n31531;
    input n31529;
    input n31527;
    input n31599;
    output n37231;
    output n37369;
    
    wire clk32MHz /* synthesis SET_AS_NETWORK=clk32MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(34[6:14])
    
    wire n28889, n2199, n2225, n28890, n28777, n1403, n1433, n28778, 
        n1503, n1404, n28776, n2299, n2200, n28888, n2300, n2201, 
        n28887, n1504, n1405, n28775, \neo_pixel_transmitter.done_N_670 , 
        n32930, n1505, n1406, n28774, n2301, n2202, n28886, n1506, 
        n1407, n28773, n2302, n2203, n28885;
    wire [31:0]n51;
    
    wire n2303, n2204, n28884, n1507, n1408, n28772, n2304, n2205, 
        n28883, n1508, n1409, n38231, n28771, n2305, n2206, n28882, 
        n3182, n3083, n3116, n29103, n3183, n3084, n29102, n2306, 
        n2207, n28881, n1509, n3184, n3085, n29101, n2307, n2208, 
        n28880, n24, n27957;
    wire [31:0]one_wire_N_613;
    
    wire n1400, n1301, n1334, n28770, n3185, n3086, n29100, n2308, 
        n2209, n38230, n28879, n3186, n3087, n29099, n2309, n3187, 
        n3088, n29098, n2192, n2093, n2126, n28878, n2193, n2094, 
        n28877, n3188, n3089, n29097, n2194, n2095, n28876, n3189, 
        n3090, n29096, n3190, n3091, n29095, n2195, n2096, n28875, 
        n2196, n2097, n28874, n3191, n3092, n29094, n27958, n30, 
        n27956, n2197, n2098, n28873, n3192, n3093, n29093, n27846, 
        n2198, n2099, n28872, n27955, n3193, n3094, n29092, n1401, 
        n1302, n28769, n1402, n1303, n28768, n3194, n3095, n29091, 
        n1109, n24968, n1105, n1104, n1106, n1108, n12, n1103, 
        n1107, n1136, n3195, n3096, n29090, n1235, n38236, n2100, 
        n28871, n27854, n16103, n25098, n4_c, n21929, n21937, 
        n2101, n28870, n1304, n28767, n1205, n1207, n1202, n1206, 
        n14_adj_4629, n1208, n1209, n9, n1203, n1204, n2103, n18, 
        n2109, n25002, n2108, n30_adj_4630, n28, n38235, n1730, 
        n38245, n2105, n2102, n29, n2798, n2804, n2791, n2795, 
        n40, n2796, n2793, n2788, n2808, n38, n2789, n2800, 
        n2803, n2805, n39, n2107, n2104, n2106, n27, n2792, 
        n2787, n2801, n2799, n37, n22, n27954, n2786, n2797, 
        n34, n2794, n2806, n2807, n2790, n42, n1895, n1902, 
        n1899, n1897, n26, n1907, n1909, n19, n1908, n1900, 
        n16_adj_4632, n1904, n1901, n1906, n1898, n24_adj_4633, 
        n46, n2802, n2809, n33, n1905, n1903, n28_adj_4634, n1896, 
        n1928, n2819, n2918, n38243, n1699, n1709, n17_adj_4635, 
        n1698, n1707, n1703, n1705, n21, n1305, n28766, n1704, 
        n1701, n1708, n20_c, n1702, n1697, n24_adj_4636, n3196, 
        n3097, n29089, n28869, n1306, n28765, n1700, n1706, n2324, 
        n38253, n1307, n28764, n1829, n38244, n1308, n28763, n1309, 
        n28762, n28761, n28760, n28759, n3197, n3098, n29088, 
        n28758, n2027, n38241, n28868, n28757, n1608, n1606, n1604, 
        n1603, n20_adj_4638, n1602, n1609, n13_adj_4639, n1598, 
        n1600, n18_adj_4640, n1605, n1599, n22_adj_4641, n28756, 
        n28755, n3198, n3099, n29087, n28867, n28754, n28753, 
        n28752, n14_adj_4643, n12_adj_4644, n28751, n28750, n16_adj_4645, 
        n3199, n3100, n29086, n1601, n1607, n1631, n28749, n28748, 
        n28866, n38237, n28747, n4_adj_4647, n1037, n28746, n1005, 
        n28745, n28865, n3200, n3101, n29085, n1006, n28744, n3201, 
        n3102, n29084, n3202, n3103, n29083, n25_adj_4648, n27953, 
        n1007, n28743, n28864, n3203, n3104, n29082, n3204, n3105, 
        n29081, n1008, n28742, n1009, n38239, n28741;
    wire [31:0]n971;
    
    wire n905, n28740, n3205, n3106, n29080, n3206, n3107, n29079, 
        n28863, n3207, n3108, n29078, n38234, n28862, n3208, n3109, 
        n38233, n29077, n906, n28739, n3209, n33675, n28738, n2984, 
        n3017, n29076, n17391, n28737, n2292, n22_adj_4652, n30_adj_4653, 
        n14852, n28736, n2294, n2297, n34_adj_4654, n2291, n32, 
        n2985, n29075, n2298, n2295, n33_adj_4655, n2986, n29074, 
        n2296, n2293, n31, n1994, n28861, n1995, n28860, n1996, 
        n28859, n2987, n29073, n1997, n28858, n23_adj_4657, n27952, 
        n1998, n28857, n2988, n29072, n6, n2989, n29071, n2990, 
        n29070, n1999, n28856, n27_adj_4659, n27951, n2991, n29069, 
        n2000, n28855, n2001, n28854, n2992, n29068, n2002, n28853, 
        n27950, n27949, n708, n30176, n33673, n2993, n29067, n2994, 
        n29066, n2995, n29065, n2003, n28852, n2004, n28851, n2996, 
        n29064, n27855, n2005, n28850, n36, n46_adj_4660, n21_adj_4661, 
        n36_adj_4662, n2006, n28849, n2997, n29063, n2007, n28848, 
        n14844, n60, n838, n2423, n38252, n27948, n6_adj_4663, 
        n27947, n2998, n29062, n2999, n29061, n7_adj_4664, n27946, 
        n27945, n3000, n29060, n42_adj_4665, n2008, n28847, n27874, 
        n3001, n29059, n3002, n29058, n1809, n25012, n1807, n1801, 
        n18_adj_4667, n32_adj_4668, n44, n50, n48, n49, n2009, 
        n28846, n1802, n1798, n1808, n1804, n24_adj_4669, n1800, 
        n1803, n1805, n22_adj_4670, n1797, n1806, n26_adj_4671, 
        n1796, n1799, n26_adj_4672, n28_adj_4673, n37_adj_4674, n29_adj_4675, 
        n8, n7_adj_4676, n28845, n47, n3003, n29057, n28844, n3004, 
        n29056, n38242, n28843;
    wire [31:0]n133;
    
    wire n30_adj_4677, n48_adj_4678, n34639, n4_adj_4679, n46_adj_4680, 
        n47_adj_4681, n45, n3005, n29055, n27873, n27944, n3006, 
        n29054, n35357, n26_adj_4683, n27943, n28842, n3007, n29053, 
        n27942, n28841, n44_adj_4686, n3008, n29052, n28840, n28839, 
        n3009, n38240, n29051, n28838, n28837, n27941, n43, n54, 
        n49_adj_4690, n37295, n28836, n2885, n29050, n28835, n2886, 
        n29049, n27940, n4_adj_4692, n2887, n29048, n28834, n2888, 
        n29047, n28833, n27872, n2889, n29046, n28832, n2890, 
        n29045, n2891, n29044, n28831, n2892, n29043, n2893, n29042, 
        n28830, n2894, n29041, n28829, n28828, n2895, n29040, 
        n2896, n29039, n28827, n27853, n2897, n29038, n18_adj_4697, 
        n2403, n2409, n27_adj_4698, n2390, n2391, n2397, n2394, 
        n33_adj_4699, n28_adj_4700, n2392, n2405, n2400, n2398, 
        n32_adj_4701, n2396, n2402, n2408, n2399, n31_adj_4702, 
        n26_adj_4703, n2393, n2406, n2395, n2407, n35, n2404, 
        n2401, n37_adj_4704, n2522, n38251, n2902, n2909, n28_adj_4705, 
        n2900, n2906, n2908, n40_adj_4706, n27_adj_4707, n25_adj_4708, 
        n38_adj_4709, n38247, n2907, n2904, n43_adj_4710, n2898, 
        n2903, n42_adj_4711, n40_adj_4712, n44_adj_4713, n42_adj_4714, 
        n2905, n41, n2901, n2899, n45_adj_4715, n43_adj_4716, n41_adj_4717, 
        n38_adj_4718, n47_adj_4719, n46_adj_4720, n50_adj_4721, n37_adj_4722, 
        n2491, n2504, n24_adj_4723, n2496, n2505, n2500, n2499, 
        n34_adj_4724, n2497, n2509, n22_adj_4725, n2490, n2494, 
        n38_adj_4726, n2501, n2502, n2506, n2492, n36_adj_4727, 
        n2495, n2498, n2493, n37_adj_4728, n2507, n2508, n2503, 
        n2489, n35_adj_4729, n2621, n38249, n1500, n1501, n18_adj_4730, 
        n1502, n1499, n20_adj_4731, n15_adj_4732, n1532, n38250, 
        n2591, n2608, n2601, n2605, n36_adj_4733, n2606, n2609, 
        n25_adj_4734, n2593, n2596, n2600, n2590, n34_adj_4735, 
        n2594, n2589, n40_adj_4736, n2602, n2588, n2604, n2607, 
        n38_adj_4737, n2598, n2603, n39_adj_4738, n2592, n2597, 
        n2595, n2599, n37_adj_4739, n28826, n28825, n29037, n28824, 
        n29036, n28823, n29035, n28822, n28821, n29034, n28820, 
        n29033, n28819, n29032, n28818, n29031, n2720, n38248, 
        n28817, n29030, n28816, n29029, n28815, n29028, n28814, 
        n29027, n28813, n28812, n29026, n28811, n28810, n29025, 
        n29024, n28809, n29023, n28808, n29022, n28807, n29021, 
        n28806, n27871, n29020, n28805, n28804, n29019, n28803, 
        n28802, n29018, n29017, n28801, n37325, n37323, n28_adj_4740, 
        n29016, n28800, n35059, \neo_pixel_transmitter.done_N_676 , 
        n807, n28799, n29015, n28798, n29014, n28797, n27847, 
        n27852, n27870, n29013, n28796, n2693, n2704, n28_adj_4742, 
        n2699, n2706, n2694, n2691, n38_adj_4743, n2709, n24956, 
        n2701, n2696, n2697, n36_adj_4744, n2700, n2705, n42_adj_4745, 
        n2702, n2690, n2689, n2708, n40_adj_4746, n2687, n2703, 
        n2695, n41_adj_4747, n2688, n2698, n2692, n2707, n39_adj_4748, 
        n29012, n28795, n28794, n24998, n16_adj_4749, n29011, n29010, 
        n29009, n29008, n29007, n29006, n38246;
    wire [3:0]state_3__N_462;
    
    wire n27869, n29005, n14_adj_4750, n13_adj_4751, n24860, n34_adj_4752, 
        n23_adj_4753, n22_adj_4754, n38_adj_4755, n36_adj_4756, n37_adj_4757, 
        n29004, n35_adj_4758, n24890, n9_adj_4759, n4_adj_4760, n37779, 
        n36317, n14_adj_4761, n29003, n17_adj_4762, n27868, n27867, 
        n29002, n32854, n27866, n17243, n29001, n29000, n28999, 
        n28998, n28997, n28996, n28995, n28994, n28993, n28992, 
        n28_adj_4763, n32_adj_4764, n30_adj_4765, n31_adj_4766, n29_adj_4767, 
        n28991, n27845, n28990, n28989, n28988, n28987, n28986, 
        n28985, n28984, n28983, n28982, n28981, n28980, n27865, 
        n28979, n28978, n28977, n28976, n28975, n28974, n28465, 
        n28464, n28973, n28972, n28463, n28971, n28462, n27851, 
        n28461, n28460, n28970, n28459, n27864, n28969, n28968, 
        n28458, n28457, n28779, n28967, n28456, n28966, n28780, 
        n28455, n28965, n28454, n27970, n28453, n28964, n28452, 
        n27863, n27844, n28451, n28450, n27850, n28963, n28781, 
        n28449, n28448, n28447, n28446, n28782, n28962, n28445, 
        n28444, n28443, n28961, n28442, n28441, n28960, n28440, 
        n28439, n28438, n28437, n28959, n28436, n28958, n28435, 
        n28957, n27862, n28956, n28955, n28954, n28953, n2_adj_4768, 
        n28952, n28951, n28950, n28949, n28948, n28947, n28946, 
        n28945, n28944, n28943, n28942, n27969, n28941, n28793, 
        n28940, n28792, n28939, n28938, n28791, n28937, n28790, 
        n28936, n28789, n28788, n28787, n28935, n27968, n28934, 
        n28786, n28933, n28785, n28784, n28932, n27861, n27967, 
        n28783, n27849, n28931, n28930, n28929, n28928, n28927, 
        n27848, n27860, n28926, n27966, n28925, n28924, n27965, 
        n28923, n28922, n27964, n27963, n27859, n28921, n27858, 
        n28920, n27962, n28919, n27857, n28918, n28917, n27856, 
        n28916, n28915, n28914, n28913, n28912, n28911, n28910, 
        n28909, n36426, n28908, n27961, n28907, n28906, n28905, 
        n28904, n28903, n28902, n28901, n28900, n28899, n27960, 
        n28898, n27959, n36434, n6_adj_4769, n28897, n28896, n28895, 
        n28894, n28893, n28892, n28891;
    
    SB_CARRY mod_5_add_1540_13 (.CI(n28889), .I0(n2199), .I1(n2225), .CO(n28890));
    SB_CARRY mod_5_add_1004_9 (.CI(n28777), .I0(n1403), .I1(n1433), .CO(n28778));
    SB_LUT4 mod_5_add_1004_8_lut (.I0(n1404), .I1(n1404), .I2(n1433), 
            .I3(n28776), .O(n1503)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1004_8_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1540_12_lut (.I0(n2200), .I1(n2200), .I2(n2225), 
            .I3(n28888), .O(n2299)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_12_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1004_8 (.CI(n28776), .I0(n1404), .I1(n1433), .CO(n28777));
    SB_CARRY mod_5_add_1540_12 (.CI(n28888), .I0(n2200), .I1(n2225), .CO(n28889));
    SB_LUT4 mod_5_add_1540_11_lut (.I0(n2201), .I1(n2201), .I2(n2225), 
            .I3(n28887), .O(n2300)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_11_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1004_7_lut (.I0(n1405), .I1(n1405), .I2(n1433), 
            .I3(n28775), .O(n1504)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1004_7_lut.LUT_INIT = 16'hCA3A;
    SB_DFFE \neo_pixel_transmitter.done_104  (.Q(\neo_pixel_transmitter.done ), 
            .C(clk32MHz), .E(n32930), .D(\neo_pixel_transmitter.done_N_670 ));   // verilog/neopixel.v(35[12] 117[6])
    SB_CARRY mod_5_add_1004_7 (.CI(n28775), .I0(n1405), .I1(n1433), .CO(n28776));
    SB_CARRY mod_5_add_1540_11 (.CI(n28887), .I0(n2201), .I1(n2225), .CO(n28888));
    SB_LUT4 mod_5_add_1004_6_lut (.I0(n1406), .I1(n1406), .I2(n1433), 
            .I3(n28774), .O(n1505)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1004_6_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1004_6 (.CI(n28774), .I0(n1406), .I1(n1433), .CO(n28775));
    SB_LUT4 mod_5_add_1540_10_lut (.I0(n2202), .I1(n2202), .I2(n2225), 
            .I3(n28886), .O(n2301)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_10_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1004_5_lut (.I0(n1407), .I1(n1407), .I2(n1433), 
            .I3(n28773), .O(n1506)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1004_5_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1004_5 (.CI(n28773), .I0(n1407), .I1(n1433), .CO(n28774));
    SB_CARRY mod_5_add_1540_10 (.CI(n28886), .I0(n2202), .I1(n2225), .CO(n28887));
    SB_LUT4 mod_5_add_1540_9_lut (.I0(n2203), .I1(n2203), .I2(n2225), 
            .I3(n28885), .O(n2302)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_9_lut.LUT_INIT = 16'hCA3A;
    SB_DFFE bit_ctr_i0_i31 (.Q(bit_ctr[31]), .C(clk32MHz), .E(VCC_net), 
            .D(n31521));   // verilog/neopixel.v(35[12] 117[6])
    SB_CARRY mod_5_add_1540_9 (.CI(n28885), .I0(n2203), .I1(n2225), .CO(n28886));
    SB_LUT4 sub_14_inv_0_i17_1_lut (.I0(\neo_pixel_transmitter.t0 [16]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n51[16]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i17_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mod_5_add_1540_8_lut (.I0(n2204), .I1(n2204), .I2(n2225), 
            .I3(n28884), .O(n2303)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_8_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1004_4_lut (.I0(n1408), .I1(n1408), .I2(n1433), 
            .I3(n28772), .O(n1507)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1004_4_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1540_8 (.CI(n28884), .I0(n2204), .I1(n2225), .CO(n28885));
    SB_LUT4 mod_5_add_1540_7_lut (.I0(n2205), .I1(n2205), .I2(n2225), 
            .I3(n28883), .O(n2304)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_7_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1004_4 (.CI(n28772), .I0(n1408), .I1(n1433), .CO(n28773));
    SB_LUT4 mod_5_add_1004_3_lut (.I0(n1409), .I1(n1409), .I2(n38231), 
            .I3(n28771), .O(n1508)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1004_3_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1540_7 (.CI(n28883), .I0(n2205), .I1(n2225), .CO(n28884));
    SB_LUT4 mod_5_add_1540_6_lut (.I0(n2206), .I1(n2206), .I2(n2225), 
            .I3(n28882), .O(n2305)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_6_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_2143_29_lut (.I0(n3083), .I1(n3083), .I2(n3116), 
            .I3(n29103), .O(n3182)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_29_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1540_6 (.CI(n28882), .I0(n2206), .I1(n2225), .CO(n28883));
    SB_CARRY mod_5_add_1004_3 (.CI(n28771), .I0(n1409), .I1(n38231), .CO(n28772));
    SB_LUT4 mod_5_add_2143_28_lut (.I0(n3084), .I1(n3084), .I2(n3116), 
            .I3(n29102), .O(n3183)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_28_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2143_28 (.CI(n29102), .I0(n3084), .I1(n3116), .CO(n29103));
    SB_LUT4 mod_5_add_1540_5_lut (.I0(n2207), .I1(n2207), .I2(n2225), 
            .I3(n28881), .O(n2306)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_5_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1004_2_lut (.I0(bit_ctr[21]), .I1(bit_ctr[21]), .I2(n38231), 
            .I3(VCC_net), .O(n1509)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1004_2_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 mod_5_add_2143_27_lut (.I0(n3085), .I1(n3085), .I2(n3116), 
            .I3(n29101), .O(n3184)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_27_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1540_5 (.CI(n28881), .I0(n2207), .I1(n2225), .CO(n28882));
    SB_CARRY mod_5_add_2143_27 (.CI(n29101), .I0(n3085), .I1(n3116), .CO(n29102));
    SB_LUT4 mod_5_add_1540_4_lut (.I0(n2208), .I1(n2208), .I2(n2225), 
            .I3(n28880), .O(n2307)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_4_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1004_2 (.CI(VCC_net), .I0(bit_ctr[21]), .I1(n38231), 
            .CO(n28771));
    SB_CARRY mod_5_add_1540_4 (.CI(n28880), .I0(n2208), .I1(n2225), .CO(n28881));
    SB_LUT4 sub_14_add_2_20_lut (.I0(one_wire_N_613[16]), .I1(timer[18]), 
            .I2(n51[18]), .I3(n27957), .O(n24)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_20_lut.LUT_INIT = 16'hebbe;
    SB_LUT4 mod_5_add_937_11_lut (.I0(n1301), .I1(n1301), .I2(n1334), 
            .I3(n28770), .O(n1400)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_937_11_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_2143_26_lut (.I0(n3086), .I1(n3086), .I2(n3116), 
            .I3(n29100), .O(n3185)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_26_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1540_3_lut (.I0(n2209), .I1(n2209), .I2(n38230), 
            .I3(n28879), .O(n2308)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_3_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_2143_26 (.CI(n29100), .I0(n3086), .I1(n3116), .CO(n29101));
    SB_CARRY mod_5_add_1540_3 (.CI(n28879), .I0(n2209), .I1(n38230), .CO(n28880));
    SB_LUT4 mod_5_add_2143_25_lut (.I0(n3087), .I1(n3087), .I2(n3116), 
            .I3(n29099), .O(n3186)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_25_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2143_25 (.CI(n29099), .I0(n3087), .I1(n3116), .CO(n29100));
    SB_LUT4 mod_5_add_1540_2_lut (.I0(bit_ctr[13]), .I1(bit_ctr[13]), .I2(n38230), 
            .I3(VCC_net), .O(n2309)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_2_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1540_2 (.CI(VCC_net), .I0(bit_ctr[13]), .I1(n38230), 
            .CO(n28879));
    SB_LUT4 mod_5_add_2143_24_lut (.I0(n3088), .I1(n3088), .I2(n3116), 
            .I3(n29098), .O(n3187)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_24_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1473_19_lut (.I0(n2093), .I1(n2093), .I2(n2126), 
            .I3(n28878), .O(n2192)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_19_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2143_24 (.CI(n29098), .I0(n3088), .I1(n3116), .CO(n29099));
    SB_LUT4 mod_5_add_1473_18_lut (.I0(n2094), .I1(n2094), .I2(n2126), 
            .I3(n28877), .O(n2193)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_18_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_2143_23_lut (.I0(n3089), .I1(n3089), .I2(n3116), 
            .I3(n29097), .O(n3188)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_23_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1473_18 (.CI(n28877), .I0(n2094), .I1(n2126), .CO(n28878));
    SB_CARRY mod_5_add_2143_23 (.CI(n29097), .I0(n3089), .I1(n3116), .CO(n29098));
    SB_LUT4 mod_5_add_1473_17_lut (.I0(n2095), .I1(n2095), .I2(n2126), 
            .I3(n28876), .O(n2194)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_17_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_2143_22_lut (.I0(n3090), .I1(n3090), .I2(n3116), 
            .I3(n29096), .O(n3189)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_22_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1473_17 (.CI(n28876), .I0(n2095), .I1(n2126), .CO(n28877));
    SB_CARRY mod_5_add_2143_22 (.CI(n29096), .I0(n3090), .I1(n3116), .CO(n29097));
    SB_LUT4 mod_5_add_2143_21_lut (.I0(n3091), .I1(n3091), .I2(n3116), 
            .I3(n29095), .O(n3190)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_21_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1473_16_lut (.I0(n2096), .I1(n2096), .I2(n2126), 
            .I3(n28875), .O(n2195)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_16_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1473_16 (.CI(n28875), .I0(n2096), .I1(n2126), .CO(n28876));
    SB_CARRY mod_5_add_2143_21 (.CI(n29095), .I0(n3091), .I1(n3116), .CO(n29096));
    SB_LUT4 mod_5_add_1473_15_lut (.I0(n2097), .I1(n2097), .I2(n2126), 
            .I3(n28874), .O(n2196)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_15_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_2143_20_lut (.I0(n3092), .I1(n3092), .I2(n3116), 
            .I3(n29094), .O(n3191)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_20_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1473_15 (.CI(n28874), .I0(n2097), .I1(n2126), .CO(n28875));
    SB_CARRY sub_14_add_2_20 (.CI(n27957), .I0(timer[18]), .I1(n51[18]), 
            .CO(n27958));
    SB_LUT4 sub_14_add_2_19_lut (.I0(one_wire_N_613[23]), .I1(timer[17]), 
            .I2(n51[17]), .I3(n27956), .O(n30)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_19_lut.LUT_INIT = 16'hebbe;
    SB_CARRY mod_5_add_2143_20 (.CI(n29094), .I0(n3092), .I1(n3116), .CO(n29095));
    SB_LUT4 mod_5_add_1473_14_lut (.I0(n2098), .I1(n2098), .I2(n2126), 
            .I3(n28873), .O(n2197)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_14_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY sub_14_add_2_19 (.CI(n27956), .I0(timer[17]), .I1(n51[17]), 
            .CO(n27957));
    SB_LUT4 mod_5_add_2143_19_lut (.I0(n3093), .I1(n3093), .I2(n3116), 
            .I3(n29093), .O(n3192)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_19_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1473_14 (.CI(n28873), .I0(n2098), .I1(n2126), .CO(n28874));
    SB_LUT4 add_21_5_lut (.I0(n1), .I1(bit_ctr[3]), .I2(GND_net), .I3(n27846), 
            .O(n37232)) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_5_lut.LUT_INIT = 16'h8228;
    SB_CARRY mod_5_add_2143_19 (.CI(n29093), .I0(n3093), .I1(n3116), .CO(n29094));
    SB_LUT4 mod_5_add_1473_13_lut (.I0(n2099), .I1(n2099), .I2(n2126), 
            .I3(n28872), .O(n2198)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_13_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 sub_14_add_2_18_lut (.I0(GND_net), .I1(timer[16]), .I2(n51[16]), 
            .I3(n27955), .O(one_wire_N_613[16])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1473_13 (.CI(n28872), .I0(n2099), .I1(n2126), .CO(n28873));
    SB_LUT4 mod_5_add_2143_18_lut (.I0(n3094), .I1(n3094), .I2(n3116), 
            .I3(n29092), .O(n3193)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_18_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_937_10_lut (.I0(n1302), .I1(n1302), .I2(n1334), 
            .I3(n28769), .O(n1401)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_937_10_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_937_10 (.CI(n28769), .I0(n1302), .I1(n1334), .CO(n28770));
    SB_LUT4 mod_5_add_937_9_lut (.I0(n1303), .I1(n1303), .I2(n1334), .I3(n28768), 
            .O(n1402)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_937_9_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_937_9 (.CI(n28768), .I0(n1303), .I1(n1334), .CO(n28769));
    SB_CARRY mod_5_add_2143_18 (.CI(n29092), .I0(n3094), .I1(n3116), .CO(n29093));
    SB_LUT4 mod_5_add_2143_17_lut (.I0(n3095), .I1(n3095), .I2(n3116), 
            .I3(n29091), .O(n3194)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_17_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 sub_14_inv_0_i18_1_lut (.I0(\neo_pixel_transmitter.t0 [17]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n51[17]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i18_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i20146_2_lut (.I0(bit_ctr[24]), .I1(n1109), .I2(GND_net), 
            .I3(GND_net), .O(n24968));
    defparam i20146_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i5_4_lut (.I0(n1105), .I1(n1104), .I2(n1106), .I3(n1108), 
            .O(n12));
    defparam i5_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i6_4_lut (.I0(n1103), .I1(n12), .I2(n1107), .I3(n24968), 
            .O(n1136));
    defparam i6_4_lut.LUT_INIT = 16'hfffe;
    SB_CARRY mod_5_add_2143_17 (.CI(n29091), .I0(n3095), .I1(n3116), .CO(n29092));
    SB_LUT4 mod_5_add_2143_16_lut (.I0(n3096), .I1(n3096), .I2(n3116), 
            .I3(n29090), .O(n3195)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_16_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i31556_1_lut (.I0(n1235), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n38236));
    defparam i31556_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mod_5_add_1473_12_lut (.I0(n2100), .I1(n2100), .I2(n2126), 
            .I3(n28871), .O(n2199)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_12_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY sub_14_add_2_18 (.CI(n27955), .I0(timer[16]), .I1(n51[16]), 
            .CO(n27956));
    SB_CARRY mod_5_add_2143_16 (.CI(n29090), .I0(n3096), .I1(n3116), .CO(n29091));
    SB_CARRY mod_5_add_1473_12 (.CI(n28871), .I0(n2100), .I1(n2126), .CO(n28872));
    SB_LUT4 add_21_13_lut (.I0(n1), .I1(bit_ctr[11]), .I2(GND_net), .I3(n27854), 
            .O(n37224)) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_13_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i20273_4_lut (.I0(one_wire_N_613[11]), .I1(n16103), .I2(one_wire_N_613[9]), 
            .I3(one_wire_N_613[10]), .O(n25098));
    defparam i20273_4_lut.LUT_INIT = 16'heeec;
    SB_LUT4 i1_2_lut (.I0(n25098), .I1(\neo_pixel_transmitter.done ), .I2(GND_net), 
            .I3(GND_net), .O(n4_c));   // verilog/neopixel.v(36[4] 116[11])
    defparam i1_2_lut.LUT_INIT = 16'hdddd;
    SB_LUT4 i17117_3_lut (.I0(n21929), .I1(n21937), .I2(\state[0] ), .I3(GND_net), 
            .O(n7));   // verilog/neopixel.v(16[20:25])
    defparam i17117_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 sub_14_inv_0_i20_1_lut (.I0(\neo_pixel_transmitter.t0 [19]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n51[19]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i20_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mod_5_add_1473_11_lut (.I0(n2101), .I1(n2101), .I2(n2126), 
            .I3(n28870), .O(n2200)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_11_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i1_4_lut (.I0(\state[0] ), .I1(n4), .I2(n4_c), .I3(\state[1] ), 
            .O(n17229));
    defparam i1_4_lut.LUT_INIT = 16'hafcc;
    SB_LUT4 i12_3_lut (.I0(n4), .I1(n35088), .I2(\state[1] ), .I3(GND_net), 
            .O(n17500));   // verilog/neopixel.v(35[12] 117[6])
    defparam i12_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 mod_5_add_937_8_lut (.I0(n1304), .I1(n1304), .I2(n1334), .I3(n28767), 
            .O(n1403)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_937_8_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i6_4_lut_adj_1473 (.I0(n1205), .I1(n1207), .I2(n1202), .I3(n1206), 
            .O(n14_adj_4629));
    defparam i6_4_lut_adj_1473.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_3_lut (.I0(bit_ctr[23]), .I1(n1208), .I2(n1209), .I3(GND_net), 
            .O(n9));
    defparam i1_3_lut.LUT_INIT = 16'hecec;
    SB_LUT4 i7_4_lut (.I0(n9), .I1(n14_adj_4629), .I2(n1203), .I3(n1204), 
            .O(n1235));
    defparam i7_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_adj_1474 (.I0(n2103), .I1(n2097), .I2(GND_net), .I3(GND_net), 
            .O(n18));
    defparam i1_2_lut_adj_1474.LUT_INIT = 16'heeee;
    SB_LUT4 i20180_2_lut (.I0(bit_ctr[14]), .I1(n2109), .I2(GND_net), 
            .I3(GND_net), .O(n25002));
    defparam i20180_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i13_4_lut (.I0(n2093), .I1(n2108), .I2(n2100), .I3(n18), 
            .O(n30_adj_4630));
    defparam i13_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i11_4_lut (.I0(n2098), .I1(n25002), .I2(n2094), .I3(n2099), 
            .O(n28));
    defparam i11_4_lut.LUT_INIT = 16'hfffe;
    SB_CARRY mod_5_add_937_8 (.CI(n28767), .I0(n1304), .I1(n1334), .CO(n28768));
    SB_LUT4 i31555_1_lut (.I0(n1334), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n38235));
    defparam i31555_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i31565_1_lut (.I0(n1730), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n38245));
    defparam i31565_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i12_4_lut (.I0(n2105), .I1(n2096), .I2(n2095), .I3(n2102), 
            .O(n29));
    defparam i12_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i16_4_lut (.I0(n2798), .I1(n2804), .I2(n2791), .I3(n2795), 
            .O(n40));
    defparam i16_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i14_4_lut (.I0(n2796), .I1(n2793), .I2(n2788), .I3(n2808), 
            .O(n38));
    defparam i14_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i15_4_lut (.I0(n2789), .I1(n2800), .I2(n2803), .I3(n2805), 
            .O(n39));
    defparam i15_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i10_4_lut (.I0(n2101), .I1(n2107), .I2(n2104), .I3(n2106), 
            .O(n27));
    defparam i10_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i16_4_lut_adj_1475 (.I0(n27), .I1(n29), .I2(n28), .I3(n30_adj_4630), 
            .O(n2126));
    defparam i16_4_lut_adj_1475.LUT_INIT = 16'hfffe;
    SB_LUT4 i13_4_lut_adj_1476 (.I0(n2792), .I1(n2787), .I2(n2801), .I3(n2799), 
            .O(n37));
    defparam i13_4_lut_adj_1476.LUT_INIT = 16'hfffe;
    SB_CARRY mod_5_add_1473_11 (.CI(n28870), .I0(n2101), .I1(n2126), .CO(n28871));
    SB_LUT4 sub_14_add_2_17_lut (.I0(one_wire_N_613[22]), .I1(timer[15]), 
            .I2(n51[15]), .I3(n27954), .O(n22)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_17_lut.LUT_INIT = 16'hebbe;
    SB_LUT4 i10_2_lut (.I0(n2786), .I1(n2797), .I2(GND_net), .I3(GND_net), 
            .O(n34));
    defparam i10_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i18_4_lut (.I0(n2794), .I1(n2806), .I2(n2807), .I3(n2790), 
            .O(n42));
    defparam i18_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i11_4_lut_adj_1477 (.I0(n1895), .I1(n1902), .I2(n1899), .I3(n1897), 
            .O(n26));
    defparam i11_4_lut_adj_1477.LUT_INIT = 16'hfffe;
    SB_LUT4 i4_3_lut (.I0(n1907), .I1(bit_ctr[16]), .I2(n1909), .I3(GND_net), 
            .O(n19));
    defparam i4_3_lut.LUT_INIT = 16'heaea;
    SB_LUT4 i1_2_lut_adj_1478 (.I0(n1908), .I1(n1900), .I2(GND_net), .I3(GND_net), 
            .O(n16_adj_4632));
    defparam i1_2_lut_adj_1478.LUT_INIT = 16'heeee;
    SB_LUT4 i9_4_lut (.I0(n1904), .I1(n1901), .I2(n1906), .I3(n1898), 
            .O(n24_adj_4633));
    defparam i9_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i22_4_lut (.I0(n37), .I1(n39), .I2(n38), .I3(n40), .O(n46));
    defparam i22_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i9_3_lut (.I0(bit_ctr[7]), .I1(n2802), .I2(n2809), .I3(GND_net), 
            .O(n33));
    defparam i9_3_lut.LUT_INIT = 16'hecec;
    SB_LUT4 i13_4_lut_adj_1479 (.I0(n19), .I1(n26), .I2(n1905), .I3(n1903), 
            .O(n28_adj_4634));
    defparam i13_4_lut_adj_1479.LUT_INIT = 16'hfffe;
    SB_LUT4 i14_4_lut_adj_1480 (.I0(n1896), .I1(n28_adj_4634), .I2(n24_adj_4633), 
            .I3(n16_adj_4632), .O(n1928));
    defparam i14_4_lut_adj_1480.LUT_INIT = 16'hfffe;
    SB_LUT4 i23_4_lut (.I0(n33), .I1(n46), .I2(n42), .I3(n34), .O(n2819));
    defparam i23_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i31563_1_lut (.I0(n2918), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n38243));
    defparam i31563_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i4_3_lut_adj_1481 (.I0(bit_ctr[18]), .I1(n1699), .I2(n1709), 
            .I3(GND_net), .O(n17_adj_4635));
    defparam i4_3_lut_adj_1481.LUT_INIT = 16'hecec;
    SB_LUT4 i8_4_lut (.I0(n1698), .I1(n1707), .I2(n1703), .I3(n1705), 
            .O(n21));
    defparam i8_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 mod_5_add_937_7_lut (.I0(n1305), .I1(n1305), .I2(n1334), .I3(n28766), 
            .O(n1404)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_937_7_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i7_3_lut (.I0(n1704), .I1(n1701), .I2(n1708), .I3(GND_net), 
            .O(n20_c));
    defparam i7_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i11_4_lut_adj_1482 (.I0(n21), .I1(n17_adj_4635), .I2(n1702), 
            .I3(n1697), .O(n24_adj_4636));
    defparam i11_4_lut_adj_1482.LUT_INIT = 16'hfffe;
    SB_LUT4 mod_5_add_2143_15_lut (.I0(n3097), .I1(n3097), .I2(n3116), 
            .I3(n29089), .O(n3196)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_15_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1473_10_lut (.I0(n2102), .I1(n2102), .I2(n2126), 
            .I3(n28869), .O(n2201)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_10_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_937_7 (.CI(n28766), .I0(n1305), .I1(n1334), .CO(n28767));
    SB_LUT4 mod_5_add_937_6_lut (.I0(n1306), .I1(n1306), .I2(n1334), .I3(n28765), 
            .O(n1405)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_937_6_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_937_6 (.CI(n28765), .I0(n1306), .I1(n1334), .CO(n28766));
    SB_LUT4 i12_4_lut_adj_1483 (.I0(n1700), .I1(n24_adj_4636), .I2(n20_c), 
            .I3(n1706), .O(n1730));
    defparam i12_4_lut_adj_1483.LUT_INIT = 16'hfffe;
    SB_LUT4 sub_14_inv_0_i16_1_lut (.I0(\neo_pixel_transmitter.t0 [15]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n51[15]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i16_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i31573_1_lut (.I0(n2324), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n38253));
    defparam i31573_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mod_5_add_937_5_lut (.I0(n1307), .I1(n1307), .I2(n1334), .I3(n28764), 
            .O(n1406)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_937_5_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_937_5 (.CI(n28764), .I0(n1307), .I1(n1334), .CO(n28765));
    SB_LUT4 i31564_1_lut (.I0(n1829), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n38244));
    defparam i31564_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mod_5_add_937_4_lut (.I0(n1308), .I1(n1308), .I2(n1334), .I3(n28763), 
            .O(n1407)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_937_4_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_937_4 (.CI(n28763), .I0(n1308), .I1(n1334), .CO(n28764));
    SB_LUT4 mod_5_add_937_3_lut (.I0(n1309), .I1(n1309), .I2(n38235), 
            .I3(n28762), .O(n1408)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_937_3_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_937_3 (.CI(n28762), .I0(n1309), .I1(n38235), .CO(n28763));
    SB_LUT4 mod_5_add_937_2_lut (.I0(bit_ctr[22]), .I1(bit_ctr[22]), .I2(n38235), 
            .I3(VCC_net), .O(n1409)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_937_2_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_937_2 (.CI(VCC_net), .I0(bit_ctr[22]), .I1(n38235), 
            .CO(n28762));
    SB_LUT4 mod_5_add_870_10_lut (.I0(n1202), .I1(n1202), .I2(n1235), 
            .I3(n28761), .O(n1301)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_870_10_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_870_9_lut (.I0(n1203), .I1(n1203), .I2(n1235), .I3(n28760), 
            .O(n1302)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_870_9_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_870_9 (.CI(n28760), .I0(n1203), .I1(n1235), .CO(n28761));
    SB_CARRY mod_5_add_2143_15 (.CI(n29089), .I0(n3097), .I1(n3116), .CO(n29090));
    SB_LUT4 sub_14_inv_0_i21_1_lut (.I0(\neo_pixel_transmitter.t0 [20]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n51[20]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i21_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mod_5_add_870_8_lut (.I0(n1204), .I1(n1204), .I2(n1235), .I3(n28759), 
            .O(n1303)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_870_8_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_870_8 (.CI(n28759), .I0(n1204), .I1(n1235), .CO(n28760));
    SB_LUT4 mod_5_add_2143_14_lut (.I0(n3098), .I1(n3098), .I2(n3116), 
            .I3(n29088), .O(n3197)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_14_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_870_7_lut (.I0(n1205), .I1(n1205), .I2(n1235), .I3(n28758), 
            .O(n1304)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_870_7_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2143_14 (.CI(n29088), .I0(n3098), .I1(n3116), .CO(n29089));
    SB_LUT4 i31561_1_lut (.I0(n2027), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n38241));
    defparam i31561_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY mod_5_add_1473_10 (.CI(n28869), .I0(n2102), .I1(n2126), .CO(n28870));
    SB_LUT4 sub_14_inv_0_i22_1_lut (.I0(\neo_pixel_transmitter.t0 [21]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n51[21]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i22_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mod_5_add_1473_9_lut (.I0(n2103), .I1(n2103), .I2(n2126), 
            .I3(n28868), .O(n2202)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_9_lut.LUT_INIT = 16'hCA3A;
    SB_DFFE state_i1 (.Q(\state[1] ), .C(clk32MHz), .E(VCC_net), .D(n17567));   // verilog/neopixel.v(35[12] 117[6])
    SB_CARRY mod_5_add_870_7 (.CI(n28758), .I0(n1205), .I1(n1235), .CO(n28759));
    SB_LUT4 mod_5_add_870_6_lut (.I0(n1206), .I1(n1206), .I2(n1235), .I3(n28757), 
            .O(n1305)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_870_6_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_870_6 (.CI(n28757), .I0(n1206), .I1(n1235), .CO(n28758));
    SB_LUT4 i8_4_lut_adj_1484 (.I0(n1608), .I1(n1606), .I2(n1604), .I3(n1603), 
            .O(n20_adj_4638));
    defparam i8_4_lut_adj_1484.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_3_lut_adj_1485 (.I0(bit_ctr[19]), .I1(n1602), .I2(n1609), 
            .I3(GND_net), .O(n13_adj_4639));
    defparam i1_3_lut_adj_1485.LUT_INIT = 16'hecec;
    SB_LUT4 i6_2_lut (.I0(n1598), .I1(n1600), .I2(GND_net), .I3(GND_net), 
            .O(n18_adj_4640));
    defparam i6_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i10_4_lut_adj_1486 (.I0(n13_adj_4639), .I1(n20_adj_4638), .I2(n1605), 
            .I3(n1599), .O(n22_adj_4641));
    defparam i10_4_lut_adj_1486.LUT_INIT = 16'hfffe;
    SB_LUT4 sub_14_inv_0_i7_1_lut (.I0(\neo_pixel_transmitter.t0 [6]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n51[6]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mod_5_add_870_5_lut (.I0(n1207), .I1(n1207), .I2(n1235), .I3(n28756), 
            .O(n1306)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_870_5_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_870_5 (.CI(n28756), .I0(n1207), .I1(n1235), .CO(n28757));
    SB_LUT4 mod_5_add_870_4_lut (.I0(n1208), .I1(n1208), .I2(n1235), .I3(n28755), 
            .O(n1307)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_870_4_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i31550_1_lut (.I0(n2225), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n38230));
    defparam i31550_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mod_5_add_2143_13_lut (.I0(n3099), .I1(n3099), .I2(n3116), 
            .I3(n29087), .O(n3198)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_13_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1473_9 (.CI(n28868), .I0(n2103), .I1(n2126), .CO(n28869));
    SB_CARRY sub_14_add_2_17 (.CI(n27954), .I0(timer[15]), .I1(n51[15]), 
            .CO(n27955));
    SB_CARRY mod_5_add_870_4 (.CI(n28755), .I0(n1208), .I1(n1235), .CO(n28756));
    SB_CARRY mod_5_add_2143_13 (.CI(n29087), .I0(n3099), .I1(n3116), .CO(n29088));
    SB_LUT4 mod_5_add_1473_8_lut (.I0(n2104), .I1(n2104), .I2(n2126), 
            .I3(n28867), .O(n2203)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_8_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_870_3_lut (.I0(n1209), .I1(n1209), .I2(n38236), 
            .I3(n28754), .O(n1308)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_870_3_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_870_3 (.CI(n28754), .I0(n1209), .I1(n38236), .CO(n28755));
    SB_LUT4 mod_5_add_870_2_lut (.I0(bit_ctr[23]), .I1(bit_ctr[23]), .I2(n38236), 
            .I3(VCC_net), .O(n1309)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_870_2_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_870_2 (.CI(VCC_net), .I0(bit_ctr[23]), .I1(n38236), 
            .CO(n28754));
    SB_LUT4 mod_5_add_803_9_lut (.I0(n1103), .I1(n1103), .I2(n1136), .I3(n28753), 
            .O(n1202)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_803_9_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1473_8 (.CI(n28867), .I0(n2104), .I1(n2126), .CO(n28868));
    SB_LUT4 mod_5_add_803_8_lut (.I0(n1104), .I1(n1104), .I2(n1136), .I3(n28752), 
            .O(n1203)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_803_8_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_803_8 (.CI(n28752), .I0(n1104), .I1(n1136), .CO(n28753));
    SB_LUT4 i5_3_lut (.I0(n1308), .I1(n1304), .I2(n1305), .I3(GND_net), 
            .O(n14_adj_4643));
    defparam i5_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i3_2_lut (.I0(n1306), .I1(n1307), .I2(GND_net), .I3(GND_net), 
            .O(n12_adj_4644));
    defparam i3_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 mod_5_add_803_7_lut (.I0(n1105), .I1(n1105), .I2(n1136), .I3(n28751), 
            .O(n1204)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_803_7_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_803_7 (.CI(n28751), .I0(n1105), .I1(n1136), .CO(n28752));
    SB_LUT4 mod_5_add_803_6_lut (.I0(n1106), .I1(n1106), .I2(n1136), .I3(n28750), 
            .O(n1205)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_803_6_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i7_4_lut_adj_1487 (.I0(n1303), .I1(n14_adj_4643), .I2(bit_ctr[22]), 
            .I3(n1309), .O(n16_adj_4645));
    defparam i7_4_lut_adj_1487.LUT_INIT = 16'hfeee;
    SB_LUT4 i8_4_lut_adj_1488 (.I0(n1301), .I1(n16_adj_4645), .I2(n12_adj_4644), 
            .I3(n1302), .O(n1334));
    defparam i8_4_lut_adj_1488.LUT_INIT = 16'hfffe;
    SB_LUT4 sub_14_inv_0_i19_1_lut (.I0(\neo_pixel_transmitter.t0 [18]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n51[18]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i19_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mod_5_add_2143_12_lut (.I0(n3100), .I1(n3100), .I2(n3116), 
            .I3(n29086), .O(n3199)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_12_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_803_6 (.CI(n28750), .I0(n1106), .I1(n1136), .CO(n28751));
    SB_CARRY mod_5_add_2143_12 (.CI(n29086), .I0(n3100), .I1(n3116), .CO(n29087));
    SB_LUT4 sub_14_inv_0_i23_1_lut (.I0(\neo_pixel_transmitter.t0 [22]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n51[22]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i23_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i11_4_lut_adj_1489 (.I0(n1601), .I1(n22_adj_4641), .I2(n18_adj_4640), 
            .I3(n1607), .O(n1631));
    defparam i11_4_lut_adj_1489.LUT_INIT = 16'hfffe;
    SB_LUT4 mod_5_add_803_5_lut (.I0(n1107), .I1(n1107), .I2(n1136), .I3(n28749), 
            .O(n1206)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_803_5_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_803_5 (.CI(n28749), .I0(n1107), .I1(n1136), .CO(n28750));
    SB_LUT4 mod_5_add_803_4_lut (.I0(n1108), .I1(n1108), .I2(n1136), .I3(n28748), 
            .O(n1207)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_803_4_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1473_7_lut (.I0(n2105), .I1(n2105), .I2(n2126), 
            .I3(n28866), .O(n2204)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_7_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_803_4 (.CI(n28748), .I0(n1108), .I1(n1136), .CO(n28749));
    SB_LUT4 mod_5_add_803_3_lut (.I0(n1109), .I1(n1109), .I2(n38237), 
            .I3(n28747), .O(n1208)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_803_3_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_803_3 (.CI(n28747), .I0(n1109), .I1(n38237), .CO(n28748));
    SB_LUT4 mod_5_add_803_2_lut (.I0(bit_ctr[24]), .I1(bit_ctr[24]), .I2(n38237), 
            .I3(VCC_net), .O(n1209)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_803_2_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_803_2 (.CI(VCC_net), .I0(bit_ctr[24]), .I1(n38237), 
            .CO(n28747));
    SB_LUT4 sub_14_inv_0_i8_1_lut (.I0(\neo_pixel_transmitter.t0 [7]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n51[7]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i8_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY mod_5_add_1473_7 (.CI(n28866), .I0(n2105), .I1(n2126), .CO(n28867));
    SB_LUT4 mod_5_add_736_8_lut (.I0(n4_adj_4647), .I1(n4_adj_4647), .I2(n1037), 
            .I3(n28746), .O(n1103)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_736_8_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_736_7_lut (.I0(n1005), .I1(n1005), .I2(n1037), .I3(n28745), 
            .O(n1104)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_736_7_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1473_6_lut (.I0(n2106), .I1(n2106), .I2(n2126), 
            .I3(n28865), .O(n2205)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_6_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_2143_11_lut (.I0(n3101), .I1(n3101), .I2(n3116), 
            .I3(n29085), .O(n3200)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_11_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2143_11 (.CI(n29085), .I0(n3101), .I1(n3116), .CO(n29086));
    SB_CARRY mod_5_add_736_7 (.CI(n28745), .I0(n1005), .I1(n1037), .CO(n28746));
    SB_LUT4 mod_5_add_736_6_lut (.I0(n1006), .I1(n1006), .I2(n1037), .I3(n28744), 
            .O(n1105)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_736_6_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 sub_14_inv_0_i9_1_lut (.I0(\neo_pixel_transmitter.t0 [8]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n51[8]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i9_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mod_5_add_2143_10_lut (.I0(n3102), .I1(n3102), .I2(n3116), 
            .I3(n29084), .O(n3201)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_10_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2143_10 (.CI(n29084), .I0(n3102), .I1(n3116), .CO(n29085));
    SB_LUT4 mod_5_add_2143_9_lut (.I0(n3103), .I1(n3103), .I2(n3116), 
            .I3(n29083), .O(n3202)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_9_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2143_9 (.CI(n29083), .I0(n3103), .I1(n3116), .CO(n29084));
    SB_CARRY mod_5_add_1473_6 (.CI(n28865), .I0(n2106), .I1(n2126), .CO(n28866));
    SB_LUT4 sub_14_add_2_16_lut (.I0(one_wire_N_613[19]), .I1(timer[14]), 
            .I2(n51[14]), .I3(n27953), .O(n25_adj_4648)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_16_lut.LUT_INIT = 16'hebbe;
    SB_CARRY mod_5_add_736_6 (.CI(n28744), .I0(n1006), .I1(n1037), .CO(n28745));
    SB_LUT4 mod_5_add_736_5_lut (.I0(n1007), .I1(n1007), .I2(n1037), .I3(n28743), 
            .O(n1106)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_736_5_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1473_5_lut (.I0(n2107), .I1(n2107), .I2(n2126), 
            .I3(n28864), .O(n2206)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_5_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_2143_8_lut (.I0(n3104), .I1(n3104), .I2(n3116), 
            .I3(n29082), .O(n3203)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_8_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2143_8 (.CI(n29082), .I0(n3104), .I1(n3116), .CO(n29083));
    SB_CARRY mod_5_add_736_5 (.CI(n28743), .I0(n1007), .I1(n1037), .CO(n28744));
    SB_CARRY sub_14_add_2_16 (.CI(n27953), .I0(timer[14]), .I1(n51[14]), 
            .CO(n27954));
    SB_LUT4 mod_5_add_2143_7_lut (.I0(n3105), .I1(n3105), .I2(n3116), 
            .I3(n29081), .O(n3204)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_7_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1473_5 (.CI(n28864), .I0(n2107), .I1(n2126), .CO(n28865));
    SB_CARRY mod_5_add_2143_7 (.CI(n29081), .I0(n3105), .I1(n3116), .CO(n29082));
    SB_LUT4 mod_5_add_736_4_lut (.I0(n1008), .I1(n1008), .I2(n1037), .I3(n28742), 
            .O(n1107)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_736_4_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_736_4 (.CI(n28742), .I0(n1008), .I1(n1037), .CO(n28743));
    SB_LUT4 mod_5_add_736_3_lut (.I0(n1009), .I1(n1009), .I2(n38239), 
            .I3(n28741), .O(n1108)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_736_3_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_736_3 (.CI(n28741), .I0(n1009), .I1(n38239), .CO(n28742));
    SB_LUT4 mod_5_add_736_2_lut (.I0(bit_ctr[25]), .I1(bit_ctr[25]), .I2(n38239), 
            .I3(VCC_net), .O(n1109)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_736_2_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_736_2 (.CI(VCC_net), .I0(bit_ctr[25]), .I1(n38239), 
            .CO(n28741));
    SB_LUT4 mod_5_add_669_7_lut (.I0(GND_net), .I1(n905), .I2(VCC_net), 
            .I3(n28740), .O(n971[31])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_669_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_14_inv_0_i10_1_lut (.I0(\neo_pixel_transmitter.t0 [9]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n51[9]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i10_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mod_5_add_2143_6_lut (.I0(n3106), .I1(n3106), .I2(n3116), 
            .I3(n29080), .O(n3205)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_6_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2143_6 (.CI(n29080), .I0(n3106), .I1(n3116), .CO(n29081));
    SB_LUT4 mod_5_add_2143_5_lut (.I0(n3107), .I1(n3107), .I2(n3116), 
            .I3(n29079), .O(n3206)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_5_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1473_4_lut (.I0(n2108), .I1(n2108), .I2(n2126), 
            .I3(n28863), .O(n2207)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_4_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2143_5 (.CI(n29079), .I0(n3107), .I1(n3116), .CO(n29080));
    SB_CARRY mod_5_add_1473_4 (.CI(n28863), .I0(n2108), .I1(n2126), .CO(n28864));
    SB_LUT4 mod_5_add_2143_4_lut (.I0(n3108), .I1(n3108), .I2(n3116), 
            .I3(n29078), .O(n3207)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_4_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1473_3_lut (.I0(n2109), .I1(n2109), .I2(n38234), 
            .I3(n28862), .O(n2208)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_3_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_2143_4 (.CI(n29078), .I0(n3108), .I1(n3116), .CO(n29079));
    SB_LUT4 mod_5_add_2143_3_lut (.I0(n3109), .I1(n3109), .I2(n38233), 
            .I3(n29077), .O(n3208)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_3_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 mod_5_add_669_6_lut (.I0(GND_net), .I1(n906), .I2(VCC_net), 
            .I3(n28739), .O(n971[30])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_669_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_2143_3 (.CI(n29077), .I0(n3109), .I1(n38233), .CO(n29078));
    SB_LUT4 mod_5_add_2143_2_lut (.I0(bit_ctr[4]), .I1(bit_ctr[4]), .I2(n38233), 
            .I3(VCC_net), .O(n3209)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_2_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1473_3 (.CI(n28862), .I0(n2109), .I1(n38234), .CO(n28863));
    SB_CARRY mod_5_add_669_6 (.CI(n28739), .I0(n906), .I1(VCC_net), .CO(n28740));
    SB_LUT4 mod_5_add_669_5_lut (.I0(GND_net), .I1(n33675), .I2(VCC_net), 
            .I3(n28738), .O(n971[29])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_669_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_2143_2 (.CI(VCC_net), .I0(bit_ctr[4]), .I1(n38233), 
            .CO(n29077));
    SB_LUT4 mod_5_add_1473_2_lut (.I0(bit_ctr[14]), .I1(bit_ctr[14]), .I2(n38234), 
            .I3(VCC_net), .O(n2209)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_2_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_669_5 (.CI(n28738), .I0(n33675), .I1(VCC_net), 
            .CO(n28739));
    SB_LUT4 mod_5_add_2076_28_lut (.I0(n2984), .I1(n2984), .I2(n3017), 
            .I3(n29076), .O(n3083)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_28_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_669_4_lut (.I0(GND_net), .I1(n17391), .I2(VCC_net), 
            .I3(n28737), .O(n971[28])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_669_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_14_inv_0_i11_1_lut (.I0(\neo_pixel_transmitter.t0 [10]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n51[10]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i11_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i12_1_lut (.I0(\neo_pixel_transmitter.t0 [11]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n51[11]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i12_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i3_2_lut_adj_1490 (.I0(n2302), .I1(n2292), .I2(GND_net), .I3(GND_net), 
            .O(n22_adj_4652));
    defparam i3_2_lut_adj_1490.LUT_INIT = 16'heeee;
    SB_CARRY mod_5_add_669_4 (.CI(n28737), .I0(n17391), .I1(VCC_net), 
            .CO(n28738));
    SB_LUT4 i11_4_lut_adj_1491 (.I0(bit_ctr[12]), .I1(n22_adj_4652), .I2(n2299), 
            .I3(n2309), .O(n30_adj_4653));
    defparam i11_4_lut_adj_1491.LUT_INIT = 16'hfefc;
    SB_LUT4 mod_5_add_669_3_lut (.I0(GND_net), .I1(n14852), .I2(GND_net), 
            .I3(n28736), .O(n971[27])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_669_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i15_4_lut_adj_1492 (.I0(n2294), .I1(n30_adj_4653), .I2(n2306), 
            .I3(n2297), .O(n34_adj_4654));
    defparam i15_4_lut_adj_1492.LUT_INIT = 16'hfffe;
    SB_LUT4 i13_4_lut_adj_1493 (.I0(n2301), .I1(n2307), .I2(n2291), .I3(n2305), 
            .O(n32));
    defparam i13_4_lut_adj_1493.LUT_INIT = 16'hfffe;
    SB_CARRY mod_5_add_1473_2 (.CI(VCC_net), .I0(bit_ctr[14]), .I1(n38234), 
            .CO(n28862));
    SB_LUT4 mod_5_add_2076_27_lut (.I0(n2985), .I1(n2985), .I2(n3017), 
            .I3(n29075), .O(n3084)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_27_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i14_4_lut_adj_1494 (.I0(n2298), .I1(n2295), .I2(n2304), .I3(n2300), 
            .O(n33_adj_4655));
    defparam i14_4_lut_adj_1494.LUT_INIT = 16'hfffe;
    SB_CARRY mod_5_add_669_3 (.CI(n28736), .I0(n14852), .I1(GND_net), 
            .CO(n28737));
    SB_CARRY mod_5_add_2076_27 (.CI(n29075), .I0(n2985), .I1(n3017), .CO(n29076));
    SB_LUT4 mod_5_add_2076_26_lut (.I0(n2986), .I1(n2986), .I2(n3017), 
            .I3(n29074), .O(n3085)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_26_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i12_4_lut_adj_1495 (.I0(n2308), .I1(n2296), .I2(n2303), .I3(n2293), 
            .O(n31));
    defparam i12_4_lut_adj_1495.LUT_INIT = 16'hfffe;
    SB_LUT4 mod_5_add_1406_18_lut (.I0(n1994), .I1(n1994), .I2(n2027), 
            .I3(n28861), .O(n2093)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_18_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i18_4_lut_adj_1496 (.I0(n31), .I1(n33_adj_4655), .I2(n32), 
            .I3(n34_adj_4654), .O(n2324));
    defparam i18_4_lut_adj_1496.LUT_INIT = 16'hfffe;
    SB_LUT4 mod_5_add_669_2_lut (.I0(GND_net), .I1(bit_ctr[26]), .I2(GND_net), 
            .I3(VCC_net), .O(n971[26])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_669_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_669_2 (.CI(VCC_net), .I0(bit_ctr[26]), .I1(GND_net), 
            .CO(n28736));
    SB_LUT4 mod_5_add_1406_17_lut (.I0(n1995), .I1(n1995), .I2(n2027), 
            .I3(n28860), .O(n2094)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_17_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1406_17 (.CI(n28860), .I0(n1995), .I1(n2027), .CO(n28861));
    SB_LUT4 mod_5_add_1406_16_lut (.I0(n1996), .I1(n1996), .I2(n2027), 
            .I3(n28859), .O(n2095)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_16_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1406_16 (.CI(n28859), .I0(n1996), .I1(n2027), .CO(n28860));
    SB_CARRY mod_5_add_2076_26 (.CI(n29074), .I0(n2986), .I1(n3017), .CO(n29075));
    SB_LUT4 mod_5_add_2076_25_lut (.I0(n2987), .I1(n2987), .I2(n3017), 
            .I3(n29073), .O(n3086)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_25_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1406_15_lut (.I0(n1997), .I1(n1997), .I2(n2027), 
            .I3(n28858), .O(n2096)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_15_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 sub_14_inv_0_i13_1_lut (.I0(\neo_pixel_transmitter.t0 [12]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n51[12]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i13_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY mod_5_add_1406_15 (.CI(n28858), .I0(n1997), .I1(n2027), .CO(n28859));
    SB_LUT4 sub_14_add_2_15_lut (.I0(one_wire_N_613[20]), .I1(timer[13]), 
            .I2(n51[13]), .I3(n27952), .O(n23_adj_4657)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_15_lut.LUT_INIT = 16'hebbe;
    SB_CARRY mod_5_add_2076_25 (.CI(n29073), .I0(n2987), .I1(n3017), .CO(n29074));
    SB_LUT4 mod_5_add_1406_14_lut (.I0(n1998), .I1(n1998), .I2(n2027), 
            .I3(n28857), .O(n2097)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_14_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_2076_24_lut (.I0(n2988), .I1(n2988), .I2(n3017), 
            .I3(n29072), .O(n3087)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_24_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2076_24 (.CI(n29072), .I0(n2988), .I1(n3017), .CO(n29073));
    SB_LUT4 i1_2_lut_adj_1497 (.I0(one_wire_N_613[10]), .I1(one_wire_N_613[11]), 
            .I2(GND_net), .I3(GND_net), .O(n6));   // verilog/neopixel.v(104[14:39])
    defparam i1_2_lut_adj_1497.LUT_INIT = 16'heeee;
    SB_LUT4 sub_14_inv_0_i14_1_lut (.I0(\neo_pixel_transmitter.t0 [13]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n51[13]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i14_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY mod_5_add_1406_14 (.CI(n28857), .I0(n1998), .I1(n2027), .CO(n28858));
    SB_LUT4 mod_5_add_2076_23_lut (.I0(n2989), .I1(n2989), .I2(n3017), 
            .I3(n29071), .O(n3088)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_23_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2076_23 (.CI(n29071), .I0(n2989), .I1(n3017), .CO(n29072));
    SB_LUT4 mod_5_add_2076_22_lut (.I0(n2990), .I1(n2990), .I2(n3017), 
            .I3(n29070), .O(n3089)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_22_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1406_13_lut (.I0(n1999), .I1(n1999), .I2(n2027), 
            .I3(n28856), .O(n2098)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_13_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY sub_14_add_2_15 (.CI(n27952), .I0(timer[13]), .I1(n51[13]), 
            .CO(n27953));
    SB_LUT4 sub_14_add_2_14_lut (.I0(one_wire_N_613[25]), .I1(timer[12]), 
            .I2(n51[12]), .I3(n27951), .O(n27_adj_4659)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_14_lut.LUT_INIT = 16'hebbe;
    SB_CARRY mod_5_add_2076_22 (.CI(n29070), .I0(n2990), .I1(n3017), .CO(n29071));
    SB_LUT4 mod_5_add_2076_21_lut (.I0(n2991), .I1(n2991), .I2(n3017), 
            .I3(n29069), .O(n3090)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_21_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2076_21 (.CI(n29069), .I0(n2991), .I1(n3017), .CO(n29070));
    SB_CARRY mod_5_add_1406_13 (.CI(n28856), .I0(n1999), .I1(n2027), .CO(n28857));
    SB_LUT4 mod_5_add_1406_12_lut (.I0(n2000), .I1(n2000), .I2(n2027), 
            .I3(n28855), .O(n2099)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_12_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1406_12 (.CI(n28855), .I0(n2000), .I1(n2027), .CO(n28856));
    SB_LUT4 mod_5_add_1406_11_lut (.I0(n2001), .I1(n2001), .I2(n2027), 
            .I3(n28854), .O(n2100)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_11_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_2076_20_lut (.I0(n2992), .I1(n2992), .I2(n3017), 
            .I3(n29068), .O(n3091)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_20_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2076_20 (.CI(n29068), .I0(n2992), .I1(n3017), .CO(n29069));
    SB_CARRY mod_5_add_1406_11 (.CI(n28854), .I0(n2001), .I1(n2027), .CO(n28855));
    SB_CARRY sub_14_add_2_14 (.CI(n27951), .I0(timer[12]), .I1(n51[12]), 
            .CO(n27952));
    SB_LUT4 mod_5_add_1406_10_lut (.I0(n2002), .I1(n2002), .I2(n2027), 
            .I3(n28853), .O(n2101)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_10_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 sub_14_add_2_13_lut (.I0(GND_net), .I1(timer[11]), .I2(n51[11]), 
            .I3(n27950), .O(one_wire_N_613[11])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_14_add_2_13 (.CI(n27950), .I0(timer[11]), .I1(n51[11]), 
            .CO(n27951));
    SB_LUT4 sub_14_add_2_12_lut (.I0(GND_net), .I1(timer[10]), .I2(n51[10]), 
            .I3(n27949), .O(one_wire_N_613[10])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i30948_3_lut_4_lut_3_lut (.I0(n708), .I1(n30176), .I2(bit_ctr[28]), 
            .I3(GND_net), .O(n33673));   // verilog/neopixel.v(22[26:36])
    defparam i30948_3_lut_4_lut_3_lut.LUT_INIT = 16'h2c2c;
    SB_CARRY sub_14_add_2_12 (.CI(n27949), .I0(timer[10]), .I1(n51[10]), 
            .CO(n27950));
    SB_CARRY mod_5_add_1406_10 (.CI(n28853), .I0(n2002), .I1(n2027), .CO(n28854));
    SB_LUT4 mod_5_add_2076_19_lut (.I0(n2993), .I1(n2993), .I2(n3017), 
            .I3(n29067), .O(n3092)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_19_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2076_19 (.CI(n29067), .I0(n2993), .I1(n3017), .CO(n29068));
    SB_LUT4 mod_5_add_2076_18_lut (.I0(n2994), .I1(n2994), .I2(n3017), 
            .I3(n29066), .O(n3093)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_18_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i12_3_lut_4_lut_3_lut (.I0(bit_ctr[30]), .I1(bit_ctr[31]), .I2(bit_ctr[29]), 
            .I3(GND_net), .O(n708));   // verilog/neopixel.v(22[26:36])
    defparam i12_3_lut_4_lut_3_lut.LUT_INIT = 16'h4242;
    SB_CARRY mod_5_add_2076_18 (.CI(n29066), .I0(n2994), .I1(n3017), .CO(n29067));
    SB_LUT4 i1_3_lut_3_lut_4_lut_3_lut (.I0(bit_ctr[30]), .I1(bit_ctr[31]), 
            .I2(bit_ctr[29]), .I3(GND_net), .O(n30176));   // verilog/neopixel.v(22[26:36])
    defparam i1_3_lut_3_lut_4_lut_3_lut.LUT_INIT = 16'h9494;
    SB_LUT4 mod_5_add_2076_17_lut (.I0(n2995), .I1(n2995), .I2(n3017), 
            .I3(n29065), .O(n3094)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_17_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2076_17 (.CI(n29065), .I0(n2995), .I1(n3017), .CO(n29066));
    SB_LUT4 mod_5_add_1406_9_lut (.I0(n2003), .I1(n2003), .I2(n2027), 
            .I3(n28852), .O(n2102)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_9_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1406_9 (.CI(n28852), .I0(n2003), .I1(n2027), .CO(n28853));
    SB_LUT4 mod_5_add_1406_8_lut (.I0(n2004), .I1(n2004), .I2(n2027), 
            .I3(n28851), .O(n2103)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_8_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_2076_16_lut (.I0(n2996), .I1(n2996), .I2(n3017), 
            .I3(n29064), .O(n3095)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_16_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY add_21_13 (.CI(n27854), .I0(bit_ctr[11]), .I1(GND_net), .CO(n27855));
    SB_CARRY mod_5_add_1406_8 (.CI(n28851), .I0(n2004), .I1(n2027), .CO(n28852));
    SB_LUT4 mod_5_add_1406_7_lut (.I0(n2005), .I1(n2005), .I2(n2027), 
            .I3(n28850), .O(n2104)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_7_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i9_3_lut_adj_1498 (.I0(bit_ctr[4]), .I1(n3107), .I2(n3109), 
            .I3(GND_net), .O(n36));
    defparam i9_3_lut_adj_1498.LUT_INIT = 16'hecec;
    SB_LUT4 i19_4_lut (.I0(n3086), .I1(n3102), .I2(n3094), .I3(n3106), 
            .O(n46_adj_4660));
    defparam i19_4_lut.LUT_INIT = 16'hfffe;
    SB_CARRY mod_5_add_1406_7 (.CI(n28850), .I0(n2005), .I1(n2027), .CO(n28851));
    SB_LUT4 i16_4_lut_adj_1499 (.I0(n21_adj_4661), .I1(n23_adj_4657), .I2(n22), 
            .I3(n24), .O(n36_adj_4662));   // verilog/neopixel.v(104[14:39])
    defparam i16_4_lut_adj_1499.LUT_INIT = 16'hfffe;
    SB_LUT4 mod_5_add_1406_6_lut (.I0(n2006), .I1(n2006), .I2(n2027), 
            .I3(n28849), .O(n2105)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_6_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2076_16 (.CI(n29064), .I0(n2996), .I1(n3017), .CO(n29065));
    SB_CARRY mod_5_add_1406_6 (.CI(n28849), .I0(n2006), .I1(n2027), .CO(n28850));
    SB_LUT4 mod_5_add_2076_15_lut (.I0(n2997), .I1(n2997), .I2(n3017), 
            .I3(n29063), .O(n3096)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_15_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1406_5_lut (.I0(n2007), .I1(n2007), .I2(n2027), 
            .I3(n28848), .O(n2106)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_5_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i3559_2_lut_3_lut (.I0(n14844), .I1(bit_ctr[27]), .I2(n33673), 
            .I3(GND_net), .O(n60));   // verilog/neopixel.v(22[26:36])
    defparam i3559_2_lut_3_lut.LUT_INIT = 16'hf4f4;
    SB_LUT4 mod_5_i606_3_lut_4_lut (.I0(n14844), .I1(bit_ctr[27]), .I2(n838), 
            .I3(n33673), .O(n33675));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i606_3_lut_4_lut.LUT_INIT = 16'hf40b;
    SB_LUT4 i31572_1_lut (.I0(n2423), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n38252));
    defparam i31572_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY mod_5_add_2076_15 (.CI(n29063), .I0(n2997), .I1(n3017), .CO(n29064));
    SB_LUT4 sub_14_add_2_11_lut (.I0(GND_net), .I1(timer[9]), .I2(n51[9]), 
            .I3(n27948), .O(one_wire_N_613[9])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_14_add_2_11 (.CI(n27948), .I0(timer[9]), .I1(n51[9]), 
            .CO(n27949));
    SB_LUT4 sub_14_add_2_10_lut (.I0(one_wire_N_613[9]), .I1(timer[8]), 
            .I2(n51[8]), .I3(n27947), .O(n6_adj_4663)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_10_lut.LUT_INIT = 16'hebbe;
    SB_LUT4 mod_5_add_2076_14_lut (.I0(n2998), .I1(n2998), .I2(n3017), 
            .I3(n29062), .O(n3097)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_14_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2076_14 (.CI(n29062), .I0(n2998), .I1(n3017), .CO(n29063));
    SB_CARRY sub_14_add_2_10 (.CI(n27947), .I0(timer[8]), .I1(n51[8]), 
            .CO(n27948));
    SB_LUT4 mod_5_add_2076_13_lut (.I0(n2999), .I1(n2999), .I2(n3017), 
            .I3(n29061), .O(n3098)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_13_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 sub_14_add_2_9_lut (.I0(one_wire_N_613[6]), .I1(timer[7]), .I2(n51[7]), 
            .I3(n27946), .O(n7_adj_4664)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_9_lut.LUT_INIT = 16'hebbe;
    SB_CARRY sub_14_add_2_9 (.CI(n27946), .I0(timer[7]), .I1(n51[7]), 
            .CO(n27947));
    SB_CARRY mod_5_add_2076_13 (.CI(n29061), .I0(n2999), .I1(n3017), .CO(n29062));
    SB_LUT4 sub_14_add_2_8_lut (.I0(GND_net), .I1(timer[6]), .I2(n51[6]), 
            .I3(n27945), .O(one_wire_N_613[6])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_2076_12_lut (.I0(n3000), .I1(n3000), .I2(n3017), 
            .I3(n29060), .O(n3099)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_12_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i15_4_lut_adj_1500 (.I0(n3095), .I1(n3089), .I2(n3092), .I3(n3096), 
            .O(n42_adj_4665));
    defparam i15_4_lut_adj_1500.LUT_INIT = 16'hfffe;
    SB_CARRY mod_5_add_1406_5 (.CI(n28848), .I0(n2007), .I1(n2027), .CO(n28849));
    SB_LUT4 mod_5_add_1406_4_lut (.I0(n2008), .I1(n2008), .I2(n2027), 
            .I3(n28847), .O(n2107)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_4_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1406_4 (.CI(n28847), .I0(n2008), .I1(n2027), .CO(n28848));
    SB_CARRY mod_5_add_2076_12 (.CI(n29060), .I0(n3000), .I1(n3017), .CO(n29061));
    SB_LUT4 add_21_33_lut (.I0(n1), .I1(bit_ctr[31]), .I2(GND_net), .I3(n27874), 
            .O(n37244)) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_33_lut.LUT_INIT = 16'h8228;
    SB_LUT4 mod_5_add_2076_11_lut (.I0(n3001), .I1(n3001), .I2(n3017), 
            .I3(n29059), .O(n3100)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_11_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2076_11 (.CI(n29059), .I0(n3001), .I1(n3017), .CO(n29060));
    SB_LUT4 mod_5_add_2076_10_lut (.I0(n3002), .I1(n3002), .I2(n3017), 
            .I3(n29058), .O(n3101)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_10_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 sub_14_inv_0_i1_1_lut (.I0(\neo_pixel_transmitter.t0 [0]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n51[0]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i1_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i20190_2_lut (.I0(bit_ctr[17]), .I1(n1809), .I2(GND_net), 
            .I3(GND_net), .O(n25012));
    defparam i20190_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i4_2_lut (.I0(n1807), .I1(n1801), .I2(GND_net), .I3(GND_net), 
            .O(n18_adj_4667));
    defparam i4_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i5_2_lut (.I0(n3085), .I1(n3083), .I2(GND_net), .I3(GND_net), 
            .O(n32_adj_4668));
    defparam i5_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i17_4_lut (.I0(n3091), .I1(n3108), .I2(n3105), .I3(n3101), 
            .O(n44));
    defparam i17_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i23_4_lut_adj_1501 (.I0(n3099), .I1(n46_adj_4660), .I2(n36), 
            .I3(n3100), .O(n50));
    defparam i23_4_lut_adj_1501.LUT_INIT = 16'hfffe;
    SB_LUT4 i21_4_lut (.I0(n3090), .I1(n42_adj_4665), .I2(n3098), .I3(n3093), 
            .O(n48));
    defparam i21_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i22_4_lut_adj_1502 (.I0(n3097), .I1(n44), .I2(n32_adj_4668), 
            .I3(n3084), .O(n49));
    defparam i22_4_lut_adj_1502.LUT_INIT = 16'hfffe;
    SB_LUT4 mod_5_add_1406_3_lut (.I0(n2009), .I1(n2009), .I2(n38241), 
            .I3(n28846), .O(n2108)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_3_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1406_3 (.CI(n28846), .I0(n2009), .I1(n38241), .CO(n28847));
    SB_LUT4 i10_4_lut_adj_1503 (.I0(n1802), .I1(n1798), .I2(n1808), .I3(n1804), 
            .O(n24_adj_4669));
    defparam i10_4_lut_adj_1503.LUT_INIT = 16'hfffe;
    SB_LUT4 i8_4_lut_adj_1504 (.I0(n1800), .I1(n1803), .I2(n25012), .I3(n1805), 
            .O(n22_adj_4670));
    defparam i8_4_lut_adj_1504.LUT_INIT = 16'hfffe;
    SB_LUT4 i12_4_lut_adj_1505 (.I0(n1797), .I1(n24_adj_4669), .I2(n18_adj_4667), 
            .I3(n1806), .O(n26_adj_4671));
    defparam i12_4_lut_adj_1505.LUT_INIT = 16'hfffe;
    SB_LUT4 i13_4_lut_adj_1506 (.I0(n1796), .I1(n26_adj_4671), .I2(n22_adj_4670), 
            .I3(n1799), .O(n1829));
    defparam i13_4_lut_adj_1506.LUT_INIT = 16'hfffe;
    SB_LUT4 mod_5_add_1406_2_lut (.I0(bit_ctr[15]), .I1(bit_ctr[15]), .I2(n38241), 
            .I3(VCC_net), .O(n2109)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_2_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1406_2 (.CI(VCC_net), .I0(bit_ctr[15]), .I1(n38241), 
            .CO(n28846));
    SB_LUT4 i17_4_lut_adj_1507 (.I0(n25_adj_4648), .I1(n27_adj_4659), .I2(n26_adj_4672), 
            .I3(n28_adj_4673), .O(n37_adj_4674));   // verilog/neopixel.v(104[14:39])
    defparam i17_4_lut_adj_1507.LUT_INIT = 16'hfffe;
    SB_LUT4 i19_4_lut_adj_1508 (.I0(n37_adj_4674), .I1(n29_adj_4675), .I2(n36_adj_4662), 
            .I3(n30), .O(n16103));   // verilog/neopixel.v(104[14:39])
    defparam i19_4_lut_adj_1508.LUT_INIT = 16'hfffe;
    SB_CARRY mod_5_add_2076_10 (.CI(n29058), .I0(n3002), .I1(n3017), .CO(n29059));
    SB_LUT4 i4_2_lut_adj_1509 (.I0(n7_adj_4664), .I1(n8), .I2(GND_net), 
            .I3(GND_net), .O(n7_adj_4676));   // verilog/neopixel.v(104[14:39])
    defparam i4_2_lut_adj_1509.LUT_INIT = 16'heeee;
    SB_LUT4 mod_5_add_1339_17_lut (.I0(n1895), .I1(n1895), .I2(n1928), 
            .I3(n28845), .O(n1994)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_17_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY sub_14_add_2_8 (.CI(n27945), .I0(timer[6]), .I1(n51[6]), 
            .CO(n27946));
    SB_LUT4 i20_4_lut (.I0(n3104), .I1(n3088), .I2(n3087), .I3(n3103), 
            .O(n47));
    defparam i20_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 mod_5_add_2076_9_lut (.I0(n3003), .I1(n3003), .I2(n3017), 
            .I3(n29057), .O(n3102)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_9_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i26_4_lut (.I0(n47), .I1(n49), .I2(n48), .I3(n50), .O(n3116));
    defparam i26_4_lut.LUT_INIT = 16'hfffe;
    SB_CARRY mod_5_add_2076_9 (.CI(n29057), .I0(n3003), .I1(n3017), .CO(n29058));
    SB_LUT4 mod_5_add_1339_16_lut (.I0(n1896), .I1(n1896), .I2(n1928), 
            .I3(n28844), .O(n1995)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_16_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_2076_8_lut (.I0(n3004), .I1(n3004), .I2(n3017), 
            .I3(n29056), .O(n3103)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_8_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1339_16 (.CI(n28844), .I0(n1896), .I1(n1928), .CO(n28845));
    SB_LUT4 i31562_1_lut (.I0(n1928), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n38242));
    defparam i31562_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mod_5_add_1339_15_lut (.I0(n1897), .I1(n1897), .I2(n1928), 
            .I3(n28843), .O(n1996)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_15_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2076_8 (.CI(n29056), .I0(n3004), .I1(n3017), .CO(n29057));
    SB_DFF timer_1524__i0 (.Q(timer[0]), .C(clk32MHz), .D(n133[0]));   // verilog/neopixel.v(12[12:21])
    SB_LUT4 i31551_1_lut (.I0(n1433), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n38231));
    defparam i31551_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i2_2_lut (.I0(bit_ctr[12]), .I1(bit_ctr[29]), .I2(GND_net), 
            .I3(GND_net), .O(n30_adj_4677));
    defparam i2_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i20_4_lut_adj_1510 (.I0(bit_ctr[8]), .I1(bit_ctr[9]), .I2(bit_ctr[27]), 
            .I3(bit_ctr[28]), .O(n48_adj_4678));
    defparam i20_4_lut_adj_1510.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_3_lut_adj_1511 (.I0(n34639), .I1(n7_adj_4676), .I2(one_wire_N_613[3]), 
            .I3(GND_net), .O(n4_adj_4679));
    defparam i1_3_lut_adj_1511.LUT_INIT = 16'hecec;
    SB_LUT4 i18_4_lut_adj_1512 (.I0(bit_ctr[18]), .I1(bit_ctr[15]), .I2(bit_ctr[13]), 
            .I3(bit_ctr[22]), .O(n46_adj_4680));
    defparam i18_4_lut_adj_1512.LUT_INIT = 16'hfffe;
    SB_LUT4 i19_4_lut_adj_1513 (.I0(bit_ctr[25]), .I1(bit_ctr[26]), .I2(bit_ctr[19]), 
            .I3(bit_ctr[14]), .O(n47_adj_4681));
    defparam i19_4_lut_adj_1513.LUT_INIT = 16'hfffe;
    SB_LUT4 i17_4_lut_adj_1514 (.I0(bit_ctr[6]), .I1(bit_ctr[10]), .I2(bit_ctr[30]), 
            .I3(bit_ctr[23]), .O(n45));
    defparam i17_4_lut_adj_1514.LUT_INIT = 16'hfffe;
    SB_LUT4 mod_5_add_2076_7_lut (.I0(n3005), .I1(n3005), .I2(n3017), 
            .I3(n29055), .O(n3104)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_7_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1339_15 (.CI(n28843), .I0(n1897), .I1(n1928), .CO(n28844));
    SB_LUT4 add_21_32_lut (.I0(n1), .I1(bit_ctr[30]), .I2(GND_net), .I3(n27873), 
            .O(n37260)) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_32_lut.LUT_INIT = 16'h8228;
    SB_LUT4 sub_14_add_2_7_lut (.I0(n6_adj_4663), .I1(timer[5]), .I2(n51[5]), 
            .I3(n27944), .O(n8)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_7_lut.LUT_INIT = 16'hebbe;
    SB_LUT4 i27110_4_lut (.I0(n16103), .I1(n6), .I2(one_wire_N_613[4]), 
            .I3(n4_adj_4679), .O(n21937));
    defparam i27110_4_lut.LUT_INIT = 16'hfffe;
    SB_CARRY mod_5_add_2076_7 (.CI(n29055), .I0(n3005), .I1(n3017), .CO(n29056));
    SB_LUT4 mod_5_add_2076_6_lut (.I0(n3006), .I1(n3006), .I2(n3017), 
            .I3(n29054), .O(n3105)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_6_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i2_3_lut (.I0(one_wire_N_613[4]), .I1(one_wire_N_613[2]), .I2(one_wire_N_613[3]), 
            .I3(GND_net), .O(n35357));   // verilog/neopixel.v(6[16:24])
    defparam i2_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 i3_4_lut (.I0(n16103), .I1(n35357), .I2(n7_adj_4676), .I3(n6), 
            .O(n21929));   // verilog/neopixel.v(104[14:39])
    defparam i3_4_lut.LUT_INIT = 16'hfffe;
    SB_CARRY mod_5_add_2076_6 (.CI(n29054), .I0(n3006), .I1(n3017), .CO(n29055));
    SB_LUT4 i1_4_lut_adj_1515 (.I0(n21929), .I1(n21937), .I2(\neo_pixel_transmitter.done ), 
            .I3(\state[0] ), .O(n26_adj_4683));
    defparam i1_4_lut_adj_1515.LUT_INIT = 16'h3553;
    SB_CARRY sub_14_add_2_7 (.CI(n27944), .I0(timer[5]), .I1(n51[5]), 
            .CO(n27945));
    SB_LUT4 sub_14_add_2_6_lut (.I0(GND_net), .I1(timer[4]), .I2(n51[4]), 
            .I3(n27943), .O(one_wire_N_613[4])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_1339_14_lut (.I0(n1898), .I1(n1898), .I2(n1928), 
            .I3(n28842), .O(n1997)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_14_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_2076_5_lut (.I0(n3007), .I1(n3007), .I2(n3017), 
            .I3(n29053), .O(n3106)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_5_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1339_14 (.CI(n28842), .I0(n1898), .I1(n1928), .CO(n28843));
    SB_LUT4 sub_14_inv_0_i24_1_lut (.I0(\neo_pixel_transmitter.t0 [23]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n51[23]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i24_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY sub_14_add_2_6 (.CI(n27943), .I0(timer[4]), .I1(n51[4]), 
            .CO(n27944));
    SB_LUT4 sub_14_add_2_5_lut (.I0(GND_net), .I1(timer[3]), .I2(n51[3]), 
            .I3(n27942), .O(one_wire_N_613[3])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_1339_13_lut (.I0(n1899), .I1(n1899), .I2(n1928), 
            .I3(n28841), .O(n1998)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_13_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1339_13 (.CI(n28841), .I0(n1899), .I1(n1928), .CO(n28842));
    SB_LUT4 i16_4_lut_adj_1516 (.I0(bit_ctr[17]), .I1(bit_ctr[5]), .I2(bit_ctr[24]), 
            .I3(bit_ctr[7]), .O(n44_adj_4686));
    defparam i16_4_lut_adj_1516.LUT_INIT = 16'hfffe;
    SB_CARRY mod_5_add_2076_5 (.CI(n29053), .I0(n3007), .I1(n3017), .CO(n29054));
    SB_CARRY add_21_32 (.CI(n27873), .I0(bit_ctr[30]), .I1(GND_net), .CO(n27874));
    SB_LUT4 mod_5_add_2076_4_lut (.I0(n3008), .I1(n3008), .I2(n3017), 
            .I3(n29052), .O(n3107)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_4_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1339_12_lut (.I0(n1900), .I1(n1900), .I2(n1928), 
            .I3(n28840), .O(n1999)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_12_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2076_4 (.CI(n29052), .I0(n3008), .I1(n3017), .CO(n29053));
    SB_CARRY mod_5_add_1339_12 (.CI(n28840), .I0(n1900), .I1(n1928), .CO(n28841));
    SB_LUT4 mod_5_add_1339_11_lut (.I0(n1901), .I1(n1901), .I2(n1928), 
            .I3(n28839), .O(n2000)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_11_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 sub_14_inv_0_i25_1_lut (.I0(\neo_pixel_transmitter.t0 [24]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n51[24]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i25_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i26_1_lut (.I0(\neo_pixel_transmitter.t0 [25]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n51[25]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i26_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY sub_14_add_2_5 (.CI(n27942), .I0(timer[3]), .I1(n51[3]), 
            .CO(n27943));
    SB_LUT4 i17162_3_lut (.I0(start), .I1(\neo_pixel_transmitter.done ), 
            .I2(\state[1] ), .I3(GND_net), .O(\neo_pixel_transmitter.done_N_670 ));   // verilog/neopixel.v(16[20:25])
    defparam i17162_3_lut.LUT_INIT = 16'hc1c1;
    SB_CARRY mod_5_add_1339_11 (.CI(n28839), .I0(n1901), .I1(n1928), .CO(n28840));
    SB_LUT4 mod_5_add_2076_3_lut (.I0(n3009), .I1(n3009), .I2(n38240), 
            .I3(n29051), .O(n3108)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_3_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 mod_5_add_1339_10_lut (.I0(n1902), .I1(n1902), .I2(n1928), 
            .I3(n28838), .O(n2001)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_10_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2076_3 (.CI(n29051), .I0(n3009), .I1(n38240), .CO(n29052));
    SB_CARRY mod_5_add_1339_10 (.CI(n28838), .I0(n1902), .I1(n1928), .CO(n28839));
    SB_LUT4 mod_5_add_2076_2_lut (.I0(bit_ctr[5]), .I1(bit_ctr[5]), .I2(n38240), 
            .I3(VCC_net), .O(n3109)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_2_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 mod_5_add_1339_9_lut (.I0(n1903), .I1(n1903), .I2(n1928), 
            .I3(n28837), .O(n2002)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_9_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 sub_14_add_2_4_lut (.I0(GND_net), .I1(timer[2]), .I2(n51[2]), 
            .I3(n27941), .O(one_wire_N_613[2])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1339_9 (.CI(n28837), .I0(n1903), .I1(n1928), .CO(n28838));
    SB_LUT4 i15_4_lut_adj_1517 (.I0(bit_ctr[3]), .I1(n30_adj_4677), .I2(bit_ctr[21]), 
            .I3(bit_ctr[4]), .O(n43));
    defparam i15_4_lut_adj_1517.LUT_INIT = 16'hfefc;
    SB_LUT4 i26_4_lut_adj_1518 (.I0(n45), .I1(n47_adj_4681), .I2(n46_adj_4680), 
            .I3(n48_adj_4678), .O(n54));
    defparam i26_4_lut_adj_1518.LUT_INIT = 16'hfffe;
    SB_LUT4 i21_4_lut_adj_1519 (.I0(bit_ctr[16]), .I1(bit_ctr[11]), .I2(bit_ctr[31]), 
            .I3(bit_ctr[20]), .O(n49_adj_4690));
    defparam i21_4_lut_adj_1519.LUT_INIT = 16'hfffe;
    SB_LUT4 i27_4_lut (.I0(n49_adj_4690), .I1(n54), .I2(n43), .I3(n44_adj_4686), 
            .O(\state_3__N_462[1] ));
    defparam i27_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i30764_2_lut (.I0(start), .I1(\neo_pixel_transmitter.done ), 
            .I2(GND_net), .I3(GND_net), .O(n37295));
    defparam i30764_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i13_4_lut_adj_1520 (.I0(n37295), .I1(\state_3__N_462[1] ), .I2(\state[1] ), 
            .I3(n21937), .O(n5));
    defparam i13_4_lut_adj_1520.LUT_INIT = 16'hcac0;
    SB_CARRY sub_14_add_2_4 (.CI(n27941), .I0(timer[2]), .I1(n51[2]), 
            .CO(n27942));
    SB_CARRY mod_5_add_2076_2 (.CI(VCC_net), .I0(bit_ctr[5]), .I1(n38240), 
            .CO(n29051));
    SB_LUT4 mod_5_add_1339_8_lut (.I0(n1904), .I1(n1904), .I2(n1928), 
            .I3(n28836), .O(n2003)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_8_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_2009_27_lut (.I0(n2885), .I1(n2885), .I2(n2918), 
            .I3(n29050), .O(n2984)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_27_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1339_8 (.CI(n28836), .I0(n1904), .I1(n1928), .CO(n28837));
    SB_LUT4 i13_4_lut_adj_1521 (.I0(n1460), .I1(n5), .I2(\state[0] ), 
            .I3(\state[1] ), .O(n33701));   // verilog/neopixel.v(16[20:25])
    defparam i13_4_lut_adj_1521.LUT_INIT = 16'h3f3a;
    SB_LUT4 mod_5_add_1339_7_lut (.I0(n1905), .I1(n1905), .I2(n1928), 
            .I3(n28835), .O(n2004)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_7_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_2009_26_lut (.I0(n2886), .I1(n2886), .I2(n2918), 
            .I3(n29049), .O(n2985)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_26_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 sub_14_add_2_3_lut (.I0(n4_adj_4692), .I1(timer[1]), .I2(n51[1]), 
            .I3(n27940), .O(n34639)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_3_lut.LUT_INIT = 16'hebbe;
    SB_CARRY mod_5_add_2009_26 (.CI(n29049), .I0(n2886), .I1(n2918), .CO(n29050));
    SB_LUT4 mod_5_add_2009_25_lut (.I0(n2887), .I1(n2887), .I2(n2918), 
            .I3(n29048), .O(n2986)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_25_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1339_7 (.CI(n28835), .I0(n1905), .I1(n1928), .CO(n28836));
    SB_CARRY mod_5_add_2009_25 (.CI(n29048), .I0(n2887), .I1(n2918), .CO(n29049));
    SB_LUT4 mod_5_add_1339_6_lut (.I0(n1906), .I1(n1906), .I2(n1928), 
            .I3(n28834), .O(n2005)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_6_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_2009_24_lut (.I0(n2888), .I1(n2888), .I2(n2918), 
            .I3(n29047), .O(n2987)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_24_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1339_6 (.CI(n28834), .I0(n1906), .I1(n1928), .CO(n28835));
    SB_CARRY mod_5_add_2009_24 (.CI(n29047), .I0(n2888), .I1(n2918), .CO(n29048));
    SB_LUT4 mod_5_add_1339_5_lut (.I0(n1907), .I1(n1907), .I2(n1928), 
            .I3(n28833), .O(n2006)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_5_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 add_21_31_lut (.I0(n1), .I1(bit_ctr[29]), .I2(GND_net), .I3(n27872), 
            .O(n37261)) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_31_lut.LUT_INIT = 16'h8228;
    SB_LUT4 mod_5_add_2009_23_lut (.I0(n2889), .I1(n2889), .I2(n2918), 
            .I3(n29046), .O(n2988)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_23_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1339_5 (.CI(n28833), .I0(n1907), .I1(n1928), .CO(n28834));
    SB_CARRY mod_5_add_2009_23 (.CI(n29046), .I0(n2889), .I1(n2918), .CO(n29047));
    SB_LUT4 mod_5_add_1339_4_lut (.I0(n1908), .I1(n1908), .I2(n1928), 
            .I3(n28832), .O(n2007)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_4_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_2009_22_lut (.I0(n2890), .I1(n2890), .I2(n2918), 
            .I3(n29045), .O(n2989)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_22_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1339_4 (.CI(n28832), .I0(n1908), .I1(n1928), .CO(n28833));
    SB_CARRY mod_5_add_2009_22 (.CI(n29045), .I0(n2890), .I1(n2918), .CO(n29046));
    SB_CARRY sub_14_add_2_3 (.CI(n27940), .I0(timer[1]), .I1(n51[1]), 
            .CO(n27941));
    SB_LUT4 mod_5_add_2009_21_lut (.I0(n2891), .I1(n2891), .I2(n2918), 
            .I3(n29044), .O(n2990)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_21_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2009_21 (.CI(n29044), .I0(n2891), .I1(n2918), .CO(n29045));
    SB_LUT4 mod_5_add_1339_3_lut (.I0(n1909), .I1(n1909), .I2(n38242), 
            .I3(n28831), .O(n2008)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_3_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 mod_5_add_2009_20_lut (.I0(n2892), .I1(n2892), .I2(n2918), 
            .I3(n29043), .O(n2991)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_20_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1339_3 (.CI(n28831), .I0(n1909), .I1(n38242), .CO(n28832));
    SB_LUT4 mod_5_add_1339_2_lut (.I0(bit_ctr[16]), .I1(bit_ctr[16]), .I2(n38242), 
            .I3(VCC_net), .O(n2009)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_2_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_2009_20 (.CI(n29043), .I0(n2892), .I1(n2918), .CO(n29044));
    SB_LUT4 mod_5_add_2009_19_lut (.I0(n2893), .I1(n2893), .I2(n2918), 
            .I3(n29042), .O(n2992)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_19_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1339_2 (.CI(VCC_net), .I0(bit_ctr[16]), .I1(n38242), 
            .CO(n28831));
    SB_LUT4 mod_5_add_1272_16_lut (.I0(n1796), .I1(n1796), .I2(n1829), 
            .I3(n28830), .O(n1895)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_16_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2009_19 (.CI(n29042), .I0(n2893), .I1(n2918), .CO(n29043));
    SB_LUT4 sub_14_add_2_2_lut (.I0(one_wire_N_613[2]), .I1(timer[0]), .I2(n51[0]), 
            .I3(VCC_net), .O(n4_adj_4692)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_2_lut.LUT_INIT = 16'hebbe;
    SB_LUT4 mod_5_add_2009_18_lut (.I0(n2894), .I1(n2894), .I2(n2918), 
            .I3(n29041), .O(n2993)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_18_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1272_15_lut (.I0(n1797), .I1(n1797), .I2(n1829), 
            .I3(n28829), .O(n1896)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_15_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1272_15 (.CI(n28829), .I0(n1797), .I1(n1829), .CO(n28830));
    SB_CARRY mod_5_add_2009_18 (.CI(n29041), .I0(n2894), .I1(n2918), .CO(n29042));
    SB_LUT4 mod_5_add_1272_14_lut (.I0(n1798), .I1(n1798), .I2(n1829), 
            .I3(n28828), .O(n1897)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_14_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY sub_14_add_2_2 (.CI(VCC_net), .I0(timer[0]), .I1(n51[0]), 
            .CO(n27940));
    SB_CARRY mod_5_add_1272_14 (.CI(n28828), .I0(n1798), .I1(n1829), .CO(n28829));
    SB_LUT4 mod_5_add_2009_17_lut (.I0(n2895), .I1(n2895), .I2(n2918), 
            .I3(n29040), .O(n2994)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_17_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2009_17 (.CI(n29040), .I0(n2895), .I1(n2918), .CO(n29041));
    SB_LUT4 mod_5_add_2009_16_lut (.I0(n2896), .I1(n2896), .I2(n2918), 
            .I3(n29039), .O(n2995)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_16_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1272_13_lut (.I0(n1799), .I1(n1799), .I2(n1829), 
            .I3(n28827), .O(n1898)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_13_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 sub_14_inv_0_i27_1_lut (.I0(\neo_pixel_transmitter.t0 [26]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n51[26]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i27_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_21_31 (.CI(n27872), .I0(bit_ctr[29]), .I1(GND_net), .CO(n27873));
    SB_CARRY mod_5_add_2009_16 (.CI(n29039), .I0(n2896), .I1(n2918), .CO(n29040));
    SB_CARRY mod_5_add_1272_13 (.CI(n28827), .I0(n1799), .I1(n1829), .CO(n28828));
    SB_LUT4 add_21_12_lut (.I0(n1), .I1(bit_ctr[10]), .I2(GND_net), .I3(n27853), 
            .O(n37225)) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_12_lut.LUT_INIT = 16'h8228;
    SB_LUT4 mod_5_add_2009_15_lut (.I0(n2897), .I1(n2897), .I2(n2918), 
            .I3(n29038), .O(n2996)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_15_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 sub_14_inv_0_i28_1_lut (.I0(\neo_pixel_transmitter.t0 [27]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n51[27]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i28_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i2_1_lut (.I0(\neo_pixel_transmitter.t0 [1]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n51[1]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i29_1_lut (.I0(\neo_pixel_transmitter.t0 [28]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n51[28]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i29_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i30_1_lut (.I0(\neo_pixel_transmitter.t0 [29]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n51[29]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i30_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i2_2_lut_adj_1522 (.I0(n1998), .I1(n2004), .I2(GND_net), .I3(GND_net), 
            .O(n18_adj_4697));
    defparam i2_2_lut_adj_1522.LUT_INIT = 16'heeee;
    SB_LUT4 i7_3_lut_adj_1523 (.I0(bit_ctr[11]), .I1(n2403), .I2(n2409), 
            .I3(GND_net), .O(n27_adj_4698));
    defparam i7_3_lut_adj_1523.LUT_INIT = 16'hecec;
    SB_LUT4 i13_4_lut_adj_1524 (.I0(n2390), .I1(n2391), .I2(n2397), .I3(n2394), 
            .O(n33_adj_4699));
    defparam i13_4_lut_adj_1524.LUT_INIT = 16'hfffe;
    SB_LUT4 i12_4_lut_adj_1525 (.I0(n2003), .I1(n1999), .I2(n1996), .I3(n2007), 
            .O(n28_adj_4700));
    defparam i12_4_lut_adj_1525.LUT_INIT = 16'hfffe;
    SB_LUT4 i12_4_lut_adj_1526 (.I0(n2392), .I1(n2405), .I2(n2400), .I3(n2398), 
            .O(n32_adj_4701));
    defparam i12_4_lut_adj_1526.LUT_INIT = 16'hfffe;
    SB_LUT4 i11_4_lut_adj_1527 (.I0(n2396), .I1(n2402), .I2(n2408), .I3(n2399), 
            .O(n31_adj_4702));
    defparam i11_4_lut_adj_1527.LUT_INIT = 16'hfffe;
    SB_LUT4 i10_4_lut_adj_1528 (.I0(n1997), .I1(n2005), .I2(n2000), .I3(n2002), 
            .O(n26_adj_4703));
    defparam i10_4_lut_adj_1528.LUT_INIT = 16'hfffe;
    SB_LUT4 i15_4_lut_adj_1529 (.I0(n2393), .I1(n2406), .I2(n2395), .I3(n2407), 
            .O(n35));
    defparam i15_4_lut_adj_1529.LUT_INIT = 16'hfffe;
    SB_LUT4 i17_4_lut_adj_1530 (.I0(n33_adj_4699), .I1(n27_adj_4698), .I2(n2404), 
            .I3(n2401), .O(n37_adj_4704));
    defparam i17_4_lut_adj_1530.LUT_INIT = 16'hfffe;
    SB_LUT4 i19_4_lut_adj_1531 (.I0(n37_adj_4704), .I1(n35), .I2(n31_adj_4702), 
            .I3(n32_adj_4701), .O(n2423));
    defparam i19_4_lut_adj_1531.LUT_INIT = 16'hfffe;
    SB_LUT4 i31571_1_lut (.I0(n2522), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n38251));
    defparam i31571_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i3_3_lut (.I0(bit_ctr[6]), .I1(n2902), .I2(n2909), .I3(GND_net), 
            .O(n28_adj_4705));
    defparam i3_3_lut.LUT_INIT = 16'hecec;
    SB_LUT4 i15_4_lut_adj_1532 (.I0(n2900), .I1(n2892), .I2(n2906), .I3(n2908), 
            .O(n40_adj_4706));
    defparam i15_4_lut_adj_1532.LUT_INIT = 16'hfffe;
    SB_LUT4 i11_4_lut_adj_1533 (.I0(n2001), .I1(n2008), .I2(n1994), .I3(n1995), 
            .O(n27_adj_4707));
    defparam i11_4_lut_adj_1533.LUT_INIT = 16'hfffe;
    SB_LUT4 i9_4_lut_adj_1534 (.I0(bit_ctr[15]), .I1(n18_adj_4697), .I2(n2006), 
            .I3(n2009), .O(n25_adj_4708));
    defparam i9_4_lut_adj_1534.LUT_INIT = 16'hfefc;
    SB_LUT4 i15_4_lut_adj_1535 (.I0(n25_adj_4708), .I1(n27_adj_4707), .I2(n26_adj_4703), 
            .I3(n28_adj_4700), .O(n2027));
    defparam i15_4_lut_adj_1535.LUT_INIT = 16'hfffe;
    SB_LUT4 i13_3_lut (.I0(n2895), .I1(n2887), .I2(n2891), .I3(GND_net), 
            .O(n38_adj_4709));
    defparam i13_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i31567_1_lut (.I0(n1631), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n38247));
    defparam i31567_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i18_4_lut_adj_1536 (.I0(n2907), .I1(n2889), .I2(n2890), .I3(n2904), 
            .O(n43_adj_4710));
    defparam i18_4_lut_adj_1536.LUT_INIT = 16'hfffe;
    SB_LUT4 sub_14_inv_0_i31_1_lut (.I0(\neo_pixel_transmitter.t0 [30]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n51[30]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i31_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i17_4_lut_adj_1537 (.I0(n2886), .I1(n2898), .I2(n2894), .I3(n2903), 
            .O(n42_adj_4711));
    defparam i17_4_lut_adj_1537.LUT_INIT = 16'hfffe;
    SB_LUT4 i14_4_lut_adj_1538 (.I0(n3004), .I1(n2989), .I2(n2990), .I3(n3007), 
            .O(n40_adj_4712));
    defparam i14_4_lut_adj_1538.LUT_INIT = 16'hfffe;
    SB_LUT4 i18_4_lut_adj_1539 (.I0(n3006), .I1(n2984), .I2(n2988), .I3(n2986), 
            .O(n44_adj_4713));
    defparam i18_4_lut_adj_1539.LUT_INIT = 16'hfffe;
    SB_LUT4 i16_4_lut_adj_1540 (.I0(n3008), .I1(n3003), .I2(n2994), .I3(n3002), 
            .O(n42_adj_4714));
    defparam i16_4_lut_adj_1540.LUT_INIT = 16'hfffe;
    SB_LUT4 i16_4_lut_adj_1541 (.I0(n2905), .I1(n2885), .I2(n2888), .I3(n2893), 
            .O(n41));
    defparam i16_4_lut_adj_1541.LUT_INIT = 16'hfffe;
    SB_LUT4 i20_4_lut_adj_1542 (.I0(n2901), .I1(n40_adj_4706), .I2(n28_adj_4705), 
            .I3(n2899), .O(n45_adj_4715));
    defparam i20_4_lut_adj_1542.LUT_INIT = 16'hfffe;
    SB_LUT4 i17_4_lut_adj_1543 (.I0(n2999), .I1(n3000), .I2(n2992), .I3(n2997), 
            .O(n43_adj_4716));
    defparam i17_4_lut_adj_1543.LUT_INIT = 16'hfffe;
    SB_LUT4 i15_4_lut_adj_1544 (.I0(n2996), .I1(n2985), .I2(n2995), .I3(n2987), 
            .O(n41_adj_4717));
    defparam i15_4_lut_adj_1544.LUT_INIT = 16'hfffe;
    SB_LUT4 i12_2_lut (.I0(n3001), .I1(n2993), .I2(GND_net), .I3(GND_net), 
            .O(n38_adj_4718));
    defparam i12_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i22_4_lut_adj_1545 (.I0(n43_adj_4710), .I1(n2896), .I2(n38_adj_4709), 
            .I3(n2897), .O(n47_adj_4719));
    defparam i22_4_lut_adj_1545.LUT_INIT = 16'hfffe;
    SB_LUT4 i20_3_lut (.I0(n2998), .I1(n40_adj_4712), .I2(n2991), .I3(GND_net), 
            .O(n46_adj_4720));
    defparam i20_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i24_4_lut (.I0(n47_adj_4719), .I1(n45_adj_4715), .I2(n41), 
            .I3(n42_adj_4711), .O(n2918));
    defparam i24_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i24_4_lut_adj_1546 (.I0(n41_adj_4717), .I1(n43_adj_4716), .I2(n42_adj_4714), 
            .I3(n44_adj_4713), .O(n50_adj_4721));
    defparam i24_4_lut_adj_1546.LUT_INIT = 16'hfffe;
    SB_LUT4 i11_3_lut (.I0(n3005), .I1(bit_ctr[5]), .I2(n3009), .I3(GND_net), 
            .O(n37_adj_4722));
    defparam i11_3_lut.LUT_INIT = 16'heaea;
    SB_LUT4 i25_4_lut (.I0(n37_adj_4722), .I1(n50_adj_4721), .I2(n46_adj_4720), 
            .I3(n38_adj_4718), .O(n3017));
    defparam i25_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i3_2_lut_adj_1547 (.I0(n2491), .I1(n2504), .I2(GND_net), .I3(GND_net), 
            .O(n24_adj_4723));
    defparam i3_2_lut_adj_1547.LUT_INIT = 16'heeee;
    SB_LUT4 i13_4_lut_adj_1548 (.I0(n2496), .I1(n2505), .I2(n2500), .I3(n2499), 
            .O(n34_adj_4724));
    defparam i13_4_lut_adj_1548.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_3_lut_adj_1549 (.I0(bit_ctr[10]), .I1(n2497), .I2(n2509), 
            .I3(GND_net), .O(n22_adj_4725));
    defparam i1_3_lut_adj_1549.LUT_INIT = 16'hecec;
    SB_LUT4 i17_4_lut_adj_1550 (.I0(n2490), .I1(n34_adj_4724), .I2(n24_adj_4723), 
            .I3(n2494), .O(n38_adj_4726));
    defparam i17_4_lut_adj_1550.LUT_INIT = 16'hfffe;
    SB_LUT4 i15_4_lut_adj_1551 (.I0(n2501), .I1(n2502), .I2(n2506), .I3(n2492), 
            .O(n36_adj_4727));
    defparam i15_4_lut_adj_1551.LUT_INIT = 16'hfffe;
    SB_LUT4 i16_4_lut_adj_1552 (.I0(n2495), .I1(n2498), .I2(n2493), .I3(n22_adj_4725), 
            .O(n37_adj_4728));
    defparam i16_4_lut_adj_1552.LUT_INIT = 16'hfffe;
    SB_LUT4 i14_4_lut_adj_1553 (.I0(n2507), .I1(n2508), .I2(n2503), .I3(n2489), 
            .O(n35_adj_4729));
    defparam i14_4_lut_adj_1553.LUT_INIT = 16'hfffe;
    SB_LUT4 i20_4_lut_adj_1554 (.I0(n35_adj_4729), .I1(n37_adj_4728), .I2(n36_adj_4727), 
            .I3(n38_adj_4726), .O(n2522));
    defparam i20_4_lut_adj_1554.LUT_INIT = 16'hfffe;
    SB_LUT4 i31569_1_lut (.I0(n2621), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n38249));
    defparam i31569_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i3_1_lut (.I0(\neo_pixel_transmitter.t0 [2]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n51[2]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i7_4_lut_adj_1555 (.I0(n1506), .I1(n1503), .I2(n1500), .I3(n1501), 
            .O(n18_adj_4730));
    defparam i7_4_lut_adj_1555.LUT_INIT = 16'hfffe;
    SB_LUT4 i9_4_lut_adj_1556 (.I0(n1504), .I1(n18_adj_4730), .I2(n1502), 
            .I3(n1499), .O(n20_adj_4731));
    defparam i9_4_lut_adj_1556.LUT_INIT = 16'hfffe;
    SB_LUT4 i4_3_lut_adj_1557 (.I0(bit_ctr[20]), .I1(n1505), .I2(n1509), 
            .I3(GND_net), .O(n15_adj_4732));
    defparam i4_3_lut_adj_1557.LUT_INIT = 16'hecec;
    SB_LUT4 i10_4_lut_adj_1558 (.I0(n15_adj_4732), .I1(n20_adj_4731), .I2(n1508), 
            .I3(n1507), .O(n1532));
    defparam i10_4_lut_adj_1558.LUT_INIT = 16'hfffe;
    SB_LUT4 i31570_1_lut (.I0(n1532), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n38250));
    defparam i31570_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i32_1_lut (.I0(\neo_pixel_transmitter.t0 [31]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n51[31]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i32_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i14_4_lut_adj_1559 (.I0(n2591), .I1(n2608), .I2(n2601), .I3(n2605), 
            .O(n36_adj_4733));
    defparam i14_4_lut_adj_1559.LUT_INIT = 16'hfffe;
    SB_LUT4 i3_3_lut_adj_1560 (.I0(n2606), .I1(bit_ctr[9]), .I2(n2609), 
            .I3(GND_net), .O(n25_adj_4734));
    defparam i3_3_lut_adj_1560.LUT_INIT = 16'heaea;
    SB_LUT4 i12_4_lut_adj_1561 (.I0(n2593), .I1(n2596), .I2(n2600), .I3(n2590), 
            .O(n34_adj_4735));
    defparam i12_4_lut_adj_1561.LUT_INIT = 16'hfffe;
    SB_LUT4 i18_4_lut_adj_1562 (.I0(n25_adj_4734), .I1(n36_adj_4733), .I2(n2594), 
            .I3(n2589), .O(n40_adj_4736));
    defparam i18_4_lut_adj_1562.LUT_INIT = 16'hfffe;
    SB_LUT4 i16_4_lut_adj_1563 (.I0(n2602), .I1(n2588), .I2(n2604), .I3(n2607), 
            .O(n38_adj_4737));
    defparam i16_4_lut_adj_1563.LUT_INIT = 16'hfffe;
    SB_LUT4 i31553_1_lut (.I0(n3116), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n38233));
    defparam i31553_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i17_3_lut (.I0(n2598), .I1(n34_adj_4735), .I2(n2603), .I3(GND_net), 
            .O(n39_adj_4738));
    defparam i17_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i15_4_lut_adj_1564 (.I0(n2592), .I1(n2597), .I2(n2595), .I3(n2599), 
            .O(n37_adj_4739));
    defparam i15_4_lut_adj_1564.LUT_INIT = 16'hfffe;
    SB_LUT4 mod_5_add_1272_12_lut (.I0(n1800), .I1(n1800), .I2(n1829), 
            .I3(n28826), .O(n1899)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_12_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i21_4_lut_adj_1565 (.I0(n37_adj_4739), .I1(n39_adj_4738), .I2(n38_adj_4737), 
            .I3(n40_adj_4736), .O(n2621));
    defparam i21_4_lut_adj_1565.LUT_INIT = 16'hfffe;
    SB_CARRY mod_5_add_1272_12 (.CI(n28826), .I0(n1800), .I1(n1829), .CO(n28827));
    SB_CARRY mod_5_add_2009_15 (.CI(n29038), .I0(n2897), .I1(n2918), .CO(n29039));
    SB_LUT4 mod_5_add_1272_11_lut (.I0(n1801), .I1(n1801), .I2(n1829), 
            .I3(n28825), .O(n1900)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_11_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1272_11 (.CI(n28825), .I0(n1801), .I1(n1829), .CO(n28826));
    SB_LUT4 mod_5_add_2009_14_lut (.I0(n2898), .I1(n2898), .I2(n2918), 
            .I3(n29037), .O(n2997)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_14_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1272_10_lut (.I0(n1802), .I1(n1802), .I2(n1829), 
            .I3(n28824), .O(n1901)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_10_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2009_14 (.CI(n29037), .I0(n2898), .I1(n2918), .CO(n29038));
    SB_CARRY mod_5_add_1272_10 (.CI(n28824), .I0(n1802), .I1(n1829), .CO(n28825));
    SB_LUT4 mod_5_add_2009_13_lut (.I0(n2899), .I1(n2899), .I2(n2918), 
            .I3(n29036), .O(n2998)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_13_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1272_9_lut (.I0(n1803), .I1(n1803), .I2(n1829), 
            .I3(n28823), .O(n1902)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_9_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2009_13 (.CI(n29036), .I0(n2899), .I1(n2918), .CO(n29037));
    SB_CARRY mod_5_add_1272_9 (.CI(n28823), .I0(n1803), .I1(n1829), .CO(n28824));
    SB_LUT4 mod_5_add_2009_12_lut (.I0(n2900), .I1(n2900), .I2(n2918), 
            .I3(n29035), .O(n2999)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_12_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1272_8_lut (.I0(n1804), .I1(n1804), .I2(n1829), 
            .I3(n28822), .O(n1903)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_8_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1272_8 (.CI(n28822), .I0(n1804), .I1(n1829), .CO(n28823));
    SB_LUT4 mod_5_add_1272_7_lut (.I0(n1805), .I1(n1805), .I2(n1829), 
            .I3(n28821), .O(n1904)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_7_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1272_7 (.CI(n28821), .I0(n1805), .I1(n1829), .CO(n28822));
    SB_CARRY mod_5_add_2009_12 (.CI(n29035), .I0(n2900), .I1(n2918), .CO(n29036));
    SB_LUT4 mod_5_add_2009_11_lut (.I0(n2901), .I1(n2901), .I2(n2918), 
            .I3(n29034), .O(n3000)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_11_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2009_11 (.CI(n29034), .I0(n2901), .I1(n2918), .CO(n29035));
    SB_LUT4 mod_5_add_1272_6_lut (.I0(n1806), .I1(n1806), .I2(n1829), 
            .I3(n28820), .O(n1905)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_6_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_2009_10_lut (.I0(n2902), .I1(n2902), .I2(n2918), 
            .I3(n29033), .O(n3001)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_10_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2009_10 (.CI(n29033), .I0(n2902), .I1(n2918), .CO(n29034));
    SB_CARRY mod_5_add_1272_6 (.CI(n28820), .I0(n1806), .I1(n1829), .CO(n28821));
    SB_LUT4 mod_5_add_1272_5_lut (.I0(n1807), .I1(n1807), .I2(n1829), 
            .I3(n28819), .O(n1906)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_5_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_2009_9_lut (.I0(n2903), .I1(n2903), .I2(n2918), 
            .I3(n29032), .O(n3002)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_9_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2009_9 (.CI(n29032), .I0(n2903), .I1(n2918), .CO(n29033));
    SB_CARRY mod_5_add_1272_5 (.CI(n28819), .I0(n1807), .I1(n1829), .CO(n28820));
    SB_LUT4 mod_5_add_1272_4_lut (.I0(n1808), .I1(n1808), .I2(n1829), 
            .I3(n28818), .O(n1907)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_4_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_2009_8_lut (.I0(n2904), .I1(n2904), .I2(n2918), 
            .I3(n29031), .O(n3003)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_8_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2009_8 (.CI(n29031), .I0(n2904), .I1(n2918), .CO(n29032));
    SB_LUT4 i31568_1_lut (.I0(n2720), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n38248));
    defparam i31568_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY mod_5_add_1272_4 (.CI(n28818), .I0(n1808), .I1(n1829), .CO(n28819));
    SB_LUT4 mod_5_add_1272_3_lut (.I0(n1809), .I1(n1809), .I2(n38244), 
            .I3(n28817), .O(n1908)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_3_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 mod_5_add_2009_7_lut (.I0(n2905), .I1(n2905), .I2(n2918), 
            .I3(n29030), .O(n3004)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_7_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1272_3 (.CI(n28817), .I0(n1809), .I1(n38244), .CO(n28818));
    SB_LUT4 mod_5_add_1272_2_lut (.I0(bit_ctr[17]), .I1(bit_ctr[17]), .I2(n38244), 
            .I3(VCC_net), .O(n1909)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_2_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_2009_7 (.CI(n29030), .I0(n2905), .I1(n2918), .CO(n29031));
    SB_CARRY mod_5_add_1272_2 (.CI(VCC_net), .I0(bit_ctr[17]), .I1(n38244), 
            .CO(n28817));
    SB_LUT4 mod_5_add_1205_15_lut (.I0(n1697), .I1(n1697), .I2(n1730), 
            .I3(n28816), .O(n1796)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1205_15_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_2009_6_lut (.I0(n2906), .I1(n2906), .I2(n2918), 
            .I3(n29029), .O(n3005)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_6_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1205_14_lut (.I0(n1698), .I1(n1698), .I2(n1730), 
            .I3(n28815), .O(n1797)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1205_14_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2009_6 (.CI(n29029), .I0(n2906), .I1(n2918), .CO(n29030));
    SB_CARRY mod_5_add_1205_14 (.CI(n28815), .I0(n1698), .I1(n1730), .CO(n28816));
    SB_LUT4 mod_5_add_2009_5_lut (.I0(n2907), .I1(n2907), .I2(n2918), 
            .I3(n29028), .O(n3006)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_5_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1205_13_lut (.I0(n1699), .I1(n1699), .I2(n1730), 
            .I3(n28814), .O(n1798)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1205_13_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2009_5 (.CI(n29028), .I0(n2907), .I1(n2918), .CO(n29029));
    SB_CARRY mod_5_add_1205_13 (.CI(n28814), .I0(n1699), .I1(n1730), .CO(n28815));
    SB_LUT4 mod_5_add_2009_4_lut (.I0(n2908), .I1(n2908), .I2(n2918), 
            .I3(n29027), .O(n3007)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_4_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1205_12_lut (.I0(n1700), .I1(n1700), .I2(n1730), 
            .I3(n28813), .O(n1799)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1205_12_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1205_12 (.CI(n28813), .I0(n1700), .I1(n1730), .CO(n28814));
    SB_CARRY mod_5_add_2009_4 (.CI(n29027), .I0(n2908), .I1(n2918), .CO(n29028));
    SB_LUT4 mod_5_add_1205_11_lut (.I0(n1701), .I1(n1701), .I2(n1730), 
            .I3(n28812), .O(n1800)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1205_11_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_2009_3_lut (.I0(n2909), .I1(n2909), .I2(n38243), 
            .I3(n29026), .O(n3008)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_3_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1205_11 (.CI(n28812), .I0(n1701), .I1(n1730), .CO(n28813));
    SB_CARRY mod_5_add_2009_3 (.CI(n29026), .I0(n2909), .I1(n38243), .CO(n29027));
    SB_LUT4 mod_5_add_2009_2_lut (.I0(bit_ctr[6]), .I1(bit_ctr[6]), .I2(n38243), 
            .I3(VCC_net), .O(n3009)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_2_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 mod_5_add_1205_10_lut (.I0(n1702), .I1(n1702), .I2(n1730), 
            .I3(n28811), .O(n1801)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1205_10_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1205_10 (.CI(n28811), .I0(n1702), .I1(n1730), .CO(n28812));
    SB_CARRY mod_5_add_2009_2 (.CI(VCC_net), .I0(bit_ctr[6]), .I1(n38243), 
            .CO(n29026));
    SB_LUT4 mod_5_add_1205_9_lut (.I0(n1703), .I1(n1703), .I2(n1730), 
            .I3(n28810), .O(n1802)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1205_9_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1942_26_lut (.I0(n2786), .I1(n2786), .I2(n2819), 
            .I3(n29025), .O(n2885)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_26_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1205_9 (.CI(n28810), .I0(n1703), .I1(n1730), .CO(n28811));
    SB_LUT4 mod_5_add_1942_25_lut (.I0(n2787), .I1(n2787), .I2(n2819), 
            .I3(n29024), .O(n2886)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_25_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1205_8_lut (.I0(n1704), .I1(n1704), .I2(n1730), 
            .I3(n28809), .O(n1803)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1205_8_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1942_25 (.CI(n29024), .I0(n2787), .I1(n2819), .CO(n29025));
    SB_CARRY mod_5_add_1205_8 (.CI(n28809), .I0(n1704), .I1(n1730), .CO(n28810));
    SB_LUT4 mod_5_add_1942_24_lut (.I0(n2788), .I1(n2788), .I2(n2819), 
            .I3(n29023), .O(n2887)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_24_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1205_7_lut (.I0(n1705), .I1(n1705), .I2(n1730), 
            .I3(n28808), .O(n1804)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1205_7_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1942_24 (.CI(n29023), .I0(n2788), .I1(n2819), .CO(n29024));
    SB_LUT4 mod_5_add_1942_23_lut (.I0(n2789), .I1(n2789), .I2(n2819), 
            .I3(n29022), .O(n2888)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_23_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1205_7 (.CI(n28808), .I0(n1705), .I1(n1730), .CO(n28809));
    SB_LUT4 mod_5_add_1205_6_lut (.I0(n1706), .I1(n1706), .I2(n1730), 
            .I3(n28807), .O(n1805)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1205_6_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1942_23 (.CI(n29022), .I0(n2789), .I1(n2819), .CO(n29023));
    SB_CARRY mod_5_add_1205_6 (.CI(n28807), .I0(n1706), .I1(n1730), .CO(n28808));
    SB_LUT4 mod_5_add_1942_22_lut (.I0(n2790), .I1(n2790), .I2(n2819), 
            .I3(n29021), .O(n2889)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_22_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1205_5_lut (.I0(n1707), .I1(n1707), .I2(n1730), 
            .I3(n28806), .O(n1806)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1205_5_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 add_21_30_lut (.I0(n1), .I1(bit_ctr[28]), .I2(GND_net), .I3(n27871), 
            .O(n37262)) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_30_lut.LUT_INIT = 16'h8228;
    SB_CARRY mod_5_add_1942_22 (.CI(n29021), .I0(n2790), .I1(n2819), .CO(n29022));
    SB_CARRY mod_5_add_1205_5 (.CI(n28806), .I0(n1707), .I1(n1730), .CO(n28807));
    SB_LUT4 mod_5_add_1942_21_lut (.I0(n2791), .I1(n2791), .I2(n2819), 
            .I3(n29020), .O(n2890)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_21_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1205_4_lut (.I0(n1708), .I1(n1708), .I2(n1730), 
            .I3(n28805), .O(n1807)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1205_4_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY add_21_12 (.CI(n27853), .I0(bit_ctr[10]), .I1(GND_net), .CO(n27854));
    SB_CARRY mod_5_add_1942_21 (.CI(n29020), .I0(n2791), .I1(n2819), .CO(n29021));
    SB_CARRY mod_5_add_1205_4 (.CI(n28805), .I0(n1708), .I1(n1730), .CO(n28806));
    SB_LUT4 mod_5_add_1205_3_lut (.I0(n1709), .I1(n1709), .I2(n38245), 
            .I3(n28804), .O(n1808)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1205_3_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 mod_5_add_1942_20_lut (.I0(n2792), .I1(n2792), .I2(n2819), 
            .I3(n29019), .O(n2891)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_20_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i31554_1_lut (.I0(n2126), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n38234));
    defparam i31554_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i31559_1_lut (.I0(n1037), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n38239));
    defparam i31559_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY mod_5_add_1205_3 (.CI(n28804), .I0(n1709), .I1(n38245), .CO(n28805));
    SB_LUT4 mod_5_add_1205_2_lut (.I0(bit_ctr[18]), .I1(bit_ctr[18]), .I2(n38245), 
            .I3(VCC_net), .O(n1809)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1205_2_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY add_21_30 (.CI(n27871), .I0(bit_ctr[28]), .I1(GND_net), .CO(n27872));
    SB_CARRY mod_5_add_1205_2 (.CI(VCC_net), .I0(bit_ctr[18]), .I1(n38245), 
            .CO(n28804));
    SB_CARRY mod_5_add_1942_20 (.CI(n29019), .I0(n2792), .I1(n2819), .CO(n29020));
    SB_LUT4 i31560_1_lut (.I0(n3017), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n38240));
    defparam i31560_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mod_5_add_1138_14_lut (.I0(n1598), .I1(n1598), .I2(n1631), 
            .I3(n28803), .O(n1697)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1138_14_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1138_13_lut (.I0(n1599), .I1(n1599), .I2(n1631), 
            .I3(n28802), .O(n1698)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1138_13_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1942_19_lut (.I0(n2793), .I1(n2793), .I2(n2819), 
            .I3(n29018), .O(n2892)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_19_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1942_19 (.CI(n29018), .I0(n2793), .I1(n2819), .CO(n29019));
    SB_LUT4 mod_5_add_1942_18_lut (.I0(n2794), .I1(n2794), .I2(n2819), 
            .I3(n29017), .O(n2893)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_18_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1138_13 (.CI(n28802), .I0(n1599), .I1(n1631), .CO(n28803));
    SB_LUT4 mod_5_add_1138_12_lut (.I0(n1600), .I1(n1600), .I2(n1631), 
            .I3(n28801), .O(n1699)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1138_12_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1942_18 (.CI(n29017), .I0(n2794), .I1(n2819), .CO(n29018));
    SB_LUT4 i30885_2_lut (.I0(n21937), .I1(\neo_pixel_transmitter.done ), 
            .I2(GND_net), .I3(GND_net), .O(n37325));
    defparam i30885_2_lut.LUT_INIT = 16'hdddd;
    SB_LUT4 i42_4_lut (.I0(n37325), .I1(n37323), .I2(\state[0] ), .I3(n1460), 
            .O(n28_adj_4740));
    defparam i42_4_lut.LUT_INIT = 16'hcac0;
    SB_LUT4 i1_3_lut_adj_1566 (.I0(\state[1] ), .I1(start), .I2(n28_adj_4740), 
            .I3(GND_net), .O(n20));
    defparam i1_3_lut_adj_1566.LUT_INIT = 16'hbaba;
    SB_CARRY mod_5_add_1138_12 (.CI(n28801), .I0(n1600), .I1(n1631), .CO(n28802));
    SB_LUT4 mod_5_add_1942_17_lut (.I0(n2795), .I1(n2795), .I2(n2819), 
            .I3(n29016), .O(n2894)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_17_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1138_11_lut (.I0(n1601), .I1(n1601), .I2(n1631), 
            .I3(n28800), .O(n1700)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1138_11_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1138_11 (.CI(n28800), .I0(n1601), .I1(n1631), .CO(n28801));
    SB_LUT4 sub_14_inv_0_i4_1_lut (.I0(\neo_pixel_transmitter.t0 [3]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n51[3]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i2_3_lut_adj_1567 (.I0(\state[0] ), .I1(\neo_pixel_transmitter.done ), 
            .I2(n25098), .I3(GND_net), .O(n35059));
    defparam i2_3_lut_adj_1567.LUT_INIT = 16'hfefe;
    SB_LUT4 i3_1_lut (.I0(\neo_pixel_transmitter.done ), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(\neo_pixel_transmitter.done_N_676 ));   // verilog/neopixel.v(35[12] 117[6])
    defparam i3_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mod_5_i538_3_lut_4_lut_3_lut_4_lut (.I0(n708), .I1(n30176), 
            .I2(bit_ctr[28]), .I3(GND_net), .O(n807));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i538_3_lut_4_lut_3_lut_4_lut.LUT_INIT = 16'h8080;
    SB_LUT4 mod_5_add_1138_10_lut (.I0(n1602), .I1(n1602), .I2(n1631), 
            .I3(n28799), .O(n1701)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1138_10_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1138_10 (.CI(n28799), .I0(n1602), .I1(n1631), .CO(n28800));
    SB_CARRY mod_5_add_1942_17 (.CI(n29016), .I0(n2795), .I1(n2819), .CO(n29017));
    SB_LUT4 mod_5_add_1942_16_lut (.I0(n2796), .I1(n2796), .I2(n2819), 
            .I3(n29015), .O(n2895)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_16_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1942_16 (.CI(n29015), .I0(n2796), .I1(n2819), .CO(n29016));
    SB_LUT4 mod_5_add_1138_9_lut (.I0(n1603), .I1(n1603), .I2(n1631), 
            .I3(n28798), .O(n1702)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1138_9_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1942_15_lut (.I0(n2797), .I1(n2797), .I2(n2819), 
            .I3(n29014), .O(n2896)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_15_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1942_15 (.CI(n29014), .I0(n2797), .I1(n2819), .CO(n29015));
    SB_CARRY mod_5_add_1138_9 (.CI(n28798), .I0(n1603), .I1(n1631), .CO(n28799));
    SB_LUT4 mod_5_add_1138_8_lut (.I0(n1604), .I1(n1604), .I2(n1631), 
            .I3(n28797), .O(n1703)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1138_8_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY add_21_5 (.CI(n27846), .I0(bit_ctr[3]), .I1(GND_net), .CO(n27847));
    SB_LUT4 add_21_11_lut (.I0(n1), .I1(bit_ctr[9]), .I2(GND_net), .I3(n27852), 
            .O(n37226)) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_11_lut.LUT_INIT = 16'h8228;
    SB_LUT4 add_21_29_lut (.I0(n1), .I1(bit_ctr[27]), .I2(GND_net), .I3(n27870), 
            .O(n37263)) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_29_lut.LUT_INIT = 16'h8228;
    SB_CARRY mod_5_add_1138_8 (.CI(n28797), .I0(n1604), .I1(n1631), .CO(n28798));
    SB_LUT4 mod_5_add_1942_14_lut (.I0(n2798), .I1(n2798), .I2(n2819), 
            .I3(n29013), .O(n2897)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_14_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1138_7_lut (.I0(n1605), .I1(n1605), .I2(n1631), 
            .I3(n28796), .O(n1704)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1138_7_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i1_2_lut_3_lut_4_lut_4_lut (.I0(n708), .I1(n30176), .I2(bit_ctr[28]), 
            .I3(GND_net), .O(n14844));   // verilog/neopixel.v(22[26:36])
    defparam i1_2_lut_3_lut_4_lut_4_lut.LUT_INIT = 16'he5e5;
    SB_LUT4 sub_14_inv_0_i5_1_lut (.I0(\neo_pixel_transmitter.t0 [4]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n51[4]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_21_29 (.CI(n27870), .I0(bit_ctr[27]), .I1(GND_net), .CO(n27871));
    SB_LUT4 i5_2_lut_adj_1568 (.I0(n2693), .I1(n2704), .I2(GND_net), .I3(GND_net), 
            .O(n28_adj_4742));
    defparam i5_2_lut_adj_1568.LUT_INIT = 16'heeee;
    SB_LUT4 i15_4_lut_adj_1569 (.I0(n2699), .I1(n2706), .I2(n2694), .I3(n2691), 
            .O(n38_adj_4743));
    defparam i15_4_lut_adj_1569.LUT_INIT = 16'hfffe;
    SB_LUT4 i20134_2_lut (.I0(bit_ctr[8]), .I1(n2709), .I2(GND_net), .I3(GND_net), 
            .O(n24956));
    defparam i20134_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i13_4_lut_adj_1570 (.I0(n2701), .I1(n2696), .I2(n2697), .I3(n24956), 
            .O(n36_adj_4744));
    defparam i13_4_lut_adj_1570.LUT_INIT = 16'hfffe;
    SB_LUT4 i19_4_lut_adj_1571 (.I0(n2700), .I1(n38_adj_4743), .I2(n28_adj_4742), 
            .I3(n2705), .O(n42_adj_4745));
    defparam i19_4_lut_adj_1571.LUT_INIT = 16'hfffe;
    SB_LUT4 i17_4_lut_adj_1572 (.I0(n2702), .I1(n2690), .I2(n2689), .I3(n2708), 
            .O(n40_adj_4746));
    defparam i17_4_lut_adj_1572.LUT_INIT = 16'hfffe;
    SB_LUT4 i18_4_lut_adj_1573 (.I0(n2687), .I1(n36_adj_4744), .I2(n2703), 
            .I3(n2695), .O(n41_adj_4747));
    defparam i18_4_lut_adj_1573.LUT_INIT = 16'hfffe;
    SB_LUT4 i16_4_lut_adj_1574 (.I0(n2688), .I1(n2698), .I2(n2692), .I3(n2707), 
            .O(n39_adj_4748));
    defparam i16_4_lut_adj_1574.LUT_INIT = 16'hfffe;
    SB_LUT4 i22_4_lut_adj_1575 (.I0(n39_adj_4748), .I1(n41_adj_4747), .I2(n40_adj_4746), 
            .I3(n42_adj_4745), .O(n2720));
    defparam i22_4_lut_adj_1575.LUT_INIT = 16'hfffe;
    SB_CARRY mod_5_add_1942_14 (.CI(n29013), .I0(n2798), .I1(n2819), .CO(n29014));
    SB_CARRY mod_5_add_1138_7 (.CI(n28796), .I0(n1605), .I1(n1631), .CO(n28797));
    SB_LUT4 mod_5_add_1942_13_lut (.I0(n2799), .I1(n2799), .I2(n2819), 
            .I3(n29012), .O(n2898)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_13_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1138_6_lut (.I0(n1606), .I1(n1606), .I2(n1631), 
            .I3(n28795), .O(n1705)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1138_6_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1138_6 (.CI(n28795), .I0(n1606), .I1(n1631), .CO(n28796));
    SB_LUT4 mod_5_add_1138_5_lut (.I0(n1607), .I1(n1607), .I2(n1631), 
            .I3(n28794), .O(n1706)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1138_5_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i20176_2_lut (.I0(bit_ctr[21]), .I1(n1409), .I2(GND_net), 
            .I3(GND_net), .O(n24998));
    defparam i20176_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i6_4_lut_adj_1576 (.I0(n1405), .I1(n24998), .I2(n1403), .I3(n1406), 
            .O(n16_adj_4749));
    defparam i6_4_lut_adj_1576.LUT_INIT = 16'hfffe;
    SB_LUT4 mod_5_add_1004_9_lut (.I0(n1403), .I1(n1403), .I2(n1433), 
            .I3(n28777), .O(n1502)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1004_9_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1942_13 (.CI(n29012), .I0(n2799), .I1(n2819), .CO(n29013));
    SB_LUT4 mod_5_add_1942_12_lut (.I0(n2800), .I1(n2800), .I2(n2819), 
            .I3(n29011), .O(n2899)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_12_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1942_12 (.CI(n29011), .I0(n2800), .I1(n2819), .CO(n29012));
    SB_LUT4 mod_5_add_1942_11_lut (.I0(n2801), .I1(n2801), .I2(n2819), 
            .I3(n29010), .O(n2900)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_11_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1942_11 (.CI(n29010), .I0(n2801), .I1(n2819), .CO(n29011));
    SB_LUT4 mod_5_add_1942_10_lut (.I0(n2802), .I1(n2802), .I2(n2819), 
            .I3(n29009), .O(n2901)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_10_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1942_10 (.CI(n29009), .I0(n2802), .I1(n2819), .CO(n29010));
    SB_LUT4 mod_5_add_1942_9_lut (.I0(n2803), .I1(n2803), .I2(n2819), 
            .I3(n29008), .O(n2902)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_9_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1942_9 (.CI(n29008), .I0(n2803), .I1(n2819), .CO(n29009));
    SB_LUT4 mod_5_add_1942_8_lut (.I0(n2804), .I1(n2804), .I2(n2819), 
            .I3(n29007), .O(n2903)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_8_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1942_8 (.CI(n29007), .I0(n2804), .I1(n2819), .CO(n29008));
    SB_LUT4 mod_5_add_1942_7_lut (.I0(n2805), .I1(n2805), .I2(n2819), 
            .I3(n29006), .O(n2904)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_7_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i31566_1_lut (.I0(n2819), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n38246));
    defparam i31566_1_lut.LUT_INIT = 16'h5555;
    SB_DFFESS state_i0 (.Q(\state[0] ), .C(clk32MHz), .E(n17229), .D(state_3__N_462[0]), 
            .S(n17500));   // verilog/neopixel.v(35[12] 117[6])
    SB_LUT4 add_21_28_lut (.I0(n1), .I1(bit_ctr[26]), .I2(GND_net), .I3(n27869), 
            .O(n37304)) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_28_lut.LUT_INIT = 16'h8228;
    SB_CARRY mod_5_add_1942_7 (.CI(n29006), .I0(n2805), .I1(n2819), .CO(n29007));
    SB_LUT4 mod_5_add_1942_6_lut (.I0(n2806), .I1(n2806), .I2(n2819), 
            .I3(n29005), .O(n2905)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_6_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i6_4_lut_adj_1577 (.I0(n3185), .I1(n3200), .I2(n3192), .I3(n3182), 
            .O(n14_adj_4750));
    defparam i6_4_lut_adj_1577.LUT_INIT = 16'hfffe;
    SB_LUT4 i5_4_lut_adj_1578 (.I0(n3193), .I1(n3201), .I2(n3184), .I3(n3190), 
            .O(n13_adj_4751));
    defparam i5_4_lut_adj_1578.LUT_INIT = 16'hfffe;
    SB_LUT4 i20039_2_lut (.I0(bit_ctr[3]), .I1(n3209), .I2(GND_net), .I3(GND_net), 
            .O(n24860));
    defparam i20039_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i13_4_lut_adj_1579 (.I0(n3196), .I1(n3186), .I2(n24860), .I3(n3202), 
            .O(n34_adj_4752));
    defparam i13_4_lut_adj_1579.LUT_INIT = 16'hfffe;
    SB_LUT4 i2_3_lut_adj_1580 (.I0(n13_adj_4751), .I1(n3206), .I2(n14_adj_4750), 
            .I3(GND_net), .O(n23_adj_4753));
    defparam i2_3_lut_adj_1580.LUT_INIT = 16'hfefe;
    SB_LUT4 i1_2_lut_adj_1581 (.I0(n3198), .I1(n3189), .I2(GND_net), .I3(GND_net), 
            .O(n22_adj_4754));
    defparam i1_2_lut_adj_1581.LUT_INIT = 16'heeee;
    SB_LUT4 i17_4_lut_adj_1582 (.I0(n23_adj_4753), .I1(n34_adj_4752), .I2(n3197), 
            .I3(n3199), .O(n38_adj_4755));
    defparam i17_4_lut_adj_1582.LUT_INIT = 16'hfffe;
    SB_LUT4 i15_4_lut_adj_1583 (.I0(n3203), .I1(n3204), .I2(n3195), .I3(n3191), 
            .O(n36_adj_4756));
    defparam i15_4_lut_adj_1583.LUT_INIT = 16'hfffe;
    SB_LUT4 i16_4_lut_adj_1584 (.I0(n3183), .I1(n3208), .I2(n3188), .I3(n22_adj_4754), 
            .O(n37_adj_4757));
    defparam i16_4_lut_adj_1584.LUT_INIT = 16'hfffe;
    SB_CARRY mod_5_add_1942_6 (.CI(n29005), .I0(n2806), .I1(n2819), .CO(n29006));
    SB_LUT4 mod_5_add_1942_5_lut (.I0(n2807), .I1(n2807), .I2(n2819), 
            .I3(n29004), .O(n2906)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_5_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i14_4_lut_adj_1585 (.I0(n3205), .I1(n3207), .I2(n3187), .I3(n3194), 
            .O(n35_adj_4758));
    defparam i14_4_lut_adj_1585.LUT_INIT = 16'hfffe;
    SB_LUT4 i20_4_lut_adj_1586 (.I0(n35_adj_4758), .I1(n37_adj_4757), .I2(n36_adj_4756), 
            .I3(n38_adj_4755), .O(n24890));
    defparam i20_4_lut_adj_1586.LUT_INIT = 16'hfffe;
    SB_CARRY mod_5_add_1942_5 (.CI(n29004), .I0(n2807), .I1(n2819), .CO(n29005));
    SB_LUT4 color_bit_I_0_i9_3_lut (.I0(\color[10] ), .I1(\color[11] ), 
            .I2(bit_ctr[0]), .I3(GND_net), .O(n9_adj_4759));   // verilog/neopixel.v(22[26:36])
    defparam color_bit_I_0_i9_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_adj_1587 (.I0(\color[12] ), .I1(bit_ctr[0]), .I2(GND_net), 
            .I3(GND_net), .O(n4_adj_4760));
    defparam i1_2_lut_adj_1587.LUT_INIT = 16'h2222;
    SB_LUT4 i31097_4_lut (.I0(\color[9] ), .I1(n9_adj_4759), .I2(bit_ctr[1]), 
            .I3(bit_ctr[0]), .O(n37779));   // verilog/neopixel.v(22[26:36])
    defparam i31097_4_lut.LUT_INIT = 16'hcac0;
    SB_LUT4 i29720_4_lut (.I0(n3209), .I1(\state_3__N_462[1] ), .I2(bit_ctr[3]), 
            .I3(n24890), .O(n36317));
    defparam i29720_4_lut.LUT_INIT = 16'hdeee;
    SB_LUT4 color_bit_I_0_i14_4_lut (.I0(n37779), .I1(bit_ctr[1]), .I2(bit_ctr[2]), 
            .I3(n4_adj_4760), .O(n14_adj_4761));   // verilog/neopixel.v(22[26:36])
    defparam color_bit_I_0_i14_4_lut.LUT_INIT = 16'h3a0a;
    SB_CARRY add_21_28 (.CI(n27869), .I0(bit_ctr[26]), .I1(GND_net), .CO(n27870));
    SB_LUT4 mod_5_add_1942_4_lut (.I0(n2808), .I1(n2808), .I2(n2819), 
            .I3(n29003), .O(n2907)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_4_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i3_4_lut_adj_1588 (.I0(n14_adj_4761), .I1(n36317), .I2(bit_ctr[3]), 
            .I3(n24890), .O(state_3__N_462[0]));   // verilog/neopixel.v(40[18] 45[12])
    defparam i3_4_lut_adj_1588.LUT_INIT = 16'h0220;
    SB_CARRY mod_5_add_1942_4 (.CI(n29003), .I0(n2808), .I1(n2819), .CO(n29004));
    SB_LUT4 i7_4_lut_adj_1589 (.I0(n1402), .I1(n1404), .I2(n1400), .I3(n1407), 
            .O(n17_adj_4762));
    defparam i7_4_lut_adj_1589.LUT_INIT = 16'hfffe;
    SB_LUT4 i9_4_lut_adj_1590 (.I0(n17_adj_4762), .I1(n1408), .I2(n16_adj_4749), 
            .I3(n1401), .O(n1433));
    defparam i9_4_lut_adj_1590.LUT_INIT = 16'hfffe;
    SB_LUT4 add_21_27_lut (.I0(n1), .I1(bit_ctr[25]), .I2(GND_net), .I3(n27868), 
            .O(n37308)) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_27_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_21_27 (.CI(n27868), .I0(bit_ctr[25]), .I1(GND_net), .CO(n27869));
    SB_LUT4 add_21_26_lut (.I0(n1), .I1(bit_ctr[24]), .I2(GND_net), .I3(n27867), 
            .O(n37309)) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_26_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_21_26 (.CI(n27867), .I0(bit_ctr[24]), .I1(GND_net), .CO(n27868));
    SB_LUT4 mod_5_add_1942_3_lut (.I0(n2809), .I1(n2809), .I2(n38246), 
            .I3(n29002), .O(n2908)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_3_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1942_3 (.CI(n29002), .I0(n2809), .I1(n38246), .CO(n29003));
    SB_LUT4 i1_2_lut_4_lut (.I0(\state[1] ), .I1(\state[0] ), .I2(\neo_pixel_transmitter.done ), 
            .I3(n25098), .O(n32854));   // verilog/neopixel.v(35[12] 117[6])
    defparam i1_2_lut_4_lut.LUT_INIT = 16'h0002;
    SB_LUT4 add_21_25_lut (.I0(n1), .I1(bit_ctr[23]), .I2(GND_net), .I3(n27866), 
            .O(n37330)) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_25_lut.LUT_INIT = 16'h8228;
    SB_LUT4 mod_5_add_1942_2_lut (.I0(bit_ctr[7]), .I1(bit_ctr[7]), .I2(n38246), 
            .I3(VCC_net), .O(n2909)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_2_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1942_2 (.CI(VCC_net), .I0(bit_ctr[7]), .I1(n38246), 
            .CO(n29002));
    SB_LUT4 i43_3_lut_4_lut (.I0(start), .I1(n26_adj_4683), .I2(\state[1] ), 
            .I3(n35059), .O(n17243));
    defparam i43_3_lut_4_lut.LUT_INIT = 16'h04f4;
    SB_LUT4 mod_5_add_1875_25_lut (.I0(n2687), .I1(n2687), .I2(n2720), 
            .I3(n29001), .O(n2786)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_25_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1875_24_lut (.I0(n2688), .I1(n2688), .I2(n2720), 
            .I3(n29000), .O(n2787)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_24_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i31522_2_lut_3_lut (.I0(start), .I1(n26_adj_4683), .I2(\state[1] ), 
            .I3(GND_net), .O(n32930));
    defparam i31522_2_lut_3_lut.LUT_INIT = 16'hfbfb;
    SB_CARRY mod_5_add_1875_24 (.CI(n29000), .I0(n2688), .I1(n2720), .CO(n29001));
    SB_LUT4 mod_5_add_1875_23_lut (.I0(n2689), .I1(n2689), .I2(n2720), 
            .I3(n28999), .O(n2788)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_23_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1875_23 (.CI(n28999), .I0(n2689), .I1(n2720), .CO(n29000));
    SB_LUT4 mod_5_add_1875_22_lut (.I0(n2690), .I1(n2690), .I2(n2720), 
            .I3(n28998), .O(n2789)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_22_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 sub_14_inv_0_i6_1_lut (.I0(\neo_pixel_transmitter.t0 [5]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n51[5]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY mod_5_add_1875_22 (.CI(n28998), .I0(n2690), .I1(n2720), .CO(n28999));
    SB_LUT4 mod_5_add_1875_21_lut (.I0(n2691), .I1(n2691), .I2(n2720), 
            .I3(n28997), .O(n2790)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_21_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1875_21 (.CI(n28997), .I0(n2691), .I1(n2720), .CO(n28998));
    SB_LUT4 mod_5_add_1875_20_lut (.I0(n2692), .I1(n2692), .I2(n2720), 
            .I3(n28996), .O(n2791)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_20_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1875_20 (.CI(n28996), .I0(n2692), .I1(n2720), .CO(n28997));
    SB_LUT4 mod_5_add_1875_19_lut (.I0(n2693), .I1(n2693), .I2(n2720), 
            .I3(n28995), .O(n2792)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_19_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1875_19 (.CI(n28995), .I0(n2693), .I1(n2720), .CO(n28996));
    SB_LUT4 mod_5_add_1875_18_lut (.I0(n2694), .I1(n2694), .I2(n2720), 
            .I3(n28994), .O(n2793)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_18_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1875_18 (.CI(n28994), .I0(n2694), .I1(n2720), .CO(n28995));
    SB_LUT4 mod_5_add_1875_17_lut (.I0(n2695), .I1(n2695), .I2(n2720), 
            .I3(n28993), .O(n2794)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_17_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1875_17 (.CI(n28993), .I0(n2695), .I1(n2720), .CO(n28994));
    SB_LUT4 mod_5_add_1875_16_lut (.I0(n2696), .I1(n2696), .I2(n2720), 
            .I3(n28992), .O(n2795)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_16_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1875_16 (.CI(n28992), .I0(n2696), .I1(n2720), .CO(n28993));
    SB_CARRY add_21_25 (.CI(n27866), .I0(bit_ctr[23]), .I1(GND_net), .CO(n27867));
    SB_LUT4 i10_4_lut_adj_1591 (.I0(n2193), .I1(n2194), .I2(n2206), .I3(n2204), 
            .O(n28_adj_4763));
    defparam i10_4_lut_adj_1591.LUT_INIT = 16'hfffe;
    SB_LUT4 i14_4_lut_adj_1592 (.I0(n2203), .I1(n28_adj_4763), .I2(bit_ctr[13]), 
            .I3(n2209), .O(n32_adj_4764));
    defparam i14_4_lut_adj_1592.LUT_INIT = 16'hfeee;
    SB_LUT4 i12_4_lut_adj_1593 (.I0(n2208), .I1(n2201), .I2(n2192), .I3(n2196), 
            .O(n30_adj_4765));
    defparam i12_4_lut_adj_1593.LUT_INIT = 16'hfffe;
    SB_LUT4 i13_4_lut_adj_1594 (.I0(n2195), .I1(n2207), .I2(n2205), .I3(n2199), 
            .O(n31_adj_4766));
    defparam i13_4_lut_adj_1594.LUT_INIT = 16'hfffe;
    SB_LUT4 i11_4_lut_adj_1595 (.I0(n2202), .I1(n2197), .I2(n2198), .I3(n2200), 
            .O(n29_adj_4767));
    defparam i11_4_lut_adj_1595.LUT_INIT = 16'hfffe;
    SB_DFFESR one_wire_108 (.Q(PIN_8_c), .C(clk32MHz), .E(n17243), .D(\neo_pixel_transmitter.done_N_676 ), 
            .R(n32854));   // verilog/neopixel.v(35[12] 117[6])
    SB_LUT4 i19658_2_lut_3_lut (.I0(start), .I1(\neo_pixel_transmitter.done ), 
            .I2(n21929), .I3(GND_net), .O(n1460));   // verilog/neopixel.v(79[18] 99[12])
    defparam i19658_2_lut_3_lut.LUT_INIT = 16'hbfbf;
    SB_LUT4 mod_5_add_1875_15_lut (.I0(n2697), .I1(n2697), .I2(n2720), 
            .I3(n28991), .O(n2796)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_15_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i30866_4_lut_4_lut (.I0(start), .I1(\neo_pixel_transmitter.done ), 
            .I2(n21937), .I3(n21929), .O(n37323));   // verilog/neopixel.v(79[18] 99[12])
    defparam i30866_4_lut_4_lut.LUT_INIT = 16'h8cbf;
    SB_LUT4 add_21_4_lut (.I0(n1), .I1(bit_ctr[2]), .I2(GND_net), .I3(n27845), 
            .O(n37251)) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_4_lut.LUT_INIT = 16'h8228;
    SB_CARRY mod_5_add_1875_15 (.CI(n28991), .I0(n2697), .I1(n2720), .CO(n28992));
    SB_LUT4 mod_5_add_1875_14_lut (.I0(n2698), .I1(n2698), .I2(n2720), 
            .I3(n28990), .O(n2797)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_14_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY add_21_11 (.CI(n27852), .I0(bit_ctr[9]), .I1(GND_net), .CO(n27853));
    SB_CARRY mod_5_add_1875_14 (.CI(n28990), .I0(n2698), .I1(n2720), .CO(n28991));
    SB_LUT4 mod_5_add_1875_13_lut (.I0(n2699), .I1(n2699), .I2(n2720), 
            .I3(n28989), .O(n2798)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_13_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1875_13 (.CI(n28989), .I0(n2699), .I1(n2720), .CO(n28990));
    SB_LUT4 mod_5_add_1875_12_lut (.I0(n2700), .I1(n2700), .I2(n2720), 
            .I3(n28988), .O(n2799)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_12_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i17_4_lut_adj_1596 (.I0(n29_adj_4767), .I1(n31_adj_4766), .I2(n30_adj_4765), 
            .I3(n32_adj_4764), .O(n2225));
    defparam i17_4_lut_adj_1596.LUT_INIT = 16'hfffe;
    SB_CARRY mod_5_add_1875_12 (.CI(n28988), .I0(n2700), .I1(n2720), .CO(n28989));
    SB_LUT4 mod_5_add_1875_11_lut (.I0(n2701), .I1(n2701), .I2(n2720), 
            .I3(n28987), .O(n2800)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_11_lut.LUT_INIT = 16'hCA3A;
    SB_DFF timer_1524__i1 (.Q(timer[1]), .C(clk32MHz), .D(n133[1]));   // verilog/neopixel.v(12[12:21])
    SB_CARRY mod_5_add_1875_11 (.CI(n28987), .I0(n2701), .I1(n2720), .CO(n28988));
    SB_LUT4 mod_5_add_1875_10_lut (.I0(n2702), .I1(n2702), .I2(n2720), 
            .I3(n28986), .O(n2801)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_10_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1875_10 (.CI(n28986), .I0(n2702), .I1(n2720), .CO(n28987));
    SB_LUT4 mod_5_add_1875_9_lut (.I0(n2703), .I1(n2703), .I2(n2720), 
            .I3(n28985), .O(n2802)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_9_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1875_9 (.CI(n28985), .I0(n2703), .I1(n2720), .CO(n28986));
    SB_LUT4 mod_5_add_1875_8_lut (.I0(n2704), .I1(n2704), .I2(n2720), 
            .I3(n28984), .O(n2803)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_8_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1875_8 (.CI(n28984), .I0(n2704), .I1(n2720), .CO(n28985));
    SB_LUT4 mod_5_add_1875_7_lut (.I0(n2705), .I1(n2705), .I2(n2720), 
            .I3(n28983), .O(n2804)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_7_lut.LUT_INIT = 16'hCA3A;
    SB_DFF timer_1524__i2 (.Q(timer[2]), .C(clk32MHz), .D(n133[2]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1524__i3 (.Q(timer[3]), .C(clk32MHz), .D(n133[3]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1524__i4 (.Q(timer[4]), .C(clk32MHz), .D(n133[4]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1524__i5 (.Q(timer[5]), .C(clk32MHz), .D(n133[5]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1524__i6 (.Q(timer[6]), .C(clk32MHz), .D(n133[6]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1524__i7 (.Q(timer[7]), .C(clk32MHz), .D(n133[7]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1524__i8 (.Q(timer[8]), .C(clk32MHz), .D(n133[8]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1524__i9 (.Q(timer[9]), .C(clk32MHz), .D(n133[9]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1524__i10 (.Q(timer[10]), .C(clk32MHz), .D(n133[10]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1524__i11 (.Q(timer[11]), .C(clk32MHz), .D(n133[11]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1524__i12 (.Q(timer[12]), .C(clk32MHz), .D(n133[12]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1524__i13 (.Q(timer[13]), .C(clk32MHz), .D(n133[13]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1524__i14 (.Q(timer[14]), .C(clk32MHz), .D(n133[14]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1524__i15 (.Q(timer[15]), .C(clk32MHz), .D(n133[15]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1524__i16 (.Q(timer[16]), .C(clk32MHz), .D(n133[16]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1524__i17 (.Q(timer[17]), .C(clk32MHz), .D(n133[17]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1524__i18 (.Q(timer[18]), .C(clk32MHz), .D(n133[18]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1524__i19 (.Q(timer[19]), .C(clk32MHz), .D(n133[19]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1524__i20 (.Q(timer[20]), .C(clk32MHz), .D(n133[20]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1524__i21 (.Q(timer[21]), .C(clk32MHz), .D(n133[21]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1524__i22 (.Q(timer[22]), .C(clk32MHz), .D(n133[22]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1524__i23 (.Q(timer[23]), .C(clk32MHz), .D(n133[23]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1524__i24 (.Q(timer[24]), .C(clk32MHz), .D(n133[24]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1524__i25 (.Q(timer[25]), .C(clk32MHz), .D(n133[25]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1524__i26 (.Q(timer[26]), .C(clk32MHz), .D(n133[26]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1524__i27 (.Q(timer[27]), .C(clk32MHz), .D(n133[27]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1524__i28 (.Q(timer[28]), .C(clk32MHz), .D(n133[28]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1524__i29 (.Q(timer[29]), .C(clk32MHz), .D(n133[29]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1524__i30 (.Q(timer[30]), .C(clk32MHz), .D(n133[30]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1524__i31 (.Q(timer[31]), .C(clk32MHz), .D(n133[31]));   // verilog/neopixel.v(12[12:21])
    SB_DFF \neo_pixel_transmitter.t0_i0_i0  (.Q(\neo_pixel_transmitter.t0 [0]), 
           .C(clk32MHz), .D(n17546));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i31  (.Q(\neo_pixel_transmitter.t0 [31]), 
           .C(clk32MHz), .D(n17767));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i30  (.Q(\neo_pixel_transmitter.t0 [30]), 
           .C(clk32MHz), .D(n17766));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i29  (.Q(\neo_pixel_transmitter.t0 [29]), 
           .C(clk32MHz), .D(n17765));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i28  (.Q(\neo_pixel_transmitter.t0 [28]), 
           .C(clk32MHz), .D(n17764));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i27  (.Q(\neo_pixel_transmitter.t0 [27]), 
           .C(clk32MHz), .D(n17763));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i26  (.Q(\neo_pixel_transmitter.t0 [26]), 
           .C(clk32MHz), .D(n17762));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i25  (.Q(\neo_pixel_transmitter.t0 [25]), 
           .C(clk32MHz), .D(n17761));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i24  (.Q(\neo_pixel_transmitter.t0 [24]), 
           .C(clk32MHz), .D(n17760));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i23  (.Q(\neo_pixel_transmitter.t0 [23]), 
           .C(clk32MHz), .D(n17759));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i22  (.Q(\neo_pixel_transmitter.t0 [22]), 
           .C(clk32MHz), .D(n17758));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i21  (.Q(\neo_pixel_transmitter.t0 [21]), 
           .C(clk32MHz), .D(n17757));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i20  (.Q(\neo_pixel_transmitter.t0 [20]), 
           .C(clk32MHz), .D(n17756));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i19  (.Q(\neo_pixel_transmitter.t0 [19]), 
           .C(clk32MHz), .D(n17755));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i18  (.Q(\neo_pixel_transmitter.t0 [18]), 
           .C(clk32MHz), .D(n17754));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i17  (.Q(\neo_pixel_transmitter.t0 [17]), 
           .C(clk32MHz), .D(n17753));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i16  (.Q(\neo_pixel_transmitter.t0 [16]), 
           .C(clk32MHz), .D(n17752));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i15  (.Q(\neo_pixel_transmitter.t0 [15]), 
           .C(clk32MHz), .D(n17751));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i14  (.Q(\neo_pixel_transmitter.t0 [14]), 
           .C(clk32MHz), .D(n17750));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i13  (.Q(\neo_pixel_transmitter.t0 [13]), 
           .C(clk32MHz), .D(n17749));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i12  (.Q(\neo_pixel_transmitter.t0 [12]), 
           .C(clk32MHz), .D(n17748));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i11  (.Q(\neo_pixel_transmitter.t0 [11]), 
           .C(clk32MHz), .D(n17747));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i10  (.Q(\neo_pixel_transmitter.t0 [10]), 
           .C(clk32MHz), .D(n17746));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i9  (.Q(\neo_pixel_transmitter.t0 [9]), 
           .C(clk32MHz), .D(n17745));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i8  (.Q(\neo_pixel_transmitter.t0 [8]), 
           .C(clk32MHz), .D(n17744));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i7  (.Q(\neo_pixel_transmitter.t0 [7]), 
           .C(clk32MHz), .D(n17743));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i6  (.Q(\neo_pixel_transmitter.t0 [6]), 
           .C(clk32MHz), .D(n17742));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i5  (.Q(\neo_pixel_transmitter.t0 [5]), 
           .C(clk32MHz), .D(n17741));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i4  (.Q(\neo_pixel_transmitter.t0 [4]), 
           .C(clk32MHz), .D(n17740));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i3  (.Q(\neo_pixel_transmitter.t0 [3]), 
           .C(clk32MHz), .D(n17739));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i2  (.Q(\neo_pixel_transmitter.t0 [2]), 
           .C(clk32MHz), .D(n17738));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i1  (.Q(\neo_pixel_transmitter.t0 [1]), 
           .C(clk32MHz), .D(n17737));   // verilog/neopixel.v(35[12] 117[6])
    SB_CARRY mod_5_add_1875_7 (.CI(n28983), .I0(n2705), .I1(n2720), .CO(n28984));
    SB_LUT4 mod_5_add_1875_6_lut (.I0(n2706), .I1(n2706), .I2(n2720), 
            .I3(n28982), .O(n2805)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_6_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1875_6 (.CI(n28982), .I0(n2706), .I1(n2720), .CO(n28983));
    SB_LUT4 mod_5_add_1875_5_lut (.I0(n2707), .I1(n2707), .I2(n2720), 
            .I3(n28981), .O(n2806)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_5_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1875_5 (.CI(n28981), .I0(n2707), .I1(n2720), .CO(n28982));
    SB_LUT4 mod_5_add_1875_4_lut (.I0(n2708), .I1(n2708), .I2(n2720), 
            .I3(n28980), .O(n2807)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_4_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1875_4 (.CI(n28980), .I0(n2708), .I1(n2720), .CO(n28981));
    SB_LUT4 add_21_24_lut (.I0(n1), .I1(bit_ctr[22]), .I2(GND_net), .I3(n27865), 
            .O(n37335)) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_24_lut.LUT_INIT = 16'h8228;
    SB_LUT4 mod_5_add_1875_3_lut (.I0(n2709), .I1(n2709), .I2(n38248), 
            .I3(n28979), .O(n2808)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_3_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1875_3 (.CI(n28979), .I0(n2709), .I1(n38248), .CO(n28980));
    SB_LUT4 mod_5_add_1875_2_lut (.I0(bit_ctr[8]), .I1(bit_ctr[8]), .I2(n38248), 
            .I3(VCC_net), .O(n2809)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_2_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY add_21_24 (.CI(n27865), .I0(bit_ctr[22]), .I1(GND_net), .CO(n27866));
    SB_CARRY mod_5_add_1875_2 (.CI(VCC_net), .I0(bit_ctr[8]), .I1(n38248), 
            .CO(n28979));
    SB_LUT4 mod_5_add_1808_24_lut (.I0(n2588), .I1(n2588), .I2(n2621), 
            .I3(n28978), .O(n2687)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_24_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1808_23_lut (.I0(n2589), .I1(n2589), .I2(n2621), 
            .I3(n28977), .O(n2688)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_23_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1808_23 (.CI(n28977), .I0(n2589), .I1(n2621), .CO(n28978));
    SB_LUT4 mod_5_add_1808_22_lut (.I0(n2590), .I1(n2590), .I2(n2621), 
            .I3(n28976), .O(n2689)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_22_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1808_22 (.CI(n28976), .I0(n2590), .I1(n2621), .CO(n28977));
    SB_CARRY add_21_4 (.CI(n27845), .I0(bit_ctr[2]), .I1(GND_net), .CO(n27846));
    SB_LUT4 mod_5_add_1808_21_lut (.I0(n2591), .I1(n2591), .I2(n2621), 
            .I3(n28975), .O(n2690)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_21_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1808_21 (.CI(n28975), .I0(n2591), .I1(n2621), .CO(n28976));
    SB_LUT4 mod_5_add_1808_20_lut (.I0(n2592), .I1(n2592), .I2(n2621), 
            .I3(n28974), .O(n2691)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_20_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 timer_1524_add_4_33_lut (.I0(GND_net), .I1(GND_net), .I2(timer[31]), 
            .I3(n28465), .O(n133[31])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1524_add_4_33_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 timer_1524_add_4_32_lut (.I0(GND_net), .I1(GND_net), .I2(timer[30]), 
            .I3(n28464), .O(n133[30])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1524_add_4_32_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1808_20 (.CI(n28974), .I0(n2592), .I1(n2621), .CO(n28975));
    SB_LUT4 mod_5_add_1808_19_lut (.I0(n2593), .I1(n2593), .I2(n2621), 
            .I3(n28973), .O(n2692)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_19_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1808_19 (.CI(n28973), .I0(n2593), .I1(n2621), .CO(n28974));
    SB_LUT4 mod_5_add_1808_18_lut (.I0(n2594), .I1(n2594), .I2(n2621), 
            .I3(n28972), .O(n2693)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_18_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1808_18 (.CI(n28972), .I0(n2594), .I1(n2621), .CO(n28973));
    SB_CARRY timer_1524_add_4_32 (.CI(n28464), .I0(GND_net), .I1(timer[30]), 
            .CO(n28465));
    SB_LUT4 timer_1524_add_4_31_lut (.I0(GND_net), .I1(GND_net), .I2(timer[29]), 
            .I3(n28463), .O(n133[29])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1524_add_4_31_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1524_add_4_31 (.CI(n28463), .I0(GND_net), .I1(timer[29]), 
            .CO(n28464));
    SB_LUT4 mod_5_add_1808_17_lut (.I0(n2595), .I1(n2595), .I2(n2621), 
            .I3(n28971), .O(n2694)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_17_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 timer_1524_add_4_30_lut (.I0(GND_net), .I1(GND_net), .I2(timer[28]), 
            .I3(n28462), .O(n133[28])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1524_add_4_30_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1524_add_4_30 (.CI(n28462), .I0(GND_net), .I1(timer[28]), 
            .CO(n28463));
    SB_LUT4 add_21_10_lut (.I0(n1), .I1(bit_ctr[8]), .I2(GND_net), .I3(n27851), 
            .O(n37227)) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_10_lut.LUT_INIT = 16'h8228;
    SB_LUT4 timer_1524_add_4_29_lut (.I0(GND_net), .I1(GND_net), .I2(timer[27]), 
            .I3(n28461), .O(n133[27])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1524_add_4_29_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1808_17 (.CI(n28971), .I0(n2595), .I1(n2621), .CO(n28972));
    SB_CARRY timer_1524_add_4_29 (.CI(n28461), .I0(GND_net), .I1(timer[27]), 
            .CO(n28462));
    SB_LUT4 timer_1524_add_4_28_lut (.I0(GND_net), .I1(GND_net), .I2(timer[26]), 
            .I3(n28460), .O(n133[26])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1524_add_4_28_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1524_add_4_28 (.CI(n28460), .I0(GND_net), .I1(timer[26]), 
            .CO(n28461));
    SB_LUT4 mod_5_add_1808_16_lut (.I0(n2596), .I1(n2596), .I2(n2621), 
            .I3(n28970), .O(n2695)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_16_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1808_16 (.CI(n28970), .I0(n2596), .I1(n2621), .CO(n28971));
    SB_LUT4 timer_1524_add_4_27_lut (.I0(GND_net), .I1(GND_net), .I2(timer[25]), 
            .I3(n28459), .O(n133[25])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1524_add_4_27_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_21_23_lut (.I0(n1), .I1(bit_ctr[21]), .I2(GND_net), .I3(n27864), 
            .O(n37359)) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_23_lut.LUT_INIT = 16'h8228;
    SB_CARRY timer_1524_add_4_27 (.CI(n28459), .I0(GND_net), .I1(timer[25]), 
            .CO(n28460));
    SB_LUT4 mod_5_add_1808_15_lut (.I0(n2597), .I1(n2597), .I2(n2621), 
            .I3(n28969), .O(n2696)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_15_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1808_15 (.CI(n28969), .I0(n2597), .I1(n2621), .CO(n28970));
    SB_LUT4 mod_5_add_1808_14_lut (.I0(n2598), .I1(n2598), .I2(n2621), 
            .I3(n28968), .O(n2697)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_14_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1808_14 (.CI(n28968), .I0(n2598), .I1(n2621), .CO(n28969));
    SB_LUT4 timer_1524_add_4_26_lut (.I0(GND_net), .I1(GND_net), .I2(timer[24]), 
            .I3(n28458), .O(n133[24])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1524_add_4_26_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1524_add_4_26 (.CI(n28458), .I0(GND_net), .I1(timer[24]), 
            .CO(n28459));
    SB_LUT4 timer_1524_add_4_25_lut (.I0(GND_net), .I1(GND_net), .I2(timer[23]), 
            .I3(n28457), .O(n133[23])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1524_add_4_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1524_add_4_25 (.CI(n28457), .I0(GND_net), .I1(timer[23]), 
            .CO(n28458));
    SB_CARRY mod_5_add_1004_10 (.CI(n28778), .I0(n1402), .I1(n1433), .CO(n28779));
    SB_LUT4 mod_5_add_1808_13_lut (.I0(n2599), .I1(n2599), .I2(n2621), 
            .I3(n28967), .O(n2698)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_13_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY add_21_10 (.CI(n27851), .I0(bit_ctr[8]), .I1(GND_net), .CO(n27852));
    SB_LUT4 timer_1524_add_4_24_lut (.I0(GND_net), .I1(GND_net), .I2(timer[22]), 
            .I3(n28456), .O(n133[22])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1524_add_4_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1808_13 (.CI(n28967), .I0(n2599), .I1(n2621), .CO(n28968));
    SB_LUT4 mod_5_add_1004_10_lut (.I0(n1402), .I1(n1402), .I2(n1433), 
            .I3(n28778), .O(n1501)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1004_10_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1808_12_lut (.I0(n2600), .I1(n2600), .I2(n2621), 
            .I3(n28966), .O(n2699)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_12_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1004_11 (.CI(n28779), .I0(n1401), .I1(n1433), .CO(n28780));
    SB_CARRY timer_1524_add_4_24 (.CI(n28456), .I0(GND_net), .I1(timer[22]), 
            .CO(n28457));
    SB_LUT4 timer_1524_add_4_23_lut (.I0(GND_net), .I1(GND_net), .I2(timer[21]), 
            .I3(n28455), .O(n133[21])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1524_add_4_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1808_12 (.CI(n28966), .I0(n2600), .I1(n2621), .CO(n28967));
    SB_CARRY add_21_23 (.CI(n27864), .I0(bit_ctr[21]), .I1(GND_net), .CO(n27865));
    SB_LUT4 mod_5_add_1808_11_lut (.I0(n2601), .I1(n2601), .I2(n2621), 
            .I3(n28965), .O(n2700)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_11_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY timer_1524_add_4_23 (.CI(n28455), .I0(GND_net), .I1(timer[21]), 
            .CO(n28456));
    SB_LUT4 timer_1524_add_4_22_lut (.I0(GND_net), .I1(GND_net), .I2(timer[20]), 
            .I3(n28454), .O(n133[20])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1524_add_4_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1524_add_4_22 (.CI(n28454), .I0(GND_net), .I1(timer[20]), 
            .CO(n28455));
    SB_LUT4 sub_14_add_2_33_lut (.I0(one_wire_N_613[21]), .I1(timer[31]), 
            .I2(n51[31]), .I3(n27970), .O(n29_adj_4675)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_33_lut.LUT_INIT = 16'hebbe;
    SB_LUT4 timer_1524_add_4_21_lut (.I0(GND_net), .I1(GND_net), .I2(timer[19]), 
            .I3(n28453), .O(n133[19])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1524_add_4_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1808_11 (.CI(n28965), .I0(n2601), .I1(n2621), .CO(n28966));
    SB_CARRY timer_1524_add_4_21 (.CI(n28453), .I0(GND_net), .I1(timer[19]), 
            .CO(n28454));
    SB_LUT4 mod_5_add_1808_10_lut (.I0(n2602), .I1(n2602), .I2(n2621), 
            .I3(n28964), .O(n2701)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_10_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1004_11_lut (.I0(n1401), .I1(n1401), .I2(n1433), 
            .I3(n28779), .O(n1500)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1004_11_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 timer_1524_add_4_20_lut (.I0(GND_net), .I1(GND_net), .I2(timer[18]), 
            .I3(n28452), .O(n133[18])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1524_add_4_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1524_add_4_20 (.CI(n28452), .I0(GND_net), .I1(timer[18]), 
            .CO(n28453));
    SB_CARRY mod_5_add_1808_10 (.CI(n28964), .I0(n2602), .I1(n2621), .CO(n28965));
    SB_LUT4 add_21_22_lut (.I0(n1), .I1(bit_ctr[20]), .I2(GND_net), .I3(n27863), 
            .O(n37360)) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_22_lut.LUT_INIT = 16'h8228;
    SB_LUT4 mod_5_add_1004_12_lut (.I0(n1400), .I1(n1400), .I2(n1433), 
            .I3(n28780), .O(n1499)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1004_12_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 add_21_3_lut (.I0(n1), .I1(bit_ctr[1]), .I2(GND_net), .I3(n27844), 
            .O(n37241)) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_3_lut.LUT_INIT = 16'h8228;
    SB_LUT4 timer_1524_add_4_19_lut (.I0(GND_net), .I1(GND_net), .I2(timer[17]), 
            .I3(n28451), .O(n133[17])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1524_add_4_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1524_add_4_19 (.CI(n28451), .I0(GND_net), .I1(timer[17]), 
            .CO(n28452));
    SB_LUT4 timer_1524_add_4_18_lut (.I0(GND_net), .I1(GND_net), .I2(timer[16]), 
            .I3(n28450), .O(n133[16])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1524_add_4_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_21_9_lut (.I0(n1), .I1(bit_ctr[7]), .I2(GND_net), .I3(n27850), 
            .O(n37228)) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_9_lut.LUT_INIT = 16'h8228;
    SB_LUT4 mod_5_add_1808_9_lut (.I0(n2603), .I1(n2603), .I2(n2621), 
            .I3(n28963), .O(n2702)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_9_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1071_2 (.CI(VCC_net), .I0(bit_ctr[20]), .I1(n38250), 
            .CO(n28781));
    SB_LUT4 mod_5_add_1071_2_lut (.I0(bit_ctr[20]), .I1(bit_ctr[20]), .I2(n38250), 
            .I3(VCC_net), .O(n1609)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1071_2_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY timer_1524_add_4_18 (.CI(n28450), .I0(GND_net), .I1(timer[16]), 
            .CO(n28451));
    SB_CARRY mod_5_add_1808_9 (.CI(n28963), .I0(n2603), .I1(n2621), .CO(n28964));
    SB_LUT4 timer_1524_add_4_17_lut (.I0(GND_net), .I1(GND_net), .I2(timer[15]), 
            .I3(n28449), .O(n133[15])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1524_add_4_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1524_add_4_17 (.CI(n28449), .I0(GND_net), .I1(timer[15]), 
            .CO(n28450));
    SB_LUT4 timer_1524_add_4_16_lut (.I0(GND_net), .I1(GND_net), .I2(timer[14]), 
            .I3(n28448), .O(n133[14])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1524_add_4_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1524_add_4_16 (.CI(n28448), .I0(GND_net), .I1(timer[14]), 
            .CO(n28449));
    SB_LUT4 timer_1524_add_4_15_lut (.I0(GND_net), .I1(GND_net), .I2(timer[13]), 
            .I3(n28447), .O(n133[13])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1524_add_4_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1524_add_4_15 (.CI(n28447), .I0(GND_net), .I1(timer[13]), 
            .CO(n28448));
    SB_LUT4 timer_1524_add_4_14_lut (.I0(GND_net), .I1(GND_net), .I2(timer[12]), 
            .I3(n28446), .O(n133[12])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1524_add_4_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1071_3 (.CI(n28781), .I0(n1509), .I1(n38250), .CO(n28782));
    SB_LUT4 mod_5_add_1808_8_lut (.I0(n2604), .I1(n2604), .I2(n2621), 
            .I3(n28962), .O(n2703)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_8_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY timer_1524_add_4_14 (.CI(n28446), .I0(GND_net), .I1(timer[12]), 
            .CO(n28447));
    SB_LUT4 timer_1524_add_4_13_lut (.I0(GND_net), .I1(GND_net), .I2(timer[11]), 
            .I3(n28445), .O(n133[11])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1524_add_4_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1524_add_4_13 (.CI(n28445), .I0(GND_net), .I1(timer[11]), 
            .CO(n28446));
    SB_CARRY mod_5_add_1808_8 (.CI(n28962), .I0(n2604), .I1(n2621), .CO(n28963));
    SB_CARRY add_21_9 (.CI(n27850), .I0(bit_ctr[7]), .I1(GND_net), .CO(n27851));
    SB_CARRY mod_5_add_1138_5 (.CI(n28794), .I0(n1607), .I1(n1631), .CO(n28795));
    SB_LUT4 timer_1524_add_4_12_lut (.I0(GND_net), .I1(GND_net), .I2(timer[10]), 
            .I3(n28444), .O(n133[10])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1524_add_4_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1524_add_4_12 (.CI(n28444), .I0(GND_net), .I1(timer[10]), 
            .CO(n28445));
    SB_LUT4 timer_1524_add_4_11_lut (.I0(GND_net), .I1(GND_net), .I2(timer[9]), 
            .I3(n28443), .O(n133[9])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1524_add_4_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1524_add_4_11 (.CI(n28443), .I0(GND_net), .I1(timer[9]), 
            .CO(n28444));
    SB_LUT4 mod_5_add_1808_7_lut (.I0(n2605), .I1(n2605), .I2(n2621), 
            .I3(n28961), .O(n2704)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_7_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1808_7 (.CI(n28961), .I0(n2605), .I1(n2621), .CO(n28962));
    SB_LUT4 timer_1524_add_4_10_lut (.I0(GND_net), .I1(GND_net), .I2(timer[8]), 
            .I3(n28442), .O(n133[8])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1524_add_4_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1524_add_4_10 (.CI(n28442), .I0(GND_net), .I1(timer[8]), 
            .CO(n28443));
    SB_LUT4 timer_1524_add_4_9_lut (.I0(GND_net), .I1(GND_net), .I2(timer[7]), 
            .I3(n28441), .O(n133[7])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1524_add_4_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1524_add_4_9 (.CI(n28441), .I0(GND_net), .I1(timer[7]), 
            .CO(n28442));
    SB_LUT4 mod_5_add_1808_6_lut (.I0(n2606), .I1(n2606), .I2(n2621), 
            .I3(n28960), .O(n2705)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_6_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 timer_1524_add_4_8_lut (.I0(GND_net), .I1(GND_net), .I2(timer[6]), 
            .I3(n28440), .O(n133[6])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1524_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1524_add_4_8 (.CI(n28440), .I0(GND_net), .I1(timer[6]), 
            .CO(n28441));
    SB_CARRY add_21_22 (.CI(n27863), .I0(bit_ctr[20]), .I1(GND_net), .CO(n27864));
    SB_LUT4 timer_1524_add_4_7_lut (.I0(GND_net), .I1(GND_net), .I2(timer[5]), 
            .I3(n28439), .O(n133[5])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1524_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1524_add_4_7 (.CI(n28439), .I0(GND_net), .I1(timer[5]), 
            .CO(n28440));
    SB_LUT4 timer_1524_add_4_6_lut (.I0(GND_net), .I1(GND_net), .I2(timer[4]), 
            .I3(n28438), .O(n133[4])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1524_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1808_6 (.CI(n28960), .I0(n2606), .I1(n2621), .CO(n28961));
    SB_CARRY timer_1524_add_4_6 (.CI(n28438), .I0(GND_net), .I1(timer[4]), 
            .CO(n28439));
    SB_LUT4 timer_1524_add_4_5_lut (.I0(GND_net), .I1(GND_net), .I2(timer[3]), 
            .I3(n28437), .O(n133[3])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1524_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1524_add_4_5 (.CI(n28437), .I0(GND_net), .I1(timer[3]), 
            .CO(n28438));
    SB_LUT4 mod_5_add_1808_5_lut (.I0(n2607), .I1(n2607), .I2(n2621), 
            .I3(n28959), .O(n2706)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_5_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 timer_1524_add_4_4_lut (.I0(GND_net), .I1(GND_net), .I2(timer[2]), 
            .I3(n28436), .O(n133[2])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1524_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1808_5 (.CI(n28959), .I0(n2607), .I1(n2621), .CO(n28960));
    SB_LUT4 mod_5_add_1808_4_lut (.I0(n2608), .I1(n2608), .I2(n2621), 
            .I3(n28958), .O(n2707)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_4_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY timer_1524_add_4_4 (.CI(n28436), .I0(GND_net), .I1(timer[2]), 
            .CO(n28437));
    SB_LUT4 timer_1524_add_4_3_lut (.I0(GND_net), .I1(GND_net), .I2(timer[1]), 
            .I3(n28435), .O(n133[1])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1524_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1524_add_4_3 (.CI(n28435), .I0(GND_net), .I1(timer[1]), 
            .CO(n28436));
    SB_LUT4 timer_1524_add_4_2_lut (.I0(GND_net), .I1(GND_net), .I2(timer[0]), 
            .I3(VCC_net), .O(n133[0])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1524_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1524_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(timer[0]), 
            .CO(n28435));
    SB_CARRY mod_5_add_1808_4 (.CI(n28958), .I0(n2608), .I1(n2621), .CO(n28959));
    SB_LUT4 mod_5_add_1808_3_lut (.I0(n2609), .I1(n2609), .I2(n38249), 
            .I3(n28957), .O(n2708)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_3_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 add_21_21_lut (.I0(n1), .I1(bit_ctr[19]), .I2(GND_net), .I3(n27862), 
            .O(n37361)) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_21_lut.LUT_INIT = 16'h8228;
    SB_CARRY mod_5_add_1808_3 (.CI(n28957), .I0(n2609), .I1(n38249), .CO(n28958));
    SB_LUT4 mod_5_add_1808_2_lut (.I0(bit_ctr[9]), .I1(bit_ctr[9]), .I2(n38249), 
            .I3(VCC_net), .O(n2709)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_2_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1808_2 (.CI(VCC_net), .I0(bit_ctr[9]), .I1(n38249), 
            .CO(n28957));
    SB_LUT4 mod_5_add_1741_23_lut (.I0(n2489), .I1(n2489), .I2(n2522), 
            .I3(n28956), .O(n2588)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_23_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1741_22_lut (.I0(n2490), .I1(n2490), .I2(n2522), 
            .I3(n28955), .O(n2589)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_22_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1741_22 (.CI(n28955), .I0(n2490), .I1(n2522), .CO(n28956));
    SB_LUT4 mod_5_add_1741_21_lut (.I0(n2491), .I1(n2491), .I2(n2522), 
            .I3(n28954), .O(n2590)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_21_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1741_21 (.CI(n28954), .I0(n2491), .I1(n2522), .CO(n28955));
    SB_LUT4 mod_5_add_1741_20_lut (.I0(n2492), .I1(n2492), .I2(n2522), 
            .I3(n28953), .O(n2591)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_20_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1741_20 (.CI(n28953), .I0(n2492), .I1(n2522), .CO(n28954));
    SB_LUT4 i31527_2_lut (.I0(n2_adj_4768), .I1(n971[28]), .I2(GND_net), 
            .I3(GND_net), .O(n1007));   // verilog/neopixel.v(22[26:36])
    defparam i31527_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 mod_5_add_1741_19_lut (.I0(n2493), .I1(n2493), .I2(n2522), 
            .I3(n28952), .O(n2592)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_19_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 sub_14_inv_0_i15_1_lut (.I0(\neo_pixel_transmitter.t0 [14]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n51[14]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i15_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY mod_5_add_1741_19 (.CI(n28952), .I0(n2493), .I1(n2522), .CO(n28953));
    SB_LUT4 mod_5_add_1741_18_lut (.I0(n2494), .I1(n2494), .I2(n2522), 
            .I3(n28951), .O(n2593)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_18_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1741_18 (.CI(n28951), .I0(n2494), .I1(n2522), .CO(n28952));
    SB_LUT4 mod_5_add_1741_17_lut (.I0(n2495), .I1(n2495), .I2(n2522), 
            .I3(n28950), .O(n2594)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_17_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1741_17 (.CI(n28950), .I0(n2495), .I1(n2522), .CO(n28951));
    SB_LUT4 mod_5_add_1741_16_lut (.I0(n2496), .I1(n2496), .I2(n2522), 
            .I3(n28949), .O(n2595)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_16_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1741_16 (.CI(n28949), .I0(n2496), .I1(n2522), .CO(n28950));
    SB_LUT4 mod_5_add_1741_15_lut (.I0(n2497), .I1(n2497), .I2(n2522), 
            .I3(n28948), .O(n2596)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_15_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1741_15 (.CI(n28948), .I0(n2497), .I1(n2522), .CO(n28949));
    SB_LUT4 mod_5_add_1741_14_lut (.I0(n2498), .I1(n2498), .I2(n2522), 
            .I3(n28947), .O(n2597)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_14_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1741_14 (.CI(n28947), .I0(n2498), .I1(n2522), .CO(n28948));
    SB_LUT4 mod_5_add_1741_13_lut (.I0(n2499), .I1(n2499), .I2(n2522), 
            .I3(n28946), .O(n2598)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_13_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1741_13 (.CI(n28946), .I0(n2499), .I1(n2522), .CO(n28947));
    SB_LUT4 mod_5_add_1741_12_lut (.I0(n2500), .I1(n2500), .I2(n2522), 
            .I3(n28945), .O(n2599)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_12_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1741_12 (.CI(n28945), .I0(n2500), .I1(n2522), .CO(n28946));
    SB_LUT4 mod_5_add_1741_11_lut (.I0(n2501), .I1(n2501), .I2(n2522), 
            .I3(n28944), .O(n2600)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_11_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1741_11 (.CI(n28944), .I0(n2501), .I1(n2522), .CO(n28945));
    SB_LUT4 mod_5_add_1741_10_lut (.I0(n2502), .I1(n2502), .I2(n2522), 
            .I3(n28943), .O(n2601)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_10_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1741_10 (.CI(n28943), .I0(n2502), .I1(n2522), .CO(n28944));
    SB_LUT4 mod_5_add_1741_9_lut (.I0(n2503), .I1(n2503), .I2(n2522), 
            .I3(n28942), .O(n2602)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_9_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i31529_2_lut (.I0(n2_adj_4768), .I1(n971[29]), .I2(GND_net), 
            .I3(GND_net), .O(n1006));   // verilog/neopixel.v(22[26:36])
    defparam i31529_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 sub_14_add_2_32_lut (.I0(one_wire_N_613[29]), .I1(timer[30]), 
            .I2(n51[30]), .I3(n27969), .O(n28_adj_4673)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_32_lut.LUT_INIT = 16'hebbe;
    SB_CARRY mod_5_add_1741_9 (.CI(n28942), .I0(n2503), .I1(n2522), .CO(n28943));
    SB_LUT4 mod_5_add_1741_8_lut (.I0(n2504), .I1(n2504), .I2(n2522), 
            .I3(n28941), .O(n2603)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_8_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1138_4_lut (.I0(n1608), .I1(n1608), .I2(n1631), 
            .I3(n28793), .O(n1707)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1138_4_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1741_8 (.CI(n28941), .I0(n2504), .I1(n2522), .CO(n28942));
    SB_LUT4 mod_5_add_1741_7_lut (.I0(n2505), .I1(n2505), .I2(n2522), 
            .I3(n28940), .O(n2604)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_7_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1138_4 (.CI(n28793), .I0(n1608), .I1(n1631), .CO(n28794));
    SB_LUT4 mod_5_add_1138_3_lut (.I0(n1609), .I1(n1609), .I2(n38247), 
            .I3(n28792), .O(n1708)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1138_3_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1741_7 (.CI(n28940), .I0(n2505), .I1(n2522), .CO(n28941));
    SB_CARRY mod_5_add_1138_3 (.CI(n28792), .I0(n1609), .I1(n38247), .CO(n28793));
    SB_LUT4 mod_5_add_1741_6_lut (.I0(n2506), .I1(n2506), .I2(n2522), 
            .I3(n28939), .O(n2605)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_6_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1138_2_lut (.I0(bit_ctr[19]), .I1(bit_ctr[19]), .I2(n38247), 
            .I3(VCC_net), .O(n1709)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1138_2_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1741_6 (.CI(n28939), .I0(n2506), .I1(n2522), .CO(n28940));
    SB_CARRY mod_5_add_1138_2 (.CI(VCC_net), .I0(bit_ctr[19]), .I1(n38247), 
            .CO(n28792));
    SB_LUT4 mod_5_add_1741_5_lut (.I0(n2507), .I1(n2507), .I2(n2522), 
            .I3(n28938), .O(n2606)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_5_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1071_13_lut (.I0(n1499), .I1(n1499), .I2(n1532), 
            .I3(n28791), .O(n1598)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1071_13_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1741_5 (.CI(n28938), .I0(n2507), .I1(n2522), .CO(n28939));
    SB_LUT4 mod_5_add_1741_4_lut (.I0(n2508), .I1(n2508), .I2(n2522), 
            .I3(n28937), .O(n2607)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_4_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1071_12_lut (.I0(n1500), .I1(n1500), .I2(n1532), 
            .I3(n28790), .O(n1599)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1071_12_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1741_4 (.CI(n28937), .I0(n2508), .I1(n2522), .CO(n28938));
    SB_LUT4 mod_5_add_1741_3_lut (.I0(n2509), .I1(n2509), .I2(n38251), 
            .I3(n28936), .O(n2608)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_3_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1071_12 (.CI(n28790), .I0(n1500), .I1(n1532), .CO(n28791));
    SB_LUT4 mod_5_add_1071_11_lut (.I0(n1501), .I1(n1501), .I2(n1532), 
            .I3(n28789), .O(n1600)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1071_11_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1741_3 (.CI(n28936), .I0(n2509), .I1(n38251), .CO(n28937));
    SB_CARRY mod_5_add_1071_11 (.CI(n28789), .I0(n1501), .I1(n1532), .CO(n28790));
    SB_LUT4 mod_5_add_1741_2_lut (.I0(bit_ctr[10]), .I1(bit_ctr[10]), .I2(n38251), 
            .I3(VCC_net), .O(n2609)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_2_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 mod_5_add_1071_10_lut (.I0(n1502), .I1(n1502), .I2(n1532), 
            .I3(n28788), .O(n1601)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1071_10_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_i672_3_lut (.I0(n906), .I1(n971[30]), .I2(n2_adj_4768), 
            .I3(GND_net), .O(n1005));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i672_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY mod_5_add_1741_2 (.CI(VCC_net), .I0(bit_ctr[10]), .I1(n38251), 
            .CO(n28936));
    SB_CARRY mod_5_add_1071_10 (.CI(n28788), .I0(n1502), .I1(n1532), .CO(n28789));
    SB_LUT4 mod_5_add_1071_9_lut (.I0(n1503), .I1(n1503), .I2(n1532), 
            .I3(n28787), .O(n1602)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1071_9_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1674_22_lut (.I0(n2390), .I1(n2390), .I2(n2423), 
            .I3(n28935), .O(n2489)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_22_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY sub_14_add_2_32 (.CI(n27969), .I0(timer[30]), .I1(n51[30]), 
            .CO(n27970));
    SB_LUT4 sub_14_add_2_31_lut (.I0(GND_net), .I1(timer[29]), .I2(n51[29]), 
            .I3(n27968), .O(one_wire_N_613[29])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_31_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_1674_21_lut (.I0(n2391), .I1(n2391), .I2(n2423), 
            .I3(n28934), .O(n2490)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_21_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1674_21 (.CI(n28934), .I0(n2391), .I1(n2423), .CO(n28935));
    SB_CARRY mod_5_add_1071_9 (.CI(n28787), .I0(n1503), .I1(n1532), .CO(n28788));
    SB_LUT4 mod_5_add_1071_8_lut (.I0(n1504), .I1(n1504), .I2(n1532), 
            .I3(n28786), .O(n1603)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1071_8_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1071_8 (.CI(n28786), .I0(n1504), .I1(n1532), .CO(n28787));
    SB_CARRY add_21_21 (.CI(n27862), .I0(bit_ctr[19]), .I1(GND_net), .CO(n27863));
    SB_LUT4 mod_5_add_1674_20_lut (.I0(n2392), .I1(n2392), .I2(n2423), 
            .I3(n28933), .O(n2491)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_20_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i30947_3_lut (.I0(n14844), .I1(bit_ctr[27]), .I2(n838), .I3(GND_net), 
            .O(n17391));
    defparam i30947_3_lut.LUT_INIT = 16'h5959;
    SB_LUT4 mod_5_add_1071_7_lut (.I0(n1505), .I1(n1505), .I2(n1532), 
            .I3(n28785), .O(n1604)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1071_7_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1071_7 (.CI(n28785), .I0(n1505), .I1(n1532), .CO(n28786));
    SB_CARRY mod_5_add_1674_20 (.CI(n28933), .I0(n2392), .I1(n2423), .CO(n28934));
    SB_LUT4 mod_5_add_1071_6_lut (.I0(n1506), .I1(n1506), .I2(n1532), 
            .I3(n28784), .O(n1605)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1071_6_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1674_19_lut (.I0(n2393), .I1(n2393), .I2(n2423), 
            .I3(n28932), .O(n2492)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_19_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 add_21_20_lut (.I0(n1), .I1(bit_ctr[18]), .I2(GND_net), .I3(n27861), 
            .O(n37362)) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_20_lut.LUT_INIT = 16'h8228;
    SB_CARRY sub_14_add_2_31 (.CI(n27968), .I0(timer[29]), .I1(n51[29]), 
            .CO(n27969));
    SB_LUT4 sub_14_add_2_30_lut (.I0(one_wire_N_613[24]), .I1(timer[28]), 
            .I2(n51[28]), .I3(n27967), .O(n26_adj_4672)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_30_lut.LUT_INIT = 16'hebbe;
    SB_CARRY mod_5_add_1071_6 (.CI(n28784), .I0(n1506), .I1(n1532), .CO(n28785));
    SB_LUT4 mod_5_add_1071_5_lut (.I0(n1507), .I1(n1507), .I2(n1532), 
            .I3(n28783), .O(n1606)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1071_5_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 add_21_8_lut (.I0(n1), .I1(bit_ctr[6]), .I2(GND_net), .I3(n27849), 
            .O(n37229)) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_8_lut.LUT_INIT = 16'h8228;
    SB_CARRY mod_5_add_1071_5 (.CI(n28783), .I0(n1507), .I1(n1532), .CO(n28784));
    SB_LUT4 mod_5_add_1071_4_lut (.I0(n1508), .I1(n1508), .I2(n1532), 
            .I3(n28782), .O(n1607)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1071_4_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i2_2_lut_3_lut (.I0(\state[0] ), .I1(n25098), .I2(\neo_pixel_transmitter.done ), 
            .I3(GND_net), .O(n35088));   // verilog/neopixel.v(36[4] 116[11])
    defparam i2_2_lut_3_lut.LUT_INIT = 16'hfbfb;
    SB_CARRY mod_5_add_1674_19 (.CI(n28932), .I0(n2393), .I1(n2423), .CO(n28933));
    SB_CARRY mod_5_add_1071_4 (.CI(n28782), .I0(n1508), .I1(n1532), .CO(n28783));
    SB_LUT4 mod_5_add_1071_3_lut (.I0(n1509), .I1(n1509), .I2(n38250), 
            .I3(n28781), .O(n1608)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1071_3_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY add_21_20 (.CI(n27861), .I0(bit_ctr[18]), .I1(GND_net), .CO(n27862));
    SB_LUT4 mod_5_add_1674_18_lut (.I0(n2394), .I1(n2394), .I2(n2423), 
            .I3(n28931), .O(n2493)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_18_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1674_18 (.CI(n28931), .I0(n2394), .I1(n2423), .CO(n28932));
    SB_LUT4 mod_5_add_1674_17_lut (.I0(n2395), .I1(n2395), .I2(n2423), 
            .I3(n28930), .O(n2494)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_17_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1674_17 (.CI(n28930), .I0(n2395), .I1(n2423), .CO(n28931));
    SB_LUT4 mod_5_add_1674_16_lut (.I0(n2396), .I1(n2396), .I2(n2423), 
            .I3(n28929), .O(n2495)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_16_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1674_16 (.CI(n28929), .I0(n2396), .I1(n2423), .CO(n28930));
    SB_CARRY add_21_3 (.CI(n27844), .I0(bit_ctr[1]), .I1(GND_net), .CO(n27845));
    SB_LUT4 mod_5_add_1674_15_lut (.I0(n2397), .I1(n2397), .I2(n2423), 
            .I3(n28928), .O(n2496)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_15_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY sub_14_add_2_30 (.CI(n27967), .I0(timer[28]), .I1(n51[28]), 
            .CO(n27968));
    SB_CARRY mod_5_add_1674_15 (.CI(n28928), .I0(n2397), .I1(n2423), .CO(n28929));
    SB_LUT4 mod_5_add_1674_14_lut (.I0(n2398), .I1(n2398), .I2(n2423), 
            .I3(n28927), .O(n2497)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_14_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY add_21_8 (.CI(n27849), .I0(bit_ctr[6]), .I1(GND_net), .CO(n27850));
    SB_LUT4 add_21_7_lut (.I0(n1), .I1(bit_ctr[5]), .I2(GND_net), .I3(n27848), 
            .O(n37230)) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_7_lut.LUT_INIT = 16'h8228;
    SB_LUT4 add_21_19_lut (.I0(n1), .I1(bit_ctr[17]), .I2(GND_net), .I3(n27860), 
            .O(n37245)) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_19_lut.LUT_INIT = 16'h8228;
    SB_CARRY mod_5_add_1674_14 (.CI(n28927), .I0(n2398), .I1(n2423), .CO(n28928));
    SB_CARRY add_21_19 (.CI(n27860), .I0(bit_ctr[17]), .I1(GND_net), .CO(n27861));
    SB_LUT4 mod_5_add_1674_13_lut (.I0(n2399), .I1(n2399), .I2(n2423), 
            .I3(n28926), .O(n2498)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_13_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1674_13 (.CI(n28926), .I0(n2399), .I1(n2423), .CO(n28927));
    SB_LUT4 sub_14_add_2_29_lut (.I0(one_wire_N_613[26]), .I1(timer[27]), 
            .I2(n51[27]), .I3(n27966), .O(n21_adj_4661)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_29_lut.LUT_INIT = 16'hebbe;
    SB_LUT4 mod_5_add_1674_12_lut (.I0(n2400), .I1(n2400), .I2(n2423), 
            .I3(n28925), .O(n2499)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_12_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1674_12 (.CI(n28925), .I0(n2400), .I1(n2423), .CO(n28926));
    SB_LUT4 mod_5_add_1674_11_lut (.I0(n2401), .I1(n2401), .I2(n2423), 
            .I3(n28924), .O(n2500)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_11_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1674_11 (.CI(n28924), .I0(n2401), .I1(n2423), .CO(n28925));
    SB_CARRY sub_14_add_2_29 (.CI(n27966), .I0(timer[27]), .I1(n51[27]), 
            .CO(n27967));
    SB_LUT4 sub_14_add_2_28_lut (.I0(GND_net), .I1(timer[26]), .I2(n51[26]), 
            .I3(n27965), .O(one_wire_N_613[26])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_28_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_1674_10_lut (.I0(n2402), .I1(n2402), .I2(n2423), 
            .I3(n28923), .O(n2501)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_10_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY sub_14_add_2_28 (.CI(n27965), .I0(timer[26]), .I1(n51[26]), 
            .CO(n27966));
    SB_CARRY mod_5_add_1674_10 (.CI(n28923), .I0(n2402), .I1(n2423), .CO(n28924));
    SB_LUT4 i3_4_lut_4_lut (.I0(n33673), .I1(n14844), .I2(n807), .I3(bit_ctr[27]), 
            .O(n838));
    defparam i3_4_lut_4_lut.LUT_INIT = 16'h0405;
    SB_LUT4 mod_5_add_1674_9_lut (.I0(n2403), .I1(n2403), .I2(n2423), 
            .I3(n28922), .O(n2502)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_9_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 sub_14_add_2_27_lut (.I0(GND_net), .I1(timer[25]), .I2(n51[25]), 
            .I3(n27964), .O(one_wire_N_613[25])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_27_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1674_9 (.CI(n28922), .I0(n2403), .I1(n2423), .CO(n28923));
    SB_CARRY sub_14_add_2_27 (.CI(n27964), .I0(timer[25]), .I1(n51[25]), 
            .CO(n27965));
    SB_LUT4 sub_14_add_2_26_lut (.I0(GND_net), .I1(timer[24]), .I2(n51[24]), 
            .I3(n27963), .O(one_wire_N_613[24])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_26_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_21_18_lut (.I0(n1), .I1(bit_ctr[16]), .I2(GND_net), .I3(n27859), 
            .O(n37363)) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_18_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_21_18 (.CI(n27859), .I0(bit_ctr[16]), .I1(GND_net), .CO(n27860));
    SB_CARRY sub_14_add_2_26 (.CI(n27963), .I0(timer[24]), .I1(n51[24]), 
            .CO(n27964));
    SB_LUT4 mod_5_add_1674_8_lut (.I0(n2404), .I1(n2404), .I2(n2423), 
            .I3(n28921), .O(n2503)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_8_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1674_8 (.CI(n28921), .I0(n2404), .I1(n2423), .CO(n28922));
    SB_LUT4 add_21_17_lut (.I0(n1), .I1(bit_ctr[15]), .I2(GND_net), .I3(n27858), 
            .O(n37364)) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_17_lut.LUT_INIT = 16'h8228;
    SB_LUT4 mod_5_add_1674_7_lut (.I0(n2405), .I1(n2405), .I2(n2423), 
            .I3(n28920), .O(n2504)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_7_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1674_7 (.CI(n28920), .I0(n2405), .I1(n2423), .CO(n28921));
    SB_LUT4 sub_14_add_2_25_lut (.I0(GND_net), .I1(timer[23]), .I2(n51[23]), 
            .I3(n27962), .O(one_wire_N_613[23])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_1674_6_lut (.I0(n2406), .I1(n2406), .I2(n2423), 
            .I3(n28919), .O(n2505)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_6_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1674_6 (.CI(n28919), .I0(n2406), .I1(n2423), .CO(n28920));
    SB_DFF bit_ctr_i0_i0 (.Q(bit_ctr[0]), .C(clk32MHz), .D(n31591));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF bit_ctr_i0_i30 (.Q(bit_ctr[30]), .C(clk32MHz), .D(n31589));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF bit_ctr_i0_i29 (.Q(bit_ctr[29]), .C(clk32MHz), .D(n31587));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF bit_ctr_i0_i28 (.Q(bit_ctr[28]), .C(clk32MHz), .D(n31585));   // verilog/neopixel.v(35[12] 117[6])
    SB_CARRY add_21_17 (.CI(n27858), .I0(bit_ctr[15]), .I1(GND_net), .CO(n27859));
    SB_LUT4 add_21_2_lut (.I0(n1), .I1(bit_ctr[0]), .I2(GND_net), .I3(VCC_net), 
            .O(n37252)) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_2_lut.LUT_INIT = 16'h8228;
    SB_DFF bit_ctr_i0_i27 (.Q(bit_ctr[27]), .C(clk32MHz), .D(n31583));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF bit_ctr_i0_i26 (.Q(bit_ctr[26]), .C(clk32MHz), .D(n31577));   // verilog/neopixel.v(35[12] 117[6])
    SB_LUT4 add_21_16_lut (.I0(n1), .I1(bit_ctr[14]), .I2(GND_net), .I3(n27857), 
            .O(n37365)) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_16_lut.LUT_INIT = 16'h8228;
    SB_DFF bit_ctr_i0_i25 (.Q(bit_ctr[25]), .C(clk32MHz), .D(n31575));   // verilog/neopixel.v(35[12] 117[6])
    SB_LUT4 mod_5_add_1674_5_lut (.I0(n2407), .I1(n2407), .I2(n2423), 
            .I3(n28918), .O(n2506)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_5_lut.LUT_INIT = 16'hCA3A;
    SB_DFF bit_ctr_i0_i24 (.Q(bit_ctr[24]), .C(clk32MHz), .D(n31573));   // verilog/neopixel.v(35[12] 117[6])
    SB_CARRY mod_5_add_1674_5 (.CI(n28918), .I0(n2407), .I1(n2423), .CO(n28919));
    SB_DFF bit_ctr_i0_i23 (.Q(bit_ctr[23]), .C(clk32MHz), .D(n31571));   // verilog/neopixel.v(35[12] 117[6])
    SB_LUT4 mod_5_add_1674_4_lut (.I0(n2408), .I1(n2408), .I2(n2423), 
            .I3(n28917), .O(n2507)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_4_lut.LUT_INIT = 16'hCA3A;
    SB_DFF bit_ctr_i0_i22 (.Q(bit_ctr[22]), .C(clk32MHz), .D(n31569));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF bit_ctr_i0_i21 (.Q(bit_ctr[21]), .C(clk32MHz), .D(n31567));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF bit_ctr_i0_i20 (.Q(bit_ctr[20]), .C(clk32MHz), .D(n31565));   // verilog/neopixel.v(35[12] 117[6])
    SB_CARRY add_21_16 (.CI(n27857), .I0(bit_ctr[14]), .I1(GND_net), .CO(n27858));
    SB_DFF bit_ctr_i0_i19 (.Q(bit_ctr[19]), .C(clk32MHz), .D(n31563));   // verilog/neopixel.v(35[12] 117[6])
    SB_CARRY mod_5_add_1674_4 (.CI(n28917), .I0(n2408), .I1(n2423), .CO(n28918));
    SB_DFF bit_ctr_i0_i18 (.Q(bit_ctr[18]), .C(clk32MHz), .D(n31561));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF bit_ctr_i0_i17 (.Q(bit_ctr[17]), .C(clk32MHz), .D(n31559));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF bit_ctr_i0_i16 (.Q(bit_ctr[16]), .C(clk32MHz), .D(n31557));   // verilog/neopixel.v(35[12] 117[6])
    SB_LUT4 add_21_15_lut (.I0(n1), .I1(bit_ctr[13]), .I2(GND_net), .I3(n27856), 
            .O(n37368)) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_15_lut.LUT_INIT = 16'h8228;
    SB_DFF bit_ctr_i0_i15 (.Q(bit_ctr[15]), .C(clk32MHz), .D(n31555));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF bit_ctr_i0_i14 (.Q(bit_ctr[14]), .C(clk32MHz), .D(n31553));   // verilog/neopixel.v(35[12] 117[6])
    SB_LUT4 mod_5_i605_3_lut (.I0(n807), .I1(n60), .I2(n838), .I3(GND_net), 
            .O(n906));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i605_3_lut.LUT_INIT = 16'ha9a9;
    SB_DFF bit_ctr_i0_i13 (.Q(bit_ctr[13]), .C(clk32MHz), .D(n31551));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF bit_ctr_i0_i12 (.Q(bit_ctr[12]), .C(clk32MHz), .D(n31549));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF bit_ctr_i0_i11 (.Q(bit_ctr[11]), .C(clk32MHz), .D(n31547));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF bit_ctr_i0_i10 (.Q(bit_ctr[10]), .C(clk32MHz), .D(n31545));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF bit_ctr_i0_i9 (.Q(bit_ctr[9]), .C(clk32MHz), .D(n31543));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF bit_ctr_i0_i8 (.Q(bit_ctr[8]), .C(clk32MHz), .D(n31541));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF bit_ctr_i0_i7 (.Q(bit_ctr[7]), .C(clk32MHz), .D(n31539));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF bit_ctr_i0_i6 (.Q(bit_ctr[6]), .C(clk32MHz), .D(n31537));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF bit_ctr_i0_i5 (.Q(bit_ctr[5]), .C(clk32MHz), .D(n31535));   // verilog/neopixel.v(35[12] 117[6])
    SB_LUT4 mod_5_add_1674_3_lut (.I0(n2409), .I1(n2409), .I2(n38252), 
            .I3(n28916), .O(n2508)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_3_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1674_3 (.CI(n28916), .I0(n2409), .I1(n38252), .CO(n28917));
    SB_LUT4 mod_5_add_1674_2_lut (.I0(bit_ctr[11]), .I1(bit_ctr[11]), .I2(n38252), 
            .I3(VCC_net), .O(n2509)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_2_lut.LUT_INIT = 16'hA3AC;
    SB_DFF bit_ctr_i0_i4 (.Q(bit_ctr[4]), .C(clk32MHz), .D(n31533));   // verilog/neopixel.v(35[12] 117[6])
    SB_CARRY mod_5_add_1674_2 (.CI(VCC_net), .I0(bit_ctr[11]), .I1(n38252), 
            .CO(n28916));
    SB_DFF bit_ctr_i0_i3 (.Q(bit_ctr[3]), .C(clk32MHz), .D(n31531));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF bit_ctr_i0_i2 (.Q(bit_ctr[2]), .C(clk32MHz), .D(n31529));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF bit_ctr_i0_i1 (.Q(bit_ctr[1]), .C(clk32MHz), .D(n31527));   // verilog/neopixel.v(35[12] 117[6])
    SB_LUT4 mod_5_add_1607_21_lut (.I0(n2291), .I1(n2291), .I2(n2324), 
            .I3(n28915), .O(n2390)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_21_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1607_20_lut (.I0(n2292), .I1(n2292), .I2(n2324), 
            .I3(n28914), .O(n2391)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_20_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_i604_4_lut (.I0(n807), .I1(n838), .I2(n60), .I3(GND_net), 
            .O(n905));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i604_4_lut.LUT_INIT = 16'h0101;
    SB_CARRY add_21_15 (.CI(n27856), .I0(bit_ctr[13]), .I1(GND_net), .CO(n27857));
    SB_CARRY mod_5_add_1607_20 (.CI(n28914), .I0(n2292), .I1(n2324), .CO(n28915));
    SB_CARRY add_21_7 (.CI(n27848), .I0(bit_ctr[5]), .I1(GND_net), .CO(n27849));
    SB_LUT4 mod_5_add_1607_19_lut (.I0(n2293), .I1(n2293), .I2(n2324), 
            .I3(n28913), .O(n2392)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_19_lut.LUT_INIT = 16'hCA3A;
    SB_DFFE start_103 (.Q(start), .C(clk32MHz), .E(VCC_net), .D(n31599));   // verilog/neopixel.v(35[12] 117[6])
    SB_CARRY mod_5_add_1607_19 (.CI(n28913), .I0(n2293), .I1(n2324), .CO(n28914));
    SB_LUT4 mod_5_add_1607_18_lut (.I0(n2294), .I1(n2294), .I2(n2324), 
            .I3(n28912), .O(n2393)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_18_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1607_18 (.CI(n28912), .I0(n2294), .I1(n2324), .CO(n28913));
    SB_LUT4 mod_5_add_1607_17_lut (.I0(n2295), .I1(n2295), .I2(n2324), 
            .I3(n28911), .O(n2394)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_17_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1607_17 (.CI(n28911), .I0(n2295), .I1(n2324), .CO(n28912));
    SB_CARRY sub_14_add_2_25 (.CI(n27962), .I0(timer[23]), .I1(n51[23]), 
            .CO(n27963));
    SB_LUT4 mod_5_add_1607_16_lut (.I0(n2296), .I1(n2296), .I2(n2324), 
            .I3(n28910), .O(n2395)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_16_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1607_16 (.CI(n28910), .I0(n2296), .I1(n2324), .CO(n28911));
    SB_LUT4 mod_5_add_1607_15_lut (.I0(n2297), .I1(n2297), .I2(n2324), 
            .I3(n28909), .O(n2396)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_15_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i29823_3_lut (.I0(n905), .I1(n906), .I2(n33675), .I3(GND_net), 
            .O(n36426));
    defparam i29823_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i4_4_lut (.I0(n17391), .I1(n36426), .I2(bit_ctr[26]), .I3(n14852), 
            .O(n2_adj_4768));
    defparam i4_4_lut.LUT_INIT = 16'h0111;
    SB_CARRY mod_5_add_1607_15 (.CI(n28909), .I0(n2297), .I1(n2324), .CO(n28910));
    SB_CARRY add_21_2 (.CI(VCC_net), .I0(bit_ctr[0]), .I1(GND_net), .CO(n27844));
    SB_LUT4 mod_5_add_1607_14_lut (.I0(n2298), .I1(n2298), .I2(n2324), 
            .I3(n28908), .O(n2397)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_14_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i1_2_lut_adj_1597 (.I0(bit_ctr[27]), .I1(n838), .I2(GND_net), 
            .I3(GND_net), .O(n14852));
    defparam i1_2_lut_adj_1597.LUT_INIT = 16'h9999;
    SB_CARRY mod_5_add_1607_14 (.CI(n28908), .I0(n2298), .I1(n2324), .CO(n28909));
    SB_LUT4 mod_5_i676_3_lut (.I0(bit_ctr[26]), .I1(n971[26]), .I2(n2_adj_4768), 
            .I3(GND_net), .O(n1009));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i676_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 sub_14_add_2_24_lut (.I0(GND_net), .I1(timer[22]), .I2(n51[22]), 
            .I3(n27961), .O(one_wire_N_613[22])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_1607_13_lut (.I0(n2299), .I1(n2299), .I2(n2324), 
            .I3(n28907), .O(n2398)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_13_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1607_13 (.CI(n28907), .I0(n2299), .I1(n2324), .CO(n28908));
    SB_LUT4 add_21_6_lut (.I0(n1), .I1(bit_ctr[4]), .I2(GND_net), .I3(n27847), 
            .O(n37231)) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_6_lut.LUT_INIT = 16'h8228;
    SB_LUT4 mod_5_add_1607_12_lut (.I0(n2300), .I1(n2300), .I2(n2324), 
            .I3(n28906), .O(n2399)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_12_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1607_12 (.CI(n28906), .I0(n2300), .I1(n2324), .CO(n28907));
    SB_LUT4 mod_5_add_1607_11_lut (.I0(n2301), .I1(n2301), .I2(n2324), 
            .I3(n28905), .O(n2400)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_11_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1607_11 (.CI(n28905), .I0(n2301), .I1(n2324), .CO(n28906));
    SB_CARRY sub_14_add_2_24 (.CI(n27961), .I0(timer[22]), .I1(n51[22]), 
            .CO(n27962));
    SB_LUT4 mod_5_add_1607_10_lut (.I0(n2302), .I1(n2302), .I2(n2324), 
            .I3(n28904), .O(n2401)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_10_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1607_10 (.CI(n28904), .I0(n2302), .I1(n2324), .CO(n28905));
    SB_LUT4 mod_5_add_1607_9_lut (.I0(n2303), .I1(n2303), .I2(n2324), 
            .I3(n28903), .O(n2402)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_9_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1607_9 (.CI(n28903), .I0(n2303), .I1(n2324), .CO(n28904));
    SB_LUT4 mod_5_add_1607_8_lut (.I0(n2304), .I1(n2304), .I2(n2324), 
            .I3(n28902), .O(n2403)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_8_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1607_8 (.CI(n28902), .I0(n2304), .I1(n2324), .CO(n28903));
    SB_LUT4 mod_5_add_1607_7_lut (.I0(n2305), .I1(n2305), .I2(n2324), 
            .I3(n28901), .O(n2404)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_7_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1607_7 (.CI(n28901), .I0(n2305), .I1(n2324), .CO(n28902));
    SB_CARRY add_21_6 (.CI(n27847), .I0(bit_ctr[4]), .I1(GND_net), .CO(n27848));
    SB_LUT4 mod_5_add_1607_6_lut (.I0(n2306), .I1(n2306), .I2(n2324), 
            .I3(n28900), .O(n2405)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_6_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1607_6 (.CI(n28900), .I0(n2306), .I1(n2324), .CO(n28901));
    SB_LUT4 mod_5_add_1607_5_lut (.I0(n2307), .I1(n2307), .I2(n2324), 
            .I3(n28899), .O(n2406)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_5_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 sub_14_add_2_23_lut (.I0(GND_net), .I1(timer[21]), .I2(n51[21]), 
            .I3(n27960), .O(one_wire_N_613[21])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_i675_3_lut (.I0(n14852), .I1(n971[27]), .I2(n2_adj_4768), 
            .I3(GND_net), .O(n1008));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i675_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY mod_5_add_1607_5 (.CI(n28899), .I0(n2307), .I1(n2324), .CO(n28900));
    SB_CARRY sub_14_add_2_23 (.CI(n27960), .I0(timer[21]), .I1(n51[21]), 
            .CO(n27961));
    SB_LUT4 mod_5_add_1607_4_lut (.I0(n2308), .I1(n2308), .I2(n2324), 
            .I3(n28898), .O(n2407)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_4_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 sub_14_add_2_22_lut (.I0(GND_net), .I1(timer[20]), .I2(n51[20]), 
            .I3(n27959), .O(one_wire_N_613[20])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i29829_3_lut (.I0(n971[28]), .I1(n971[31]), .I2(n971[29]), 
            .I3(GND_net), .O(n36434));
    defparam i29829_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i2_3_lut_adj_1598 (.I0(n1008), .I1(bit_ctr[25]), .I2(n1009), 
            .I3(GND_net), .O(n6_adj_4769));
    defparam i2_3_lut_adj_1598.LUT_INIT = 16'heaea;
    SB_LUT4 i3_4_lut_adj_1599 (.I0(n2_adj_4768), .I1(n6_adj_4769), .I2(n1005), 
            .I3(n36434), .O(n1037));
    defparam i3_4_lut_adj_1599.LUT_INIT = 16'hfdfc;
    SB_LUT4 i31483_2_lut (.I0(n2_adj_4768), .I1(n971[31]), .I2(GND_net), 
            .I3(GND_net), .O(n4_adj_4647));   // verilog/neopixel.v(22[26:36])
    defparam i31483_2_lut.LUT_INIT = 16'h4444;
    SB_CARRY mod_5_add_1607_4 (.CI(n28898), .I0(n2308), .I1(n2324), .CO(n28899));
    SB_LUT4 mod_5_add_1607_3_lut (.I0(n2309), .I1(n2309), .I2(n38253), 
            .I3(n28897), .O(n2408)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_3_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1607_3 (.CI(n28897), .I0(n2309), .I1(n38253), .CO(n28898));
    SB_LUT4 mod_5_add_1607_2_lut (.I0(bit_ctr[12]), .I1(bit_ctr[12]), .I2(n38253), 
            .I3(VCC_net), .O(n2409)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_2_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1607_2 (.CI(VCC_net), .I0(bit_ctr[12]), .I1(n38253), 
            .CO(n28897));
    SB_LUT4 mod_5_add_1540_20_lut (.I0(n2192), .I1(n2192), .I2(n2225), 
            .I3(n28896), .O(n2291)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_20_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1540_19_lut (.I0(n2193), .I1(n2193), .I2(n2225), 
            .I3(n28895), .O(n2292)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_19_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i31557_1_lut (.I0(n1136), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n38237));
    defparam i31557_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY mod_5_add_1540_19 (.CI(n28895), .I0(n2193), .I1(n2225), .CO(n28896));
    SB_LUT4 mod_5_add_1540_18_lut (.I0(n2194), .I1(n2194), .I2(n2225), 
            .I3(n28894), .O(n2293)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_18_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY sub_14_add_2_22 (.CI(n27959), .I0(timer[20]), .I1(n51[20]), 
            .CO(n27960));
    SB_LUT4 add_21_14_lut (.I0(n1), .I1(bit_ctr[12]), .I2(GND_net), .I3(n27855), 
            .O(n37369)) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_14_lut.LUT_INIT = 16'h8228;
    SB_CARRY mod_5_add_1540_18 (.CI(n28894), .I0(n2194), .I1(n2225), .CO(n28895));
    SB_LUT4 mod_5_add_1540_17_lut (.I0(n2195), .I1(n2195), .I2(n2225), 
            .I3(n28893), .O(n2294)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_17_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1540_17 (.CI(n28893), .I0(n2195), .I1(n2225), .CO(n28894));
    SB_LUT4 mod_5_add_1540_16_lut (.I0(n2196), .I1(n2196), .I2(n2225), 
            .I3(n28892), .O(n2295)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_16_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1540_16 (.CI(n28892), .I0(n2196), .I1(n2225), .CO(n28893));
    SB_LUT4 sub_14_add_2_21_lut (.I0(GND_net), .I1(timer[19]), .I2(n51[19]), 
            .I3(n27958), .O(one_wire_N_613[19])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_21_14 (.CI(n27855), .I0(bit_ctr[12]), .I1(GND_net), .CO(n27856));
    SB_LUT4 mod_5_add_1540_15_lut (.I0(n2197), .I1(n2197), .I2(n2225), 
            .I3(n28891), .O(n2296)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_15_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY sub_14_add_2_21 (.CI(n27958), .I0(timer[19]), .I1(n51[19]), 
            .CO(n27959));
    SB_CARRY mod_5_add_1540_15 (.CI(n28891), .I0(n2197), .I1(n2225), .CO(n28892));
    SB_LUT4 mod_5_add_1540_14_lut (.I0(n2198), .I1(n2198), .I2(n2225), 
            .I3(n28890), .O(n2297)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_14_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1540_14 (.CI(n28890), .I0(n2198), .I1(n2225), .CO(n28891));
    SB_LUT4 mod_5_add_1540_13_lut (.I0(n2199), .I1(n2199), .I2(n2225), 
            .I3(n28889), .O(n2298)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_13_lut.LUT_INIT = 16'hCA3A;
    
endmodule
//
// Verilog Description of module pll32MHz
//

module pll32MHz (GND_net, CLK_c, VCC_net, clk32MHz) /* synthesis lattice_noprune=1, syn_preserve=0, syn_module_defined=1, syn_noprune=0 */ ;
    input GND_net;
    input CLK_c;
    input VCC_net;
    output clk32MHz;
    
    wire CLK_c /* synthesis SET_AS_NETWORK=CLK_c, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(3[9:12])
    wire clk32MHz /* synthesis SET_AS_NETWORK=clk32MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(34[6:14])
    
    SB_PLL40_CORE pll32MHz_inst (.REFERENCECLK(CLK_c), .PLLOUTGLOBAL(clk32MHz), 
            .BYPASS(GND_net), .RESETB(VCC_net)) /* synthesis lattice_noprune=1, syn_instantiated=1, LSE_LINE_FILE_ID=49, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=35, LSE_RLINE=38, syn_preserve=0 */ ;   // verilog/TinyFPGA_B.v(35[10] 38[2])
    defparam pll32MHz_inst.FEEDBACK_PATH = "PHASE_AND_DELAY";
    defparam pll32MHz_inst.DELAY_ADJUSTMENT_MODE_FEEDBACK = "FIXED";
    defparam pll32MHz_inst.DELAY_ADJUSTMENT_MODE_RELATIVE = "FIXED";
    defparam pll32MHz_inst.SHIFTREG_DIV_MODE = 2'b00;
    defparam pll32MHz_inst.FDA_FEEDBACK = 4'b0000;
    defparam pll32MHz_inst.FDA_RELATIVE = 4'b0000;
    defparam pll32MHz_inst.PLLOUT_SELECT = "SHIFTREG_0deg";
    defparam pll32MHz_inst.DIVR = 4'b0000;
    defparam pll32MHz_inst.DIVF = 7'b0000001;
    defparam pll32MHz_inst.DIVQ = 3'b011;
    defparam pll32MHz_inst.FILTER_RANGE = 3'b001;
    defparam pll32MHz_inst.ENABLE_ICEGATE = 1'b0;
    defparam pll32MHz_inst.TEST_MODE = 1'b0;
    defparam pll32MHz_inst.EXTERNAL_DIVIDE_FACTOR = 1;
    
endmodule
//
// Verilog Description of module coms
//

module coms (\data_in_frame[10] , clk32MHz, \data_out_frame[11] , \data_out_frame[9] , 
            GND_net, \data_in_frame[8] , \data_out_frame[6] , rx_data, 
            \data_in_frame[5] , \data_out_frame[8] , \data_out_frame[12] , 
            \data_out_frame[7] , n18202, PWMLimit, n18203, n18204, 
            n18205, n18206, n18207, n18208, n18194, n18195, n18196, 
            n18197, n18198, n18199, n34206, n38508, n18200, n18201, 
            n18186, n18187, n18188, n18189, n18190, n18191, n18192, 
            n18193, \data_in_frame[13] , \data_out_frame[5] , \data_in_frame[12] , 
            \data_in_frame[4] , n34066, \data_in_frame[3] , n4997, n4998, 
            n4999, \data_out_frame[13] , n5000, n5001, \data_out_frame[10] , 
            n5002, n5003, \data_in_frame[2] , n5004, n5005, n5006, 
            \data_out_frame[16] , n5007, n5008, \data_out_frame[18] , 
            n5009, n24786, \data_out_frame[15] , n5010, \data_out_frame[20] , 
            n5011, \data_in_frame[17] , \data_in_frame[1] , n5012, n5013, 
            n5014, n5015, n5016, n5017, n5018, n35492, n5019, 
            n18025, n18024, n18023, n18022, n18021, n18020, \data_in[1] , 
            rx_data_ready, byte_transmit_counter, \data_out_frame[17] , 
            \data_out_frame[19] , \r_SM_Main_2__N_3458[0] , n18019, n18018, 
            \data_in_frame[11] , n18010, control_mode, n18009, n18008, 
            n18007, n18006, n18005, n18004, n18003, \data_out_frame[23][6] , 
            n18002, n18001, n18000, n17999, n17998, n17997, n17996, 
            n17995, n17994, n17993, \data_in[2] , n17992, n17991, 
            n17990, n13724, n17989, n16158, n16154, n3893, n3007, 
            \data_out_frame[14] , n17988, n17987, n17986, n17985, 
            n17984, n17983, \data_in_frame[9] , n17982, n17981, n17980, 
            n17979, n17978, n17977, n17976, n17975, n17974, n17973, 
            n17972, n17971, \data_in[0][6] , n17970, n17969, n17968, 
            n17967, n17966, n17965, n17964, n17963, n17962, n17961, 
            n17960, n17959, n17958, n17957, n17956, n33657, \data_in[3][0] , 
            \data_in[0][3] , \data_in[0][1] , \data_in[0][5] , \data_in[3][2] , 
            \data_in[3][7] , n17955, n17954, n17953, n17952, n17951, 
            n17950, n17949, n17948, n17947, n17946, n17945, n17944, 
            n17943, n17942, n17941, n17940, n17939, n17938, n17937, 
            n17936, n17935, n17934, n17933, n17932, n17931, n17930, 
            n17929, n17928, n17927, n17926, n17925, n17924, n17923, 
            n17922, n17921, n17920, n17919, n17918, n17917, n17916, 
            n17915, n17914, n17913, n17912, n17911, n17910, n17909, 
            n17908, n17907, n17906, n17905, n17904, n17903, n17902, 
            n17901, n17900, n17899, n17898, n17897, n17896, n17895, 
            n17894, n17893, n17892, n17891, n17890, \data_in[3][6] , 
            n17889, n17888, \data_in[0][7] , n17887, n17886, n17885, 
            n17884, n17883, n17882, n17881, n17880, n17879, n17878, 
            n17877, n17876, n17875, n17874, setpoint, n17873, n17872, 
            n17871, n17870, n17869, n17868, n17867, n17866, n17865, 
            n17864, n17863, n17862, n17861, n17860, n17859, n17858, 
            n17857, n17856, n17855, n17854, n17853, n17852, n17851, 
            \Ki[15] , n17850, \Ki[14] , n17849, \Ki[13] , n17848, 
            \Ki[12] , n17847, \Ki[11] , n17846, \Ki[10] , n17845, 
            \Ki[9] , n17844, \Ki[8] , n17843, \Ki[7] , n17842, \Ki[6] , 
            n17841, \Ki[5] , n17840, \Ki[4] , n17839, \Ki[3] , n63, 
            n17838, \Ki[2] , n17837, \Ki[1] , n17836, \Kp[15] , 
            n17835, \Kp[14] , n17834, \Kp[13] , n17833, \Kp[12] , 
            n17832, \Kp[11] , n17831, \Kp[10] , \data_in[0][0] , \data_in[0][4] , 
            \data_in[3][4] , n17830, \Kp[9] , n17829, \Kp[8] , n17828, 
            \Kp[7] , n17827, \Kp[6] , n17826, \Kp[5] , n17825, \Kp[4] , 
            n17824, \Kp[3] , n17823, \Kp[2] , n17822, \Kp[1] , n17821, 
            n17820, n17818, n17816, n17814, n17813, n17812, n17810, 
            n17808, n17806, n33228, n737, \FRAME_MATCHER.state_31__N_2566[1] , 
            n4996, n5, n16159, n2958, n32962, n32941, n32957, 
            n5439, n17308, PIN_11_c, n17805, n4, n17804, n17803, 
            n17802, n17801, n17800, n17799, n17798, n17797, n17796, 
            n17795, n17794, n17793, n17791, n17790, IntegralLimit, 
            n17789, n17788, n17787, n17786, n17785, n17784, n17783, 
            n17782, n17781, n17780, n17779, n17778, LED_c, n17777, 
            n17776, n17527, n18153, n18152, n18151, n18150, n18149, 
            n18089, n17775, n17774, n18088, n17656, n25050, n17659, 
            n18087, n18086, n18085, n17662, n17665, n18084, n18083, 
            n18082, n17668, n18148, n18147, n17550, n17773, n17772, 
            n17771, n17770, n17769, n17768, n17671, n17674, n8014, 
            tx_transmit_N_3355, n16157, n34531, n18146, \FRAME_MATCHER.state_31__N_2566[2] , 
            n17696, n17694, n17693, n17692, \Ki[0] , n17691, \Kp[0] , 
            n17690, n17658, n17661, n17664, n17667, n17670, n17673, 
            n17676, n17731, \r_SM_Main[2] , r_Bit_Index, n17362, n17534, 
            n5600, \r_Clock_Count[6] , \r_Clock_Count[7] , \r_Clock_Count[8] , 
            \r_Clock_Count[0] , \r_Clock_Count[3] , n313, n314, n315, 
            n316, \r_Clock_Count[5] , tx_active, n5478, n318, n321, 
            VCC_net, tx_o, tx_enable, n17559, n18278, n17652, n17655, 
            n17708, n17713, n17728, n17549, n17553, n25112, \r_SM_Main[1] , 
            n18260, r_Rx_Data, n37332, PIN_13_N_105, \r_SM_Main[2]_adj_3 , 
            n33769, n17681, r_Bit_Index_adj_10, n5578, n24193, n4_adj_7, 
            n4_adj_8, n16148, n25070, n1, n37333, n17701, n17689, 
            n17688, n17687, n17686, n17685, n17684, n17683, n16143, 
            n17679, n17682, n17735, n4_adj_9) /* synthesis lattice_noprune=1, syn_preserve=0, syn_module_defined=1, syn_noprune=0 */ ;
    output [7:0]\data_in_frame[10] ;
    input clk32MHz;
    output [7:0]\data_out_frame[11] ;
    output [7:0]\data_out_frame[9] ;
    input GND_net;
    output [7:0]\data_in_frame[8] ;
    output [7:0]\data_out_frame[6] ;
    output [7:0]rx_data;
    output [7:0]\data_in_frame[5] ;
    output [7:0]\data_out_frame[8] ;
    output [7:0]\data_out_frame[12] ;
    output [7:0]\data_out_frame[7] ;
    input n18202;
    output [23:0]PWMLimit;
    input n18203;
    input n18204;
    input n18205;
    input n18206;
    input n18207;
    input n18208;
    input n18194;
    input n18195;
    input n18196;
    input n18197;
    input n18198;
    input n18199;
    input n34206;
    input n38508;
    input n18200;
    input n18201;
    input n18186;
    input n18187;
    input n18188;
    input n18189;
    input n18190;
    input n18191;
    input n18192;
    input n18193;
    output [7:0]\data_in_frame[13] ;
    output [7:0]\data_out_frame[5] ;
    output [7:0]\data_in_frame[12] ;
    output [7:0]\data_in_frame[4] ;
    output n34066;
    output [7:0]\data_in_frame[3] ;
    output n4997;
    output n4998;
    output n4999;
    output [7:0]\data_out_frame[13] ;
    output n5000;
    output n5001;
    output [7:0]\data_out_frame[10] ;
    output n5002;
    output n5003;
    output [7:0]\data_in_frame[2] ;
    output n5004;
    output n5005;
    output n5006;
    output [7:0]\data_out_frame[16] ;
    output n5007;
    output n5008;
    output [7:0]\data_out_frame[18] ;
    output n5009;
    output n24786;
    output [7:0]\data_out_frame[15] ;
    output n5010;
    output [7:0]\data_out_frame[20] ;
    output n5011;
    output [7:0]\data_in_frame[17] ;
    output [7:0]\data_in_frame[1] ;
    output n5012;
    output n5013;
    output n5014;
    output n5015;
    output n5016;
    output n5017;
    output n5018;
    output n35492;
    output n5019;
    input n18025;
    input n18024;
    input n18023;
    input n18022;
    input n18021;
    input n18020;
    output [7:0]\data_in[1] ;
    output rx_data_ready;
    output [7:0]byte_transmit_counter;
    output [7:0]\data_out_frame[17] ;
    output [7:0]\data_out_frame[19] ;
    output \r_SM_Main_2__N_3458[0] ;
    input n18019;
    input n18018;
    output [7:0]\data_in_frame[11] ;
    input n18010;
    output [7:0]control_mode;
    input n18009;
    input n18008;
    input n18007;
    input n18006;
    input n18005;
    input n18004;
    input n18003;
    output \data_out_frame[23][6] ;
    input n18002;
    input n18001;
    input n18000;
    input n17999;
    input n17998;
    input n17997;
    input n17996;
    input n17995;
    input n17994;
    input n17993;
    output [7:0]\data_in[2] ;
    input n17992;
    input n17991;
    input n17990;
    output n13724;
    input n17989;
    output n16158;
    output n16154;
    output n3893;
    output n3007;
    output [7:0]\data_out_frame[14] ;
    input n17988;
    input n17987;
    input n17986;
    input n17985;
    input n17984;
    input n17983;
    output [7:0]\data_in_frame[9] ;
    input n17982;
    input n17981;
    input n17980;
    input n17979;
    input n17978;
    input n17977;
    input n17976;
    input n17975;
    input n17974;
    input n17973;
    input n17972;
    input n17971;
    output \data_in[0][6] ;
    input n17970;
    input n17969;
    input n17968;
    input n17967;
    input n17966;
    input n17965;
    input n17964;
    input n17963;
    input n17962;
    input n17961;
    input n17960;
    input n17959;
    input n17958;
    input n17957;
    input n17956;
    output n33657;
    output \data_in[3][0] ;
    output \data_in[0][3] ;
    output \data_in[0][1] ;
    output \data_in[0][5] ;
    output \data_in[3][2] ;
    output \data_in[3][7] ;
    input n17955;
    input n17954;
    input n17953;
    input n17952;
    input n17951;
    input n17950;
    input n17949;
    input n17948;
    input n17947;
    input n17946;
    input n17945;
    input n17944;
    input n17943;
    input n17942;
    input n17941;
    input n17940;
    input n17939;
    input n17938;
    input n17937;
    input n17936;
    input n17935;
    input n17934;
    input n17933;
    input n17932;
    input n17931;
    input n17930;
    input n17929;
    input n17928;
    input n17927;
    input n17926;
    input n17925;
    input n17924;
    input n17923;
    input n17922;
    input n17921;
    input n17920;
    input n17919;
    input n17918;
    input n17917;
    input n17916;
    input n17915;
    input n17914;
    input n17913;
    input n17912;
    input n17911;
    input n17910;
    input n17909;
    input n17908;
    input n17907;
    input n17906;
    input n17905;
    input n17904;
    input n17903;
    input n17902;
    input n17901;
    input n17900;
    input n17899;
    input n17898;
    input n17897;
    input n17896;
    input n17895;
    input n17894;
    input n17893;
    input n17892;
    input n17891;
    input n17890;
    output \data_in[3][6] ;
    input n17889;
    input n17888;
    output \data_in[0][7] ;
    input n17887;
    input n17886;
    input n17885;
    input n17884;
    input n17883;
    input n17882;
    input n17881;
    input n17880;
    input n17879;
    input n17878;
    input n17877;
    input n17876;
    input n17875;
    input n17874;
    output [23:0]setpoint;
    input n17873;
    input n17872;
    input n17871;
    input n17870;
    input n17869;
    input n17868;
    input n17867;
    input n17866;
    input n17865;
    input n17864;
    input n17863;
    input n17862;
    input n17861;
    input n17860;
    input n17859;
    input n17858;
    input n17857;
    input n17856;
    input n17855;
    input n17854;
    input n17853;
    input n17852;
    input n17851;
    output \Ki[15] ;
    input n17850;
    output \Ki[14] ;
    input n17849;
    output \Ki[13] ;
    input n17848;
    output \Ki[12] ;
    input n17847;
    output \Ki[11] ;
    input n17846;
    output \Ki[10] ;
    input n17845;
    output \Ki[9] ;
    input n17844;
    output \Ki[8] ;
    input n17843;
    output \Ki[7] ;
    input n17842;
    output \Ki[6] ;
    input n17841;
    output \Ki[5] ;
    input n17840;
    output \Ki[4] ;
    input n17839;
    output \Ki[3] ;
    output n63;
    input n17838;
    output \Ki[2] ;
    input n17837;
    output \Ki[1] ;
    input n17836;
    output \Kp[15] ;
    input n17835;
    output \Kp[14] ;
    input n17834;
    output \Kp[13] ;
    input n17833;
    output \Kp[12] ;
    input n17832;
    output \Kp[11] ;
    input n17831;
    output \Kp[10] ;
    output \data_in[0][0] ;
    output \data_in[0][4] ;
    output \data_in[3][4] ;
    input n17830;
    output \Kp[9] ;
    input n17829;
    output \Kp[8] ;
    input n17828;
    output \Kp[7] ;
    input n17827;
    output \Kp[6] ;
    input n17826;
    output \Kp[5] ;
    input n17825;
    output \Kp[4] ;
    input n17824;
    output \Kp[3] ;
    input n17823;
    output \Kp[2] ;
    input n17822;
    output \Kp[1] ;
    input n17821;
    input n17820;
    input n17818;
    input n17816;
    input n17814;
    input n17813;
    input n17812;
    input n17810;
    input n17808;
    input n17806;
    output n33228;
    output n737;
    output \FRAME_MATCHER.state_31__N_2566[1] ;
    output n4996;
    input n5;
    output n16159;
    output n2958;
    output n32962;
    output n32941;
    output n32957;
    output n5439;
    output n17308;
    output PIN_11_c;
    input n17805;
    output n4;
    input n17804;
    input n17803;
    input n17802;
    input n17801;
    input n17800;
    input n17799;
    input n17798;
    input n17797;
    input n17796;
    input n17795;
    input n17794;
    input n17793;
    input n17791;
    input n17790;
    output [23:0]IntegralLimit;
    input n17789;
    input n17788;
    input n17787;
    input n17786;
    input n17785;
    input n17784;
    input n17783;
    input n17782;
    input n17781;
    input n17780;
    input n17779;
    input n17778;
    output LED_c;
    input n17777;
    input n17776;
    output n17527;
    input n18153;
    input n18152;
    input n18151;
    input n18150;
    input n18149;
    input n18089;
    input n17775;
    input n17774;
    input n18088;
    output n17656;
    output n25050;
    output n17659;
    input n18087;
    input n18086;
    input n18085;
    output n17662;
    output n17665;
    input n18084;
    input n18083;
    input n18082;
    output n17668;
    input n18148;
    input n18147;
    input n17550;
    input n17773;
    input n17772;
    input n17771;
    input n17770;
    input n17769;
    input n17768;
    output n17671;
    output n17674;
    output n8014;
    output tx_transmit_N_3355;
    output n16157;
    output n34531;
    input n18146;
    output \FRAME_MATCHER.state_31__N_2566[2] ;
    input n17696;
    input n17694;
    input n17693;
    input n17692;
    output \Ki[0] ;
    input n17691;
    output \Kp[0] ;
    input n17690;
    input n17658;
    input n17661;
    input n17664;
    input n17667;
    input n17670;
    input n17673;
    input n17676;
    input n17731;
    output \r_SM_Main[2] ;
    output [2:0]r_Bit_Index;
    output n17362;
    output n17534;
    output n5600;
    output \r_Clock_Count[6] ;
    output \r_Clock_Count[7] ;
    output \r_Clock_Count[8] ;
    output \r_Clock_Count[0] ;
    output \r_Clock_Count[3] ;
    output n313;
    output n314;
    output n315;
    output n316;
    output \r_Clock_Count[5] ;
    output tx_active;
    output n5478;
    output n318;
    output n321;
    input VCC_net;
    output tx_o;
    output tx_enable;
    input n17559;
    input n18278;
    input n17652;
    input n17655;
    input n17708;
    input n17713;
    input n17728;
    input n17549;
    input n17553;
    input n25112;
    output \r_SM_Main[1] ;
    input n18260;
    output r_Rx_Data;
    output n37332;
    input PIN_13_N_105;
    output \r_SM_Main[2]_adj_3 ;
    output n33769;
    output n17681;
    output [2:0]r_Bit_Index_adj_10;
    output n5578;
    output n24193;
    output n4_adj_7;
    output n4_adj_8;
    output n16148;
    output n25070;
    output n1;
    output n37333;
    input n17701;
    input n17689;
    input n17688;
    input n17687;
    input n17686;
    input n17685;
    input n17684;
    input n17683;
    output n16143;
    input n17679;
    input n17682;
    input n17735;
    output n4_adj_9;
    
    wire clk32MHz /* synthesis SET_AS_NETWORK=clk32MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(34[6:14])
    wire LED_c /* synthesis SET_AS_NETWORK=LED_c, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(4[10:13])
    
    wire n14, n10, n32982, n16413, n18168;
    wire [7:0]\data_in_frame[19] ;   // verilog/coms.v(95[12:25])
    wire [7:0]\data_in_frame[14] ;   // verilog/coms.v(95[12:25])
    
    wire n16314;
    wire [7:0]\data_in_frame[15] ;   // verilog/coms.v(95[12:25])
    
    wire n33310, n17068, n18076, n18167, n33546, n16229, n1270, 
        n14_adj_4339, n18166, n18165, n9, n33381, n30857, n18164, 
        n18163, n18162, n18161;
    wire [7:0]\data_in_frame[18] ;   // verilog/coms.v(95[12:25])
    
    wire n18160, n18159, n8, n32959, n18051, n18075, n18074, n18137, 
        n2;
    wire [31:0]\FRAME_MATCHER.i ;   // verilog/coms.v(114[11:12])
    
    wire n3, n18124, n27910, n27911, n2_adj_4340, n27909, n2290, 
        n33107, n1301, n16672, n16163, n16687, n16880, n16525, 
        n33313, n6, n33066, n16304, n33427, n33115, n16548, n30801, 
        n16521, n18073;
    wire [7:0]\data_in_frame[7] ;   // verilog/coms.v(95[12:25])
    
    wire n18183;
    wire [7:0]\data_in_frame[21] ;   // verilog/coms.v(95[12:25])
    
    wire n18184;
    wire [31:0]\FRAME_MATCHER.state ;   // verilog/coms.v(111[11:16])
    
    wire n18072, n18071, n18070, n18169, n18069, n18068, n18185, 
        n18181, n18182, n18179, n18180, n18177;
    wire [7:0]\data_in_frame[20] ;   // verilog/coms.v(95[12:25])
    
    wire n18178, n18175, n18176, n18173, n18174, n18067, n18170, 
        n18171, n18172, n18066, n18123, n18122, n18121, n18120, 
        n18119, n18118, n18117, n18136, n18065;
    wire [7:0]\data_in_frame[6] ;   // verilog/coms.v(95[12:25])
    
    wire n18064, n18063, n18062, n18061, n18060, n18059, n18058, 
        n18057, n18056, n18055, n18054, n18053, n18052, n18116, 
        n33330, n33127, n33508, n18050, n18115, n18049, n18114, 
        n18048, n18047, n18046, n18045, n18113, n18112, n1251, 
        n6_adj_4341, n33241, n15783, n1254, n33265, n13947, n31, 
        n16162, n4995, n18111, n33073, n33204, n33256, n16946, 
        n33540, n32, n22, n31287, n36, n33494, n33253, n33287, 
        n34, n16545, n35, n33610, n33, n31223, n10_adj_4342, n34521, 
        n16676, n31188, n6_adj_4343, n33303, n30451, n13554, n25118, 
        n33773, n16195, n16000, n8_adj_4344, n7, n5069;
    wire [0:0]n3693;
    
    wire n33520, n33060, n14_adj_4345, n10_adj_4346, n16711, n34672, 
        n33789, n35075, n33201, n33020, n33371, n16647, n42, n34894, 
        n35045, n4_c, n18044, n33634, n33636, n31_adj_4347, Kp_23__N_993, 
        n15, n16791, Kp_23__N_996, n21, n31230, n30217, n28, n6_adj_4348, 
        n16722, n16380, n16834, n26, n16335, Kp_23__N_1046, n27, 
        n16608, n31002, n16765, n16384, n25;
    wire [7:0]\data_in_frame[0] ;   // verilog/coms.v(95[12:25])
    
    wire n14_adj_4349, n9_adj_4350, n6_adj_4351, n6_adj_4352, n18043, 
        n18042, n18041, n18040, n18039, n18038, n18037, n18036, 
        n18035, n18034, n18033, n18032, n18031, n18030, n18029, 
        n18028, n18027, n18026, n18110, n33186, n34651, n8_adj_4353, 
        n18109, n33279, n33483, n10_adj_4354, n18108, n18135;
    wire [7:0]\data_in[0] ;   // verilog/coms.v(94[12:19])
    
    wire n17792, n8_adj_4355;
    wire [7:0]byte_transmit_counter_c;   // verilog/coms.v(101[12:33])
    
    wire n6_adj_4356, n18134, n5_c, n37177, n7_adj_4357, n38438, 
        n38444, n14_adj_4358, n6_adj_4359, n5_adj_4360, n7_adj_4361, 
        n18133, n38348, n38450, n14_adj_4362, n6_adj_4363, n5_adj_4364, 
        n7_adj_4365, n38342, n38456, n14_adj_4366, n16, n17;
    wire [7:0]\data_out_frame[23] ;   // verilog/coms.v(96[12:26])
    
    wire n37271, n37270, n33238, n34170, n16233, n30694, n6_adj_4367, 
        n5_adj_4368, n24810, n34514;
    wire [7:0]\data_in_frame[16] ;   // verilog/coms.v(95[12:25])
    
    wire n31184, n33464, n7_adj_4369, \FRAME_MATCHER.rx_data_ready_prev , 
        n38330, n38462, n14_adj_4370, n18107, Kp_23__N_1183, n34073, 
        n37536, n14_adj_4371, n10_adj_4372, n5_adj_4373, n33323, n33583, 
        n8_adj_4374, n33076, n5034, n33781, n13, n11, n16930, 
        n34659, n18132, n33247, n33471, n12, n7_adj_4375, n18106, 
        n33385, n33350, n33526, n33250, n12_adj_4376, n18017, n18016, 
        n18015, n18014, n38324, n38318, n14_adj_4377, n16_adj_4378, 
        n17_adj_4379, n33604, n33104, n37531, n17157, n33316, n10_adj_4380, 
        n15795, n33269, n35077, n33445, n10_adj_4381, n5_adj_4382, 
        Kp_23__N_1026, n7_adj_4383, n32994, n32937, n38372, n38288, 
        n14_adj_4384, n33532, n16_adj_4385, n18013, n18012, n18011, 
        n18125, n33217, n11_adj_4386, n33409, n33607, n33036, n17_adj_4387, 
        n18105, n33354, n15781, n16740, n9_adj_4388, n12_adj_4389, 
        n32271, n37837, n5_adj_4390, n7_adj_4391, n38366, n38294, 
        n14_adj_4392, n32219, n32221, n6_adj_4393, n5_adj_4394, n7_adj_4395, 
        n32223, n33155, n38354, n38312, n14_adj_4396, n33335, n31196, 
        n32225, n18131, n32227, n32161, n33474, n10_adj_4397, n32181, 
        n33010, n16447, n161, n32229, n32231, n32233, n32235, 
        n10_adj_4398, n33142, n33357, n32149, n32237, n33397;
    wire [7:0]\data_in[3] ;   // verilog/coms.v(94[12:19])
    
    wire n17807, n32239, n16466, n31228, n17809, n36323, n30, 
        n17811, n32855, n28_adj_4399, n29, n27_adj_4400;
    wire [31:0]\FRAME_MATCHER.state_31__N_2630 ;
    
    wire n18130, n33403, n16951, n16299, n1_c, n4_adj_4401, n7_adj_4402, 
        n33406, n33306, n16161, n36418, n32241, n17815, n33178, 
        n17817, n136, n4_adj_4403, n8_adj_4404, n17819, n10_adj_4405, 
        n34982, n18129, n30241, n33388, n6_adj_4406, n33054, n6_adj_4407, 
        n18128, n33292, n17126, n8_adj_4408, n33503, n35487, n17169, 
        n33003, n33529, n6_adj_4409, n33063, n33616, n33552, n32989, 
        n4_adj_4410, n24185, n22566, n42_adj_4411, n30769, n16661, 
        n31295, n4_adj_4412, n33013, n33589, n33377, n33622, n10_adj_4413, 
        n33488, n31265, n14_adj_4414, n10_adj_4415, n33439, n16975, 
        n33514, n33145, n16746, n32952, n16153, n10_adj_4416, n31298, 
        n10_adj_4417, n16114, n15973, n14_adj_4418, n16108, n15_adj_4419, 
        n18, n16_adj_4420, n16097, n20, n33158, n16570, n16906, 
        n6_adj_4421, n33189, n10_adj_4422, n33164, n33543, n22_adj_4423, 
        n20_adj_4424, n98, n53, n6_adj_4425, n16_adj_4426, n24, 
        n16090, n32109, n16350, n34236, n158, n16_adj_4427, n17_adj_4428, 
        n22269, n35535, n16319, n12_adj_4429, n3_adj_4430, n32183, 
        n12_adj_4431, n31163, n33195, n1999, n35212, n33570, n14584, 
        n33262, n32979, n34522, n16679, n33087, n16795, n15982, 
        n35262, n35254, n24089, n31190, n33168, n33169, n14531, 
        n6_adj_4432, n6_adj_4433, n31225, n33549, n33338, n33511, 
        n30360, n67, n34726, n6_adj_4434, n30231, n8_adj_4435, n33368, 
        n16536, n6_adj_4436, n31249, n33223, n10_adj_4437, n10_adj_4438, 
        n14_adj_4439, n30192, n16291, n37292, n37291, n10_adj_4440, 
        n16_adj_4441, n16_adj_4442, n17_adj_4443, n17_adj_4444, n136_adj_4445, 
        n33017, n33430, n34266, n5_adj_4446, n34116, n33564, n6_adj_4447, 
        n33171, n14_adj_4448, n8_adj_4449, n12_adj_4450, n13_adj_4451, 
        n34664, n11_adj_4452, n42_adj_4453, n18079, n18104, n40, 
        n28_adj_4454, n32_adj_4455, n33523, n33598, n33477, n33042, 
        n33586, n33344, n33457, n8_adj_4456, n41, n34691, n39, 
        n38, n37, n16404, n33619, n33210, n30_adj_4457, n48, n10_adj_4458, 
        n33207, n33631, n10_adj_4459, Kp_23__N_843, n7_adj_4460, n33505, 
        n17072, n34_adj_4461, n4_adj_4462, n8_adj_4463, n17695, n12_adj_4464, 
        n30339, n43, n33573, n33451, n32_adj_4465, n4_adj_4466, 
        n33148, n33023, n33_adj_4467, n31_adj_4468, n31178, n18098, 
        n18099, n18100, n36430, n30968, n16477, n1981, n18101, 
        n22275, n36422, n10599;
    wire [31:0]n92;
    
    wire n1337, n4_adj_4469, n32976, n35602, n18102, n4_adj_4471, 
        n34351, n18103, n37283, n37282, n18080, n6_adj_4472, n16954, 
        n16726, n17135, n9_adj_4473, n33558, n18081, n18077, n18078, 
        n34996, n33057, n16998, n33442, n28_adj_4474, n26_adj_4475, 
        n33576, n33069, n27_adj_4476, n32985, n25_adj_4477, n33175, 
        n38459, n38453, n38447, n38441, n38435, n38258, n37290, 
        n38423;
    wire [7:0]tx_data;   // verilog/coms.v(104[13:20])
    
    wire n38264, n37281, n38417, n16_adj_4478, n17_adj_4479, n37280, 
        n37279, n38270, n37278, n38411, n38276, n37275, n38405, 
        n38282, n37272, n38399, n38393, n37807, n37269, n38387, 
        n38306, n37266, n38381, n38336, n37257, n38375, n38369, 
        n38363, n16_adj_4480, n17_adj_4481, n33424, n33436, n25_adj_4482, 
        n31209, n30_adj_4483, n2_adj_4484, n27939, n3_adj_4485, n37277, 
        n34_adj_4486, n29_adj_4487, n37276, n16_adj_4488, n17_adj_4489, 
        n17_adj_4490, n21_adj_4491, n2_adj_4492, n27938, n2_adj_4493, 
        n27937, n2_adj_4494, n27936, n2_adj_4495, n3_adj_4496, n2_adj_4497, 
        n3_adj_4498, n2_adj_4499, n3_adj_4500, n2_adj_4501, n3_adj_4502, 
        n2_adj_4503, n3_adj_4504, n2_adj_4505, n3_adj_4506, n2_adj_4507, 
        n3_adj_4508, n2_adj_4509, n3_adj_4510, n2_adj_4511, n3_adj_4512, 
        n2_adj_4513, n3_adj_4514, n2_adj_4515, n3_adj_4516, n2_adj_4517, 
        n3_adj_4518, n2_adj_4519, n3_adj_4520, n2_adj_4521, n3_adj_4522, 
        n2_adj_4523, n3_adj_4524, n2_adj_4525, n3_adj_4526, n2_adj_4527, 
        n3_adj_4528, n2_adj_4529, n3_adj_4530, n2_adj_4531, n3_adj_4532, 
        n2_adj_4533, n3_adj_4534, n2_adj_4535, n3_adj_4536, n2_adj_4537, 
        n3_adj_4538, n2_adj_4539, n3_adj_4540, n2_adj_4541, n3_adj_4542, 
        n2_adj_4543, n3_adj_4544, n2_adj_4545, n3_adj_4546, n3_adj_4547, 
        n3_adj_4548, n3_adj_4549, n3_adj_4550, n33202, n34730, n24_adj_4551, 
        n20_adj_4552, n35248, n33421, n6_adj_4553, n28_adj_4554, n34864, 
        n34374, n34501, n34502, n34130;
    wire [7:0]\data_out_frame[24] ;   // verilog/coms.v(96[12:26])
    
    wire n34495, n32999, n33480, n5_adj_4555, n24102, n24819, n32277, 
        n32279, n7_adj_4556, n8_adj_4557, n24104, n24821, n24106, 
        n32113, n24108, n32117, n32281, n32283, n32285, n32287, 
        n32289, n32291, n24110, n24823, n32275, n32185, n24112, 
        n24825, n32293, n32295, n29601, n29605, n32297, n32299, 
        n32301, n32171, n29611, n32273, n32173, n29609, n32175, 
        n29613, n32179, n29607, n32_adj_4558, n30_adj_4559, n31_adj_4560, 
        n33467, n29_adj_4561, n18138, n18139, n18140, n33198, n18141, 
        n33273, n18142, n30899, n33081, n16855, n20_adj_4562, n33259, 
        n33039, n19, n33045, n21_adj_4563, n33613, n10_adj_4564, 
        n18143, n18144, n6_adj_4565, n9_adj_4566, n30900, n33500, 
        n18145, n33183, n4_adj_4567, n33567, n16_adj_4569, n31235, 
        n27935, n16347, n16_adj_4570, n17_adj_4571, n37274, n37273, 
        n18154, n18155, n18156, n18157, n33580, n33448, n17_adj_4572, 
        n16_adj_4573, n33244, n17_adj_4574, n37268, n37267, n17081, 
        n19_adj_4575, n33374, n33094, n31257, Kp_23__N_1662, n33595, 
        n33628, n33394, n18158, n27934, n38351, n18097, n18096, 
        n18095, n18094, n18093, n17449, n27933, n18092, n27932, 
        n18091, n6_adj_4576, n31204, n31168, n16292, n33121, n16262, 
        n16_adj_4577, n20_adj_4578, n33000, n19_adj_4579, n33555, 
        n33118, n21_adj_4580, n33537, n17_adj_4581, n27931, n34934, 
        Kp_23__N_860, n10_adj_4582, n38345, n38339, n37258, n37259, 
        n38333, n17_adj_4583, n16_adj_4584, n38327, n38321, n38315, 
        n33517, n16862, n33110, n18_adj_4585, n27930, n27929, n16248, 
        n33414, n16242, n33192, n33341, n20_adj_4586, n27928, n33151, 
        n6_adj_4587, n16840, n16_adj_4588, n6_adj_4589, n6_adj_4590, 
        n6_adj_4591, n30930, n17132, n33090, n17042, n18090, n7_adj_4592, 
        n30438, n31219, n27927, n35345, n16626, n33232, n33320, 
        n38309, n16816, n33625, n10_adj_4593, n33298, n16435, n30805, 
        Kp_23__N_1453, n33235, n12_adj_4594, n17036, n12_adj_4595, 
        n27926, n28024, n28023, n14_adj_4596, n15_adj_4597, n33491, 
        n22_adj_4598, n32_adj_4599, n35349, n36_adj_4600, n34_adj_4601, 
        n35_adj_4602, n33_adj_4603, n16080, n18127, n10_adj_4604, 
        n14_adj_4605, n10_adj_4606, n27925, n28022, n38303, n33601, 
        n10_adj_4607, n33220, n28021, n12_adj_4608, n27924, n28020, 
        n16399, n27923, n38291, n38285, n27922, n38279, n16418, 
        n35410, n28019, n14758, n16780, n6_adj_4609, n50, n38273, 
        n17111, n57, n54, n52, n28018, n18126, n38267, n27921, 
        n53_adj_4610, n33454, n51, n56, n62, n33592, n55, n118, 
        n63_adj_4611, n27920, n1502, n16392, n16620, n6_adj_4612, 
        n27919, n17182, n34605, n38261, n27918, n27917, n27916, 
        n27915, n23, n22_adj_4613, n26_adj_4614, n38255, n27914, 
        n10_adj_4615, n27913, n33295, n14_adj_4616, n17004, n16179, 
        n12_adj_4617, n27912, n12_adj_4618, n33007;
    
    SB_LUT4 i7_4_lut (.I0(\data_in_frame[10] [5]), .I1(n14), .I2(n10), 
            .I3(n32982), .O(n16413));   // verilog/coms.v(72[16:42])
    defparam i7_4_lut.LUT_INIT = 16'h6996;
    SB_DFF data_in_frame_0__i159 (.Q(\data_in_frame[19] [6]), .C(clk32MHz), 
           .D(n18168));   // verilog/coms.v(126[12] 293[6])
    SB_LUT4 i3_4_lut (.I0(\data_in_frame[14] [7]), .I1(n16314), .I2(\data_in_frame[14] [6]), 
            .I3(\data_in_frame[15] [0]), .O(n33310));
    defparam i3_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut (.I0(\data_out_frame[11] [4]), .I1(\data_out_frame[9] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n17068));
    defparam i1_2_lut.LUT_INIT = 16'h6666;
    SB_DFF data_in_frame_0__i67 (.Q(\data_in_frame[8] [2]), .C(clk32MHz), 
           .D(n18076));   // verilog/coms.v(126[12] 293[6])
    SB_DFF data_in_frame_0__i158 (.Q(\data_in_frame[19] [5]), .C(clk32MHz), 
           .D(n18167));   // verilog/coms.v(126[12] 293[6])
    SB_LUT4 i6_4_lut (.I0(n33546), .I1(n16229), .I2(\data_out_frame[6] [4]), 
            .I3(n1270), .O(n14_adj_4339));   // verilog/coms.v(70[16:27])
    defparam i6_4_lut.LUT_INIT = 16'h6996;
    SB_DFF data_in_frame_0__i157 (.Q(\data_in_frame[19] [4]), .C(clk32MHz), 
           .D(n18166));   // verilog/coms.v(126[12] 293[6])
    SB_DFF data_in_frame_0__i156 (.Q(\data_in_frame[19] [3]), .C(clk32MHz), 
           .D(n18165));   // verilog/coms.v(126[12] 293[6])
    SB_LUT4 i1_3_lut (.I0(\data_out_frame[6] [1]), .I1(\data_out_frame[6] [3]), 
            .I2(\data_out_frame[6] [2]), .I3(GND_net), .O(n9));   // verilog/coms.v(70[16:27])
    defparam i1_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 i7_4_lut_adj_877 (.I0(n9), .I1(n14_adj_4339), .I2(n33381), 
            .I3(\data_out_frame[6] [5]), .O(n30857));   // verilog/coms.v(70[16:27])
    defparam i7_4_lut_adj_877.LUT_INIT = 16'h6996;
    SB_DFF data_in_frame_0__i155 (.Q(\data_in_frame[19] [2]), .C(clk32MHz), 
           .D(n18164));   // verilog/coms.v(126[12] 293[6])
    SB_DFF data_in_frame_0__i154 (.Q(\data_in_frame[19] [1]), .C(clk32MHz), 
           .D(n18163));   // verilog/coms.v(126[12] 293[6])
    SB_DFF data_in_frame_0__i153 (.Q(\data_in_frame[19] [0]), .C(clk32MHz), 
           .D(n18162));   // verilog/coms.v(126[12] 293[6])
    SB_DFF data_in_frame_0__i152 (.Q(\data_in_frame[18] [7]), .C(clk32MHz), 
           .D(n18161));   // verilog/coms.v(126[12] 293[6])
    SB_DFF data_in_frame_0__i151 (.Q(\data_in_frame[18] [6]), .C(clk32MHz), 
           .D(n18160));   // verilog/coms.v(126[12] 293[6])
    SB_DFF data_in_frame_0__i150 (.Q(\data_in_frame[18] [5]), .C(clk32MHz), 
           .D(n18159));   // verilog/coms.v(126[12] 293[6])
    SB_LUT4 i13222_3_lut_4_lut (.I0(n8), .I1(n32959), .I2(rx_data[1]), 
            .I3(\data_in_frame[5] [1]), .O(n18051));
    defparam i13222_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF data_in_frame_0__i66 (.Q(\data_in_frame[8] [1]), .C(clk32MHz), 
           .D(n18075));   // verilog/coms.v(126[12] 293[6])
    SB_DFF data_in_frame_0__i65 (.Q(\data_in_frame[8] [0]), .C(clk32MHz), 
           .D(n18074));   // verilog/coms.v(126[12] 293[6])
    SB_DFF data_in_frame_0__i128 (.Q(\data_in_frame[15] [7]), .C(clk32MHz), 
           .D(n18137));   // verilog/coms.v(126[12] 293[6])
    SB_DFFSS \FRAME_MATCHER.i_i0  (.Q(\FRAME_MATCHER.i [0]), .C(clk32MHz), 
            .D(n2), .S(n3));   // verilog/coms.v(126[12] 293[6])
    SB_DFF data_in_frame_0__i115 (.Q(\data_in_frame[14] [2]), .C(clk32MHz), 
           .D(n18124));   // verilog/coms.v(126[12] 293[6])
    SB_CARRY add_41_4 (.CI(n27910), .I0(\FRAME_MATCHER.i [2]), .I1(GND_net), 
            .CO(n27911));
    SB_LUT4 add_41_3_lut (.I0(n2290), .I1(\FRAME_MATCHER.i [1]), .I2(GND_net), 
            .I3(n27909), .O(n2_adj_4340)) /* synthesis syn_instantiated=1 */ ;
    defparam add_41_3_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_41_3 (.CI(n27909), .I0(\FRAME_MATCHER.i [1]), .I1(GND_net), 
            .CO(n27910));
    SB_LUT4 i1_2_lut_adj_878 (.I0(\data_out_frame[6] [6]), .I1(\data_out_frame[11] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n33107));   // verilog/coms.v(75[16:27])
    defparam i1_2_lut_adj_878.LUT_INIT = 16'h6666;
    SB_LUT4 i545_2_lut (.I0(\data_out_frame[8] [7]), .I1(\data_out_frame[8] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n1301));   // verilog/coms.v(70[16:27])
    defparam i545_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut (.I0(\data_out_frame[9] [0]), .I1(\data_out_frame[9] [2]), 
            .I2(\data_out_frame[11] [3]), .I3(GND_net), .O(n16672));
    defparam i2_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 i3_4_lut_adj_879 (.I0(n16163), .I1(n16687), .I2(n16880), .I3(n16525), 
            .O(n33313));
    defparam i3_4_lut_adj_879.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut (.I0(\data_out_frame[9] [4]), .I1(\data_out_frame[12] [0]), 
            .I2(n33313), .I3(n6), .O(n33066));   // verilog/coms.v(84[17:63])
    defparam i4_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_880 (.I0(\data_out_frame[12] [7]), .I1(n16304), 
            .I2(GND_net), .I3(GND_net), .O(n33427));   // verilog/coms.v(74[16:27])
    defparam i1_2_lut_adj_880.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_881 (.I0(\data_out_frame[9] [5]), .I1(n33115), 
            .I2(GND_net), .I3(GND_net), .O(n16548));
    defparam i1_2_lut_adj_881.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_882 (.I0(\data_out_frame[11] [7]), .I1(n33066), 
            .I2(GND_net), .I3(GND_net), .O(n30801));   // verilog/coms.v(84[17:63])
    defparam i1_2_lut_adj_882.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_883 (.I0(\data_out_frame[7] [1]), .I1(\data_out_frame[7] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n16521));
    defparam i1_2_lut_adj_883.LUT_INIT = 16'h6666;
    SB_DFF data_in_frame_0__i64 (.Q(\data_in_frame[7] [7]), .C(clk32MHz), 
           .D(n18073));   // verilog/coms.v(126[12] 293[6])
    SB_DFF PWMLimit_i0_i17 (.Q(PWMLimit[17]), .C(clk32MHz), .D(n18202));   // verilog/coms.v(126[12] 293[6])
    SB_DFF PWMLimit_i0_i18 (.Q(PWMLimit[18]), .C(clk32MHz), .D(n18203));   // verilog/coms.v(126[12] 293[6])
    SB_DFF PWMLimit_i0_i19 (.Q(PWMLimit[19]), .C(clk32MHz), .D(n18204));   // verilog/coms.v(126[12] 293[6])
    SB_DFF PWMLimit_i0_i20 (.Q(PWMLimit[20]), .C(clk32MHz), .D(n18205));   // verilog/coms.v(126[12] 293[6])
    SB_DFF PWMLimit_i0_i21 (.Q(PWMLimit[21]), .C(clk32MHz), .D(n18206));   // verilog/coms.v(126[12] 293[6])
    SB_DFF PWMLimit_i0_i22 (.Q(PWMLimit[22]), .C(clk32MHz), .D(n18207));   // verilog/coms.v(126[12] 293[6])
    SB_DFF PWMLimit_i0_i23 (.Q(PWMLimit[23]), .C(clk32MHz), .D(n18208));   // verilog/coms.v(126[12] 293[6])
    SB_DFF PWMLimit_i0_i9 (.Q(PWMLimit[9]), .C(clk32MHz), .D(n18194));   // verilog/coms.v(126[12] 293[6])
    SB_DFF PWMLimit_i0_i10 (.Q(PWMLimit[10]), .C(clk32MHz), .D(n18195));   // verilog/coms.v(126[12] 293[6])
    SB_DFF PWMLimit_i0_i11 (.Q(PWMLimit[11]), .C(clk32MHz), .D(n18196));   // verilog/coms.v(126[12] 293[6])
    SB_DFF PWMLimit_i0_i12 (.Q(PWMLimit[12]), .C(clk32MHz), .D(n18197));   // verilog/coms.v(126[12] 293[6])
    SB_DFF PWMLimit_i0_i13 (.Q(PWMLimit[13]), .C(clk32MHz), .D(n18198));   // verilog/coms.v(126[12] 293[6])
    SB_DFF PWMLimit_i0_i14 (.Q(PWMLimit[14]), .C(clk32MHz), .D(n18199));   // verilog/coms.v(126[12] 293[6])
    SB_DFF data_in_frame_0__i174 (.Q(\data_in_frame[21] [5]), .C(clk32MHz), 
           .D(n18183));   // verilog/coms.v(126[12] 293[6])
    SB_DFF data_in_frame_0__i175 (.Q(\data_in_frame[21] [6]), .C(clk32MHz), 
           .D(n18184));   // verilog/coms.v(126[12] 293[6])
    SB_DFF \FRAME_MATCHER.state_i1  (.Q(\FRAME_MATCHER.state [1]), .C(clk32MHz), 
           .D(n34206));   // verilog/coms.v(126[12] 293[6])
    SB_DFF \FRAME_MATCHER.state_i2  (.Q(\FRAME_MATCHER.state [2]), .C(clk32MHz), 
           .D(n38508));   // verilog/coms.v(126[12] 293[6])
    SB_DFF data_in_frame_0__i63 (.Q(\data_in_frame[7] [6]), .C(clk32MHz), 
           .D(n18072));   // verilog/coms.v(126[12] 293[6])
    SB_DFF data_in_frame_0__i62 (.Q(\data_in_frame[7] [5]), .C(clk32MHz), 
           .D(n18071));   // verilog/coms.v(126[12] 293[6])
    SB_DFF data_in_frame_0__i61 (.Q(\data_in_frame[7] [4]), .C(clk32MHz), 
           .D(n18070));   // verilog/coms.v(126[12] 293[6])
    SB_DFF data_in_frame_0__i160 (.Q(\data_in_frame[19] [7]), .C(clk32MHz), 
           .D(n18169));   // verilog/coms.v(126[12] 293[6])
    SB_DFF data_in_frame_0__i60 (.Q(\data_in_frame[7] [3]), .C(clk32MHz), 
           .D(n18069));   // verilog/coms.v(126[12] 293[6])
    SB_DFF data_in_frame_0__i59 (.Q(\data_in_frame[7] [2]), .C(clk32MHz), 
           .D(n18068));   // verilog/coms.v(126[12] 293[6])
    SB_DFF PWMLimit_i0_i15 (.Q(PWMLimit[15]), .C(clk32MHz), .D(n18200));   // verilog/coms.v(126[12] 293[6])
    SB_DFF PWMLimit_i0_i16 (.Q(PWMLimit[16]), .C(clk32MHz), .D(n18201));   // verilog/coms.v(126[12] 293[6])
    SB_DFF data_in_frame_0__i176 (.Q(\data_in_frame[21] [7]), .C(clk32MHz), 
           .D(n18185));   // verilog/coms.v(126[12] 293[6])
    SB_DFF PWMLimit_i0_i1 (.Q(PWMLimit[1]), .C(clk32MHz), .D(n18186));   // verilog/coms.v(126[12] 293[6])
    SB_DFF PWMLimit_i0_i2 (.Q(PWMLimit[2]), .C(clk32MHz), .D(n18187));   // verilog/coms.v(126[12] 293[6])
    SB_DFF PWMLimit_i0_i3 (.Q(PWMLimit[3]), .C(clk32MHz), .D(n18188));   // verilog/coms.v(126[12] 293[6])
    SB_DFF PWMLimit_i0_i4 (.Q(PWMLimit[4]), .C(clk32MHz), .D(n18189));   // verilog/coms.v(126[12] 293[6])
    SB_DFF PWMLimit_i0_i5 (.Q(PWMLimit[5]), .C(clk32MHz), .D(n18190));   // verilog/coms.v(126[12] 293[6])
    SB_DFF PWMLimit_i0_i6 (.Q(PWMLimit[6]), .C(clk32MHz), .D(n18191));   // verilog/coms.v(126[12] 293[6])
    SB_DFF PWMLimit_i0_i7 (.Q(PWMLimit[7]), .C(clk32MHz), .D(n18192));   // verilog/coms.v(126[12] 293[6])
    SB_DFF PWMLimit_i0_i8 (.Q(PWMLimit[8]), .C(clk32MHz), .D(n18193));   // verilog/coms.v(126[12] 293[6])
    SB_DFF data_in_frame_0__i172 (.Q(\data_in_frame[21] [3]), .C(clk32MHz), 
           .D(n18181));   // verilog/coms.v(126[12] 293[6])
    SB_DFF data_in_frame_0__i173 (.Q(\data_in_frame[21] [4]), .C(clk32MHz), 
           .D(n18182));   // verilog/coms.v(126[12] 293[6])
    SB_DFF data_in_frame_0__i170 (.Q(\data_in_frame[21] [1]), .C(clk32MHz), 
           .D(n18179));   // verilog/coms.v(126[12] 293[6])
    SB_DFF data_in_frame_0__i171 (.Q(\data_in_frame[21] [2]), .C(clk32MHz), 
           .D(n18180));   // verilog/coms.v(126[12] 293[6])
    SB_DFF data_in_frame_0__i168 (.Q(\data_in_frame[20] [7]), .C(clk32MHz), 
           .D(n18177));   // verilog/coms.v(126[12] 293[6])
    SB_DFF data_in_frame_0__i169 (.Q(\data_in_frame[21] [0]), .C(clk32MHz), 
           .D(n18178));   // verilog/coms.v(126[12] 293[6])
    SB_DFF data_in_frame_0__i166 (.Q(\data_in_frame[20] [5]), .C(clk32MHz), 
           .D(n18175));   // verilog/coms.v(126[12] 293[6])
    SB_DFF data_in_frame_0__i167 (.Q(\data_in_frame[20] [6]), .C(clk32MHz), 
           .D(n18176));   // verilog/coms.v(126[12] 293[6])
    SB_DFF data_in_frame_0__i164 (.Q(\data_in_frame[20] [3]), .C(clk32MHz), 
           .D(n18173));   // verilog/coms.v(126[12] 293[6])
    SB_DFF data_in_frame_0__i165 (.Q(\data_in_frame[20] [4]), .C(clk32MHz), 
           .D(n18174));   // verilog/coms.v(126[12] 293[6])
    SB_DFF data_in_frame_0__i58 (.Q(\data_in_frame[7] [1]), .C(clk32MHz), 
           .D(n18067));   // verilog/coms.v(126[12] 293[6])
    SB_DFF data_in_frame_0__i161 (.Q(\data_in_frame[20] [0]), .C(clk32MHz), 
           .D(n18170));   // verilog/coms.v(126[12] 293[6])
    SB_DFF data_in_frame_0__i162 (.Q(\data_in_frame[20] [1]), .C(clk32MHz), 
           .D(n18171));   // verilog/coms.v(126[12] 293[6])
    SB_DFF data_in_frame_0__i163 (.Q(\data_in_frame[20] [2]), .C(clk32MHz), 
           .D(n18172));   // verilog/coms.v(126[12] 293[6])
    SB_DFF data_in_frame_0__i57 (.Q(\data_in_frame[7] [0]), .C(clk32MHz), 
           .D(n18066));   // verilog/coms.v(126[12] 293[6])
    SB_DFF data_in_frame_0__i114 (.Q(\data_in_frame[14] [1]), .C(clk32MHz), 
           .D(n18123));   // verilog/coms.v(126[12] 293[6])
    SB_DFF data_in_frame_0__i113 (.Q(\data_in_frame[14] [0]), .C(clk32MHz), 
           .D(n18122));   // verilog/coms.v(126[12] 293[6])
    SB_DFF data_in_frame_0__i112 (.Q(\data_in_frame[13] [7]), .C(clk32MHz), 
           .D(n18121));   // verilog/coms.v(126[12] 293[6])
    SB_DFF data_in_frame_0__i111 (.Q(\data_in_frame[13] [6]), .C(clk32MHz), 
           .D(n18120));   // verilog/coms.v(126[12] 293[6])
    SB_DFF data_in_frame_0__i110 (.Q(\data_in_frame[13] [5]), .C(clk32MHz), 
           .D(n18119));   // verilog/coms.v(126[12] 293[6])
    SB_DFF data_in_frame_0__i109 (.Q(\data_in_frame[13] [4]), .C(clk32MHz), 
           .D(n18118));   // verilog/coms.v(126[12] 293[6])
    SB_DFF data_in_frame_0__i108 (.Q(\data_in_frame[13] [3]), .C(clk32MHz), 
           .D(n18117));   // verilog/coms.v(126[12] 293[6])
    SB_DFF data_in_frame_0__i127 (.Q(\data_in_frame[15] [6]), .C(clk32MHz), 
           .D(n18136));   // verilog/coms.v(126[12] 293[6])
    SB_DFF data_in_frame_0__i56 (.Q(\data_in_frame[6] [7]), .C(clk32MHz), 
           .D(n18065));   // verilog/coms.v(126[12] 293[6])
    SB_DFF data_in_frame_0__i55 (.Q(\data_in_frame[6] [6]), .C(clk32MHz), 
           .D(n18064));   // verilog/coms.v(126[12] 293[6])
    SB_DFF data_in_frame_0__i54 (.Q(\data_in_frame[6] [5]), .C(clk32MHz), 
           .D(n18063));   // verilog/coms.v(126[12] 293[6])
    SB_LUT4 i1_2_lut_adj_884 (.I0(\data_out_frame[6] [7]), .I1(\data_out_frame[6] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n16229));   // verilog/coms.v(70[16:27])
    defparam i1_2_lut_adj_884.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_885 (.I0(\data_out_frame[5] [2]), .I1(\data_out_frame[5] [0]), 
            .I2(\data_out_frame[7] [3]), .I3(GND_net), .O(n16525));
    defparam i2_3_lut_adj_885.LUT_INIT = 16'h9696;
    SB_DFF data_in_frame_0__i53 (.Q(\data_in_frame[6] [4]), .C(clk32MHz), 
           .D(n18062));   // verilog/coms.v(126[12] 293[6])
    SB_DFF data_in_frame_0__i52 (.Q(\data_in_frame[6] [3]), .C(clk32MHz), 
           .D(n18061));   // verilog/coms.v(126[12] 293[6])
    SB_DFF data_in_frame_0__i51 (.Q(\data_in_frame[6] [2]), .C(clk32MHz), 
           .D(n18060));   // verilog/coms.v(126[12] 293[6])
    SB_DFF data_in_frame_0__i50 (.Q(\data_in_frame[6] [1]), .C(clk32MHz), 
           .D(n18059));   // verilog/coms.v(126[12] 293[6])
    SB_DFF data_in_frame_0__i49 (.Q(\data_in_frame[6] [0]), .C(clk32MHz), 
           .D(n18058));   // verilog/coms.v(126[12] 293[6])
    SB_DFF data_in_frame_0__i48 (.Q(\data_in_frame[5] [7]), .C(clk32MHz), 
           .D(n18057));   // verilog/coms.v(126[12] 293[6])
    SB_DFF data_in_frame_0__i47 (.Q(\data_in_frame[5] [6]), .C(clk32MHz), 
           .D(n18056));   // verilog/coms.v(126[12] 293[6])
    SB_DFF data_in_frame_0__i46 (.Q(\data_in_frame[5] [5]), .C(clk32MHz), 
           .D(n18055));   // verilog/coms.v(126[12] 293[6])
    SB_DFF data_in_frame_0__i45 (.Q(\data_in_frame[5] [4]), .C(clk32MHz), 
           .D(n18054));   // verilog/coms.v(126[12] 293[6])
    SB_DFF data_in_frame_0__i44 (.Q(\data_in_frame[5] [3]), .C(clk32MHz), 
           .D(n18053));   // verilog/coms.v(126[12] 293[6])
    SB_DFF data_in_frame_0__i43 (.Q(\data_in_frame[5] [2]), .C(clk32MHz), 
           .D(n18052));   // verilog/coms.v(126[12] 293[6])
    SB_DFF data_in_frame_0__i42 (.Q(\data_in_frame[5] [1]), .C(clk32MHz), 
           .D(n18051));   // verilog/coms.v(126[12] 293[6])
    SB_DFF data_in_frame_0__i107 (.Q(\data_in_frame[13] [2]), .C(clk32MHz), 
           .D(n18116));   // verilog/coms.v(126[12] 293[6])
    SB_LUT4 i3_4_lut_adj_886 (.I0(\data_in_frame[10] [0]), .I1(n33330), 
            .I2(n33127), .I3(\data_in_frame[12] [2]), .O(n33508));   // verilog/coms.v(84[17:28])
    defparam i3_4_lut_adj_886.LUT_INIT = 16'h6996;
    SB_DFF data_in_frame_0__i41 (.Q(\data_in_frame[5] [0]), .C(clk32MHz), 
           .D(n18050));   // verilog/coms.v(126[12] 293[6])
    SB_DFF data_in_frame_0__i106 (.Q(\data_in_frame[13] [1]), .C(clk32MHz), 
           .D(n18115));   // verilog/coms.v(126[12] 293[6])
    SB_DFF data_in_frame_0__i40 (.Q(\data_in_frame[4] [7]), .C(clk32MHz), 
           .D(n18049));   // verilog/coms.v(126[12] 293[6])
    SB_DFF data_in_frame_0__i105 (.Q(\data_in_frame[13] [0]), .C(clk32MHz), 
           .D(n18114));   // verilog/coms.v(126[12] 293[6])
    SB_DFF data_in_frame_0__i39 (.Q(\data_in_frame[4] [6]), .C(clk32MHz), 
           .D(n18048));   // verilog/coms.v(126[12] 293[6])
    SB_DFF data_in_frame_0__i38 (.Q(\data_in_frame[4] [5]), .C(clk32MHz), 
           .D(n18047));   // verilog/coms.v(126[12] 293[6])
    SB_DFF data_in_frame_0__i37 (.Q(\data_in_frame[4] [4]), .C(clk32MHz), 
           .D(n18046));   // verilog/coms.v(126[12] 293[6])
    SB_DFF data_in_frame_0__i36 (.Q(\data_in_frame[4] [3]), .C(clk32MHz), 
           .D(n18045));   // verilog/coms.v(126[12] 293[6])
    SB_DFF data_in_frame_0__i104 (.Q(\data_in_frame[12] [7]), .C(clk32MHz), 
           .D(n18113));   // verilog/coms.v(126[12] 293[6])
    SB_DFF data_in_frame_0__i103 (.Q(\data_in_frame[12] [6]), .C(clk32MHz), 
           .D(n18112));   // verilog/coms.v(126[12] 293[6])
    SB_LUT4 i1_2_lut_adj_887 (.I0(n1251), .I1(\data_out_frame[11] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_4341));   // verilog/coms.v(75[16:43])
    defparam i1_2_lut_adj_887.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_888 (.I0(n33241), .I1(n15783), .I2(n1254), .I3(n6_adj_4341), 
            .O(n33265));   // verilog/coms.v(75[16:43])
    defparam i4_4_lut_adj_888.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_889 (.I0(n13947), .I1(n31), .I2(n16162), .I3(GND_net), 
            .O(n34066));
    defparam i2_3_lut_adj_889.LUT_INIT = 16'hfefe;
    SB_LUT4 mux_1255_i2_3_lut (.I0(\data_in_frame[19] [1]), .I1(\data_in_frame[3] [1]), 
            .I2(n4995), .I3(GND_net), .O(n4997));
    defparam mux_1255_i2_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF data_in_frame_0__i102 (.Q(\data_in_frame[12] [5]), .C(clk32MHz), 
           .D(n18111));   // verilog/coms.v(126[12] 293[6])
    SB_LUT4 mux_1255_i3_3_lut (.I0(\data_in_frame[19] [2]), .I1(\data_in_frame[3] [2]), 
            .I2(n4995), .I3(GND_net), .O(n4998));
    defparam mux_1255_i3_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_1255_i4_3_lut (.I0(\data_in_frame[19] [3]), .I1(\data_in_frame[3] [3]), 
            .I2(n4995), .I3(GND_net), .O(n4999));
    defparam mux_1255_i4_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2_3_lut_adj_890 (.I0(n33073), .I1(\data_out_frame[13] [6]), 
            .I2(\data_out_frame[13] [4]), .I3(GND_net), .O(n33204));   // verilog/coms.v(84[17:63])
    defparam i2_3_lut_adj_890.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_adj_891 (.I0(n1251), .I1(n33256), .I2(n1254), .I3(GND_net), 
            .O(n16946));   // verilog/coms.v(74[16:43])
    defparam i2_3_lut_adj_891.LUT_INIT = 16'h9696;
    SB_LUT4 mux_1255_i5_3_lut (.I0(\data_in_frame[19] [4]), .I1(\data_in_frame[3] [4]), 
            .I2(n4995), .I3(GND_net), .O(n5000));
    defparam mux_1255_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12_4_lut (.I0(n33540), .I1(n30801), .I2(n16548), .I3(n33427), 
            .O(n32));
    defparam i12_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 mux_1255_i6_3_lut (.I0(\data_in_frame[19] [5]), .I1(\data_in_frame[3] [5]), 
            .I2(n4995), .I3(GND_net), .O(n5001));
    defparam mux_1255_i6_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16_4_lut (.I0(\data_out_frame[13] [0]), .I1(n32), .I2(n22), 
            .I3(n31287), .O(n36));
    defparam i16_4_lut.LUT_INIT = 16'h9669;
    SB_LUT4 i14_4_lut (.I0(n33494), .I1(n33253), .I2(n33287), .I3(\data_out_frame[9] [4]), 
            .O(n34));
    defparam i14_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i15_4_lut (.I0(n16545), .I1(\data_out_frame[10] [4]), .I2(n30857), 
            .I3(\data_out_frame[12] [1]), .O(n35));
    defparam i15_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i13_4_lut (.I0(\data_out_frame[12] [6]), .I1(n17068), .I2(\data_out_frame[11] [1]), 
            .I3(n33610), .O(n33));
    defparam i13_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 mux_1255_i7_3_lut (.I0(\data_in_frame[19] [6]), .I1(\data_in_frame[3] [6]), 
            .I2(n4995), .I3(GND_net), .O(n5002));
    defparam mux_1255_i7_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_1255_i8_3_lut (.I0(\data_in_frame[19] [7]), .I1(\data_in_frame[3] [7]), 
            .I2(n4995), .I3(GND_net), .O(n5003));
    defparam mux_1255_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_1255_i9_3_lut (.I0(\data_in_frame[18] [0]), .I1(\data_in_frame[2] [0]), 
            .I2(n4995), .I3(GND_net), .O(n5004));
    defparam mux_1255_i9_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i19_4_lut (.I0(n33), .I1(n35), .I2(n34), .I3(n36), .O(n31223));
    defparam i19_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i13223_3_lut_4_lut (.I0(n8), .I1(n32959), .I2(rx_data[2]), 
            .I3(\data_in_frame[5] [2]), .O(n18052));
    defparam i13223_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 mux_1255_i10_3_lut (.I0(\data_in_frame[18] [1]), .I1(\data_in_frame[2] [1]), 
            .I2(n4995), .I3(GND_net), .O(n5005));
    defparam mux_1255_i10_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13224_3_lut_4_lut (.I0(n8), .I1(n32959), .I2(rx_data[3]), 
            .I3(\data_in_frame[5] [3]), .O(n18053));
    defparam i13224_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i4_4_lut_adj_892 (.I0(\data_out_frame[13] [5]), .I1(n16946), 
            .I2(\data_out_frame[11] [4]), .I3(n33204), .O(n10_adj_4342));
    defparam i4_4_lut_adj_892.LUT_INIT = 16'h6996;
    SB_LUT4 i5_3_lut (.I0(\data_out_frame[13] [7]), .I1(n10_adj_4342), .I2(n31223), 
            .I3(GND_net), .O(n34521));
    defparam i5_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 i13225_3_lut_4_lut (.I0(n8), .I1(n32959), .I2(rx_data[4]), 
            .I3(\data_in_frame[5] [4]), .O(n18054));
    defparam i13225_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13226_3_lut_4_lut (.I0(n8), .I1(n32959), .I2(rx_data[5]), 
            .I3(\data_in_frame[5] [5]), .O(n18055));
    defparam i13226_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_893 (.I0(\data_out_frame[13] [2]), .I1(\data_out_frame[13] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n16676));
    defparam i1_2_lut_adj_893.LUT_INIT = 16'h6666;
    SB_LUT4 mux_1255_i11_3_lut (.I0(\data_in_frame[18] [2]), .I1(\data_in_frame[2] [2]), 
            .I2(n4995), .I3(GND_net), .O(n5006));
    defparam mux_1255_i11_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4_4_lut_adj_894 (.I0(\data_out_frame[16] [0]), .I1(n31188), 
            .I2(\data_out_frame[13] [7]), .I3(n6_adj_4343), .O(n33303));
    defparam i4_4_lut_adj_894.LUT_INIT = 16'h6996;
    SB_LUT4 mux_1255_i12_3_lut (.I0(\data_in_frame[18] [3]), .I1(\data_in_frame[2] [3]), 
            .I2(n4995), .I3(GND_net), .O(n5007));
    defparam mux_1255_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_adj_895 (.I0(n15783), .I1(n33253), .I2(GND_net), 
            .I3(GND_net), .O(n30451));
    defparam i1_2_lut_adj_895.LUT_INIT = 16'h6666;
    SB_LUT4 mux_1255_i13_3_lut (.I0(\data_in_frame[18] [4]), .I1(\data_in_frame[2] [4]), 
            .I2(n4995), .I3(GND_net), .O(n5008));
    defparam mux_1255_i13_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_adj_896 (.I0(\FRAME_MATCHER.state [1]), .I1(\FRAME_MATCHER.state [0]), 
            .I2(GND_net), .I3(GND_net), .O(n13554));
    defparam i1_2_lut_adj_896.LUT_INIT = 16'heeee;
    SB_LUT4 i27179_4_lut (.I0(n25118), .I1(\FRAME_MATCHER.state [3]), .I2(\FRAME_MATCHER.state [2]), 
            .I3(n13554), .O(n33773));
    defparam i27179_4_lut.LUT_INIT = 16'heeea;
    SB_LUT4 i1_2_lut_adj_897 (.I0(\data_out_frame[18] [2]), .I1(\data_out_frame[18] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n16195));
    defparam i1_2_lut_adj_897.LUT_INIT = 16'h6666;
    SB_LUT4 mux_1255_i14_3_lut (.I0(\data_in_frame[18] [5]), .I1(\data_in_frame[2] [5]), 
            .I2(n4995), .I3(GND_net), .O(n5009));
    defparam mux_1255_i14_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3_3_lut (.I0(n16000), .I1(\FRAME_MATCHER.state [1]), .I2(n24786), 
            .I3(GND_net), .O(n8_adj_4344));
    defparam i3_3_lut.LUT_INIT = 16'hbfbf;
    SB_LUT4 mux_833_i1_4_lut (.I0(n7), .I1(\FRAME_MATCHER.state [3]), .I2(n5069), 
            .I3(n8_adj_4344), .O(n3693[0]));   // verilog/coms.v(144[4] 292[11])
    defparam mux_833_i1_4_lut.LUT_INIT = 16'h0c5c;
    SB_LUT4 i6_4_lut_adj_898 (.I0(n33520), .I1(\data_out_frame[13] [6]), 
            .I2(n33060), .I3(\data_out_frame[6] [6]), .O(n14_adj_4345));
    defparam i6_4_lut_adj_898.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut_adj_899 (.I0(\data_out_frame[16] [2]), .I1(n14_adj_4345), 
            .I2(n10_adj_4346), .I3(n1251), .O(n16711));
    defparam i7_4_lut_adj_899.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_900 (.I0(n30451), .I1(n33303), .I2(\data_out_frame[15] [6]), 
            .I3(n16676), .O(n34672));
    defparam i3_4_lut_adj_900.LUT_INIT = 16'h6996;
    SB_LUT4 mux_1255_i15_3_lut (.I0(\data_in_frame[18] [6]), .I1(\data_in_frame[2] [6]), 
            .I2(n4995), .I3(GND_net), .O(n5010));
    defparam mux_1255_i15_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i31535_4_lut (.I0(\FRAME_MATCHER.state [3]), .I1(n33789), .I2(\FRAME_MATCHER.state [1]), 
            .I3(n33773), .O(n35075));
    defparam i31535_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 i3_4_lut_adj_901 (.I0(\data_out_frame[20] [4]), .I1(n34672), 
            .I2(n16711), .I3(n16195), .O(n33201));
    defparam i3_4_lut_adj_901.LUT_INIT = 16'h9669;
    SB_LUT4 i2_3_lut_adj_902 (.I0(n33020), .I1(n33371), .I2(\data_out_frame[20] [6]), 
            .I3(GND_net), .O(n16647));
    defparam i2_3_lut_adj_902.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_adj_903 (.I0(\FRAME_MATCHER.state [0]), .I1(\FRAME_MATCHER.state [2]), 
            .I2(n42), .I3(GND_net), .O(n34894));
    defparam i2_3_lut_adj_903.LUT_INIT = 16'h4040;
    SB_LUT4 i1_4_lut (.I0(n5069), .I1(n33773), .I2(n34894), .I3(n35045), 
            .O(n4_c));
    defparam i1_4_lut.LUT_INIT = 16'hecee;
    SB_LUT4 mux_1255_i16_3_lut (.I0(\data_in_frame[18] [7]), .I1(\data_in_frame[2] [7]), 
            .I2(n4995), .I3(GND_net), .O(n5011));
    defparam mux_1255_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF data_in_frame_0__i35 (.Q(\data_in_frame[4] [2]), .C(clk32MHz), 
           .D(n18044));   // verilog/coms.v(126[12] 293[6])
    SB_LUT4 i31495_4_lut (.I0(n5069), .I1(\FRAME_MATCHER.state [3]), .I2(n33634), 
            .I3(n4_c), .O(n33636));
    defparam i31495_4_lut.LUT_INIT = 16'h001b;
    SB_LUT4 mux_1255_i17_3_lut (.I0(\data_in_frame[17] [0]), .I1(\data_in_frame[1] [0]), 
            .I2(n4995), .I3(GND_net), .O(n5012));
    defparam mux_1255_i17_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_1255_i18_3_lut (.I0(\data_in_frame[17] [1]), .I1(\data_in_frame[1] [1]), 
            .I2(n4995), .I3(GND_net), .O(n5013));
    defparam mux_1255_i18_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_1255_i19_3_lut (.I0(\data_in_frame[17] [2]), .I1(\data_in_frame[1] [2]), 
            .I2(n4995), .I3(GND_net), .O(n5014));
    defparam mux_1255_i19_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_1255_i20_3_lut (.I0(\data_in_frame[17] [3]), .I1(\data_in_frame[1] [3]), 
            .I2(n4995), .I3(GND_net), .O(n5015));
    defparam mux_1255_i20_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_1255_i21_3_lut (.I0(\data_in_frame[17] [4]), .I1(\data_in_frame[1] [4]), 
            .I2(n4995), .I3(GND_net), .O(n5016));
    defparam mux_1255_i21_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_1255_i22_3_lut (.I0(\data_in_frame[17] [5]), .I1(\data_in_frame[1] [5]), 
            .I2(n4995), .I3(GND_net), .O(n5017));
    defparam mux_1255_i22_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_1255_i23_3_lut (.I0(\data_in_frame[17] [6]), .I1(\data_in_frame[1] [6]), 
            .I2(n4995), .I3(GND_net), .O(n5018));
    defparam mux_1255_i23_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2_3_lut_adj_904 (.I0(n31_adj_4347), .I1(\FRAME_MATCHER.state [1]), 
            .I2(n13947), .I3(GND_net), .O(n4995));
    defparam i2_3_lut_adj_904.LUT_INIT = 16'h0404;
    SB_LUT4 equal_1520_i15_2_lut (.I0(Kp_23__N_993), .I1(\data_in_frame[4] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n15));   // verilog/coms.v(232[9:81])
    defparam equal_1520_i15_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i5_3_lut_adj_905 (.I0(n16791), .I1(Kp_23__N_996), .I2(\data_in_frame[4] [7]), 
            .I3(GND_net), .O(n21));
    defparam i5_3_lut_adj_905.LUT_INIT = 16'hbebe;
    SB_LUT4 i12_4_lut_adj_906 (.I0(n33127), .I1(n31230), .I2(n15), .I3(n30217), 
            .O(n28));
    defparam i12_4_lut_adj_906.LUT_INIT = 16'hfeff;
    SB_LUT4 i10_4_lut (.I0(n6_adj_4348), .I1(n16722), .I2(n16380), .I3(n16834), 
            .O(n26));
    defparam i10_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i11_4_lut (.I0(n21), .I1(n16335), .I2(Kp_23__N_1046), .I3(\data_in_frame[5] [7]), 
            .O(n27));
    defparam i11_4_lut.LUT_INIT = 16'hbffb;
    SB_LUT4 i9_4_lut (.I0(n16608), .I1(n31002), .I2(n16765), .I3(n16384), 
            .O(n25));
    defparam i9_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i15_4_lut_adj_907 (.I0(n25), .I1(n27), .I2(n26), .I3(n28), 
            .O(n31_adj_4347));
    defparam i15_4_lut_adj_907.LUT_INIT = 16'hfffe;
    SB_LUT4 i6_4_lut_adj_908 (.I0(\data_in_frame[0] [6]), .I1(\data_in_frame[0] [1]), 
            .I2(\data_in_frame[0] [4]), .I3(\data_in_frame[0] [2]), .O(n14_adj_4349));
    defparam i6_4_lut_adj_908.LUT_INIT = 16'hfbff;
    SB_LUT4 i1_2_lut_adj_909 (.I0(\data_in_frame[0] [3]), .I1(\data_in_frame[0] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n9_adj_4350));
    defparam i1_2_lut_adj_909.LUT_INIT = 16'heeee;
    SB_LUT4 i7_4_lut_adj_910 (.I0(n9_adj_4350), .I1(n14_adj_4349), .I2(\data_in_frame[0] [5]), 
            .I3(\data_in_frame[0] [0]), .O(n13947));
    defparam i7_4_lut_adj_910.LUT_INIT = 16'hfeff;
    SB_LUT4 i1_2_lut_adj_911 (.I0(\data_in_frame[7] [7]), .I1(n33508), .I2(GND_net), 
            .I3(GND_net), .O(n6_adj_4351));   // verilog/coms.v(84[17:28])
    defparam i1_2_lut_adj_911.LUT_INIT = 16'h6666;
    SB_LUT4 i1_4_lut_adj_912 (.I0(n13947), .I1(n31), .I2(n31_adj_4347), 
            .I3(\FRAME_MATCHER.state [1]), .O(n42));   // verilog/coms.v(111[11:16])
    defparam i1_4_lut_adj_912.LUT_INIT = 16'hfaee;
    SB_LUT4 i1_2_lut_adj_913 (.I0(n42), .I1(\FRAME_MATCHER.state [3]), .I2(GND_net), 
            .I3(GND_net), .O(n6_adj_4352));
    defparam i1_2_lut_adj_913.LUT_INIT = 16'heeee;
    SB_LUT4 i4_4_lut_adj_914 (.I0(\FRAME_MATCHER.state [0]), .I1(\FRAME_MATCHER.state [2]), 
            .I2(n25118), .I3(n6_adj_4352), .O(n35492));
    defparam i4_4_lut_adj_914.LUT_INIT = 16'hfffb;
    SB_LUT4 mux_1255_i24_3_lut (.I0(\data_in_frame[17] [7]), .I1(\data_in_frame[1] [7]), 
            .I2(n4995), .I3(GND_net), .O(n5019));
    defparam mux_1255_i24_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13227_3_lut_4_lut (.I0(n8), .I1(n32959), .I2(rx_data[6]), 
            .I3(\data_in_frame[5] [6]), .O(n18056));
    defparam i13227_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13228_3_lut_4_lut (.I0(n8), .I1(n32959), .I2(rx_data[7]), 
            .I3(\data_in_frame[5] [7]), .O(n18057));
    defparam i13228_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF data_in_frame_0__i34 (.Q(\data_in_frame[4] [1]), .C(clk32MHz), 
           .D(n18043));   // verilog/coms.v(126[12] 293[6])
    SB_DFF data_in_frame_0__i33 (.Q(\data_in_frame[4] [0]), .C(clk32MHz), 
           .D(n18042));   // verilog/coms.v(126[12] 293[6])
    SB_DFF data_in_frame_0__i32 (.Q(\data_in_frame[3] [7]), .C(clk32MHz), 
           .D(n18041));   // verilog/coms.v(126[12] 293[6])
    SB_DFF data_in_frame_0__i31 (.Q(\data_in_frame[3] [6]), .C(clk32MHz), 
           .D(n18040));   // verilog/coms.v(126[12] 293[6])
    SB_DFF data_in_frame_0__i30 (.Q(\data_in_frame[3] [5]), .C(clk32MHz), 
           .D(n18039));   // verilog/coms.v(126[12] 293[6])
    SB_DFF data_in_frame_0__i29 (.Q(\data_in_frame[3] [4]), .C(clk32MHz), 
           .D(n18038));   // verilog/coms.v(126[12] 293[6])
    SB_DFF data_in_frame_0__i28 (.Q(\data_in_frame[3] [3]), .C(clk32MHz), 
           .D(n18037));   // verilog/coms.v(126[12] 293[6])
    SB_DFF data_in_frame_0__i27 (.Q(\data_in_frame[3] [2]), .C(clk32MHz), 
           .D(n18036));   // verilog/coms.v(126[12] 293[6])
    SB_DFF data_in_frame_0__i26 (.Q(\data_in_frame[3] [1]), .C(clk32MHz), 
           .D(n18035));   // verilog/coms.v(126[12] 293[6])
    SB_DFF data_in_frame_0__i25 (.Q(\data_in_frame[3] [0]), .C(clk32MHz), 
           .D(n18034));   // verilog/coms.v(126[12] 293[6])
    SB_DFF data_in_frame_0__i24 (.Q(\data_in_frame[2] [7]), .C(clk32MHz), 
           .D(n18033));   // verilog/coms.v(126[12] 293[6])
    SB_DFF data_in_frame_0__i23 (.Q(\data_in_frame[2] [6]), .C(clk32MHz), 
           .D(n18032));   // verilog/coms.v(126[12] 293[6])
    SB_DFF data_in_frame_0__i22 (.Q(\data_in_frame[2] [5]), .C(clk32MHz), 
           .D(n18031));   // verilog/coms.v(126[12] 293[6])
    SB_DFF data_in_frame_0__i21 (.Q(\data_in_frame[2] [4]), .C(clk32MHz), 
           .D(n18030));   // verilog/coms.v(126[12] 293[6])
    SB_DFF data_in_frame_0__i20 (.Q(\data_in_frame[2] [3]), .C(clk32MHz), 
           .D(n18029));   // verilog/coms.v(126[12] 293[6])
    SB_DFF data_in_frame_0__i19 (.Q(\data_in_frame[2] [2]), .C(clk32MHz), 
           .D(n18028));   // verilog/coms.v(126[12] 293[6])
    SB_DFF data_in_frame_0__i18 (.Q(\data_in_frame[2] [1]), .C(clk32MHz), 
           .D(n18027));   // verilog/coms.v(126[12] 293[6])
    SB_DFF data_in_frame_0__i17 (.Q(\data_in_frame[2] [0]), .C(clk32MHz), 
           .D(n18026));   // verilog/coms.v(126[12] 293[6])
    SB_DFF data_in_frame_0__i16 (.Q(\data_in_frame[1] [7]), .C(clk32MHz), 
           .D(n18025));   // verilog/coms.v(126[12] 293[6])
    SB_DFF data_in_frame_0__i15 (.Q(\data_in_frame[1] [6]), .C(clk32MHz), 
           .D(n18024));   // verilog/coms.v(126[12] 293[6])
    SB_DFF data_in_frame_0__i14 (.Q(\data_in_frame[1] [5]), .C(clk32MHz), 
           .D(n18023));   // verilog/coms.v(126[12] 293[6])
    SB_DFF data_in_frame_0__i13 (.Q(\data_in_frame[1] [4]), .C(clk32MHz), 
           .D(n18022));   // verilog/coms.v(126[12] 293[6])
    SB_DFF data_in_frame_0__i12 (.Q(\data_in_frame[1] [3]), .C(clk32MHz), 
           .D(n18021));   // verilog/coms.v(126[12] 293[6])
    SB_DFF data_in_frame_0__i11 (.Q(\data_in_frame[1] [2]), .C(clk32MHz), 
           .D(n18020));   // verilog/coms.v(126[12] 293[6])
    SB_DFF data_in_frame_0__i101 (.Q(\data_in_frame[12] [4]), .C(clk32MHz), 
           .D(n18110));   // verilog/coms.v(126[12] 293[6])
    SB_LUT4 i3_4_lut_adj_915 (.I0(\data_in_frame[19] [7]), .I1(\data_in_frame[17] [7]), 
            .I2(\data_in_frame[20] [1]), .I3(n33186), .O(n34651));
    defparam i3_4_lut_adj_915.LUT_INIT = 16'h6996;
    SB_LUT4 i13213_3_lut_4_lut (.I0(n8_adj_4353), .I1(n32959), .I2(rx_data[0]), 
            .I3(\data_in_frame[4] [0]), .O(n18042));
    defparam i13213_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF data_in_frame_0__i100 (.Q(\data_in_frame[12] [3]), .C(clk32MHz), 
           .D(n18109));   // verilog/coms.v(126[12] 293[6])
    SB_LUT4 i4_4_lut_adj_916 (.I0(n33279), .I1(\data_in_frame[18] [2]), 
            .I2(\data_in_frame[20] [4]), .I3(n33483), .O(n10_adj_4354));
    defparam i4_4_lut_adj_916.LUT_INIT = 16'h6996;
    SB_DFF data_in_frame_0__i99 (.Q(\data_in_frame[12] [2]), .C(clk32MHz), 
           .D(n18108));   // verilog/coms.v(126[12] 293[6])
    SB_DFF data_in_frame_0__i126 (.Q(\data_in_frame[15] [5]), .C(clk32MHz), 
           .D(n18135));   // verilog/coms.v(126[12] 293[6])
    SB_LUT4 i17820_3_lut (.I0(\data_in[0] [2]), .I1(\data_in[1] [2]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n17792));   // verilog/coms.v(89[7:20])
    defparam i17820_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13232_3_lut_4_lut (.I0(n8_adj_4355), .I1(n32959), .I2(rx_data[3]), 
            .I3(\data_in_frame[6] [3]), .O(n18061));
    defparam i13232_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_1_i6_3_lut (.I0(\data_out_frame[5] [1]), 
            .I1(byte_transmit_counter[0]), .I2(byte_transmit_counter_c[2]), 
            .I3(GND_net), .O(n6_adj_4356));   // verilog/coms.v(105[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_1_i6_3_lut.LUT_INIT = 16'hbcbc;
    SB_DFF data_in_frame_0__i125 (.Q(\data_in_frame[15] [4]), .C(clk32MHz), 
           .D(n18134));   // verilog/coms.v(126[12] 293[6])
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_1_i5_3_lut (.I0(\data_out_frame[6] [1]), 
            .I1(\data_out_frame[7] [1]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n5_c));   // verilog/coms.v(105[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_1_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_1_i7_3_lut (.I0(n5_c), .I1(n6_adj_4356), 
            .I2(n37177), .I3(GND_net), .O(n7_adj_4357));   // verilog/coms.v(105[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_1_i7_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i2032929_i1_3_lut (.I0(n38438), .I1(n38444), .I2(byte_transmit_counter_c[2]), 
            .I3(GND_net), .O(n14_adj_4358));
    defparam i2032929_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_2_i6_4_lut (.I0(\data_out_frame[5] [2]), 
            .I1(byte_transmit_counter[0]), .I2(byte_transmit_counter_c[2]), 
            .I3(byte_transmit_counter_c[1]), .O(n6_adj_4359));   // verilog/coms.v(105[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_2_i6_4_lut.LUT_INIT = 16'hb0b3;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_2_i5_3_lut (.I0(\data_out_frame[6] [2]), 
            .I1(\data_out_frame[7] [2]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n5_adj_4360));   // verilog/coms.v(105[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_2_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_2_i7_3_lut (.I0(n5_adj_4360), 
            .I1(n6_adj_4359), .I2(n37177), .I3(GND_net), .O(n7_adj_4361));   // verilog/coms.v(105[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_2_i7_3_lut.LUT_INIT = 16'hacac;
    SB_DFF data_in_frame_0__i124 (.Q(\data_in_frame[15] [3]), .C(clk32MHz), 
           .D(n18133));   // verilog/coms.v(126[12] 293[6])
    SB_LUT4 i13214_3_lut_4_lut (.I0(n8_adj_4353), .I1(n32959), .I2(rx_data[1]), 
            .I3(\data_in_frame[4] [1]), .O(n18043));
    defparam i13214_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2033532_i1_3_lut (.I0(n38348), .I1(n38450), .I2(byte_transmit_counter_c[2]), 
            .I3(GND_net), .O(n14_adj_4362));
    defparam i2033532_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_3_i6_4_lut (.I0(\data_out_frame[5] [3]), 
            .I1(byte_transmit_counter_c[1]), .I2(byte_transmit_counter_c[2]), 
            .I3(byte_transmit_counter[0]), .O(n6_adj_4363));   // verilog/coms.v(105[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_3_i6_4_lut.LUT_INIT = 16'haf03;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_3_i5_3_lut (.I0(\data_out_frame[6] [3]), 
            .I1(\data_out_frame[7] [3]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n5_adj_4364));   // verilog/coms.v(105[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_3_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_3_i7_3_lut (.I0(n5_adj_4364), 
            .I1(n6_adj_4363), .I2(n37177), .I3(GND_net), .O(n7_adj_4365));   // verilog/coms.v(105[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_3_i7_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i2034135_i1_3_lut (.I0(n38342), .I1(n38456), .I2(byte_transmit_counter_c[2]), 
            .I3(GND_net), .O(n14_adj_4366));
    defparam i2034135_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13215_3_lut_4_lut (.I0(n8_adj_4353), .I1(n32959), .I2(rx_data[2]), 
            .I3(\data_in_frame[4] [2]), .O(n18044));
    defparam i13215_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_3_i16_3_lut (.I0(\data_out_frame[16] [3]), 
            .I1(\data_out_frame[17] [3]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n16));   // verilog/coms.v(105[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_3_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13216_3_lut_4_lut (.I0(n8_adj_4353), .I1(n32959), .I2(rx_data[3]), 
            .I3(\data_in_frame[4] [3]), .O(n18045));
    defparam i13216_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13217_3_lut_4_lut (.I0(n8_adj_4353), .I1(n32959), .I2(rx_data[4]), 
            .I3(\data_in_frame[4] [4]), .O(n18046));
    defparam i13217_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_3_i17_3_lut (.I0(\data_out_frame[18] [3]), 
            .I1(\data_out_frame[19] [3]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n17));   // verilog/coms.v(105[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_3_i17_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i30862_2_lut (.I0(\data_out_frame[23] [3]), .I1(byte_transmit_counter[0]), 
            .I2(GND_net), .I3(GND_net), .O(n37271));
    defparam i30862_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i13218_3_lut_4_lut (.I0(n8_adj_4353), .I1(n32959), .I2(rx_data[5]), 
            .I3(\data_in_frame[4] [5]), .O(n18047));
    defparam i13218_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i30838_2_lut (.I0(\data_out_frame[20] [3]), .I1(byte_transmit_counter[0]), 
            .I2(GND_net), .I3(GND_net), .O(n37270));
    defparam i30838_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i2_3_lut_adj_917 (.I0(\data_in_frame[20] [6]), .I1(n33238), 
            .I2(\data_in_frame[18] [5]), .I3(GND_net), .O(n34170));
    defparam i2_3_lut_adj_917.LUT_INIT = 16'h9696;
    SB_LUT4 i4_4_lut_adj_918 (.I0(\data_in_frame[7] [6]), .I1(n16233), .I2(\data_in_frame[8] [0]), 
            .I3(n6_adj_4351), .O(n30694));   // verilog/coms.v(84[17:28])
    defparam i4_4_lut_adj_918.LUT_INIT = 16'h6996;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_4_i6_4_lut (.I0(\data_out_frame[5] [4]), 
            .I1(byte_transmit_counter_c[1]), .I2(byte_transmit_counter_c[2]), 
            .I3(byte_transmit_counter[0]), .O(n6_adj_4367));   // verilog/coms.v(105[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_4_i6_4_lut.LUT_INIT = 16'hac03;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_4_i5_3_lut (.I0(\data_out_frame[6] [4]), 
            .I1(\data_out_frame[7] [4]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n5_adj_4368));   // verilog/coms.v(105[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_4_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_DFFSR tx_transmit_3429 (.Q(\r_SM_Main_2__N_3458[0] ), .C(clk32MHz), 
            .D(n3693[0]), .R(n33773));   // verilog/coms.v(126[12] 293[6])
    SB_LUT4 i19995_1_lut (.I0(n24810), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n2290));
    defparam i19995_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i13219_3_lut_4_lut (.I0(n8_adj_4353), .I1(n32959), .I2(rx_data[6]), 
            .I3(\data_in_frame[4] [6]), .O(n18048));
    defparam i13219_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_919 (.I0(n34514), .I1(\data_in_frame[16] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n31184));
    defparam i1_2_lut_adj_919.LUT_INIT = 16'h9999;
    SB_LUT4 i1_2_lut_adj_920 (.I0(\data_in_frame[8] [0]), .I1(\data_in_frame[12] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n33464));   // verilog/coms.v(84[17:28])
    defparam i1_2_lut_adj_920.LUT_INIT = 16'h6666;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_4_i7_3_lut (.I0(n5_adj_4368), 
            .I1(n6_adj_4367), .I2(n37177), .I3(GND_net), .O(n7_adj_4369));   // verilog/coms.v(105[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_4_i7_3_lut.LUT_INIT = 16'hacac;
    SB_DFF \FRAME_MATCHER.rx_data_ready_prev_3430  (.Q(\FRAME_MATCHER.rx_data_ready_prev ), 
           .C(clk32MHz), .D(rx_data_ready));   // verilog/coms.v(126[12] 293[6])
    SB_LUT4 i2034738_i1_3_lut (.I0(n38330), .I1(n38462), .I2(byte_transmit_counter_c[2]), 
            .I3(GND_net), .O(n14_adj_4370));
    defparam i2034738_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF data_in_frame_0__i98 (.Q(\data_in_frame[12] [1]), .C(clk32MHz), 
           .D(n18107));   // verilog/coms.v(126[12] 293[6])
    SB_LUT4 data_in_frame_7__7__I_0_2_lut (.I0(\data_in_frame[7] [7]), .I1(\data_in_frame[7] [6]), 
            .I2(GND_net), .I3(GND_net), .O(Kp_23__N_1183));   // verilog/coms.v(84[17:28])
    defparam data_in_frame_7__7__I_0_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i31492_3_lut (.I0(\FRAME_MATCHER.state [3]), .I1(n33773), .I2(n5069), 
            .I3(GND_net), .O(n34073));
    defparam i31492_3_lut.LUT_INIT = 16'h0101;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_5_i6_3_lut (.I0(\data_out_frame[5] [5]), 
            .I1(byte_transmit_counter_c[1]), .I2(byte_transmit_counter_c[2]), 
            .I3(GND_net), .O(n37536));   // verilog/coms.v(105[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_5_i6_3_lut.LUT_INIT = 16'ha3a3;
    SB_LUT4 i6_4_lut_adj_921 (.I0(n33464), .I1(\data_in_frame[6] [1]), .I2(\data_in_frame[10] [3]), 
            .I3(n16791), .O(n14_adj_4371));   // verilog/coms.v(84[17:28])
    defparam i6_4_lut_adj_921.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut_adj_922 (.I0(\data_in_frame[8] [2]), .I1(n14_adj_4371), 
            .I2(n10_adj_4372), .I3(n6_adj_4348), .O(n16314));   // verilog/coms.v(84[17:28])
    defparam i7_4_lut_adj_922.LUT_INIT = 16'h6996;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_5_i5_3_lut (.I0(\data_out_frame[6] [5]), 
            .I1(\data_out_frame[7] [5]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n5_adj_4373));   // verilog/coms.v(105[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_5_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3_3_lut_adj_923 (.I0(\data_in_frame[20] [2]), .I1(n33323), 
            .I2(n33583), .I3(GND_net), .O(n8_adj_4374));
    defparam i3_3_lut_adj_923.LUT_INIT = 16'h9696;
    SB_LUT4 i1_4_lut_adj_924 (.I0(\data_in_frame[5] [6]), .I1(\data_in_frame[1] [2]), 
            .I2(n33076), .I3(\data_in_frame[1] [4]), .O(n33127));   // verilog/coms.v(84[17:28])
    defparam i1_4_lut_adj_924.LUT_INIT = 16'h6996;
    SB_LUT4 i31541_4_lut (.I0(n33773), .I1(\FRAME_MATCHER.state [3]), .I2(n5034), 
            .I3(n5069), .O(n33781));
    defparam i31541_4_lut.LUT_INIT = 16'h5011;
    SB_LUT4 i7_4_lut_adj_925 (.I0(n13), .I1(n11), .I2(\data_in_frame[20] [7]), 
            .I3(n16930), .O(n34659));
    defparam i7_4_lut_adj_925.LUT_INIT = 16'h6996;
    SB_DFF data_in_frame_0__i123 (.Q(\data_in_frame[15] [2]), .C(clk32MHz), 
           .D(n18132));   // verilog/coms.v(126[12] 293[6])
    SB_LUT4 i4_4_lut_adj_926 (.I0(n34651), .I1(n33247), .I2(n33471), .I3(\data_in_frame[20] [3]), 
            .O(n12));
    defparam i4_4_lut_adj_926.LUT_INIT = 16'hd77d;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_5_i7_4_lut (.I0(n5_adj_4373), 
            .I1(byte_transmit_counter[0]), .I2(n37177), .I3(n37536), .O(n7_adj_4375));   // verilog/coms.v(105[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_5_i7_4_lut.LUT_INIT = 16'haca0;
    SB_DFF data_in_frame_0__i97 (.Q(\data_in_frame[12] [0]), .C(clk32MHz), 
           .D(n18106));   // verilog/coms.v(126[12] 293[6])
    SB_DFF data_in_frame_0__i10 (.Q(\data_in_frame[1] [1]), .C(clk32MHz), 
           .D(n18019));   // verilog/coms.v(126[12] 293[6])
    SB_LUT4 i2_3_lut_adj_927 (.I0(\data_in_frame[10] [5]), .I1(\data_in_frame[15] [1]), 
            .I2(\data_in_frame[14] [7]), .I3(GND_net), .O(n33385));   // verilog/coms.v(84[17:28])
    defparam i2_3_lut_adj_927.LUT_INIT = 16'h9696;
    SB_LUT4 i5_4_lut (.I0(n33350), .I1(n33526), .I2(\data_in_frame[5] [0]), 
            .I3(n33250), .O(n12_adj_4376));   // verilog/coms.v(75[16:27])
    defparam i5_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i31487_2_lut (.I0(\FRAME_MATCHER.state [1]), .I1(\FRAME_MATCHER.state [2]), 
            .I2(GND_net), .I3(GND_net), .O(n5034));   // verilog/coms.v(144[4] 292[11])
    defparam i31487_2_lut.LUT_INIT = 16'h1111;
    SB_DFF data_in_frame_0__i9 (.Q(\data_in_frame[1] [0]), .C(clk32MHz), 
           .D(n18018));   // verilog/coms.v(126[12] 293[6])
    SB_DFF data_in_frame_0__i8 (.Q(\data_in_frame[0] [7]), .C(clk32MHz), 
           .D(n18017));   // verilog/coms.v(126[12] 293[6])
    SB_DFF data_in_frame_0__i7 (.Q(\data_in_frame[0] [6]), .C(clk32MHz), 
           .D(n18016));   // verilog/coms.v(126[12] 293[6])
    SB_DFF data_in_frame_0__i6 (.Q(\data_in_frame[0] [5]), .C(clk32MHz), 
           .D(n18015));   // verilog/coms.v(126[12] 293[6])
    SB_DFF data_in_frame_0__i5 (.Q(\data_in_frame[0] [4]), .C(clk32MHz), 
           .D(n18014));   // verilog/coms.v(126[12] 293[6])
    SB_LUT4 i2035341_i1_3_lut (.I0(n38324), .I1(n38318), .I2(byte_transmit_counter_c[2]), 
            .I3(GND_net), .O(n14_adj_4377));
    defparam i2035341_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_0_i16_3_lut (.I0(\data_out_frame[16] [0]), 
            .I1(\data_out_frame[17] [0]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n16_adj_4378));   // verilog/coms.v(105[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_0_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_0_i17_3_lut (.I0(\data_out_frame[18] [0]), 
            .I1(\data_out_frame[19] [0]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n17_adj_4379));   // verilog/coms.v(105[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_0_i17_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i6_4_lut_adj_928 (.I0(\data_in_frame[1] [0]), .I1(n12_adj_4376), 
            .I2(n33604), .I3(n33104), .O(n31002));   // verilog/coms.v(75[16:27])
    defparam i6_4_lut_adj_928.LUT_INIT = 16'h6996;
    SB_LUT4 i30850_2_lut (.I0(byte_transmit_counter_c[2]), .I1(\data_out_frame[5] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n37531));   // verilog/coms.v(105[34:55])
    defparam i30850_2_lut.LUT_INIT = 16'hdddd;
    SB_LUT4 i1_2_lut_adj_929 (.I0(Kp_23__N_993), .I1(Kp_23__N_996), .I2(GND_net), 
            .I3(GND_net), .O(n17157));
    defparam i1_2_lut_adj_929.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_930 (.I0(n17157), .I1(\data_in_frame[4] [6]), .I2(n30217), 
            .I3(n33316), .O(n10_adj_4380));
    defparam i4_4_lut_adj_930.LUT_INIT = 16'h6996;
    SB_LUT4 i5_3_lut_adj_931 (.I0(n31002), .I1(n10_adj_4380), .I2(\data_in_frame[7] [2]), 
            .I3(GND_net), .O(n15795));
    defparam i5_3_lut_adj_931.LUT_INIT = 16'h9696;
    SB_LUT4 i2_4_lut (.I0(n33269), .I1(n35077), .I2(n33445), .I3(\data_in_frame[21] [2]), 
            .O(n10_adj_4381));
    defparam i2_4_lut.LUT_INIT = 16'hb77b;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_6_i5_3_lut (.I0(\data_out_frame[6] [6]), 
            .I1(\data_out_frame[7] [6]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n5_adj_4382));   // verilog/coms.v(105[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_6_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2_3_lut_adj_932 (.I0(Kp_23__N_1026), .I1(\data_in_frame[3] [0]), 
            .I2(\data_in_frame[0] [6]), .I3(GND_net), .O(n33250));
    defparam i2_3_lut_adj_932.LUT_INIT = 16'h9696;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_6_i7_4_lut (.I0(n5_adj_4382), 
            .I1(n37531), .I2(n37177), .I3(byte_transmit_counter[0]), .O(n7_adj_4383));   // verilog/coms.v(105[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_6_i7_4_lut.LUT_INIT = 16'haca0;
    SB_LUT4 i13220_3_lut_4_lut (.I0(n8_adj_4353), .I1(n32959), .I2(rx_data[7]), 
            .I3(\data_in_frame[4] [7]), .O(n18049));
    defparam i13220_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i3_4_lut_adj_933 (.I0(\data_in_frame[3] [2]), .I1(\data_in_frame[1] [0]), 
            .I2(\data_in_frame[0] [6]), .I3(\data_in_frame[1] [1]), .O(n32994));   // verilog/coms.v(77[16:27])
    defparam i3_4_lut_adj_933.LUT_INIT = 16'h6996;
    SB_LUT4 i13277_3_lut_4_lut (.I0(n8_adj_4353), .I1(n32937), .I2(rx_data[0]), 
            .I3(\data_in_frame[12] [0]), .O(n18106));
    defparam i13277_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2035944_i1_3_lut (.I0(n38372), .I1(n38288), .I2(byte_transmit_counter_c[2]), 
            .I3(GND_net), .O(n14_adj_4384));
    defparam i2035944_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2_3_lut_adj_934 (.I0(n16765), .I1(\data_in_frame[6] [1]), .I2(Kp_23__N_1046), 
            .I3(GND_net), .O(n33532));   // verilog/coms.v(71[16:41])
    defparam i2_3_lut_adj_934.LUT_INIT = 16'h9696;
    SB_LUT4 i13278_3_lut_4_lut (.I0(n8_adj_4353), .I1(n32937), .I2(rx_data[1]), 
            .I3(\data_in_frame[12] [1]), .O(n18107));
    defparam i13278_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i6_4_lut_adj_935 (.I0(\data_in_frame[6] [2]), .I1(\data_in_frame[17] [1]), 
            .I2(n33532), .I3(n33385), .O(n16_adj_4385));   // verilog/coms.v(84[17:28])
    defparam i6_4_lut_adj_935.LUT_INIT = 16'h6996;
    SB_DFF data_in_frame_0__i4 (.Q(\data_in_frame[0] [3]), .C(clk32MHz), 
           .D(n18013));   // verilog/coms.v(126[12] 293[6])
    SB_LUT4 i13279_3_lut_4_lut (.I0(n8_adj_4353), .I1(n32937), .I2(rx_data[2]), 
            .I3(\data_in_frame[12] [2]), .O(n18108));
    defparam i13279_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i30486_2_lut (.I0(byte_transmit_counter_c[2]), .I1(byte_transmit_counter_c[1]), 
            .I2(GND_net), .I3(GND_net), .O(n37177));   // verilog/coms.v(105[34:55])
    defparam i30486_2_lut.LUT_INIT = 16'h8888;
    SB_DFF data_in_frame_0__i3 (.Q(\data_in_frame[0] [2]), .C(clk32MHz), 
           .D(n18012));   // verilog/coms.v(126[12] 293[6])
    SB_DFF data_in_frame_0__i2 (.Q(\data_in_frame[0] [1]), .C(clk32MHz), 
           .D(n18011));   // verilog/coms.v(126[12] 293[6])
    SB_DFF data_in_frame_0__i116 (.Q(\data_in_frame[14] [3]), .C(clk32MHz), 
           .D(n18125));   // verilog/coms.v(126[12] 293[6])
    SB_LUT4 i3_4_lut_adj_936 (.I0(n33217), .I1(n34170), .I2(n10_adj_4354), 
            .I3(\data_in_frame[16] [2]), .O(n11_adj_4386));
    defparam i3_4_lut_adj_936.LUT_INIT = 16'hdeed;
    SB_LUT4 i7_4_lut_adj_937 (.I0(\data_in_frame[17] [2]), .I1(n33409), 
            .I2(n33607), .I3(n33036), .O(n17_adj_4387));   // verilog/coms.v(84[17:28])
    defparam i7_4_lut_adj_937.LUT_INIT = 16'h6996;
    SB_DFF data_in_frame_0__i96 (.Q(\data_in_frame[11] [7]), .C(clk32MHz), 
           .D(n18105));   // verilog/coms.v(126[12] 293[6])
    SB_LUT4 i2_3_lut_adj_938 (.I0(n32994), .I1(n33354), .I2(\data_in_frame[5] [4]), 
            .I3(GND_net), .O(n16791));
    defparam i2_3_lut_adj_938.LUT_INIT = 16'h9696;
    SB_LUT4 i9_4_lut_adj_939 (.I0(n17_adj_4387), .I1(\data_in_frame[16] [7]), 
            .I2(n16_adj_4385), .I3(\data_in_frame[14] [5]), .O(n15781));   // verilog/coms.v(84[17:28])
    defparam i9_4_lut_adj_939.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_940 (.I0(n16740), .I1(n34659), .I2(n8_adj_4374), 
            .I3(n33471), .O(n9_adj_4388));
    defparam i1_4_lut_adj_940.LUT_INIT = 16'hb77b;
    SB_LUT4 i13280_3_lut_4_lut (.I0(n8_adj_4353), .I1(n32937), .I2(rx_data[3]), 
            .I3(\data_in_frame[12] [3]), .O(n18109));
    defparam i13280_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF control_mode_i0_i7 (.Q(control_mode[7]), .C(clk32MHz), .D(n18010));   // verilog/coms.v(126[12] 293[6])
    SB_LUT4 i1_2_lut_adj_941 (.I0(\FRAME_MATCHER.state [28]), .I1(n12_adj_4389), 
            .I2(GND_net), .I3(GND_net), .O(n32271));
    defparam i1_2_lut_adj_941.LUT_INIT = 16'h8888;
    SB_LUT4 i31155_2_lut (.I0(byte_transmit_counter_c[2]), .I1(\data_out_frame[5] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n37837));   // verilog/coms.v(105[34:55])
    defparam i31155_2_lut.LUT_INIT = 16'hdddd;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_7_i5_3_lut (.I0(\data_out_frame[6] [7]), 
            .I1(\data_out_frame[7] [7]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n5_adj_4390));   // verilog/coms.v(105[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_7_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_7_i7_4_lut (.I0(n5_adj_4390), 
            .I1(n37837), .I2(n37177), .I3(byte_transmit_counter[0]), .O(n7_adj_4391));   // verilog/coms.v(105[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_7_i7_4_lut.LUT_INIT = 16'haca0;
    SB_DFF control_mode_i0_i6 (.Q(control_mode[6]), .C(clk32MHz), .D(n18009));   // verilog/coms.v(126[12] 293[6])
    SB_DFF control_mode_i0_i5 (.Q(control_mode[5]), .C(clk32MHz), .D(n18008));   // verilog/coms.v(126[12] 293[6])
    SB_DFF control_mode_i0_i4 (.Q(control_mode[4]), .C(clk32MHz), .D(n18007));   // verilog/coms.v(126[12] 293[6])
    SB_DFF control_mode_i0_i3 (.Q(control_mode[3]), .C(clk32MHz), .D(n18006));   // verilog/coms.v(126[12] 293[6])
    SB_DFF control_mode_i0_i2 (.Q(control_mode[2]), .C(clk32MHz), .D(n18005));   // verilog/coms.v(126[12] 293[6])
    SB_LUT4 i2036547_i1_3_lut (.I0(n38366), .I1(n38294), .I2(byte_transmit_counter_c[2]), 
            .I3(GND_net), .O(n14_adj_4392));
    defparam i2036547_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_adj_942 (.I0(\FRAME_MATCHER.state [26]), .I1(n12_adj_4389), 
            .I2(GND_net), .I3(GND_net), .O(n32219));
    defparam i1_2_lut_adj_942.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_943 (.I0(\FRAME_MATCHER.state [25]), .I1(n12_adj_4389), 
            .I2(GND_net), .I3(GND_net), .O(n32221));
    defparam i1_2_lut_adj_943.LUT_INIT = 16'h8888;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_0_i6_4_lut (.I0(\data_out_frame[5] [0]), 
            .I1(byte_transmit_counter[0]), .I2(byte_transmit_counter_c[2]), 
            .I3(byte_transmit_counter_c[1]), .O(n6_adj_4393));   // verilog/coms.v(105[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_0_i6_4_lut.LUT_INIT = 16'hb0bc;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_0_i5_3_lut (.I0(\data_out_frame[6] [0]), 
            .I1(\data_out_frame[7] [0]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n5_adj_4394));   // verilog/coms.v(105[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_0_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_0_i7_4_lut (.I0(n5_adj_4394), 
            .I1(n6_adj_4393), .I2(byte_transmit_counter_c[2]), .I3(byte_transmit_counter_c[1]), 
            .O(n7_adj_4395));   // verilog/coms.v(105[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_0_i7_4_lut.LUT_INIT = 16'haccc;
    SB_LUT4 i13281_3_lut_4_lut (.I0(n8_adj_4353), .I1(n32937), .I2(rx_data[4]), 
            .I3(\data_in_frame[12] [4]), .O(n18110));
    defparam i13281_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_944 (.I0(\FRAME_MATCHER.state [24]), .I1(n12_adj_4389), 
            .I2(GND_net), .I3(GND_net), .O(n32223));
    defparam i1_2_lut_adj_944.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_945 (.I0(n16608), .I1(\data_in_frame[7] [5]), .I2(GND_net), 
            .I3(GND_net), .O(n33155));
    defparam i1_2_lut_adj_945.LUT_INIT = 16'h6666;
    SB_LUT4 i2037753_i1_3_lut (.I0(n38354), .I1(n38312), .I2(byte_transmit_counter_c[2]), 
            .I3(GND_net), .O(n14_adj_4396));
    defparam i2037753_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3_4_lut_adj_946 (.I0(\data_in_frame[16] [4]), .I1(n33335), 
            .I2(n31184), .I3(\data_in_frame[19] [0]), .O(n31196));
    defparam i3_4_lut_adj_946.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_947 (.I0(\FRAME_MATCHER.state [22]), .I1(n12_adj_4389), 
            .I2(GND_net), .I3(GND_net), .O(n32225));
    defparam i1_2_lut_adj_947.LUT_INIT = 16'h8888;
    SB_DFF data_in_frame_0__i122 (.Q(\data_in_frame[15] [1]), .C(clk32MHz), 
           .D(n18131));   // verilog/coms.v(126[12] 293[6])
    SB_LUT4 i1_2_lut_adj_948 (.I0(\FRAME_MATCHER.state [21]), .I1(n12_adj_4389), 
            .I2(GND_net), .I3(GND_net), .O(n32227));
    defparam i1_2_lut_adj_948.LUT_INIT = 16'h8888;
    SB_DFF control_mode_i0_i1 (.Q(control_mode[1]), .C(clk32MHz), .D(n18004));   // verilog/coms.v(126[12] 293[6])
    SB_LUT4 i1_2_lut_adj_949 (.I0(\FRAME_MATCHER.state [19]), .I1(n12_adj_4389), 
            .I2(GND_net), .I3(GND_net), .O(n32161));   // verilog/coms.v(114[11:12])
    defparam i1_2_lut_adj_949.LUT_INIT = 16'h8888;
    SB_DFF data_out_frame_0___i191 (.Q(\data_out_frame[23][6] ), .C(clk32MHz), 
           .D(n18003));   // verilog/coms.v(126[12] 293[6])
    SB_DFF data_out_frame_0___i168 (.Q(\data_out_frame[20] [7]), .C(clk32MHz), 
           .D(n18002));   // verilog/coms.v(126[12] 293[6])
    SB_DFF data_out_frame_0___i167 (.Q(\data_out_frame[20] [6]), .C(clk32MHz), 
           .D(n18001));   // verilog/coms.v(126[12] 293[6])
    SB_DFF data_out_frame_0___i166 (.Q(\data_out_frame[20] [5]), .C(clk32MHz), 
           .D(n18000));   // verilog/coms.v(126[12] 293[6])
    SB_DFF data_out_frame_0___i165 (.Q(\data_out_frame[20] [4]), .C(clk32MHz), 
           .D(n17999));   // verilog/coms.v(126[12] 293[6])
    SB_LUT4 i4_4_lut_adj_950 (.I0(n33310), .I1(n16413), .I2(n31184), .I3(n33474), 
            .O(n10_adj_4397));
    defparam i4_4_lut_adj_950.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_adj_951 (.I0(\FRAME_MATCHER.state [18]), .I1(n12_adj_4389), 
            .I2(GND_net), .I3(GND_net), .O(n32181));
    defparam i1_2_lut_adj_951.LUT_INIT = 16'h8888;
    SB_LUT4 i2_3_lut_4_lut (.I0(\data_in_frame[6] [2]), .I1(n6_adj_4348), 
            .I2(n33010), .I3(\data_in_frame[8] [7]), .O(n16447));   // verilog/coms.v(84[17:28])
    defparam i2_3_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i13233_3_lut_4_lut (.I0(n8_adj_4355), .I1(n32959), .I2(rx_data[4]), 
            .I3(\data_in_frame[6] [4]), .O(n18062));
    defparam i13233_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 add_41_2_lut (.I0(n2290), .I1(\FRAME_MATCHER.i [0]), .I2(n161), 
            .I3(GND_net), .O(n2)) /* synthesis syn_instantiated=1 */ ;
    defparam add_41_2_lut.LUT_INIT = 16'h8228;
    SB_DFF data_out_frame_0___i164 (.Q(\data_out_frame[20] [3]), .C(clk32MHz), 
           .D(n17998));   // verilog/coms.v(126[12] 293[6])
    SB_LUT4 i1_2_lut_adj_952 (.I0(\FRAME_MATCHER.state [16]), .I1(n12_adj_4389), 
            .I2(GND_net), .I3(GND_net), .O(n32229));
    defparam i1_2_lut_adj_952.LUT_INIT = 16'h8888;
    SB_DFF data_out_frame_0___i163 (.Q(\data_out_frame[20] [2]), .C(clk32MHz), 
           .D(n17997));   // verilog/coms.v(126[12] 293[6])
    SB_LUT4 i1_2_lut_adj_953 (.I0(\FRAME_MATCHER.state [15]), .I1(n12_adj_4389), 
            .I2(GND_net), .I3(GND_net), .O(n32231));
    defparam i1_2_lut_adj_953.LUT_INIT = 16'h8888;
    SB_DFF data_out_frame_0___i162 (.Q(\data_out_frame[20] [1]), .C(clk32MHz), 
           .D(n17996));   // verilog/coms.v(126[12] 293[6])
    SB_LUT4 i1_2_lut_adj_954 (.I0(\FRAME_MATCHER.state [14]), .I1(n12_adj_4389), 
            .I2(GND_net), .I3(GND_net), .O(n32233));
    defparam i1_2_lut_adj_954.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_955 (.I0(\FRAME_MATCHER.state [13]), .I1(n12_adj_4389), 
            .I2(GND_net), .I3(GND_net), .O(n32235));
    defparam i1_2_lut_adj_955.LUT_INIT = 16'h8888;
    SB_LUT4 i5_3_lut_4_lut (.I0(\data_in_frame[6] [2]), .I1(n6_adj_4348), 
            .I2(n10_adj_4398), .I3(n33142), .O(n33357));   // verilog/coms.v(84[17:28])
    defparam i5_3_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_956 (.I0(\FRAME_MATCHER.state [12]), .I1(n12_adj_4389), 
            .I2(GND_net), .I3(GND_net), .O(n32149));
    defparam i1_2_lut_adj_956.LUT_INIT = 16'h8888;
    SB_CARRY add_41_2 (.CI(GND_net), .I0(\FRAME_MATCHER.i [0]), .I1(n161), 
            .CO(n27909));
    SB_LUT4 i1_2_lut_adj_957 (.I0(\FRAME_MATCHER.state [11]), .I1(n12_adj_4389), 
            .I2(GND_net), .I3(GND_net), .O(n32237));
    defparam i1_2_lut_adj_957.LUT_INIT = 16'h8888;
    SB_LUT4 i2_3_lut_4_lut_adj_958 (.I0(\data_in_frame[6] [2]), .I1(n6_adj_4348), 
            .I2(n16765), .I3(\data_in_frame[8] [2]), .O(n33397));   // verilog/coms.v(84[17:28])
    defparam i2_3_lut_4_lut_adj_958.LUT_INIT = 16'h6996;
    SB_DFF data_out_frame_0___i161 (.Q(\data_out_frame[20] [0]), .C(clk32MHz), 
           .D(n17995));   // verilog/coms.v(126[12] 293[6])
    SB_DFF data_out_frame_0___i160 (.Q(\data_out_frame[19] [7]), .C(clk32MHz), 
           .D(n17994));   // verilog/coms.v(126[12] 293[6])
    SB_DFF data_out_frame_0___i159 (.Q(\data_out_frame[19] [6]), .C(clk32MHz), 
           .D(n17993));   // verilog/coms.v(126[12] 293[6])
    SB_LUT4 i17819_3_lut (.I0(\data_in[2] [1]), .I1(\data_in[3] [1]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n17807));   // verilog/coms.v(89[7:20])
    defparam i17819_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF data_out_frame_0___i158 (.Q(\data_out_frame[19] [5]), .C(clk32MHz), 
           .D(n17992));   // verilog/coms.v(126[12] 293[6])
    SB_DFF data_out_frame_0___i157 (.Q(\data_out_frame[19] [4]), .C(clk32MHz), 
           .D(n17991));   // verilog/coms.v(126[12] 293[6])
    SB_DFF data_out_frame_0___i156 (.Q(\data_out_frame[19] [3]), .C(clk32MHz), 
           .D(n17990));   // verilog/coms.v(126[12] 293[6])
    SB_LUT4 i13282_3_lut_4_lut (.I0(n8_adj_4353), .I1(n32937), .I2(rx_data[5]), 
            .I3(\data_in_frame[12] [5]), .O(n18111));
    defparam i13282_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_959 (.I0(\FRAME_MATCHER.state [6]), .I1(n12_adj_4389), 
            .I2(GND_net), .I3(GND_net), .O(n32239));
    defparam i1_2_lut_adj_959.LUT_INIT = 16'h8888;
    SB_LUT4 i13283_3_lut_4_lut (.I0(n8_adj_4353), .I1(n32937), .I2(rx_data[6]), 
            .I3(\data_in_frame[12] [6]), .O(n18112));
    defparam i13283_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i5_3_lut_adj_960 (.I0(n16466), .I1(n10_adj_4397), .I2(\data_in_frame[12] [6]), 
            .I3(GND_net), .O(n31228));
    defparam i5_3_lut_adj_960.LUT_INIT = 16'h9696;
    SB_LUT4 i13284_3_lut_4_lut (.I0(n8_adj_4353), .I1(n32937), .I2(rx_data[7]), 
            .I3(\data_in_frame[12] [7]), .O(n18113));
    defparam i13284_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i17822_3_lut (.I0(\data_in[2] [3]), .I1(\data_in[3] [3]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n17809));   // verilog/coms.v(89[7:20])
    defparam i17822_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i29726_2_lut (.I0(\data_in_frame[2] [5]), .I1(\data_in_frame[2] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n36323));
    defparam i29726_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i13_4_lut_adj_961 (.I0(n36323), .I1(\data_in_frame[2] [7]), 
            .I2(\data_in_frame[2] [0]), .I3(\data_in_frame[1] [7]), .O(n30));
    defparam i13_4_lut_adj_961.LUT_INIT = 16'h0010;
    SB_LUT4 i17818_3_lut (.I0(\data_in[2] [5]), .I1(\data_in[3] [5]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n17811));   // verilog/coms.v(89[7:20])
    defparam i17818_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11_4_lut_adj_962 (.I0(n32855), .I1(\data_in_frame[2] [4]), 
            .I2(\data_in_frame[1] [4]), .I3(\data_in_frame[1] [6]), .O(n28_adj_4399));
    defparam i11_4_lut_adj_962.LUT_INIT = 16'h8000;
    SB_LUT4 i12_4_lut_adj_963 (.I0(\data_in_frame[1] [5]), .I1(\data_in_frame[1] [1]), 
            .I2(\data_in_frame[2] [2]), .I3(\data_in_frame[2] [6]), .O(n29));
    defparam i12_4_lut_adj_963.LUT_INIT = 16'h0002;
    SB_LUT4 i10_4_lut_adj_964 (.I0(\data_in_frame[1] [2]), .I1(\data_in_frame[2] [1]), 
            .I2(\data_in_frame[1] [0]), .I3(\data_in_frame[1] [3]), .O(n27_adj_4400));
    defparam i10_4_lut_adj_964.LUT_INIT = 16'h8000;
    SB_LUT4 i16_4_lut_adj_965 (.I0(n27_adj_4400), .I1(n29), .I2(n28_adj_4399), 
            .I3(n30), .O(\FRAME_MATCHER.state_31__N_2630 [3]));
    defparam i16_4_lut_adj_965.LUT_INIT = 16'h8000;
    SB_DFF data_in_frame_0__i121 (.Q(\data_in_frame[15] [0]), .C(clk32MHz), 
           .D(n18130));   // verilog/coms.v(126[12] 293[6])
    SB_LUT4 i1_2_lut_3_lut (.I0(\data_in_frame[1] [4]), .I1(\data_in_frame[1] [6]), 
            .I2(\data_in_frame[1] [0]), .I3(GND_net), .O(n33403));   // verilog/coms.v(84[17:28])
    defparam i1_2_lut_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 i3_4_lut_adj_966 (.I0(n33789), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.state [1]), .I3(\FRAME_MATCHER.state_31__N_2630 [3]), 
            .O(n13724));   // verilog/coms.v(126[12] 293[6])
    defparam i3_4_lut_adj_966.LUT_INIT = 16'h1000;
    SB_DFF data_out_frame_0___i155 (.Q(\data_out_frame[19] [2]), .C(clk32MHz), 
           .D(n17989));   // verilog/coms.v(126[12] 293[6])
    SB_LUT4 i1_2_lut_adj_967 (.I0(\data_out_frame[9] [7]), .I1(\data_out_frame[7] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n16951));
    defparam i1_2_lut_adj_967.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_3_lut_4_lut (.I0(\data_in_frame[1] [4]), .I1(\data_in_frame[1] [6]), 
            .I2(\data_in_frame[4] [0]), .I3(n16299), .O(n6_adj_4348));   // verilog/coms.v(84[17:28])
    defparam i1_2_lut_3_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_968 (.I0(n1_c), .I1(n16158), .I2(n4_adj_4401), 
            .I3(n7_adj_4402), .O(n12_adj_4389));
    defparam i1_4_lut_adj_968.LUT_INIT = 16'hbbba;
    SB_LUT4 i2_3_lut_4_lut_adj_969 (.I0(\data_in_frame[1] [4]), .I1(\data_in_frame[1] [6]), 
            .I2(\data_in_frame[0] [7]), .I3(n33406), .O(Kp_23__N_1026));   // verilog/coms.v(84[17:28])
    defparam i2_3_lut_4_lut_adj_969.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_970 (.I0(\data_out_frame[5] [2]), .I1(\data_out_frame[7] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n33306));   // verilog/coms.v(75[16:43])
    defparam i1_2_lut_adj_970.LUT_INIT = 16'h6666;
    SB_LUT4 i29815_3_lut_4_lut (.I0(n16161), .I1(n16154), .I2(n3893), 
            .I3(n3007), .O(n36418));
    defparam i29815_3_lut_4_lut.LUT_INIT = 16'hfca8;
    SB_LUT4 i3_4_lut_adj_971 (.I0(\data_out_frame[10] [1]), .I1(n33306), 
            .I2(\data_out_frame[10] [0]), .I3(\data_out_frame[12] [2]), 
            .O(n33494));
    defparam i3_4_lut_adj_971.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_972 (.I0(\FRAME_MATCHER.state [5]), .I1(n12_adj_4389), 
            .I2(GND_net), .I3(GND_net), .O(n32241));
    defparam i1_2_lut_adj_972.LUT_INIT = 16'h8888;
    SB_LUT4 i17821_3_lut (.I0(\data_in[3] [1]), .I1(rx_data[1]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n17815));   // verilog/coms.v(89[7:20])
    defparam i17821_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_adj_973 (.I0(\data_out_frame[14] [7]), .I1(\data_out_frame[17] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n33178));   // verilog/coms.v(70[16:27])
    defparam i1_2_lut_adj_973.LUT_INIT = 16'h6666;
    SB_LUT4 i17817_3_lut (.I0(\data_in[3] [3]), .I1(rx_data[3]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n17817));   // verilog/coms.v(89[7:20])
    defparam i17817_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_adj_974 (.I0(n1_c), .I1(n136), .I2(GND_net), .I3(GND_net), 
            .O(n4_adj_4403));
    defparam i1_2_lut_adj_974.LUT_INIT = 16'heeee;
    SB_LUT4 i13205_3_lut_4_lut (.I0(n8_adj_4404), .I1(n32959), .I2(rx_data[0]), 
            .I3(\data_in_frame[3] [0]), .O(n18034));
    defparam i13205_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF data_out_frame_0___i154 (.Q(\data_out_frame[19] [1]), .C(clk32MHz), 
           .D(n17988));   // verilog/coms.v(126[12] 293[6])
    SB_DFF data_out_frame_0___i153 (.Q(\data_out_frame[19] [0]), .C(clk32MHz), 
           .D(n17987));   // verilog/coms.v(126[12] 293[6])
    SB_DFF data_out_frame_0___i152 (.Q(\data_out_frame[18] [7]), .C(clk32MHz), 
           .D(n17986));   // verilog/coms.v(126[12] 293[6])
    SB_LUT4 i17823_3_lut (.I0(\data_in[3] [5]), .I1(rx_data[5]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n17819));   // verilog/coms.v(89[7:20])
    defparam i17823_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF data_out_frame_0___i151 (.Q(\data_out_frame[18] [6]), .C(clk32MHz), 
           .D(n17985));   // verilog/coms.v(126[12] 293[6])
    SB_LUT4 i5_3_lut_4_lut_adj_975 (.I0(n1251), .I1(\data_out_frame[9] [3]), 
            .I2(\data_out_frame[13] [7]), .I3(n10_adj_4405), .O(n34982));
    defparam i5_3_lut_4_lut_adj_975.LUT_INIT = 16'h6996;
    SB_DFF data_out_frame_0___i150 (.Q(\data_out_frame[18] [5]), .C(clk32MHz), 
           .D(n17984));   // verilog/coms.v(126[12] 293[6])
    SB_DFF data_out_frame_0___i149 (.Q(\data_out_frame[18] [4]), .C(clk32MHz), 
           .D(n17983));   // verilog/coms.v(126[12] 293[6])
    SB_DFF data_in_frame_0__i120 (.Q(\data_in_frame[14] [7]), .C(clk32MHz), 
           .D(n18129));   // verilog/coms.v(126[12] 293[6])
    SB_LUT4 i2_3_lut_4_lut_adj_976 (.I0(n1251), .I1(\data_out_frame[9] [3]), 
            .I2(\data_out_frame[9] [2]), .I3(n15783), .O(n30241));
    defparam i2_3_lut_4_lut_adj_976.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_977 (.I0(\data_in_frame[8] [6]), .I1(\data_in_frame[9] [0]), 
            .I2(n33388), .I3(GND_net), .O(n6_adj_4406));   // verilog/coms.v(73[16:43])
    defparam i1_2_lut_3_lut_adj_977.LUT_INIT = 16'h9696;
    SB_LUT4 i13206_3_lut_4_lut (.I0(n8_adj_4404), .I1(n32959), .I2(rx_data[1]), 
            .I3(\data_in_frame[3] [1]), .O(n18035));
    defparam i13206_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF data_out_frame_0___i148 (.Q(\data_out_frame[18] [3]), .C(clk32MHz), 
           .D(n17982));   // verilog/coms.v(126[12] 293[6])
    SB_LUT4 i1_2_lut_3_lut_adj_978 (.I0(\data_in_frame[8] [6]), .I1(\data_in_frame[9] [0]), 
            .I2(n33054), .I3(GND_net), .O(n6_adj_4407));   // verilog/coms.v(73[16:43])
    defparam i1_2_lut_3_lut_adj_978.LUT_INIT = 16'h9696;
    SB_DFF data_in_frame_0__i119 (.Q(\data_in_frame[14] [6]), .C(clk32MHz), 
           .D(n18128));   // verilog/coms.v(126[12] 293[6])
    SB_DFF data_out_frame_0___i147 (.Q(\data_out_frame[18] [2]), .C(clk32MHz), 
           .D(n17981));   // verilog/coms.v(126[12] 293[6])
    SB_LUT4 i1_2_lut_adj_979 (.I0(\data_out_frame[14] [5]), .I1(\data_out_frame[12] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n33292));   // verilog/coms.v(84[17:28])
    defparam i1_2_lut_adj_979.LUT_INIT = 16'h6666;
    SB_LUT4 i13207_3_lut_4_lut (.I0(n8_adj_4404), .I1(n32959), .I2(rx_data[2]), 
            .I3(\data_in_frame[3] [2]), .O(n18036));
    defparam i13207_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i3_3_lut_4_lut (.I0(\data_in_frame[4] [7]), .I1(\data_in_frame[4] [6]), 
            .I2(\data_in_frame[7] [2]), .I3(n17126), .O(n8_adj_4408));
    defparam i3_3_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_980 (.I0(\data_in_frame[4] [7]), .I1(\data_in_frame[4] [6]), 
            .I2(n31002), .I3(GND_net), .O(n33503));
    defparam i1_2_lut_3_lut_adj_980.LUT_INIT = 16'h9696;
    SB_LUT4 i7_4_lut_adj_981 (.I0(n9_adj_4388), .I1(n11_adj_4386), .I2(n10_adj_4381), 
            .I3(n12), .O(n35487));
    defparam i7_4_lut_adj_981.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_4_lut (.I0(\data_in_frame[9] [2]), .I1(n17169), .I2(\data_in_frame[7] [0]), 
            .I3(n33003), .O(n33529));
    defparam i1_2_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_adj_982 (.I0(\data_in_frame[9] [2]), .I1(n17169), 
            .I2(\data_in_frame[7] [0]), .I3(n31002), .O(n6_adj_4409));
    defparam i1_2_lut_4_lut_adj_982.LUT_INIT = 16'h6996;
    SB_DFF data_out_frame_0___i146 (.Q(\data_out_frame[18] [1]), .C(clk32MHz), 
           .D(n17980));   // verilog/coms.v(126[12] 293[6])
    SB_DFF data_out_frame_0___i145 (.Q(\data_out_frame[18] [0]), .C(clk32MHz), 
           .D(n17979));   // verilog/coms.v(126[12] 293[6])
    SB_LUT4 i1_2_lut_3_lut_adj_983 (.I0(\data_out_frame[12] [1]), .I1(n33063), 
            .I2(\data_out_frame[11] [7]), .I3(GND_net), .O(n33616));   // verilog/coms.v(84[17:63])
    defparam i1_2_lut_3_lut_adj_983.LUT_INIT = 16'h9696;
    SB_DFF data_out_frame_0___i144 (.Q(\data_out_frame[17] [7]), .C(clk32MHz), 
           .D(n17978));   // verilog/coms.v(126[12] 293[6])
    SB_DFF data_out_frame_0___i143 (.Q(\data_out_frame[17] [6]), .C(clk32MHz), 
           .D(n17977));   // verilog/coms.v(126[12] 293[6])
    SB_LUT4 i2_3_lut_4_lut_adj_984 (.I0(\data_out_frame[12] [1]), .I1(n33063), 
            .I2(\data_out_frame[14] [2]), .I3(n33066), .O(n33552));   // verilog/coms.v(84[17:63])
    defparam i2_3_lut_4_lut_adj_984.LUT_INIT = 16'h6996;
    SB_DFF data_out_frame_0___i142 (.Q(\data_out_frame[17] [5]), .C(clk32MHz), 
           .D(n17976));   // verilog/coms.v(126[12] 293[6])
    SB_DFF data_out_frame_0___i141 (.Q(\data_out_frame[17] [4]), .C(clk32MHz), 
           .D(n17975));   // verilog/coms.v(126[12] 293[6])
    SB_LUT4 i13234_3_lut_4_lut (.I0(n8_adj_4355), .I1(n32959), .I2(rx_data[5]), 
            .I3(\data_in_frame[6] [5]), .O(n18063));
    defparam i13234_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF data_out_frame_0___i140 (.Q(\data_out_frame[17] [3]), .C(clk32MHz), 
           .D(n17974));   // verilog/coms.v(126[12] 293[6])
    SB_DFF data_out_frame_0___i139 (.Q(\data_out_frame[17] [2]), .C(clk32MHz), 
           .D(n17973));   // verilog/coms.v(126[12] 293[6])
    SB_LUT4 i2_3_lut_4_lut_adj_985 (.I0(\data_in_frame[0] [0]), .I1(n32989), 
            .I2(\data_in_frame[2] [3]), .I3(Kp_23__N_993), .O(n33604));   // verilog/coms.v(165[9:87])
    defparam i2_3_lut_4_lut_adj_985.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_986 (.I0(\data_in_frame[0] [0]), .I1(n32989), 
            .I2(n4_adj_4410), .I3(\data_in_frame[4] [4]), .O(n16384));   // verilog/coms.v(165[9:87])
    defparam i2_3_lut_4_lut_adj_986.LUT_INIT = 16'h6996;
    SB_LUT4 i13237_3_lut_4_lut (.I0(n24185), .I1(n32959), .I2(rx_data[0]), 
            .I3(\data_in_frame[7] [0]), .O(n18066));
    defparam i13237_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i13238_3_lut_4_lut (.I0(n24185), .I1(n32959), .I2(rx_data[1]), 
            .I3(\data_in_frame[7] [1]), .O(n18067));
    defparam i13238_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF data_out_frame_0___i138 (.Q(\data_out_frame[17] [1]), .C(clk32MHz), 
           .D(n17972));   // verilog/coms.v(126[12] 293[6])
    SB_LUT4 i13239_3_lut_4_lut (.I0(n24185), .I1(n32959), .I2(rx_data[2]), 
            .I3(\data_in_frame[7] [2]), .O(n18068));
    defparam i13239_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF data_out_frame_0___i137 (.Q(\data_out_frame[17] [0]), .C(clk32MHz), 
           .D(n17971));   // verilog/coms.v(126[12] 293[6])
    SB_LUT4 i13240_3_lut_4_lut (.I0(n24185), .I1(n32959), .I2(rx_data[3]), 
            .I3(\data_in_frame[7] [3]), .O(n18069));
    defparam i13240_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i13241_3_lut_4_lut (.I0(n24185), .I1(n32959), .I2(rx_data[4]), 
            .I3(\data_in_frame[7] [4]), .O(n18070));
    defparam i13241_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1_2_lut_adj_987 (.I0(\data_in[0][6] ), .I1(n22566), .I2(GND_net), 
            .I3(GND_net), .O(n42_adj_4411));   // verilog/coms.v(94[12:19])
    defparam i1_2_lut_adj_987.LUT_INIT = 16'h2222;
    SB_DFF data_out_frame_0___i136 (.Q(\data_out_frame[16] [7]), .C(clk32MHz), 
           .D(n17970));   // verilog/coms.v(126[12] 293[6])
    SB_LUT4 i13242_3_lut_4_lut (.I0(n24185), .I1(n32959), .I2(rx_data[5]), 
            .I3(\data_in_frame[7] [5]), .O(n18071));
    defparam i13242_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF data_out_frame_0___i135 (.Q(\data_out_frame[16] [6]), .C(clk32MHz), 
           .D(n17969));   // verilog/coms.v(126[12] 293[6])
    SB_LUT4 i13243_3_lut_4_lut (.I0(n24185), .I1(n32959), .I2(rx_data[6]), 
            .I3(\data_in_frame[7] [6]), .O(n18072));
    defparam i13243_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i13244_3_lut_4_lut (.I0(n24185), .I1(n32959), .I2(rx_data[7]), 
            .I3(\data_in_frame[7] [7]), .O(n18073));
    defparam i13244_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF data_out_frame_0___i134 (.Q(\data_out_frame[16] [5]), .C(clk32MHz), 
           .D(n17968));   // verilog/coms.v(126[12] 293[6])
    SB_LUT4 i1_2_lut_3_lut_adj_988 (.I0(\data_out_frame[17] [5]), .I1(n30769), 
            .I2(n16661), .I3(GND_net), .O(n31295));
    defparam i1_2_lut_3_lut_adj_988.LUT_INIT = 16'h9696;
    SB_LUT4 i3_4_lut_adj_989 (.I0(\data_out_frame[10] [5]), .I1(n4_adj_4412), 
            .I2(n33013), .I3(\data_out_frame[6] [1]), .O(n16304));
    defparam i3_4_lut_adj_989.LUT_INIT = 16'h6996;
    SB_DFF data_out_frame_0___i133 (.Q(\data_out_frame[16] [4]), .C(clk32MHz), 
           .D(n17967));   // verilog/coms.v(126[12] 293[6])
    SB_DFF data_out_frame_0___i132 (.Q(\data_out_frame[16] [3]), .C(clk32MHz), 
           .D(n17966));   // verilog/coms.v(126[12] 293[6])
    SB_DFF data_out_frame_0___i131 (.Q(\data_out_frame[16] [2]), .C(clk32MHz), 
           .D(n17965));   // verilog/coms.v(126[12] 293[6])
    SB_LUT4 i4_4_lut_adj_990 (.I0(n33589), .I1(n33377), .I2(n1270), .I3(n33622), 
            .O(n10_adj_4413));
    defparam i4_4_lut_adj_990.LUT_INIT = 16'h6996;
    SB_DFF data_out_frame_0___i130 (.Q(\data_out_frame[16] [1]), .C(clk32MHz), 
           .D(n17964));   // verilog/coms.v(126[12] 293[6])
    SB_LUT4 i13208_3_lut_4_lut (.I0(n8_adj_4404), .I1(n32959), .I2(rx_data[3]), 
            .I3(\data_in_frame[3] [3]), .O(n18037));
    defparam i13208_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i5_3_lut_adj_991 (.I0(n33488), .I1(n10_adj_4413), .I2(\data_out_frame[10] [1]), 
            .I3(GND_net), .O(n31265));
    defparam i5_3_lut_adj_991.LUT_INIT = 16'h9696;
    SB_LUT4 i6_4_lut_adj_992 (.I0(\data_out_frame[5] [6]), .I1(n33292), 
            .I2(n33540), .I3(\data_out_frame[10] [1]), .O(n14_adj_4414));   // verilog/coms.v(84[17:28])
    defparam i6_4_lut_adj_992.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut_adj_993 (.I0(n33178), .I1(n14_adj_4414), .I2(n10_adj_4415), 
            .I3(n33546), .O(n33439));   // verilog/coms.v(84[17:28])
    defparam i7_4_lut_adj_993.LUT_INIT = 16'h6996;
    SB_DFF data_out_frame_0___i129 (.Q(\data_out_frame[16] [0]), .C(clk32MHz), 
           .D(n17963));   // verilog/coms.v(126[12] 293[6])
    SB_LUT4 i2_3_lut_4_lut_adj_994 (.I0(\data_out_frame[17] [5]), .I1(n30769), 
            .I2(n16975), .I3(\data_out_frame[20] [1]), .O(n33514));
    defparam i2_3_lut_4_lut_adj_994.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_995 (.I0(\data_out_frame[9] [6]), .I1(n33494), 
            .I2(n33145), .I3(\data_out_frame[7] [5]), .O(n16746));
    defparam i3_4_lut_adj_995.LUT_INIT = 16'h6996;
    SB_LUT4 i514_2_lut (.I0(\data_out_frame[7] [7]), .I1(\data_out_frame[7] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n1270));   // verilog/coms.v(84[17:28])
    defparam i514_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i13340_3_lut_4_lut (.I0(n8_adj_4404), .I1(n32952), .I2(rx_data[7]), 
            .I3(\data_in_frame[19] [7]), .O(n18169));
    defparam i13340_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_3_lut_adj_996 (.I0(\data_out_frame[10] [2]), .I1(\data_out_frame[8] [1]), 
            .I2(\data_out_frame[5] [4]), .I3(GND_net), .O(n33488));
    defparam i2_3_lut_adj_996.LUT_INIT = 16'h9696;
    SB_DFF data_out_frame_0___i128 (.Q(\data_out_frame[15] [7]), .C(clk32MHz), 
           .D(n17962));   // verilog/coms.v(126[12] 293[6])
    SB_DFF data_out_frame_0___i127 (.Q(\data_out_frame[15] [6]), .C(clk32MHz), 
           .D(n17961));   // verilog/coms.v(126[12] 293[6])
    SB_DFF data_out_frame_0___i126 (.Q(\data_out_frame[15] [5]), .C(clk32MHz), 
           .D(n17960));   // verilog/coms.v(126[12] 293[6])
    SB_DFF data_out_frame_0___i125 (.Q(\data_out_frame[15] [4]), .C(clk32MHz), 
           .D(n17959));   // verilog/coms.v(126[12] 293[6])
    SB_DFF data_out_frame_0___i124 (.Q(\data_out_frame[15] [3]), .C(clk32MHz), 
           .D(n17958));   // verilog/coms.v(126[12] 293[6])
    SB_DFF data_out_frame_0___i123 (.Q(\data_out_frame[15] [2]), .C(clk32MHz), 
           .D(n17957));   // verilog/coms.v(126[12] 293[6])
    SB_DFF data_out_frame_0___i122 (.Q(\data_out_frame[15] [1]), .C(clk32MHz), 
           .D(n17956));   // verilog/coms.v(126[12] 293[6])
    SB_LUT4 i2_3_lut_adj_997 (.I0(\FRAME_MATCHER.state [3]), .I1(n25118), 
            .I2(\FRAME_MATCHER.state [1]), .I3(GND_net), .O(n16153));   // verilog/coms.v(247[5:25])
    defparam i2_3_lut_adj_997.LUT_INIT = 16'hefef;
    SB_LUT4 i13333_3_lut_4_lut (.I0(n8_adj_4404), .I1(n32952), .I2(rx_data[0]), 
            .I3(\data_in_frame[19] [0]), .O(n18162));
    defparam i13333_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_3_lut_adj_998 (.I0(byte_transmit_counter_c[5]), .I1(byte_transmit_counter_c[7]), 
            .I2(byte_transmit_counter_c[6]), .I3(GND_net), .O(n16000));   // verilog/coms.v(210[11:56])
    defparam i2_3_lut_adj_998.LUT_INIT = 16'hfefe;
    SB_LUT4 i5_3_lut_4_lut_adj_999 (.I0(n33303), .I1(n10_adj_4416), .I2(\data_out_frame[18] [0]), 
            .I3(\data_out_frame[17] [6]), .O(n31298));
    defparam i5_3_lut_4_lut_adj_999.LUT_INIT = 16'h6996;
    SB_LUT4 i13209_3_lut_4_lut (.I0(n8_adj_4404), .I1(n32959), .I2(rx_data[4]), 
            .I3(\data_in_frame[3] [4]), .O(n18038));
    defparam i13209_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13210_3_lut_4_lut (.I0(n8_adj_4404), .I1(n32959), .I2(rx_data[5]), 
            .I3(\data_in_frame[3] [5]), .O(n18039));
    defparam i13210_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i19343_4_lut (.I0(n10_adj_4417), .I1(\FRAME_MATCHER.i [31]), 
            .I2(\FRAME_MATCHER.i [5]), .I3(n16114), .O(n3893));   // verilog/coms.v(252[9:58])
    defparam i19343_4_lut.LUT_INIT = 16'h3332;
    SB_LUT4 i27067_2_lut (.I0(n16154), .I1(n3893), .I2(GND_net), .I3(GND_net), 
            .O(n33657));
    defparam i27067_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i13334_3_lut_4_lut (.I0(n8_adj_4404), .I1(n32952), .I2(rx_data[1]), 
            .I3(\data_in_frame[19] [1]), .O(n18163));
    defparam i13334_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i5_3_lut_adj_1000 (.I0(\data_in[1] [4]), .I1(\data_in[3][0] ), 
            .I2(n15973), .I3(GND_net), .O(n14_adj_4418));
    defparam i5_3_lut_adj_1000.LUT_INIT = 16'hfdfd;
    SB_LUT4 i13211_3_lut_4_lut (.I0(n8_adj_4404), .I1(n32959), .I2(rx_data[6]), 
            .I3(\data_in_frame[3] [6]), .O(n18040));
    defparam i13211_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i6_4_lut_adj_1001 (.I0(\data_in[2] [4]), .I1(n16108), .I2(\data_in[2] [2]), 
            .I3(\data_in[1] [5]), .O(n15_adj_4419));
    defparam i6_4_lut_adj_1001.LUT_INIT = 16'hfffd;
    SB_LUT4 i8_4_lut (.I0(n15_adj_4419), .I1(\data_in[1] [0]), .I2(n14_adj_4418), 
            .I3(\data_in[0][3] ), .O(n22566));
    defparam i8_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i7_4_lut_adj_1002 (.I0(\data_in[1] [2]), .I1(\data_in[1] [3]), 
            .I2(\data_in[2] [5]), .I3(\data_in[1] [6]), .O(n18));
    defparam i7_4_lut_adj_1002.LUT_INIT = 16'hfeff;
    SB_LUT4 i5_2_lut (.I0(\data_in[0][1] ), .I1(\data_in[0][5] ), .I2(GND_net), 
            .I3(GND_net), .O(n16_adj_4420));
    defparam i5_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i9_4_lut_adj_1003 (.I0(\data_in[2] [6]), .I1(n18), .I2(n16097), 
            .I3(\data_in[3][2] ), .O(n20));
    defparam i9_4_lut_adj_1003.LUT_INIT = 16'hfffd;
    SB_LUT4 i10_4_lut_adj_1004 (.I0(\data_in[2] [0]), .I1(n20), .I2(n16_adj_4420), 
            .I3(\data_in[3][7] ), .O(n15973));
    defparam i10_4_lut_adj_1004.LUT_INIT = 16'hfeff;
    SB_DFF data_out_frame_0___i121 (.Q(\data_out_frame[15] [0]), .C(clk32MHz), 
           .D(n17955));   // verilog/coms.v(126[12] 293[6])
    SB_DFF data_out_frame_0___i120 (.Q(\data_out_frame[14] [7]), .C(clk32MHz), 
           .D(n17954));   // verilog/coms.v(126[12] 293[6])
    SB_DFF data_out_frame_0___i119 (.Q(\data_out_frame[14] [6]), .C(clk32MHz), 
           .D(n17953));   // verilog/coms.v(126[12] 293[6])
    SB_DFF data_out_frame_0___i118 (.Q(\data_out_frame[14] [5]), .C(clk32MHz), 
           .D(n17952));   // verilog/coms.v(126[12] 293[6])
    SB_DFF data_out_frame_0___i117 (.Q(\data_out_frame[14] [4]), .C(clk32MHz), 
           .D(n17951));   // verilog/coms.v(126[12] 293[6])
    SB_DFF data_out_frame_0___i116 (.Q(\data_out_frame[14] [3]), .C(clk32MHz), 
           .D(n17950));   // verilog/coms.v(126[12] 293[6])
    SB_DFF data_out_frame_0___i115 (.Q(\data_out_frame[14] [2]), .C(clk32MHz), 
           .D(n17949));   // verilog/coms.v(126[12] 293[6])
    SB_DFF data_out_frame_0___i114 (.Q(\data_out_frame[14] [1]), .C(clk32MHz), 
           .D(n17948));   // verilog/coms.v(126[12] 293[6])
    SB_LUT4 i1_2_lut_adj_1005 (.I0(\data_out_frame[14] [6]), .I1(\data_out_frame[17] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n33158));
    defparam i1_2_lut_adj_1005.LUT_INIT = 16'h6666;
    SB_DFF data_out_frame_0___i113 (.Q(\data_out_frame[14] [0]), .C(clk32MHz), 
           .D(n17947));   // verilog/coms.v(126[12] 293[6])
    SB_DFF data_out_frame_0___i112 (.Q(\data_out_frame[13] [7]), .C(clk32MHz), 
           .D(n17946));   // verilog/coms.v(126[12] 293[6])
    SB_DFF data_out_frame_0___i111 (.Q(\data_out_frame[13] [6]), .C(clk32MHz), 
           .D(n17945));   // verilog/coms.v(126[12] 293[6])
    SB_LUT4 i3_4_lut_adj_1006 (.I0(\data_out_frame[12] [4]), .I1(n33488), 
            .I2(n33287), .I3(n33145), .O(n16570));
    defparam i3_4_lut_adj_1006.LUT_INIT = 16'h6996;
    SB_DFF data_out_frame_0___i110 (.Q(\data_out_frame[13] [5]), .C(clk32MHz), 
           .D(n17944));   // verilog/coms.v(126[12] 293[6])
    SB_DFF data_out_frame_0___i109 (.Q(\data_out_frame[13] [4]), .C(clk32MHz), 
           .D(n17943));   // verilog/coms.v(126[12] 293[6])
    SB_DFF data_out_frame_0___i108 (.Q(\data_out_frame[13] [3]), .C(clk32MHz), 
           .D(n17942));   // verilog/coms.v(126[12] 293[6])
    SB_DFF data_out_frame_0___i107 (.Q(\data_out_frame[13] [2]), .C(clk32MHz), 
           .D(n17941));   // verilog/coms.v(126[12] 293[6])
    SB_DFF data_out_frame_0___i106 (.Q(\data_out_frame[13] [1]), .C(clk32MHz), 
           .D(n17940));   // verilog/coms.v(126[12] 293[6])
    SB_DFF data_out_frame_0___i105 (.Q(\data_out_frame[13] [0]), .C(clk32MHz), 
           .D(n17939));   // verilog/coms.v(126[12] 293[6])
    SB_DFF data_out_frame_0___i104 (.Q(\data_out_frame[12] [7]), .C(clk32MHz), 
           .D(n17938));   // verilog/coms.v(126[12] 293[6])
    SB_DFF data_out_frame_0___i103 (.Q(\data_out_frame[12] [6]), .C(clk32MHz), 
           .D(n17937));   // verilog/coms.v(126[12] 293[6])
    SB_DFF data_out_frame_0___i102 (.Q(\data_out_frame[12] [5]), .C(clk32MHz), 
           .D(n17936));   // verilog/coms.v(126[12] 293[6])
    SB_DFF data_out_frame_0___i101 (.Q(\data_out_frame[12] [4]), .C(clk32MHz), 
           .D(n17935));   // verilog/coms.v(126[12] 293[6])
    SB_DFF data_out_frame_0___i100 (.Q(\data_out_frame[12] [3]), .C(clk32MHz), 
           .D(n17934));   // verilog/coms.v(126[12] 293[6])
    SB_DFF data_out_frame_0___i99 (.Q(\data_out_frame[12] [2]), .C(clk32MHz), 
           .D(n17933));   // verilog/coms.v(126[12] 293[6])
    SB_DFF data_out_frame_0___i98 (.Q(\data_out_frame[12] [1]), .C(clk32MHz), 
           .D(n17932));   // verilog/coms.v(126[12] 293[6])
    SB_LUT4 i1_2_lut_adj_1007 (.I0(\data_out_frame[12] [5]), .I1(\data_out_frame[10] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n33610));
    defparam i1_2_lut_adj_1007.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1008 (.I0(\data_out_frame[12] [6]), .I1(\data_out_frame[15] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n16906));   // verilog/coms.v(70[16:27])
    defparam i1_2_lut_adj_1008.LUT_INIT = 16'h6666;
    SB_DFF data_out_frame_0___i97 (.Q(\data_out_frame[12] [0]), .C(clk32MHz), 
           .D(n17931));   // verilog/coms.v(126[12] 293[6])
    SB_DFF data_out_frame_0___i96 (.Q(\data_out_frame[11] [7]), .C(clk32MHz), 
           .D(n17930));   // verilog/coms.v(126[12] 293[6])
    SB_DFF data_out_frame_0___i95 (.Q(\data_out_frame[11] [6]), .C(clk32MHz), 
           .D(n17929));   // verilog/coms.v(126[12] 293[6])
    SB_DFF data_out_frame_0___i94 (.Q(\data_out_frame[11] [5]), .C(clk32MHz), 
           .D(n17928));   // verilog/coms.v(126[12] 293[6])
    SB_DFF data_out_frame_0___i93 (.Q(\data_out_frame[11] [4]), .C(clk32MHz), 
           .D(n17927));   // verilog/coms.v(126[12] 293[6])
    SB_DFF data_out_frame_0___i92 (.Q(\data_out_frame[11] [3]), .C(clk32MHz), 
           .D(n17926));   // verilog/coms.v(126[12] 293[6])
    SB_LUT4 i1_4_lut_adj_1009 (.I0(\data_in_frame[21] [0]), .I1(n35487), 
            .I2(n6_adj_4421), .I3(n33189), .O(n10_adj_4422));
    defparam i1_4_lut_adj_1009.LUT_INIT = 16'hedde;
    SB_DFF data_out_frame_0___i91 (.Q(\data_out_frame[11] [2]), .C(clk32MHz), 
           .D(n17925));   // verilog/coms.v(126[12] 293[6])
    SB_DFF data_out_frame_0___i90 (.Q(\data_out_frame[11] [1]), .C(clk32MHz), 
           .D(n17924));   // verilog/coms.v(126[12] 293[6])
    SB_LUT4 i13335_3_lut_4_lut (.I0(n8_adj_4404), .I1(n32952), .I2(rx_data[2]), 
            .I3(\data_in_frame[19] [2]), .O(n18164));
    defparam i13335_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF data_out_frame_0___i89 (.Q(\data_out_frame[11] [0]), .C(clk32MHz), 
           .D(n17923));   // verilog/coms.v(126[12] 293[6])
    SB_DFF data_out_frame_0___i88 (.Q(\data_out_frame[10] [7]), .C(clk32MHz), 
           .D(n17922));   // verilog/coms.v(126[12] 293[6])
    SB_DFF data_out_frame_0___i87 (.Q(\data_out_frame[10] [6]), .C(clk32MHz), 
           .D(n17921));   // verilog/coms.v(126[12] 293[6])
    SB_DFF data_out_frame_0___i86 (.Q(\data_out_frame[10] [5]), .C(clk32MHz), 
           .D(n17920));   // verilog/coms.v(126[12] 293[6])
    SB_DFF data_out_frame_0___i85 (.Q(\data_out_frame[10] [4]), .C(clk32MHz), 
           .D(n17919));   // verilog/coms.v(126[12] 293[6])
    SB_DFF data_out_frame_0___i84 (.Q(\data_out_frame[10] [3]), .C(clk32MHz), 
           .D(n17918));   // verilog/coms.v(126[12] 293[6])
    SB_DFF data_out_frame_0___i83 (.Q(\data_out_frame[10] [2]), .C(clk32MHz), 
           .D(n17917));   // verilog/coms.v(126[12] 293[6])
    SB_LUT4 i9_4_lut_adj_1010 (.I0(n16906), .I1(n33164), .I2(n33543), 
            .I3(\data_out_frame[8] [0]), .O(n22_adj_4423));
    defparam i9_4_lut_adj_1010.LUT_INIT = 16'h6996;
    SB_DFF data_out_frame_0___i82 (.Q(\data_out_frame[10] [1]), .C(clk32MHz), 
           .D(n17916));   // verilog/coms.v(126[12] 293[6])
    SB_DFF data_out_frame_0___i81 (.Q(\data_out_frame[10] [0]), .C(clk32MHz), 
           .D(n17915));   // verilog/coms.v(126[12] 293[6])
    SB_DFF data_out_frame_0___i80 (.Q(\data_out_frame[9] [7]), .C(clk32MHz), 
           .D(n17914));   // verilog/coms.v(126[12] 293[6])
    SB_LUT4 i7_3_lut (.I0(\data_out_frame[15] [1]), .I1(n33381), .I2(\data_out_frame[14] [6]), 
            .I3(GND_net), .O(n20_adj_4424));
    defparam i7_3_lut.LUT_INIT = 16'h9696;
    SB_DFF data_out_frame_0___i79 (.Q(\data_out_frame[9] [6]), .C(clk32MHz), 
           .D(n17913));   // verilog/coms.v(126[12] 293[6])
    SB_DFF data_out_frame_0___i78 (.Q(\data_out_frame[9] [5]), .C(clk32MHz), 
           .D(n17912));   // verilog/coms.v(126[12] 293[6])
    SB_DFF data_out_frame_0___i77 (.Q(\data_out_frame[9] [4]), .C(clk32MHz), 
           .D(n17911));   // verilog/coms.v(126[12] 293[6])
    SB_DFF data_out_frame_0___i76 (.Q(\data_out_frame[9] [3]), .C(clk32MHz), 
           .D(n17910));   // verilog/coms.v(126[12] 293[6])
    SB_DFF data_out_frame_0___i75 (.Q(\data_out_frame[9] [2]), .C(clk32MHz), 
           .D(n17909));   // verilog/coms.v(126[12] 293[6])
    SB_DFF data_out_frame_0___i74 (.Q(\data_out_frame[9] [1]), .C(clk32MHz), 
           .D(n17908));   // verilog/coms.v(126[12] 293[6])
    SB_LUT4 i1_4_lut_adj_1011 (.I0(\FRAME_MATCHER.state [3]), .I1(n98), 
            .I2(n53), .I3(n136), .O(n6_adj_4425));   // verilog/coms.v(114[11:12])
    defparam i1_4_lut_adj_1011.LUT_INIT = 16'haaa8;
    SB_DFF data_out_frame_0___i73 (.Q(\data_out_frame[9] [0]), .C(clk32MHz), 
           .D(n17907));   // verilog/coms.v(126[12] 293[6])
    SB_LUT4 i11_4_lut_adj_1012 (.I0(\data_out_frame[7] [6]), .I1(n22_adj_4423), 
            .I2(n16_adj_4426), .I3(n33610), .O(n24));
    defparam i11_4_lut_adj_1012.LUT_INIT = 16'h6996;
    SB_DFF data_out_frame_0___i72 (.Q(\data_out_frame[8] [7]), .C(clk32MHz), 
           .D(n17906));   // verilog/coms.v(126[12] 293[6])
    SB_DFF data_out_frame_0___i71 (.Q(\data_out_frame[8] [6]), .C(clk32MHz), 
           .D(n17905));   // verilog/coms.v(126[12] 293[6])
    SB_DFF data_out_frame_0___i70 (.Q(\data_out_frame[8] [5]), .C(clk32MHz), 
           .D(n17904));   // verilog/coms.v(126[12] 293[6])
    SB_DFF data_out_frame_0___i69 (.Q(\data_out_frame[8] [4]), .C(clk32MHz), 
           .D(n17903));   // verilog/coms.v(126[12] 293[6])
    SB_DFF data_out_frame_0___i68 (.Q(\data_out_frame[8] [3]), .C(clk32MHz), 
           .D(n17902));   // verilog/coms.v(126[12] 293[6])
    SB_LUT4 i1_4_lut_adj_1013 (.I0(n16153), .I1(n6_adj_4425), .I2(\FRAME_MATCHER.state_31__N_2630 [3]), 
            .I3(n16090), .O(n32109));   // verilog/coms.v(114[11:12])
    defparam i1_4_lut_adj_1013.LUT_INIT = 16'hccdc;
    SB_DFF data_out_frame_0___i67 (.Q(\data_out_frame[8] [2]), .C(clk32MHz), 
           .D(n17901));   // verilog/coms.v(126[12] 293[6])
    SB_LUT4 i12_4_lut_adj_1014 (.I0(n16350), .I1(n24), .I2(n20_adj_4424), 
            .I3(\data_out_frame[8] [1]), .O(n34236));
    defparam i12_4_lut_adj_1014.LUT_INIT = 16'h6996;
    SB_DFF data_out_frame_0___i66 (.Q(\data_out_frame[8] [1]), .C(clk32MHz), 
           .D(n17900));   // verilog/coms.v(126[12] 293[6])
    SB_DFF data_out_frame_0___i65 (.Q(\data_out_frame[8] [0]), .C(clk32MHz), 
           .D(n17899));   // verilog/coms.v(126[12] 293[6])
    SB_DFF data_out_frame_0___i64 (.Q(\data_out_frame[7] [7]), .C(clk32MHz), 
           .D(n17898));   // verilog/coms.v(126[12] 293[6])
    SB_LUT4 i1_2_lut_adj_1015 (.I0(\data_in[1] [4]), .I1(\data_in[3][0] ), 
            .I2(GND_net), .I3(GND_net), .O(n158));   // verilog/coms.v(126[12] 293[6])
    defparam i1_2_lut_adj_1015.LUT_INIT = 16'hbbbb;
    SB_DFF data_out_frame_0___i63 (.Q(\data_out_frame[7] [6]), .C(clk32MHz), 
           .D(n17897));   // verilog/coms.v(126[12] 293[6])
    SB_DFF data_out_frame_0___i62 (.Q(\data_out_frame[7] [5]), .C(clk32MHz), 
           .D(n17896));   // verilog/coms.v(126[12] 293[6])
    SB_DFF data_out_frame_0___i61 (.Q(\data_out_frame[7] [4]), .C(clk32MHz), 
           .D(n17895));   // verilog/coms.v(126[12] 293[6])
    SB_LUT4 i13336_3_lut_4_lut (.I0(n8_adj_4404), .I1(n32952), .I2(rx_data[3]), 
            .I3(\data_in_frame[19] [3]), .O(n18165));
    defparam i13336_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF data_out_frame_0___i60 (.Q(\data_out_frame[7] [3]), .C(clk32MHz), 
           .D(n17894));   // verilog/coms.v(126[12] 293[6])
    SB_DFF data_out_frame_0___i59 (.Q(\data_out_frame[7] [2]), .C(clk32MHz), 
           .D(n17893));   // verilog/coms.v(126[12] 293[6])
    SB_DFF data_out_frame_0___i58 (.Q(\data_out_frame[7] [1]), .C(clk32MHz), 
           .D(n17892));   // verilog/coms.v(126[12] 293[6])
    SB_DFF data_out_frame_0___i57 (.Q(\data_out_frame[7] [0]), .C(clk32MHz), 
           .D(n17891));   // verilog/coms.v(126[12] 293[6])
    SB_DFF data_out_frame_0___i56 (.Q(\data_out_frame[6] [7]), .C(clk32MHz), 
           .D(n17890));   // verilog/coms.v(126[12] 293[6])
    SB_LUT4 i6_4_lut_adj_1016 (.I0(\data_in[2] [3]), .I1(n15973), .I2(\data_in[3][6] ), 
            .I3(\data_in[3] [5]), .O(n16_adj_4427));
    defparam i6_4_lut_adj_1016.LUT_INIT = 16'h0200;
    SB_LUT4 i2_3_lut_adj_1017 (.I0(n16158), .I1(\FRAME_MATCHER.state [2]), 
            .I2(\FRAME_MATCHER.state [0]), .I3(GND_net), .O(n16162));   // verilog/coms.v(256[5:27])
    defparam i2_3_lut_adj_1017.LUT_INIT = 16'hfbfb;
    SB_LUT4 i7_4_lut_adj_1018 (.I0(\data_in[0] [2]), .I1(\data_in[2] [1]), 
            .I2(\data_in[3] [3]), .I3(\data_in[3] [1]), .O(n17_adj_4428));
    defparam i7_4_lut_adj_1018.LUT_INIT = 16'h8000;
    SB_DFF data_out_frame_0___i55 (.Q(\data_out_frame[6] [6]), .C(clk32MHz), 
           .D(n17889));   // verilog/coms.v(126[12] 293[6])
    SB_DFF data_out_frame_0___i54 (.Q(\data_out_frame[6] [5]), .C(clk32MHz), 
           .D(n17888));   // verilog/coms.v(126[12] 293[6])
    SB_LUT4 i9_4_lut_adj_1019 (.I0(n17_adj_4428), .I1(\data_in[0][7] ), 
            .I2(n16_adj_4427), .I3(n22269), .O(n35535));
    defparam i9_4_lut_adj_1019.LUT_INIT = 16'h0020;
    SB_DFF data_out_frame_0___i53 (.Q(\data_out_frame[6] [4]), .C(clk32MHz), 
           .D(n17887));   // verilog/coms.v(126[12] 293[6])
    SB_LUT4 i5_4_lut_adj_1020 (.I0(\data_in_frame[2] [6]), .I1(\data_in_frame[0] [4]), 
            .I2(n16319), .I3(\data_in_frame[3] [1]), .O(n12_adj_4429));   // verilog/coms.v(75[16:27])
    defparam i5_4_lut_adj_1020.LUT_INIT = 16'h6996;
    SB_LUT4 i1_3_lut_adj_1021 (.I0(\FRAME_MATCHER.state [3]), .I1(n1_c), 
            .I2(n3_adj_4430), .I3(GND_net), .O(n32183));
    defparam i1_3_lut_adj_1021.LUT_INIT = 16'ha8a8;
    SB_DFF data_out_frame_0___i52 (.Q(\data_out_frame[6] [3]), .C(clk32MHz), 
           .D(n17886));   // verilog/coms.v(126[12] 293[6])
    SB_LUT4 i5_4_lut_adj_1022 (.I0(n16746), .I1(n33439), .I2(\data_out_frame[14] [4]), 
            .I3(n31265), .O(n12_adj_4431));
    defparam i5_4_lut_adj_1022.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1023 (.I0(n31163), .I1(n33195), .I2(n1999), .I3(GND_net), 
            .O(n35212));
    defparam i2_3_lut_adj_1023.LUT_INIT = 16'h9696;
    SB_LUT4 i6_4_lut_adj_1024 (.I0(\data_out_frame[16] [6]), .I1(n12_adj_4431), 
            .I2(n33570), .I3(n16570), .O(n14584));
    defparam i6_4_lut_adj_1024.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1025 (.I0(\data_out_frame[15] [2]), .I1(\data_out_frame[11] [0]), 
            .I2(\data_out_frame[13] [1]), .I3(GND_net), .O(n33262));
    defparam i2_3_lut_adj_1025.LUT_INIT = 16'h9696;
    SB_LUT4 i13337_3_lut_4_lut (.I0(n8_adj_4404), .I1(n32952), .I2(rx_data[4]), 
            .I3(\data_in_frame[19] [4]), .O(n18166));
    defparam i13337_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_1026 (.I0(\data_out_frame[5] [4]), .I1(\data_out_frame[5] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n32979));   // verilog/coms.v(75[16:43])
    defparam i1_2_lut_adj_1026.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_1027 (.I0(\data_out_frame[20] [2]), .I1(n33201), 
            .I2(n31298), .I3(GND_net), .O(n34522));
    defparam i2_3_lut_adj_1027.LUT_INIT = 16'h6969;
    SB_LUT4 i13338_3_lut_4_lut (.I0(n8_adj_4404), .I1(n32952), .I2(rx_data[5]), 
            .I3(\data_in_frame[19] [5]), .O(n18167));
    defparam i13338_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_3_lut_adj_1028 (.I0(n16679), .I1(n33087), .I2(\data_out_frame[18] [2]), 
            .I3(GND_net), .O(n1999));
    defparam i2_3_lut_adj_1028.LUT_INIT = 16'h9696;
    SB_DFF data_out_frame_0___i51 (.Q(\data_out_frame[6] [2]), .C(clk32MHz), 
           .D(n17885));   // verilog/coms.v(126[12] 293[6])
    SB_LUT4 i13339_3_lut_4_lut (.I0(n8_adj_4404), .I1(n32952), .I2(rx_data[6]), 
            .I3(\data_in_frame[19] [6]), .O(n18168));
    defparam i13339_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF data_out_frame_0___i50 (.Q(\data_out_frame[6] [1]), .C(clk32MHz), 
           .D(n17884));   // verilog/coms.v(126[12] 293[6])
    SB_LUT4 i3_4_lut_adj_1029 (.I0(\data_out_frame[5] [7]), .I1(\data_out_frame[6] [0]), 
            .I2(n33377), .I3(n32979), .O(n33589));   // verilog/coms.v(84[17:28])
    defparam i3_4_lut_adj_1029.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1030 (.I0(\data_out_frame[5] [3]), .I1(\data_out_frame[5] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n16795));   // verilog/coms.v(84[17:28])
    defparam i1_2_lut_adj_1030.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_4_lut_adj_1031 (.I0(\FRAME_MATCHER.i [3]), .I1(\FRAME_MATCHER.i [5]), 
            .I2(n16114), .I3(\FRAME_MATCHER.i [4]), .O(n15982));   // verilog/coms.v(153[7:23])
    defparam i2_3_lut_4_lut_adj_1031.LUT_INIT = 16'hfffe;
    SB_LUT4 i2_3_lut_adj_1032 (.I0(\data_out_frame[20] [3]), .I1(n1999), 
            .I2(n35262), .I3(GND_net), .O(n35254));
    defparam i2_3_lut_adj_1032.LUT_INIT = 16'h6969;
    SB_LUT4 i2_3_lut_4_lut_adj_1033 (.I0(\FRAME_MATCHER.i [3]), .I1(\FRAME_MATCHER.i [5]), 
            .I2(\FRAME_MATCHER.i [4]), .I3(n24089), .O(n32952));   // verilog/coms.v(153[7:23])
    defparam i2_3_lut_4_lut_adj_1033.LUT_INIT = 16'hefff;
    SB_LUT4 i13212_3_lut_4_lut (.I0(n8_adj_4404), .I1(n32959), .I2(rx_data[7]), 
            .I3(\data_in_frame[3] [7]), .O(n18041));
    defparam i13212_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_1034 (.I0(n31190), .I1(n33168), .I2(GND_net), 
            .I3(GND_net), .O(n33169));
    defparam i1_2_lut_adj_1034.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1035 (.I0(\data_out_frame[5] [6]), .I1(n33381), 
            .I2(GND_net), .I3(GND_net), .O(n33377));   // verilog/coms.v(84[17:28])
    defparam i1_2_lut_adj_1035.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_3_lut_adj_1036 (.I0(\data_out_frame[11] [1]), .I1(n14531), 
            .I2(n33265), .I3(GND_net), .O(n6_adj_4432));
    defparam i1_2_lut_3_lut_adj_1036.LUT_INIT = 16'h9696;
    SB_DFF data_out_frame_0___i49 (.Q(\data_out_frame[6] [0]), .C(clk32MHz), 
           .D(n17883));   // verilog/coms.v(126[12] 293[6])
    SB_LUT4 i4_4_lut_adj_1037 (.I0(n33514), .I1(\data_out_frame[17] [6]), 
            .I2(\data_out_frame[17] [7]), .I3(n6_adj_4433), .O(n35262));   // verilog/coms.v(77[16:27])
    defparam i4_4_lut_adj_1037.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1038 (.I0(\data_out_frame[11] [1]), .I1(n14531), 
            .I2(n31225), .I3(GND_net), .O(n33549));
    defparam i1_2_lut_3_lut_adj_1038.LUT_INIT = 16'h6969;
    SB_DFF data_out_frame_0___i48 (.Q(\data_out_frame[5] [7]), .C(clk32MHz), 
           .D(n17882));   // verilog/coms.v(126[12] 293[6])
    SB_DFF data_out_frame_0___i47 (.Q(\data_out_frame[5] [6]), .C(clk32MHz), 
           .D(n17881));   // verilog/coms.v(126[12] 293[6])
    SB_LUT4 i2_3_lut_adj_1039 (.I0(n16679), .I1(n16661), .I2(\data_out_frame[19] [7]), 
            .I3(GND_net), .O(n33338));
    defparam i2_3_lut_adj_1039.LUT_INIT = 16'h9696;
    SB_LUT4 i3_4_lut_adj_1040 (.I0(\data_out_frame[17] [6]), .I1(n33511), 
            .I2(n33338), .I3(n30360), .O(n31190));
    defparam i3_4_lut_adj_1040.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1041 (.I0(\data_out_frame[5] [7]), .I1(\data_out_frame[8] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n33013));
    defparam i1_2_lut_adj_1041.LUT_INIT = 16'h6666;
    SB_DFF data_out_frame_0___i46 (.Q(\data_out_frame[5] [5]), .C(clk32MHz), 
           .D(n17880));   // verilog/coms.v(126[12] 293[6])
    SB_DFF data_out_frame_0___i45 (.Q(\data_out_frame[5] [4]), .C(clk32MHz), 
           .D(n17879));   // verilog/coms.v(126[12] 293[6])
    SB_DFF data_out_frame_0___i44 (.Q(\data_out_frame[5] [3]), .C(clk32MHz), 
           .D(n17878));   // verilog/coms.v(126[12] 293[6])
    SB_DFF data_out_frame_0___i43 (.Q(\data_out_frame[5] [2]), .C(clk32MHz), 
           .D(n17877));   // verilog/coms.v(126[12] 293[6])
    SB_DFF data_out_frame_0___i42 (.Q(\data_out_frame[5] [1]), .C(clk32MHz), 
           .D(n17876));   // verilog/coms.v(126[12] 293[6])
    SB_DFF data_out_frame_0___i41 (.Q(\data_out_frame[5] [0]), .C(clk32MHz), 
           .D(n17875));   // verilog/coms.v(126[12] 293[6])
    SB_DFF setpoint__i23 (.Q(setpoint[23]), .C(clk32MHz), .D(n17874));   // verilog/coms.v(126[12] 293[6])
    SB_DFF setpoint__i22 (.Q(setpoint[22]), .C(clk32MHz), .D(n17873));   // verilog/coms.v(126[12] 293[6])
    SB_DFF setpoint__i21 (.Q(setpoint[21]), .C(clk32MHz), .D(n17872));   // verilog/coms.v(126[12] 293[6])
    SB_DFF setpoint__i20 (.Q(setpoint[20]), .C(clk32MHz), .D(n17871));   // verilog/coms.v(126[12] 293[6])
    SB_DFF setpoint__i19 (.Q(setpoint[19]), .C(clk32MHz), .D(n17870));   // verilog/coms.v(126[12] 293[6])
    SB_DFF setpoint__i18 (.Q(setpoint[18]), .C(clk32MHz), .D(n17869));   // verilog/coms.v(126[12] 293[6])
    SB_DFF setpoint__i17 (.Q(setpoint[17]), .C(clk32MHz), .D(n17868));   // verilog/coms.v(126[12] 293[6])
    SB_DFF setpoint__i16 (.Q(setpoint[16]), .C(clk32MHz), .D(n17867));   // verilog/coms.v(126[12] 293[6])
    SB_DFF setpoint__i15 (.Q(setpoint[15]), .C(clk32MHz), .D(n17866));   // verilog/coms.v(126[12] 293[6])
    SB_DFF setpoint__i14 (.Q(setpoint[14]), .C(clk32MHz), .D(n17865));   // verilog/coms.v(126[12] 293[6])
    SB_LUT4 i1_2_lut_adj_1042 (.I0(\FRAME_MATCHER.state [0]), .I1(\FRAME_MATCHER.state [2]), 
            .I2(GND_net), .I3(GND_net), .O(n16090));   // verilog/coms.v(160[5:29])
    defparam i1_2_lut_adj_1042.LUT_INIT = 16'heeee;
    SB_DFF setpoint__i13 (.Q(setpoint[13]), .C(clk32MHz), .D(n17864));   // verilog/coms.v(126[12] 293[6])
    SB_DFF setpoint__i12 (.Q(setpoint[12]), .C(clk32MHz), .D(n17863));   // verilog/coms.v(126[12] 293[6])
    SB_DFF setpoint__i11 (.Q(setpoint[11]), .C(clk32MHz), .D(n17862));   // verilog/coms.v(126[12] 293[6])
    SB_DFF setpoint__i10 (.Q(setpoint[10]), .C(clk32MHz), .D(n17861));   // verilog/coms.v(126[12] 293[6])
    SB_DFF setpoint__i9 (.Q(setpoint[9]), .C(clk32MHz), .D(n17860));   // verilog/coms.v(126[12] 293[6])
    SB_DFF setpoint__i8 (.Q(setpoint[8]), .C(clk32MHz), .D(n17859));   // verilog/coms.v(126[12] 293[6])
    SB_DFF setpoint__i7 (.Q(setpoint[7]), .C(clk32MHz), .D(n17858));   // verilog/coms.v(126[12] 293[6])
    SB_DFF setpoint__i6 (.Q(setpoint[6]), .C(clk32MHz), .D(n17857));   // verilog/coms.v(126[12] 293[6])
    SB_DFF setpoint__i5 (.Q(setpoint[5]), .C(clk32MHz), .D(n17856));   // verilog/coms.v(126[12] 293[6])
    SB_DFF setpoint__i4 (.Q(setpoint[4]), .C(clk32MHz), .D(n17855));   // verilog/coms.v(126[12] 293[6])
    SB_DFF setpoint__i3 (.Q(setpoint[3]), .C(clk32MHz), .D(n17854));   // verilog/coms.v(126[12] 293[6])
    SB_DFF setpoint__i2 (.Q(setpoint[2]), .C(clk32MHz), .D(n17853));   // verilog/coms.v(126[12] 293[6])
    SB_DFF setpoint__i1 (.Q(setpoint[1]), .C(clk32MHz), .D(n17852));   // verilog/coms.v(126[12] 293[6])
    SB_DFF Ki_i15 (.Q(\Ki[15] ), .C(clk32MHz), .D(n17851));   // verilog/coms.v(126[12] 293[6])
    SB_DFF Ki_i14 (.Q(\Ki[14] ), .C(clk32MHz), .D(n17850));   // verilog/coms.v(126[12] 293[6])
    SB_DFF Ki_i13 (.Q(\Ki[13] ), .C(clk32MHz), .D(n17849));   // verilog/coms.v(126[12] 293[6])
    SB_DFF Ki_i12 (.Q(\Ki[12] ), .C(clk32MHz), .D(n17848));   // verilog/coms.v(126[12] 293[6])
    SB_DFF Ki_i11 (.Q(\Ki[11] ), .C(clk32MHz), .D(n17847));   // verilog/coms.v(126[12] 293[6])
    SB_LUT4 i1_2_lut_adj_1043 (.I0(\data_in[0][6] ), .I1(n22566), .I2(GND_net), 
            .I3(GND_net), .O(n67));   // verilog/coms.v(94[12:19])
    defparam i1_2_lut_adj_1043.LUT_INIT = 16'hdddd;
    SB_DFF Ki_i10 (.Q(\Ki[10] ), .C(clk32MHz), .D(n17846));   // verilog/coms.v(126[12] 293[6])
    SB_DFF Ki_i9 (.Q(\Ki[9] ), .C(clk32MHz), .D(n17845));   // verilog/coms.v(126[12] 293[6])
    SB_LUT4 i6_4_lut_adj_1044 (.I0(\data_in_frame[0] [5]), .I1(n12_adj_4429), 
            .I2(n33250), .I3(\data_in_frame[5] [2]), .O(n30217));   // verilog/coms.v(75[16:27])
    defparam i6_4_lut_adj_1044.LUT_INIT = 16'h6996;
    SB_DFF Ki_i8 (.Q(\Ki[8] ), .C(clk32MHz), .D(n17844));   // verilog/coms.v(126[12] 293[6])
    SB_DFF Ki_i7 (.Q(\Ki[7] ), .C(clk32MHz), .D(n17843));   // verilog/coms.v(126[12] 293[6])
    SB_DFF Ki_i6 (.Q(\Ki[6] ), .C(clk32MHz), .D(n17842));   // verilog/coms.v(126[12] 293[6])
    SB_DFF Ki_i5 (.Q(\Ki[5] ), .C(clk32MHz), .D(n17841));   // verilog/coms.v(126[12] 293[6])
    SB_DFF Ki_i4 (.Q(\Ki[4] ), .C(clk32MHz), .D(n17840));   // verilog/coms.v(126[12] 293[6])
    SB_DFF Ki_i3 (.Q(\Ki[3] ), .C(clk32MHz), .D(n17839));   // verilog/coms.v(126[12] 293[6])
    SB_LUT4 i2_3_lut_4_lut_adj_1045 (.I0(\FRAME_MATCHER.state [1]), .I1(n25118), 
            .I2(n16090), .I3(\FRAME_MATCHER.state [3]), .O(n63));   // verilog/coms.v(197[5:24])
    defparam i2_3_lut_4_lut_adj_1045.LUT_INIT = 16'hfeff;
    SB_LUT4 i1_2_lut_3_lut_adj_1046 (.I0(\FRAME_MATCHER.state [1]), .I1(n25118), 
            .I2(\FRAME_MATCHER.state [3]), .I3(GND_net), .O(n16158));   // verilog/coms.v(197[5:24])
    defparam i1_2_lut_3_lut_adj_1046.LUT_INIT = 16'hfefe;
    SB_LUT4 equal_134_i8_2_lut_3_lut (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(\FRAME_MATCHER.i [0]), .I3(GND_net), .O(n8_adj_4404));   // verilog/coms.v(153[7:23])
    defparam equal_134_i8_2_lut_3_lut.LUT_INIT = 16'hdfdf;
    SB_DFF Ki_i2 (.Q(\Ki[2] ), .C(clk32MHz), .D(n17838));   // verilog/coms.v(126[12] 293[6])
    SB_DFF Ki_i1 (.Q(\Ki[1] ), .C(clk32MHz), .D(n17837));   // verilog/coms.v(126[12] 293[6])
    SB_DFF Kp_i15 (.Q(\Kp[15] ), .C(clk32MHz), .D(n17836));   // verilog/coms.v(126[12] 293[6])
    SB_DFF Kp_i14 (.Q(\Kp[14] ), .C(clk32MHz), .D(n17835));   // verilog/coms.v(126[12] 293[6])
    SB_DFF Kp_i13 (.Q(\Kp[13] ), .C(clk32MHz), .D(n17834));   // verilog/coms.v(126[12] 293[6])
    SB_DFF Kp_i12 (.Q(\Kp[12] ), .C(clk32MHz), .D(n17833));   // verilog/coms.v(126[12] 293[6])
    SB_DFF Kp_i11 (.Q(\Kp[11] ), .C(clk32MHz), .D(n17832));   // verilog/coms.v(126[12] 293[6])
    SB_LUT4 i4_4_lut_adj_1047 (.I0(n34726), .I1(n14584), .I2(n30360), 
            .I3(n6_adj_4434), .O(n30231));
    defparam i4_4_lut_adj_1047.LUT_INIT = 16'h9669;
    SB_DFF Kp_i10 (.Q(\Kp[10] ), .C(clk32MHz), .D(n17831));   // verilog/coms.v(126[12] 293[6])
    SB_LUT4 equal_135_i8_2_lut_3_lut (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(\FRAME_MATCHER.i [0]), .I3(GND_net), .O(n8_adj_4435));   // verilog/coms.v(153[7:23])
    defparam equal_135_i8_2_lut_3_lut.LUT_INIT = 16'hfdfd;
    SB_LUT4 i1_2_lut_adj_1048 (.I0(\data_out_frame[6] [2]), .I1(n33368), 
            .I2(GND_net), .I3(GND_net), .O(n16536));
    defparam i1_2_lut_adj_1048.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1049 (.I0(n33287), .I1(\data_out_frame[7] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_4436));
    defparam i1_2_lut_adj_1049.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1050 (.I0(n33377), .I1(\data_out_frame[5] [4]), 
            .I2(n33543), .I3(n6_adj_4436), .O(n31249));
    defparam i4_4_lut_adj_1050.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1051 (.I0(\data_out_frame[12] [5]), .I1(n31249), 
            .I2(n33223), .I3(n16536), .O(n31287));
    defparam i3_4_lut_adj_1051.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_1052 (.I0(\data_in[1] [7]), .I1(\data_in[0][0] ), 
            .I2(\data_in[1] [1]), .I3(\data_in[0][4] ), .O(n10_adj_4437));
    defparam i4_4_lut_adj_1052.LUT_INIT = 16'hfdff;
    SB_LUT4 i5_3_lut_adj_1053 (.I0(\data_in[2] [7]), .I1(n10_adj_4437), 
            .I2(\data_in[3][4] ), .I3(GND_net), .O(n16097));
    defparam i5_3_lut_adj_1053.LUT_INIT = 16'hdfdf;
    SB_LUT4 i2_2_lut (.I0(\data_in[0] [2]), .I1(\data_in[3] [1]), .I2(GND_net), 
            .I3(GND_net), .O(n10_adj_4438));
    defparam i2_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i6_4_lut_adj_1054 (.I0(\data_in[3][6] ), .I1(\data_in[3] [3]), 
            .I2(\data_in[3] [5]), .I3(\data_in[2] [3]), .O(n14_adj_4439));
    defparam i6_4_lut_adj_1054.LUT_INIT = 16'hfffd;
    SB_LUT4 i1_2_lut_adj_1055 (.I0(n30192), .I1(n30231), .I2(GND_net), 
            .I3(GND_net), .O(n16291));
    defparam i1_2_lut_adj_1055.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1056 (.I0(\data_out_frame[6] [3]), .I1(\data_out_frame[8] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n33164));
    defparam i1_2_lut_adj_1056.LUT_INIT = 16'h6666;
    SB_LUT4 i30815_2_lut (.I0(\data_out_frame[23] [0]), .I1(byte_transmit_counter[0]), 
            .I2(GND_net), .I3(GND_net), .O(n37292));
    defparam i30815_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i30884_2_lut (.I0(\data_out_frame[20] [0]), .I1(byte_transmit_counter[0]), 
            .I2(GND_net), .I3(GND_net), .O(n37291));
    defparam i30884_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i1_2_lut_adj_1057 (.I0(\data_out_frame[8] [2]), .I1(\data_out_frame[10] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n33223));
    defparam i1_2_lut_adj_1057.LUT_INIT = 16'h6666;
    SB_LUT4 i13285_3_lut_4_lut (.I0(n8), .I1(n32937), .I2(rx_data[0]), 
            .I3(\data_in_frame[13] [0]), .O(n18114));
    defparam i13285_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i7_4_lut_adj_1058 (.I0(\data_in[0][7] ), .I1(n14_adj_4439), 
            .I2(n10_adj_4438), .I3(\data_in[2] [1]), .O(n16108));
    defparam i7_4_lut_adj_1058.LUT_INIT = 16'hfffd;
    SB_LUT4 i4_4_lut_adj_1059 (.I0(\data_in[1] [0]), .I1(\data_in[0][6] ), 
            .I2(\data_in[2] [4]), .I3(\data_in[0][3] ), .O(n10_adj_4440));
    defparam i4_4_lut_adj_1059.LUT_INIT = 16'hfdff;
    SB_LUT4 i6_4_lut_adj_1060 (.I0(\data_in[1] [6]), .I1(n16097), .I2(\data_in[3][2] ), 
            .I3(\data_in[2] [6]), .O(n16_adj_4441));
    defparam i6_4_lut_adj_1060.LUT_INIT = 16'hffef;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_7_i16_3_lut (.I0(\data_out_frame[16] [7]), 
            .I1(\data_out_frame[17] [7]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n16_adj_4442));   // verilog/coms.v(105[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_7_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_7_i17_3_lut (.I0(\data_out_frame[18] [7]), 
            .I1(\data_out_frame[19] [7]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n17_adj_4443));   // verilog/coms.v(105[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_7_i17_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i7_4_lut_adj_1061 (.I0(n16108), .I1(\data_in[2] [5]), .I2(\data_in[1] [3]), 
            .I3(\data_in[2] [0]), .O(n17_adj_4444));
    defparam i7_4_lut_adj_1061.LUT_INIT = 16'hbfff;
    SB_LUT4 i9_4_lut_adj_1062 (.I0(n17_adj_4444), .I1(\data_in[1] [2]), 
            .I2(n16_adj_4441), .I3(\data_in[0][1] ), .O(n136_adj_4445));
    defparam i9_4_lut_adj_1062.LUT_INIT = 16'hfbff;
    SB_LUT4 i13235_3_lut_4_lut (.I0(n8_adj_4355), .I1(n32959), .I2(rx_data[6]), 
            .I3(\data_in_frame[6] [6]), .O(n18064));
    defparam i13235_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_3_lut_adj_1063 (.I0(\data_out_frame[10] [6]), .I1(\data_out_frame[13] [0]), 
            .I2(\data_out_frame[12] [7]), .I3(GND_net), .O(n33017));   // verilog/coms.v(70[16:27])
    defparam i2_3_lut_adj_1063.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1064 (.I0(\data_out_frame[8] [4]), .I1(\data_out_frame[6] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n4_adj_4412));   // verilog/coms.v(73[16:27])
    defparam i1_2_lut_adj_1064.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1065 (.I0(\data_out_frame[19] [6]), .I1(\data_out_frame[20] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n33511));
    defparam i1_2_lut_adj_1065.LUT_INIT = 16'h6666;
    SB_LUT4 i2_4_lut_adj_1066 (.I0(n15781), .I1(\data_in_frame[19] [3]), 
            .I2(\data_in_frame[21] [5]), .I3(n33430), .O(n34266));
    defparam i2_4_lut_adj_1066.LUT_INIT = 16'h6996;
    SB_LUT4 i1_3_lut_adj_1067 (.I0(\data_in_frame[19] [3]), .I1(n31228), 
            .I2(n15781), .I3(GND_net), .O(n5_adj_4446));
    defparam i1_3_lut_adj_1067.LUT_INIT = 16'h9696;
    SB_LUT4 i2_4_lut_adj_1068 (.I0(n31228), .I1(n33189), .I2(n15781), 
            .I3(\data_in_frame[21] [1]), .O(n34116));
    defparam i2_4_lut_adj_1068.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1069 (.I0(n33323), .I1(\data_in_frame[19] [7]), 
            .I2(n33564), .I3(GND_net), .O(n6_adj_4447));
    defparam i2_3_lut_adj_1069.LUT_INIT = 16'h9696;
    SB_LUT4 i5_4_lut_adj_1070 (.I0(n33171), .I1(n10_adj_4422), .I2(n33430), 
            .I3(\data_in_frame[21] [6]), .O(n14_adj_4448));
    defparam i5_4_lut_adj_1070.LUT_INIT = 16'hdeed;
    SB_LUT4 i3_4_lut_adj_1071 (.I0(n34266), .I1(\data_in_frame[18] [4]), 
            .I2(n8_adj_4449), .I3(\data_in_frame[16] [1]), .O(n12_adj_4450));
    defparam i3_4_lut_adj_1071.LUT_INIT = 16'hebbe;
    SB_LUT4 i4_4_lut_adj_1072 (.I0(n34116), .I1(n5_adj_4446), .I2(\data_in_frame[19] [2]), 
            .I3(\data_in_frame[21] [4]), .O(n13_adj_4451));
    defparam i4_4_lut_adj_1072.LUT_INIT = 16'hbeeb;
    SB_LUT4 i2_4_lut_adj_1073 (.I0(\data_in_frame[20] [0]), .I1(n34664), 
            .I2(n6_adj_4447), .I3(n33186), .O(n11_adj_4452));
    defparam i2_4_lut_adj_1073.LUT_INIT = 16'hedde;
    SB_LUT4 i8_4_lut_adj_1074 (.I0(n11_adj_4452), .I1(n13_adj_4451), .I2(n12_adj_4450), 
            .I3(n14_adj_4448), .O(n31));
    defparam i8_4_lut_adj_1074.LUT_INIT = 16'hfffe;
    SB_LUT4 i13286_3_lut_4_lut (.I0(n8), .I1(n32937), .I2(rx_data[1]), 
            .I3(\data_in_frame[13] [1]), .O(n18115));
    defparam i13286_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13287_3_lut_4_lut (.I0(n8), .I1(n32937), .I2(rx_data[2]), 
            .I3(\data_in_frame[13] [2]), .O(n18116));
    defparam i13287_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_3_lut_adj_1075 (.I0(\data_in_frame[9] [6]), .I1(n30217), 
            .I2(\data_in_frame[7] [4]), .I3(GND_net), .O(n33330));
    defparam i2_3_lut_adj_1075.LUT_INIT = 16'h9696;
    SB_LUT4 i17_4_lut (.I0(\FRAME_MATCHER.i [17]), .I1(\FRAME_MATCHER.i [26]), 
            .I2(\FRAME_MATCHER.i [14]), .I3(\FRAME_MATCHER.i [23]), .O(n42_adj_4453));
    defparam i17_4_lut.LUT_INIT = 16'hfffe;
    SB_DFF data_in_frame_0__i70 (.Q(\data_in_frame[8] [5]), .C(clk32MHz), 
           .D(n18079));   // verilog/coms.v(126[12] 293[6])
    SB_DFF data_in_frame_0__i95 (.Q(\data_in_frame[11] [6]), .C(clk32MHz), 
           .D(n18104));   // verilog/coms.v(126[12] 293[6])
    SB_DFF Kp_i9 (.Q(\Kp[9] ), .C(clk32MHz), .D(n17830));   // verilog/coms.v(126[12] 293[6])
    SB_LUT4 i13288_3_lut_4_lut (.I0(n8), .I1(n32937), .I2(rx_data[3]), 
            .I3(\data_in_frame[13] [3]), .O(n18117));
    defparam i13288_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15_4_lut_adj_1076 (.I0(\FRAME_MATCHER.i [13]), .I1(\FRAME_MATCHER.i [24]), 
            .I2(\FRAME_MATCHER.i [15]), .I3(\FRAME_MATCHER.i [16]), .O(n40));
    defparam i15_4_lut_adj_1076.LUT_INIT = 16'hfffe;
    SB_LUT4 i14_3_lut_4_lut (.I0(\data_out_frame[16] [7]), .I1(\data_out_frame[16] [6]), 
            .I2(n28_adj_4454), .I3(n15783), .O(n32_adj_4455));   // verilog/coms.v(70[16:27])
    defparam i14_3_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1077 (.I0(\data_in_frame[5] [3]), .I1(n33523), 
            .I2(n32994), .I3(Kp_23__N_1026), .O(n16608));   // verilog/coms.v(69[16:69])
    defparam i3_4_lut_adj_1077.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1078 (.I0(\data_in_frame[11] [6]), .I1(\data_in_frame[14] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n33598));
    defparam i1_2_lut_adj_1078.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1079 (.I0(n33477), .I1(n33042), .I2(\data_out_frame[18] [1]), 
            .I3(n33586), .O(n10_adj_4416));
    defparam i4_4_lut_adj_1079.LUT_INIT = 16'h6996;
    SB_LUT4 i13289_3_lut_4_lut (.I0(n8), .I1(n32937), .I2(rx_data[4]), 
            .I3(\data_in_frame[13] [4]), .O(n18118));
    defparam i13289_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF Kp_i8 (.Q(\Kp[8] ), .C(clk32MHz), .D(n17829));   // verilog/coms.v(126[12] 293[6])
    SB_DFF Kp_i7 (.Q(\Kp[7] ), .C(clk32MHz), .D(n17828));   // verilog/coms.v(126[12] 293[6])
    SB_LUT4 i2_3_lut_adj_1080 (.I0(\data_out_frame[8] [6]), .I1(\data_out_frame[6] [5]), 
            .I2(n16350), .I3(GND_net), .O(n33344));
    defparam i2_3_lut_adj_1080.LUT_INIT = 16'h9696;
    SB_LUT4 i3_3_lut_adj_1081 (.I0(\data_out_frame[12] [6]), .I1(n33017), 
            .I2(n33457), .I3(GND_net), .O(n8_adj_4456));   // verilog/coms.v(70[16:27])
    defparam i3_3_lut_adj_1081.LUT_INIT = 16'h9696;
    SB_DFF Kp_i6 (.Q(\Kp[6] ), .C(clk32MHz), .D(n17827));   // verilog/coms.v(126[12] 293[6])
    SB_DFF Kp_i5 (.Q(\Kp[5] ), .C(clk32MHz), .D(n17826));   // verilog/coms.v(126[12] 293[6])
    SB_DFF Kp_i4 (.Q(\Kp[4] ), .C(clk32MHz), .D(n17825));   // verilog/coms.v(126[12] 293[6])
    SB_DFF Kp_i3 (.Q(\Kp[3] ), .C(clk32MHz), .D(n17824));   // verilog/coms.v(126[12] 293[6])
    SB_LUT4 i16_4_lut_adj_1082 (.I0(\FRAME_MATCHER.i [28]), .I1(\FRAME_MATCHER.i [12]), 
            .I2(\FRAME_MATCHER.i [11]), .I3(\FRAME_MATCHER.i [30]), .O(n41));
    defparam i16_4_lut_adj_1082.LUT_INIT = 16'hfffe;
    SB_LUT4 i2_3_lut_4_lut_adj_1083 (.I0(n34691), .I1(\data_in_frame[18] [4]), 
            .I2(\data_in_frame[16] [4]), .I3(\data_in_frame[16] [2]), .O(n33238));
    defparam i2_3_lut_4_lut_adj_1083.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_adj_1084 (.I0(\data_out_frame[20] [5]), .I1(\data_out_frame[20] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n33195));
    defparam i1_2_lut_adj_1084.LUT_INIT = 16'h6666;
    SB_LUT4 i14_4_lut_adj_1085 (.I0(\FRAME_MATCHER.i [7]), .I1(\FRAME_MATCHER.i [20]), 
            .I2(\FRAME_MATCHER.i [22]), .I3(\FRAME_MATCHER.i [25]), .O(n39));
    defparam i14_4_lut_adj_1085.LUT_INIT = 16'hfffe;
    SB_LUT4 i13290_3_lut_4_lut (.I0(n8), .I1(n32937), .I2(rx_data[5]), 
            .I3(\data_in_frame[13] [5]), .O(n18119));
    defparam i13290_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13_3_lut (.I0(\FRAME_MATCHER.i [29]), .I1(\FRAME_MATCHER.i [18]), 
            .I2(\FRAME_MATCHER.i [8]), .I3(GND_net), .O(n38));
    defparam i13_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i1_2_lut_adj_1086 (.I0(\data_out_frame[18] [0]), .I1(\data_out_frame[17] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n16975));   // verilog/coms.v(77[16:27])
    defparam i1_2_lut_adj_1086.LUT_INIT = 16'h6666;
    SB_DFF Kp_i2 (.Q(\Kp[2] ), .C(clk32MHz), .D(n17823));   // verilog/coms.v(126[12] 293[6])
    SB_LUT4 i12_2_lut (.I0(\FRAME_MATCHER.i [21]), .I1(\FRAME_MATCHER.i [10]), 
            .I2(GND_net), .I3(GND_net), .O(n37));
    defparam i12_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i1_2_lut_adj_1087 (.I0(\data_out_frame[19] [6]), .I1(\data_out_frame[19] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n16404));   // verilog/coms.v(77[16:27])
    defparam i1_2_lut_adj_1087.LUT_INIT = 16'h6666;
    SB_LUT4 i11_4_lut_adj_1088 (.I0(n33619), .I1(n16975), .I2(n33210), 
            .I3(n33549), .O(n30_adj_4457));
    defparam i11_4_lut_adj_1088.LUT_INIT = 16'h6996;
    SB_DFF Kp_i1 (.Q(\Kp[1] ), .C(clk32MHz), .D(n17822));   // verilog/coms.v(126[12] 293[6])
    SB_LUT4 i23_4_lut (.I0(n39), .I1(n41), .I2(n40), .I3(n42_adj_4453), 
            .O(n48));
    defparam i23_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_4_lut_adj_1089 (.I0(n33529), .I1(n10_adj_4458), .I2(n33207), 
            .I3(\data_in_frame[18] [3]), .O(n33279));
    defparam i1_2_lut_4_lut_adj_1089.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_1090 (.I0(n16608), .I1(\data_in_frame[11] [7]), 
            .I2(n33631), .I3(n33330), .O(n10_adj_4459));
    defparam i4_4_lut_adj_1090.LUT_INIT = 16'h6996;
    SB_LUT4 i2_2_lut_4_lut (.I0(n33529), .I1(n10_adj_4458), .I2(n33207), 
            .I3(Kp_23__N_843), .O(n7_adj_4460));
    defparam i2_2_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i5_3_lut_adj_1091 (.I0(\data_in_frame[9] [4]), .I1(n10_adj_4459), 
            .I2(n15795), .I3(GND_net), .O(n33505));
    defparam i5_3_lut_adj_1091.LUT_INIT = 16'h9696;
    SB_DFF data_in_0___i32 (.Q(\data_in[3][7] ), .C(clk32MHz), .D(n17821));   // verilog/coms.v(126[12] 293[6])
    SB_LUT4 i15_4_lut_adj_1092 (.I0(n16404), .I1(n30_adj_4457), .I2(n17072), 
            .I3(n33371), .O(n34_adj_4461));
    defparam i15_4_lut_adj_1092.LUT_INIT = 16'h6996;
    SB_DFF data_in_0___i31 (.Q(\data_in[3][6] ), .C(clk32MHz), .D(n17820));   // verilog/coms.v(126[12] 293[6])
    SB_DFF data_in_0___i30 (.Q(\data_in[3] [5]), .C(clk32MHz), .D(n17819));   // verilog/coms.v(126[12] 293[6])
    SB_DFF data_in_0___i29 (.Q(\data_in[3][4] ), .C(clk32MHz), .D(n17818));   // verilog/coms.v(126[12] 293[6])
    SB_DFF data_in_0___i28 (.Q(\data_in[3] [3]), .C(clk32MHz), .D(n17817));   // verilog/coms.v(126[12] 293[6])
    SB_DFF data_in_0___i27 (.Q(\data_in[3][2] ), .C(clk32MHz), .D(n17816));   // verilog/coms.v(126[12] 293[6])
    SB_DFF data_in_0___i26 (.Q(\data_in[3] [1]), .C(clk32MHz), .D(n17815));   // verilog/coms.v(126[12] 293[6])
    SB_LUT4 i1_4_lut_adj_1093 (.I0(n33262), .I1(n33368), .I2(n8_adj_4456), 
            .I3(n4_adj_4412), .O(n4_adj_4462));
    defparam i1_4_lut_adj_1093.LUT_INIT = 16'h6996;
    SB_LUT4 i12866_3_lut_4_lut (.I0(n8_adj_4463), .I1(n32959), .I2(rx_data[0]), 
            .I3(\data_in_frame[0] [0]), .O(n17695));
    defparam i12866_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF data_in_0___i25 (.Q(\data_in[3][0] ), .C(clk32MHz), .D(n17814));   // verilog/coms.v(126[12] 293[6])
    SB_LUT4 i5_4_lut_adj_1094 (.I0(\data_out_frame[13] [0]), .I1(n31287), 
            .I2(\data_out_frame[15] [1]), .I3(\data_out_frame[14] [7]), 
            .O(n12_adj_4464));
    defparam i5_4_lut_adj_1094.LUT_INIT = 16'h6996;
    SB_DFF data_in_0___i24 (.Q(\data_in[2] [7]), .C(clk32MHz), .D(n17813));   // verilog/coms.v(126[12] 293[6])
    SB_LUT4 i6_3_lut (.I0(n4_adj_4462), .I1(n12_adj_4464), .I2(n14531), 
            .I3(GND_net), .O(n30339));
    defparam i6_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 i13182_3_lut_4_lut (.I0(n8_adj_4463), .I1(n32959), .I2(rx_data[1]), 
            .I3(\data_in_frame[0] [1]), .O(n18011));
    defparam i13182_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13183_3_lut_4_lut (.I0(n8_adj_4463), .I1(n32959), .I2(rx_data[2]), 
            .I3(\data_in_frame[0] [2]), .O(n18012));
    defparam i13183_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i18_4_lut (.I0(\FRAME_MATCHER.i [19]), .I1(\FRAME_MATCHER.i [6]), 
            .I2(\FRAME_MATCHER.i [9]), .I3(\FRAME_MATCHER.i [27]), .O(n43));
    defparam i18_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i24_4_lut (.I0(n43), .I1(n48), .I2(n37), .I3(n38), .O(n16114));
    defparam i24_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i13184_3_lut_4_lut (.I0(n8_adj_4463), .I1(n32959), .I2(rx_data[3]), 
            .I3(\data_in_frame[0] [3]), .O(n18013));
    defparam i13184_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF data_in_0___i23 (.Q(\data_in[2] [6]), .C(clk32MHz), .D(n17812));   // verilog/coms.v(126[12] 293[6])
    SB_LUT4 i13185_3_lut_4_lut (.I0(n8_adj_4463), .I1(n32959), .I2(rx_data[4]), 
            .I3(\data_in_frame[0] [4]), .O(n18014));
    defparam i13185_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13186_3_lut_4_lut (.I0(n8_adj_4463), .I1(n32959), .I2(rx_data[5]), 
            .I3(\data_in_frame[0] [5]), .O(n18015));
    defparam i13186_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF data_in_0___i22 (.Q(\data_in[2] [5]), .C(clk32MHz), .D(n17811));   // verilog/coms.v(126[12] 293[6])
    SB_DFF data_in_0___i21 (.Q(\data_in[2] [4]), .C(clk32MHz), .D(n17810));   // verilog/coms.v(126[12] 293[6])
    SB_DFF data_in_0___i20 (.Q(\data_in[2] [3]), .C(clk32MHz), .D(n17809));   // verilog/coms.v(126[12] 293[6])
    SB_LUT4 i13_4_lut_adj_1095 (.I0(n33573), .I1(n33262), .I2(n33451), 
            .I3(n33241), .O(n32_adj_4465));
    defparam i13_4_lut_adj_1095.LUT_INIT = 16'h6996;
    SB_DFF data_in_0___i19 (.Q(\data_in[2] [2]), .C(clk32MHz), .D(n17808));   // verilog/coms.v(126[12] 293[6])
    SB_LUT4 i13187_3_lut_4_lut (.I0(n8_adj_4463), .I1(n32959), .I2(rx_data[6]), 
            .I3(\data_in_frame[0] [6]), .O(n18016));
    defparam i13187_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF data_in_0___i18 (.Q(\data_in[2] [1]), .C(clk32MHz), .D(n17807));   // verilog/coms.v(126[12] 293[6])
    SB_DFF data_in_0___i17 (.Q(\data_in[2] [0]), .C(clk32MHz), .D(n17806));   // verilog/coms.v(126[12] 293[6])
    SB_LUT4 i1_2_lut_adj_1096 (.I0(n15982), .I1(\FRAME_MATCHER.i [2]), .I2(GND_net), 
            .I3(GND_net), .O(n4_adj_4466));
    defparam i1_2_lut_adj_1096.LUT_INIT = 16'heeee;
    SB_LUT4 i14_4_lut_adj_1097 (.I0(n33148), .I1(\data_out_frame[17] [2]), 
            .I2(n33023), .I3(\data_out_frame[18] [5]), .O(n33_adj_4467));
    defparam i14_4_lut_adj_1097.LUT_INIT = 16'h6996;
    SB_LUT4 i12_4_lut_adj_1098 (.I0(n33256), .I1(\data_out_frame[17] [3]), 
            .I2(n33087), .I3(\data_out_frame[19] [4]), .O(n31_adj_4468));
    defparam i12_4_lut_adj_1098.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1099 (.I0(\data_out_frame[19] [2]), .I1(n31178), 
            .I2(GND_net), .I3(GND_net), .O(n33228));
    defparam i1_2_lut_adj_1099.LUT_INIT = 16'h6666;
    SB_LUT4 i13188_3_lut_4_lut (.I0(n8_adj_4463), .I1(n32959), .I2(rx_data[7]), 
            .I3(\data_in_frame[0] [7]), .O(n18017));
    defparam i13188_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i19361_4_lut (.I0(\FRAME_MATCHER.i [0]), .I1(\FRAME_MATCHER.i [31]), 
            .I2(n4_adj_4466), .I3(\FRAME_MATCHER.i [1]), .O(n737));   // verilog/coms.v(156[9:60])
    defparam i19361_4_lut.LUT_INIT = 16'h3230;
    SB_LUT4 i13269_3_lut_4_lut (.I0(n8_adj_4404), .I1(n32937), .I2(rx_data[0]), 
            .I3(\data_in_frame[11] [0]), .O(n18098));
    defparam i13269_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13270_3_lut_4_lut (.I0(n8_adj_4404), .I1(n32937), .I2(rx_data[1]), 
            .I3(\data_in_frame[11] [1]), .O(n18099));
    defparam i13270_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13291_3_lut_4_lut (.I0(n8), .I1(n32937), .I2(rx_data[6]), 
            .I3(\data_in_frame[13] [6]), .O(n18120));
    defparam i13291_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13271_3_lut_4_lut (.I0(n8_adj_4404), .I1(n32937), .I2(rx_data[2]), 
            .I3(\data_in_frame[11] [2]), .O(n18100));
    defparam i13271_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i29826_4_lut (.I0(\data_in_frame[0] [3]), .I1(\data_in_frame[0] [7]), 
            .I2(\data_in_frame[0] [4]), .I3(\data_in_frame[0] [5]), .O(n36430));
    defparam i29826_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i18_4_lut_adj_1100 (.I0(n31_adj_4468), .I1(n33_adj_4467), .I2(n32_adj_4465), 
            .I3(n34_adj_4461), .O(n30968));
    defparam i18_4_lut_adj_1100.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1101 (.I0(\data_out_frame[19] [7]), .I1(n16195), 
            .I2(n16477), .I3(n1981), .O(n33573));
    defparam i3_4_lut_adj_1101.LUT_INIT = 16'h6996;
    SB_LUT4 i13272_3_lut_4_lut (.I0(n8_adj_4404), .I1(n32937), .I2(rx_data[3]), 
            .I3(\data_in_frame[11] [3]), .O(n18101));
    defparam i13272_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i29819_3_lut (.I0(n22275), .I1(\data_in[3][7] ), .I2(\data_in[1] [4]), 
            .I3(GND_net), .O(n36422));
    defparam i29819_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i1_2_lut_adj_1102 (.I0(n10599), .I1(\FRAME_MATCHER.state [1]), 
            .I2(GND_net), .I3(GND_net), .O(n92[1]));   // verilog/coms.v(94[12:19])
    defparam i1_2_lut_adj_1102.LUT_INIT = 16'h8888;
    SB_LUT4 i1_4_lut_adj_1103 (.I0(\data_in[3][0] ), .I1(n92[1]), .I2(n36422), 
            .I3(\data_in[0][5] ), .O(\FRAME_MATCHER.state_31__N_2566[1] ));   // verilog/coms.v(94[12:19])
    defparam i1_4_lut_adj_1103.LUT_INIT = 16'hcecc;
    SB_LUT4 mux_1255_i1_3_lut (.I0(\data_in_frame[19] [0]), .I1(\data_in_frame[3] [0]), 
            .I2(n4995), .I3(GND_net), .O(n4996));
    defparam mux_1255_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2_3_lut_adj_1104 (.I0(n1337), .I1(\data_out_frame[15] [6]), 
            .I2(\data_out_frame[13] [4]), .I3(GND_net), .O(n33042));
    defparam i2_3_lut_adj_1104.LUT_INIT = 16'h9696;
    SB_LUT4 i2_4_lut_adj_1105 (.I0(n35535), .I1(\FRAME_MATCHER.state [0]), 
            .I2(n136_adj_4445), .I3(n4_adj_4469), .O(n32976));
    defparam i2_4_lut_adj_1105.LUT_INIT = 16'heeef;
    SB_LUT4 i13292_3_lut_4_lut (.I0(n8), .I1(n32937), .I2(rx_data[7]), 
            .I3(\data_in_frame[13] [7]), .O(n18121));
    defparam i13292_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_1106 (.I0(\data_in_frame[3] [1]), .I1(\data_in_frame[2] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n33350));   // verilog/coms.v(69[16:69])
    defparam i1_2_lut_adj_1106.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_1107 (.I0(n36418), .I1(n5), .I2(n16159), .I3(n737), 
            .O(n35602));
    defparam i3_4_lut_adj_1107.LUT_INIT = 16'hdddf;
    SB_LUT4 i13273_3_lut_4_lut (.I0(n8_adj_4404), .I1(n32937), .I2(rx_data[4]), 
            .I3(\data_in_frame[11] [4]), .O(n18102));
    defparam i13273_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_4_lut_adj_1108 (.I0(n63), .I1(n42_adj_4411), .I2(n2958), 
            .I3(n32976), .O(n4_adj_4471));   // verilog/coms.v(197[5:24])
    defparam i1_4_lut_adj_1108.LUT_INIT = 16'hf5d5;
    SB_LUT4 i2_4_lut_adj_1109 (.I0(n67), .I1(n4_adj_4471), .I2(n35602), 
            .I3(n32976), .O(n34351));   // verilog/coms.v(197[5:24])
    defparam i2_4_lut_adj_1109.LUT_INIT = 16'hfcdc;
    SB_LUT4 i13197_3_lut_4_lut (.I0(n8_adj_4435), .I1(n32959), .I2(rx_data[0]), 
            .I3(\data_in_frame[2] [0]), .O(n18026));
    defparam i13197_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13274_3_lut_4_lut (.I0(n8_adj_4404), .I1(n32937), .I2(rx_data[5]), 
            .I3(\data_in_frame[11] [5]), .O(n18103));
    defparam i13274_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i30846_2_lut (.I0(\data_out_frame[23] [7]), .I1(byte_transmit_counter[0]), 
            .I2(GND_net), .I3(GND_net), .O(n37283));
    defparam i30846_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i30844_2_lut (.I0(\data_out_frame[20] [7]), .I1(byte_transmit_counter[0]), 
            .I2(GND_net), .I3(GND_net), .O(n37282));
    defparam i30844_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i13275_3_lut_4_lut (.I0(n8_adj_4404), .I1(n32937), .I2(rx_data[6]), 
            .I3(\data_in_frame[11] [6]), .O(n18104));
    defparam i13275_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13276_3_lut_4_lut (.I0(n8_adj_4404), .I1(n32937), .I2(rx_data[7]), 
            .I3(\data_in_frame[11] [7]), .O(n18105));
    defparam i13276_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13251_3_lut_4_lut (.I0(n8_adj_4463), .I1(n32937), .I2(rx_data[6]), 
            .I3(\data_in_frame[8] [6]), .O(n18080));
    defparam i13251_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i4_4_lut_adj_1110 (.I0(\data_out_frame[9] [0]), .I1(n31188), 
            .I2(n17068), .I3(n6_adj_4472), .O(n16954));
    defparam i4_4_lut_adj_1110.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_adj_1111 (.I0(n16726), .I1(n16954), .I2(GND_net), 
            .I3(GND_net), .O(n17135));
    defparam i1_2_lut_adj_1111.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1112 (.I0(\data_in_frame[0] [0]), .I1(\data_in_frame[0] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n9_adj_4473));
    defparam i1_2_lut_adj_1112.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_1113 (.I0(\data_in_frame[3] [3]), .I1(n33558), 
            .I2(GND_net), .I3(GND_net), .O(n33526));   // verilog/coms.v(75[16:27])
    defparam i1_2_lut_adj_1113.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_1114 (.I0(n16319), .I1(n33350), .I2(\data_in_frame[0] [5]), 
            .I3(GND_net), .O(n33523));   // verilog/coms.v(69[16:69])
    defparam i2_3_lut_adj_1114.LUT_INIT = 16'h9696;
    SB_LUT4 i13252_3_lut_4_lut (.I0(n8_adj_4463), .I1(n32937), .I2(rx_data[7]), 
            .I3(\data_in_frame[8] [7]), .O(n18081));
    defparam i13252_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13248_3_lut_4_lut (.I0(n8_adj_4463), .I1(n32937), .I2(rx_data[3]), 
            .I3(\data_in_frame[8] [3]), .O(n18077));
    defparam i13248_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_1115 (.I0(\data_out_frame[13] [3]), .I1(\data_out_frame[15] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n33586));
    defparam i1_2_lut_adj_1115.LUT_INIT = 16'h6666;
    SB_LUT4 i13198_3_lut_4_lut (.I0(n8_adj_4435), .I1(n32959), .I2(rx_data[1]), 
            .I3(\data_in_frame[2] [1]), .O(n18027));
    defparam i13198_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i7_4_lut_adj_1116 (.I0(n9_adj_4473), .I1(n36430), .I2(\data_in_frame[0] [6]), 
            .I3(\data_in_frame[0] [2]), .O(n32855));
    defparam i7_4_lut_adj_1116.LUT_INIT = 16'h0200;
    SB_LUT4 i13249_3_lut_4_lut (.I0(n8_adj_4463), .I1(n32937), .I2(rx_data[4]), 
            .I3(\data_in_frame[8] [4]), .O(n18078));
    defparam i13249_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13199_3_lut_4_lut (.I0(n8_adj_4435), .I1(n32959), .I2(rx_data[2]), 
            .I3(\data_in_frame[2] [2]), .O(n18028));
    defparam i13199_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_3_lut_adj_1117 (.I0(n34996), .I1(n33210), .I2(n30451), 
            .I3(GND_net), .O(n16679));
    defparam i2_3_lut_adj_1117.LUT_INIT = 16'h6969;
    SB_LUT4 i13250_3_lut_4_lut (.I0(n8_adj_4463), .I1(n32937), .I2(rx_data[5]), 
            .I3(\data_in_frame[8] [5]), .O(n18079));
    defparam i13250_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13245_3_lut_4_lut (.I0(n8_adj_4463), .I1(n32937), .I2(rx_data[0]), 
            .I3(\data_in_frame[8] [0]), .O(n18074));
    defparam i13245_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_3_lut_adj_1118 (.I0(\data_out_frame[6] [5]), .I1(n33057), 
            .I2(\data_out_frame[10] [7]), .I3(GND_net), .O(n16998));   // verilog/coms.v(74[16:27])
    defparam i2_3_lut_adj_1118.LUT_INIT = 16'h9696;
    SB_LUT4 i13246_3_lut_4_lut (.I0(n8_adj_4463), .I1(n32937), .I2(rx_data[1]), 
            .I3(\data_in_frame[8] [1]), .O(n18075));
    defparam i13246_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_4_lut_adj_1119 (.I0(n30769), .I1(n16998), .I2(\data_out_frame[17] [4]), 
            .I3(n4_adj_4462), .O(n30360));
    defparam i2_4_lut_adj_1119.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1120 (.I0(n30360), .I1(n16679), .I2(\data_out_frame[18] [1]), 
            .I3(GND_net), .O(n33442));
    defparam i2_3_lut_adj_1120.LUT_INIT = 16'h9696;
    SB_LUT4 i12_4_lut_adj_1121 (.I0(\data_out_frame[11] [3]), .I1(\data_out_frame[16] [0]), 
            .I2(\data_out_frame[10] [6]), .I3(\data_out_frame[17] [4]), 
            .O(n28_adj_4474));
    defparam i12_4_lut_adj_1121.LUT_INIT = 16'h6996;
    SB_LUT4 i13247_3_lut_4_lut (.I0(n8_adj_4463), .I1(n32937), .I2(rx_data[2]), 
            .I3(\data_in_frame[8] [2]), .O(n18076));
    defparam i13247_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_3_lut_4_lut_adj_1122 (.I0(\FRAME_MATCHER.i [4]), .I1(\FRAME_MATCHER.i [5]), 
            .I2(\FRAME_MATCHER.i [3]), .I3(n24089), .O(n32959));   // verilog/coms.v(153[7:23])
    defparam i2_3_lut_4_lut_adj_1122.LUT_INIT = 16'hfeff;
    SB_LUT4 i10_4_lut_adj_1123 (.I0(n33457), .I1(\data_out_frame[13] [6]), 
            .I2(\data_out_frame[10] [5]), .I3(n30241), .O(n26_adj_4475));
    defparam i10_4_lut_adj_1123.LUT_INIT = 16'h6996;
    SB_LUT4 i11_4_lut_adj_1124 (.I0(n33576), .I1(\data_out_frame[15] [0]), 
            .I2(n33069), .I3(n34521), .O(n27_adj_4476));
    defparam i11_4_lut_adj_1124.LUT_INIT = 16'h9669;
    SB_LUT4 i9_4_lut_adj_1125 (.I0(\data_out_frame[12] [7]), .I1(n32985), 
            .I2(\data_out_frame[14] [0]), .I3(\data_out_frame[15] [1]), 
            .O(n25_adj_4477));
    defparam i9_4_lut_adj_1125.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_1126 (.I0(\FRAME_MATCHER.i [4]), .I1(\FRAME_MATCHER.i [5]), 
            .I2(\FRAME_MATCHER.i [3]), .I3(n24089), .O(n32937));   // verilog/coms.v(153[7:23])
    defparam i2_3_lut_4_lut_adj_1126.LUT_INIT = 16'hefff;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1127 (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(n32959), .I3(\FRAME_MATCHER.i [0]), .O(n32962));   // verilog/coms.v(153[7:23])
    defparam i1_2_lut_3_lut_4_lut_adj_1127.LUT_INIT = 16'hfeff;
    SB_LUT4 i15_4_lut_adj_1128 (.I0(n25_adj_4477), .I1(n27_adj_4476), .I2(n26_adj_4475), 
            .I3(n28_adj_4474), .O(n33619));
    defparam i15_4_lut_adj_1128.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1129 (.I0(\data_out_frame[14] [3]), .I1(\data_out_frame[16] [5]), 
            .I2(\data_out_frame[14] [4]), .I3(GND_net), .O(n33175));
    defparam i2_3_lut_adj_1129.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1130 (.I0(\data_out_frame[19] [2]), .I1(\data_out_frame[19] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n16477));
    defparam i1_2_lut_adj_1130.LUT_INIT = 16'h6666;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[14] [4]), .I2(\data_out_frame[15] [4]), 
            .I3(byte_transmit_counter_c[1]), .O(n38459));
    defparam byte_transmit_counter_0__bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_LUT4 n38459_bdd_4_lut (.I0(n38459), .I1(\data_out_frame[13] [4]), 
            .I2(\data_out_frame[12] [4]), .I3(byte_transmit_counter_c[1]), 
            .O(n38462));
    defparam n38459_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_31743 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[14] [3]), .I2(\data_out_frame[15] [3]), 
            .I3(byte_transmit_counter_c[1]), .O(n38453));
    defparam byte_transmit_counter_0__bdd_4_lut_31743.LUT_INIT = 16'he4aa;
    SB_LUT4 n38453_bdd_4_lut (.I0(n38453), .I1(\data_out_frame[13] [3]), 
            .I2(\data_out_frame[12] [3]), .I3(byte_transmit_counter_c[1]), 
            .O(n38456));
    defparam n38453_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_31738 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[14] [2]), .I2(\data_out_frame[15] [2]), 
            .I3(byte_transmit_counter_c[1]), .O(n38447));
    defparam byte_transmit_counter_0__bdd_4_lut_31738.LUT_INIT = 16'he4aa;
    SB_LUT4 n38447_bdd_4_lut (.I0(n38447), .I1(\data_out_frame[13] [2]), 
            .I2(\data_out_frame[12] [2]), .I3(byte_transmit_counter_c[1]), 
            .O(n38450));
    defparam n38447_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_31733 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[14] [1]), .I2(\data_out_frame[15] [1]), 
            .I3(byte_transmit_counter_c[1]), .O(n38441));
    defparam byte_transmit_counter_0__bdd_4_lut_31733.LUT_INIT = 16'he4aa;
    SB_LUT4 n38441_bdd_4_lut (.I0(n38441), .I1(\data_out_frame[13] [1]), 
            .I2(\data_out_frame[12] [1]), .I3(byte_transmit_counter_c[1]), 
            .O(n38444));
    defparam n38441_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_31728 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[10] [1]), .I2(\data_out_frame[11] [1]), 
            .I3(byte_transmit_counter_c[1]), .O(n38435));
    defparam byte_transmit_counter_0__bdd_4_lut_31728.LUT_INIT = 16'he4aa;
    SB_LUT4 n38435_bdd_4_lut (.I0(n38435), .I1(\data_out_frame[9] [1]), 
            .I2(\data_out_frame[8] [1]), .I3(byte_transmit_counter_c[1]), 
            .O(n38438));
    defparam n38435_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_3__bdd_4_lut (.I0(byte_transmit_counter_c[3]), 
            .I1(n38258), .I2(n37290), .I3(byte_transmit_counter_c[4]), 
            .O(n38423));
    defparam byte_transmit_counter_3__bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_LUT4 n38423_bdd_4_lut (.I0(n38423), .I1(n14_adj_4396), .I2(n7_adj_4395), 
            .I3(byte_transmit_counter_c[4]), .O(tx_data[0]));
    defparam n38423_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_3__bdd_4_lut_31714 (.I0(byte_transmit_counter_c[3]), 
            .I1(n38264), .I2(n37281), .I3(byte_transmit_counter_c[4]), 
            .O(n38417));
    defparam byte_transmit_counter_3__bdd_4_lut_31714.LUT_INIT = 16'he4aa;
    SB_LUT4 n38417_bdd_4_lut (.I0(n38417), .I1(n14_adj_4392), .I2(n7_adj_4391), 
            .I3(byte_transmit_counter_c[4]), .O(tx_data[7]));
    defparam n38417_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_6_i16_3_lut (.I0(\data_out_frame[16] [6]), 
            .I1(\data_out_frame[17] [6]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n16_adj_4478));   // verilog/coms.v(105[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_6_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1131 (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(n32937), .I3(\FRAME_MATCHER.i [0]), .O(n32941));   // verilog/coms.v(153[7:23])
    defparam i1_2_lut_3_lut_4_lut_adj_1131.LUT_INIT = 16'hfeff;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_6_i17_3_lut (.I0(\data_out_frame[18] [6]), 
            .I1(\data_out_frame[19] [6]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n17_adj_4479));   // verilog/coms.v(105[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_6_i17_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i30849_2_lut (.I0(\data_out_frame[23][6] ), .I1(byte_transmit_counter[0]), 
            .I2(GND_net), .I3(GND_net), .O(n37280));
    defparam i30849_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i30843_2_lut (.I0(\data_out_frame[20] [6]), .I1(byte_transmit_counter[0]), 
            .I2(GND_net), .I3(GND_net), .O(n37279));
    defparam i30843_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 byte_transmit_counter_3__bdd_4_lut_31709 (.I0(byte_transmit_counter_c[3]), 
            .I1(n38270), .I2(n37278), .I3(byte_transmit_counter_c[4]), 
            .O(n38411));
    defparam byte_transmit_counter_3__bdd_4_lut_31709.LUT_INIT = 16'he4aa;
    SB_LUT4 n38411_bdd_4_lut (.I0(n38411), .I1(n14_adj_4384), .I2(n7_adj_4383), 
            .I3(byte_transmit_counter_c[4]), .O(tx_data[6]));
    defparam n38411_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_3__bdd_4_lut_31704 (.I0(byte_transmit_counter_c[3]), 
            .I1(n38276), .I2(n37275), .I3(byte_transmit_counter_c[4]), 
            .O(n38405));
    defparam byte_transmit_counter_3__bdd_4_lut_31704.LUT_INIT = 16'he4aa;
    SB_LUT4 n38405_bdd_4_lut (.I0(n38405), .I1(n14_adj_4377), .I2(n7_adj_4375), 
            .I3(byte_transmit_counter_c[4]), .O(tx_data[5]));
    defparam n38405_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_3__bdd_4_lut_31699 (.I0(byte_transmit_counter_c[3]), 
            .I1(n38282), .I2(n37272), .I3(byte_transmit_counter_c[4]), 
            .O(n38399));
    defparam byte_transmit_counter_3__bdd_4_lut_31699.LUT_INIT = 16'he4aa;
    SB_LUT4 n38399_bdd_4_lut (.I0(n38399), .I1(n14_adj_4370), .I2(n7_adj_4369), 
            .I3(byte_transmit_counter_c[4]), .O(tx_data[4]));
    defparam n38399_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut (.I0(byte_transmit_counter_c[1]), 
            .I1(n37270), .I2(n37271), .I3(byte_transmit_counter_c[2]), 
            .O(n38393));
    defparam byte_transmit_counter_1__bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_LUT4 n38393_bdd_4_lut (.I0(n38393), .I1(n17), .I2(n16), .I3(byte_transmit_counter_c[2]), 
            .O(n37807));
    defparam n38393_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_3__bdd_4_lut_31694 (.I0(byte_transmit_counter_c[3]), 
            .I1(n37807), .I2(n37269), .I3(byte_transmit_counter_c[4]), 
            .O(n38387));
    defparam byte_transmit_counter_3__bdd_4_lut_31694.LUT_INIT = 16'he4aa;
    SB_LUT4 n38387_bdd_4_lut (.I0(n38387), .I1(n14_adj_4366), .I2(n7_adj_4365), 
            .I3(byte_transmit_counter_c[4]), .O(tx_data[3]));
    defparam n38387_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_3__bdd_4_lut_31684 (.I0(byte_transmit_counter_c[3]), 
            .I1(n38306), .I2(n37266), .I3(byte_transmit_counter_c[4]), 
            .O(n38381));
    defparam byte_transmit_counter_3__bdd_4_lut_31684.LUT_INIT = 16'he4aa;
    SB_LUT4 n38381_bdd_4_lut (.I0(n38381), .I1(n14_adj_4362), .I2(n7_adj_4361), 
            .I3(byte_transmit_counter_c[4]), .O(tx_data[2]));
    defparam n38381_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_3__bdd_4_lut_31679 (.I0(byte_transmit_counter_c[3]), 
            .I1(n38336), .I2(n37257), .I3(byte_transmit_counter_c[4]), 
            .O(n38375));
    defparam byte_transmit_counter_3__bdd_4_lut_31679.LUT_INIT = 16'he4aa;
    SB_LUT4 n38375_bdd_4_lut (.I0(n38375), .I1(n14_adj_4358), .I2(n7_adj_4357), 
            .I3(byte_transmit_counter_c[4]), .O(tx_data[1]));
    defparam n38375_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_31723 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[10] [6]), .I2(\data_out_frame[11] [6]), 
            .I3(byte_transmit_counter_c[1]), .O(n38369));
    defparam byte_transmit_counter_0__bdd_4_lut_31723.LUT_INIT = 16'he4aa;
    SB_LUT4 n38369_bdd_4_lut (.I0(n38369), .I1(\data_out_frame[9] [6]), 
            .I2(\data_out_frame[8] [6]), .I3(byte_transmit_counter_c[1]), 
            .O(n38372));
    defparam n38369_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_31670 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[10] [7]), .I2(\data_out_frame[11] [7]), 
            .I3(byte_transmit_counter_c[1]), .O(n38363));
    defparam byte_transmit_counter_0__bdd_4_lut_31670.LUT_INIT = 16'he4aa;
    SB_LUT4 n38363_bdd_4_lut (.I0(n38363), .I1(\data_out_frame[9] [7]), 
            .I2(\data_out_frame[8] [7]), .I3(byte_transmit_counter_c[1]), 
            .O(n38366));
    defparam n38363_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_5_i16_3_lut (.I0(\data_out_frame[16] [5]), 
            .I1(\data_out_frame[17] [5]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n16_adj_4480));   // verilog/coms.v(105[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_5_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_5_i17_3_lut (.I0(\data_out_frame[18] [5]), 
            .I1(\data_out_frame[19] [5]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n17_adj_4481));   // verilog/coms.v(105[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_5_i17_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10_4_lut_adj_1132 (.I0(\data_out_frame[15] [4]), .I1(n33424), 
            .I2(n31265), .I3(n16946), .O(n28_adj_4454));
    defparam i10_4_lut_adj_1132.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut_adj_1133 (.I0(n33175), .I1(n1337), .I2(n33436), .I3(n31265), 
            .O(n25_adj_4482));
    defparam i7_4_lut_adj_1133.LUT_INIT = 16'h9669;
    SB_LUT4 equal_121_i8_2_lut_3_lut (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(\FRAME_MATCHER.i [0]), .I3(GND_net), .O(n8_adj_4463));   // verilog/coms.v(153[7:23])
    defparam equal_121_i8_2_lut_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i12_4_lut_adj_1134 (.I0(n31209), .I1(n33292), .I2(n33619), 
            .I3(n33073), .O(n30_adj_4483));
    defparam i12_4_lut_adj_1134.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1135 (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(n32952), .I3(\FRAME_MATCHER.i [0]), .O(n32957));   // verilog/coms.v(153[7:23])
    defparam i1_2_lut_3_lut_4_lut_adj_1135.LUT_INIT = 16'hfeff;
    SB_LUT4 i2_3_lut_adj_1136 (.I0(\data_in_frame[2] [3]), .I1(\data_in_frame[0] [1]), 
            .I2(\data_in_frame[0] [2]), .I3(GND_net), .O(n4_adj_4410));   // verilog/coms.v(165[9:87])
    defparam i2_3_lut_adj_1136.LUT_INIT = 16'h9696;
    SB_LUT4 add_41_33_lut (.I0(n2290), .I1(\FRAME_MATCHER.i [31]), .I2(GND_net), 
            .I3(n27939), .O(n2_adj_4484)) /* synthesis syn_instantiated=1 */ ;
    defparam add_41_33_lut.LUT_INIT = 16'h8228;
    SB_DFFSS \FRAME_MATCHER.i_i1  (.Q(\FRAME_MATCHER.i [1]), .C(clk32MHz), 
            .D(n2_adj_4340), .S(n3_adj_4485));   // verilog/coms.v(126[12] 293[6])
    SB_LUT4 i2_3_lut_adj_1137 (.I0(n31), .I1(n32855), .I2(n16162), .I3(GND_net), 
            .O(n5439));
    defparam i2_3_lut_adj_1137.LUT_INIT = 16'h0404;
    SB_LUT4 i30854_2_lut (.I0(\data_out_frame[23] [5]), .I1(byte_transmit_counter[0]), 
            .I2(GND_net), .I3(GND_net), .O(n37277));
    defparam i30854_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i16_4_lut_adj_1138 (.I0(n25_adj_4482), .I1(n32_adj_4455), .I2(n30451), 
            .I3(\data_out_frame[15] [2]), .O(n34_adj_4486));
    defparam i16_4_lut_adj_1138.LUT_INIT = 16'h6996;
    SB_LUT4 i11_4_lut_adj_1139 (.I0(n17135), .I1(n31249), .I2(n33178), 
            .I3(n30769), .O(n29_adj_4487));
    defparam i11_4_lut_adj_1139.LUT_INIT = 16'h9669;
    SB_LUT4 i30841_2_lut (.I0(\data_out_frame[20] [5]), .I1(byte_transmit_counter[0]), 
            .I2(GND_net), .I3(GND_net), .O(n37276));
    defparam i30841_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i6_4_lut_adj_1140 (.I0(n4_adj_4410), .I1(\data_in_frame[2] [4]), 
            .I2(\data_in_frame[0] [6]), .I3(\data_in_frame[2] [2]), .O(n16_adj_4488));   // verilog/coms.v(74[16:43])
    defparam i6_4_lut_adj_1140.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut_adj_1141 (.I0(\data_in_frame[0] [0]), .I1(n33523), 
            .I2(n33526), .I3(\data_in_frame[0] [7]), .O(n17_adj_4489));   // verilog/coms.v(74[16:43])
    defparam i7_4_lut_adj_1141.LUT_INIT = 16'h6996;
    SB_DFF data_in_frame_0__i94 (.Q(\data_in_frame[11] [5]), .C(clk32MHz), 
           .D(n18103));   // verilog/coms.v(126[12] 293[6])
    SB_DFF data_in_frame_0__i93 (.Q(\data_in_frame[11] [4]), .C(clk32MHz), 
           .D(n18102));   // verilog/coms.v(126[12] 293[6])
    SB_LUT4 i4_4_lut_adj_1142 (.I0(n29_adj_4487), .I1(n33442), .I2(n34_adj_4486), 
            .I3(n30_adj_4483), .O(n17_adj_4490));
    defparam i4_4_lut_adj_1142.LUT_INIT = 16'h9669;
    SB_LUT4 i13349_3_lut_4_lut (.I0(n8), .I1(n32952), .I2(rx_data[0]), 
            .I3(\data_in_frame[21] [0]), .O(n18178));
    defparam i13349_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i8_4_lut_adj_1143 (.I0(\data_out_frame[17] [6]), .I1(\data_out_frame[17] [7]), 
            .I2(n33573), .I3(n30339), .O(n21_adj_4491));
    defparam i8_4_lut_adj_1143.LUT_INIT = 16'h6996;
    SB_DFF data_in_frame_0__i92 (.Q(\data_in_frame[11] [3]), .C(clk32MHz), 
           .D(n18101));   // verilog/coms.v(126[12] 293[6])
    SB_LUT4 add_41_32_lut (.I0(n2290), .I1(\FRAME_MATCHER.i [30]), .I2(GND_net), 
            .I3(n27938), .O(n2_adj_4492)) /* synthesis syn_instantiated=1 */ ;
    defparam add_41_32_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i13351_3_lut_4_lut (.I0(n8), .I1(n32952), .I2(rx_data[2]), 
            .I3(\data_in_frame[21] [2]), .O(n18180));
    defparam i13351_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_CARRY add_41_32 (.CI(n27938), .I0(\FRAME_MATCHER.i [30]), .I1(GND_net), 
            .CO(n27939));
    SB_LUT4 add_41_31_lut (.I0(n2290), .I1(\FRAME_MATCHER.i [29]), .I2(GND_net), 
            .I3(n27937), .O(n2_adj_4493)) /* synthesis syn_instantiated=1 */ ;
    defparam add_41_31_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_41_31 (.CI(n27937), .I0(\FRAME_MATCHER.i [29]), .I1(GND_net), 
            .CO(n27938));
    SB_LUT4 add_41_30_lut (.I0(n2290), .I1(\FRAME_MATCHER.i [28]), .I2(GND_net), 
            .I3(n27936), .O(n2_adj_4494)) /* synthesis syn_instantiated=1 */ ;
    defparam add_41_30_lut.LUT_INIT = 16'h8228;
    SB_DFFSS \FRAME_MATCHER.i_i2  (.Q(\FRAME_MATCHER.i [2]), .C(clk32MHz), 
            .D(n2_adj_4495), .S(n3_adj_4496));   // verilog/coms.v(126[12] 293[6])
    SB_LUT4 i13350_3_lut_4_lut (.I0(n8), .I1(n32952), .I2(rx_data[1]), 
            .I3(\data_in_frame[21] [1]), .O(n18179));
    defparam i13350_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13353_3_lut_4_lut (.I0(n8), .I1(n32952), .I2(rx_data[4]), 
            .I3(\data_in_frame[21] [4]), .O(n18182));
    defparam i13353_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFFSS \FRAME_MATCHER.i_i3  (.Q(\FRAME_MATCHER.i [3]), .C(clk32MHz), 
            .D(n2_adj_4497), .S(n3_adj_4498));   // verilog/coms.v(126[12] 293[6])
    SB_DFFSS \FRAME_MATCHER.i_i4  (.Q(\FRAME_MATCHER.i [4]), .C(clk32MHz), 
            .D(n2_adj_4499), .S(n3_adj_4500));   // verilog/coms.v(126[12] 293[6])
    SB_DFFSS \FRAME_MATCHER.i_i5  (.Q(\FRAME_MATCHER.i [5]), .C(clk32MHz), 
            .D(n2_adj_4501), .S(n3_adj_4502));   // verilog/coms.v(126[12] 293[6])
    SB_DFFSS \FRAME_MATCHER.i_i6  (.Q(\FRAME_MATCHER.i [6]), .C(clk32MHz), 
            .D(n2_adj_4503), .S(n3_adj_4504));   // verilog/coms.v(126[12] 293[6])
    SB_DFFSS \FRAME_MATCHER.i_i7  (.Q(\FRAME_MATCHER.i [7]), .C(clk32MHz), 
            .D(n2_adj_4505), .S(n3_adj_4506));   // verilog/coms.v(126[12] 293[6])
    SB_DFFSS \FRAME_MATCHER.i_i8  (.Q(\FRAME_MATCHER.i [8]), .C(clk32MHz), 
            .D(n2_adj_4507), .S(n3_adj_4508));   // verilog/coms.v(126[12] 293[6])
    SB_DFFSS \FRAME_MATCHER.i_i9  (.Q(\FRAME_MATCHER.i [9]), .C(clk32MHz), 
            .D(n2_adj_4509), .S(n3_adj_4510));   // verilog/coms.v(126[12] 293[6])
    SB_DFFSS \FRAME_MATCHER.i_i10  (.Q(\FRAME_MATCHER.i [10]), .C(clk32MHz), 
            .D(n2_adj_4511), .S(n3_adj_4512));   // verilog/coms.v(126[12] 293[6])
    SB_DFFSS \FRAME_MATCHER.i_i11  (.Q(\FRAME_MATCHER.i [11]), .C(clk32MHz), 
            .D(n2_adj_4513), .S(n3_adj_4514));   // verilog/coms.v(126[12] 293[6])
    SB_DFFSS \FRAME_MATCHER.i_i12  (.Q(\FRAME_MATCHER.i [12]), .C(clk32MHz), 
            .D(n2_adj_4515), .S(n3_adj_4516));   // verilog/coms.v(126[12] 293[6])
    SB_DFFSS \FRAME_MATCHER.i_i13  (.Q(\FRAME_MATCHER.i [13]), .C(clk32MHz), 
            .D(n2_adj_4517), .S(n3_adj_4518));   // verilog/coms.v(126[12] 293[6])
    SB_DFFSS \FRAME_MATCHER.i_i14  (.Q(\FRAME_MATCHER.i [14]), .C(clk32MHz), 
            .D(n2_adj_4519), .S(n3_adj_4520));   // verilog/coms.v(126[12] 293[6])
    SB_DFFSS \FRAME_MATCHER.i_i15  (.Q(\FRAME_MATCHER.i [15]), .C(clk32MHz), 
            .D(n2_adj_4521), .S(n3_adj_4522));   // verilog/coms.v(126[12] 293[6])
    SB_DFFSS \FRAME_MATCHER.i_i16  (.Q(\FRAME_MATCHER.i [16]), .C(clk32MHz), 
            .D(n2_adj_4523), .S(n3_adj_4524));   // verilog/coms.v(126[12] 293[6])
    SB_DFFSS \FRAME_MATCHER.i_i17  (.Q(\FRAME_MATCHER.i [17]), .C(clk32MHz), 
            .D(n2_adj_4525), .S(n3_adj_4526));   // verilog/coms.v(126[12] 293[6])
    SB_DFFSS \FRAME_MATCHER.i_i18  (.Q(\FRAME_MATCHER.i [18]), .C(clk32MHz), 
            .D(n2_adj_4527), .S(n3_adj_4528));   // verilog/coms.v(126[12] 293[6])
    SB_DFFSS \FRAME_MATCHER.i_i19  (.Q(\FRAME_MATCHER.i [19]), .C(clk32MHz), 
            .D(n2_adj_4529), .S(n3_adj_4530));   // verilog/coms.v(126[12] 293[6])
    SB_DFFSS \FRAME_MATCHER.i_i20  (.Q(\FRAME_MATCHER.i [20]), .C(clk32MHz), 
            .D(n2_adj_4531), .S(n3_adj_4532));   // verilog/coms.v(126[12] 293[6])
    SB_DFFSS \FRAME_MATCHER.i_i21  (.Q(\FRAME_MATCHER.i [21]), .C(clk32MHz), 
            .D(n2_adj_4533), .S(n3_adj_4534));   // verilog/coms.v(126[12] 293[6])
    SB_DFFSS \FRAME_MATCHER.i_i22  (.Q(\FRAME_MATCHER.i [22]), .C(clk32MHz), 
            .D(n2_adj_4535), .S(n3_adj_4536));   // verilog/coms.v(126[12] 293[6])
    SB_DFFSS \FRAME_MATCHER.i_i23  (.Q(\FRAME_MATCHER.i [23]), .C(clk32MHz), 
            .D(n2_adj_4537), .S(n3_adj_4538));   // verilog/coms.v(126[12] 293[6])
    SB_DFFSS \FRAME_MATCHER.i_i24  (.Q(\FRAME_MATCHER.i [24]), .C(clk32MHz), 
            .D(n2_adj_4539), .S(n3_adj_4540));   // verilog/coms.v(126[12] 293[6])
    SB_DFFSS \FRAME_MATCHER.i_i25  (.Q(\FRAME_MATCHER.i [25]), .C(clk32MHz), 
            .D(n2_adj_4541), .S(n3_adj_4542));   // verilog/coms.v(126[12] 293[6])
    SB_DFFSS \FRAME_MATCHER.i_i26  (.Q(\FRAME_MATCHER.i [26]), .C(clk32MHz), 
            .D(n2_adj_4543), .S(n3_adj_4544));   // verilog/coms.v(126[12] 293[6])
    SB_DFFSS \FRAME_MATCHER.i_i27  (.Q(\FRAME_MATCHER.i [27]), .C(clk32MHz), 
            .D(n2_adj_4545), .S(n3_adj_4546));   // verilog/coms.v(126[12] 293[6])
    SB_DFFSS \FRAME_MATCHER.i_i28  (.Q(\FRAME_MATCHER.i [28]), .C(clk32MHz), 
            .D(n2_adj_4494), .S(n3_adj_4547));   // verilog/coms.v(126[12] 293[6])
    SB_DFFSS \FRAME_MATCHER.i_i29  (.Q(\FRAME_MATCHER.i [29]), .C(clk32MHz), 
            .D(n2_adj_4493), .S(n3_adj_4548));   // verilog/coms.v(126[12] 293[6])
    SB_DFFSS \FRAME_MATCHER.i_i30  (.Q(\FRAME_MATCHER.i [30]), .C(clk32MHz), 
            .D(n2_adj_4492), .S(n3_adj_4549));   // verilog/coms.v(126[12] 293[6])
    SB_DFFSS \FRAME_MATCHER.i_i31  (.Q(\FRAME_MATCHER.i [31]), .C(clk32MHz), 
            .D(n2_adj_4484), .S(n3_adj_4550));   // verilog/coms.v(126[12] 293[6])
    SB_DFFE data_out_frame_0___i185 (.Q(\data_out_frame[23] [0]), .C(clk32MHz), 
            .E(n17308), .D(n33202));   // verilog/coms.v(126[12] 293[6])
    SB_LUT4 i13352_3_lut_4_lut (.I0(n8), .I1(n32952), .I2(rx_data[3]), 
            .I3(\data_in_frame[21] [3]), .O(n18181));
    defparam i13352_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13356_3_lut_4_lut (.I0(n8), .I1(n32952), .I2(rx_data[7]), 
            .I3(\data_in_frame[21] [7]), .O(n18185));
    defparam i13356_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_1144 (.I0(n16930), .I1(n34730), .I2(GND_net), 
            .I3(GND_net), .O(n33189));
    defparam i1_2_lut_adj_1144.LUT_INIT = 16'h9999;
    SB_LUT4 i11_4_lut_adj_1145 (.I0(n21_adj_4491), .I1(n17_adj_4490), .I2(n30968), 
            .I3(\data_out_frame[19] [5]), .O(n24_adj_4551));
    defparam i11_4_lut_adj_1145.LUT_INIT = 16'h6996;
    SB_LUT4 i12_4_lut_adj_1146 (.I0(\data_out_frame[17] [5]), .I1(n24_adj_4551), 
            .I2(n20_adj_4552), .I3(\data_out_frame[18] [4]), .O(n30192));
    defparam i12_4_lut_adj_1146.LUT_INIT = 16'h6996;
    SB_DFFE data_out_frame_0___i186 (.Q(\data_out_frame[23] [1]), .C(clk32MHz), 
            .E(n17308), .D(n35248));   // verilog/coms.v(126[12] 293[6])
    SB_LUT4 i4_4_lut_adj_1147 (.I0(n33357), .I1(n33310), .I2(n33421), 
            .I3(n6_adj_4553), .O(n33430));   // verilog/coms.v(70[16:27])
    defparam i4_4_lut_adj_1147.LUT_INIT = 16'h6996;
    SB_LUT4 i10_4_lut_adj_1148 (.I0(\data_out_frame[20] [6]), .I1(n33514), 
            .I2(n33228), .I3(\data_out_frame[19] [0]), .O(n28_adj_4554));
    defparam i10_4_lut_adj_1148.LUT_INIT = 16'h6996;
    SB_DFFE data_out_frame_0___i187 (.Q(\data_out_frame[23] [2]), .C(clk32MHz), 
            .E(n17308), .D(n34864));   // verilog/coms.v(126[12] 293[6])
    SB_DFFE data_out_frame_0___i188 (.Q(\data_out_frame[23] [3]), .C(clk32MHz), 
            .E(n17308), .D(n34374));   // verilog/coms.v(126[12] 293[6])
    SB_DFFE data_out_frame_0___i189 (.Q(\data_out_frame[23] [4]), .C(clk32MHz), 
            .E(n17308), .D(n34501));   // verilog/coms.v(126[12] 293[6])
    SB_DFFE data_out_frame_0___i190 (.Q(\data_out_frame[23] [5]), .C(clk32MHz), 
            .E(n17308), .D(n34502));   // verilog/coms.v(126[12] 293[6])
    SB_DFFE data_out_frame_0___i192 (.Q(\data_out_frame[23] [7]), .C(clk32MHz), 
            .E(n17308), .D(n34130));   // verilog/coms.v(126[12] 293[6])
    SB_DFFE data_out_frame_0___i193 (.Q(\data_out_frame[24] [0]), .C(clk32MHz), 
            .E(n17308), .D(n16291));   // verilog/coms.v(126[12] 293[6])
    SB_DFFE data_out_frame_0___i194 (.Q(\data_out_frame[24] [1]), .C(clk32MHz), 
            .E(n17308), .D(n30231));   // verilog/coms.v(126[12] 293[6])
    SB_DFFE data_out_frame_0___i195 (.Q(\data_out_frame[24] [2]), .C(clk32MHz), 
            .E(n17308), .D(n34495));   // verilog/coms.v(126[12] 293[6])
    SB_DFFE data_out_frame_0___i196 (.Q(\data_out_frame[24] [3]), .C(clk32MHz), 
            .E(n17308), .D(n32999));   // verilog/coms.v(126[12] 293[6])
    SB_DFFE data_out_frame_0___i197 (.Q(\data_out_frame[24] [4]), .C(clk32MHz), 
            .E(n17308), .D(n33169));   // verilog/coms.v(126[12] 293[6])
    SB_DFFE data_out_frame_0___i198 (.Q(\data_out_frame[24] [5]), .C(clk32MHz), 
            .E(n17308), .D(n35254));   // verilog/coms.v(126[12] 293[6])
    SB_DFFE data_out_frame_0___i199 (.Q(\data_out_frame[24] [6]), .C(clk32MHz), 
            .E(n17308), .D(n34522));   // verilog/coms.v(126[12] 293[6])
    SB_DFFE data_out_frame_0___i200 (.Q(\data_out_frame[24] [7]), .C(clk32MHz), 
            .E(n17308), .D(n35212));   // verilog/coms.v(126[12] 293[6])
    SB_DFFSS \FRAME_MATCHER.state_i3  (.Q(\FRAME_MATCHER.state [3]), .C(clk32MHz), 
            .D(n32183), .S(n32109));   // verilog/coms.v(126[12] 293[6])
    SB_LUT4 i1_2_lut_adj_1149 (.I0(\data_in_frame[19] [2]), .I1(n33269), 
            .I2(GND_net), .I3(GND_net), .O(n33480));
    defparam i1_2_lut_adj_1149.LUT_INIT = 16'h6666;
    SB_LUT4 i1_4_lut_adj_1150 (.I0(\data_in_frame[19] [7]), .I1(n16740), 
            .I2(n33564), .I3(n33171), .O(n5_adj_4555));   // verilog/coms.v(84[17:28])
    defparam i1_4_lut_adj_1150.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1151 (.I0(n5_adj_4555), .I1(n33480), .I2(\data_in_frame[19] [3]), 
            .I3(n33430), .O(n16930));   // verilog/coms.v(84[17:28])
    defparam i3_4_lut_adj_1151.LUT_INIT = 16'h6996;
    SB_DFFSS \FRAME_MATCHER.state_i4  (.Q(\FRAME_MATCHER.state [4]), .C(clk32MHz), 
            .D(n24102), .S(n24819));   // verilog/coms.v(126[12] 293[6])
    SB_DFFSS \FRAME_MATCHER.state_i5  (.Q(\FRAME_MATCHER.state [5]), .C(clk32MHz), 
            .D(n32277), .S(n32241));   // verilog/coms.v(126[12] 293[6])
    SB_DFFSS \FRAME_MATCHER.state_i6  (.Q(\FRAME_MATCHER.state [6]), .C(clk32MHz), 
            .D(n32279), .S(n32239));   // verilog/coms.v(126[12] 293[6])
    SB_DFFSS \FRAME_MATCHER.state_i7  (.Q(\FRAME_MATCHER.state [7]), .C(clk32MHz), 
            .D(n7_adj_4556), .S(n8_adj_4557));   // verilog/coms.v(126[12] 293[6])
    SB_DFFSS \FRAME_MATCHER.state_i8  (.Q(\FRAME_MATCHER.state [8]), .C(clk32MHz), 
            .D(n24104), .S(n24821));   // verilog/coms.v(126[12] 293[6])
    SB_DFFSS \FRAME_MATCHER.state_i9  (.Q(\FRAME_MATCHER.state [9]), .C(clk32MHz), 
            .D(n24106), .S(n32113));   // verilog/coms.v(126[12] 293[6])
    SB_DFFSS \FRAME_MATCHER.state_i10  (.Q(\FRAME_MATCHER.state [10]), .C(clk32MHz), 
            .D(n24108), .S(n32117));   // verilog/coms.v(126[12] 293[6])
    SB_DFFSS \FRAME_MATCHER.state_i11  (.Q(\FRAME_MATCHER.state [11]), .C(clk32MHz), 
            .D(n32281), .S(n32237));   // verilog/coms.v(126[12] 293[6])
    SB_DFFSS \FRAME_MATCHER.state_i12  (.Q(\FRAME_MATCHER.state [12]), .C(clk32MHz), 
            .D(n32283), .S(n32149));   // verilog/coms.v(126[12] 293[6])
    SB_DFFSS \FRAME_MATCHER.state_i13  (.Q(\FRAME_MATCHER.state [13]), .C(clk32MHz), 
            .D(n32285), .S(n32235));   // verilog/coms.v(126[12] 293[6])
    SB_DFFSS \FRAME_MATCHER.state_i14  (.Q(\FRAME_MATCHER.state [14]), .C(clk32MHz), 
            .D(n32287), .S(n32233));   // verilog/coms.v(126[12] 293[6])
    SB_DFFSS \FRAME_MATCHER.state_i15  (.Q(\FRAME_MATCHER.state [15]), .C(clk32MHz), 
            .D(n32289), .S(n32231));   // verilog/coms.v(126[12] 293[6])
    SB_DFFSS \FRAME_MATCHER.state_i16  (.Q(\FRAME_MATCHER.state [16]), .C(clk32MHz), 
            .D(n32291), .S(n32229));   // verilog/coms.v(126[12] 293[6])
    SB_DFFSS \FRAME_MATCHER.state_i17  (.Q(\FRAME_MATCHER.state [17]), .C(clk32MHz), 
            .D(n24110), .S(n24823));   // verilog/coms.v(126[12] 293[6])
    SB_DFFSS \FRAME_MATCHER.state_i18  (.Q(\FRAME_MATCHER.state [18]), .C(clk32MHz), 
            .D(n32275), .S(n32181));   // verilog/coms.v(126[12] 293[6])
    SB_DFFSS \FRAME_MATCHER.state_i19  (.Q(\FRAME_MATCHER.state [19]), .C(clk32MHz), 
            .D(n32185), .S(n32161));   // verilog/coms.v(126[12] 293[6])
    SB_DFFSS \FRAME_MATCHER.state_i20  (.Q(\FRAME_MATCHER.state [20]), .C(clk32MHz), 
            .D(n24112), .S(n24825));   // verilog/coms.v(126[12] 293[6])
    SB_DFFSS \FRAME_MATCHER.state_i21  (.Q(\FRAME_MATCHER.state [21]), .C(clk32MHz), 
            .D(n32293), .S(n32227));   // verilog/coms.v(126[12] 293[6])
    SB_DFFSS \FRAME_MATCHER.state_i22  (.Q(\FRAME_MATCHER.state [22]), .C(clk32MHz), 
            .D(n32295), .S(n32225));   // verilog/coms.v(126[12] 293[6])
    SB_DFFSS \FRAME_MATCHER.state_i23  (.Q(\FRAME_MATCHER.state [23]), .C(clk32MHz), 
            .D(n29601), .S(n29605));   // verilog/coms.v(126[12] 293[6])
    SB_DFFSS \FRAME_MATCHER.state_i24  (.Q(\FRAME_MATCHER.state [24]), .C(clk32MHz), 
            .D(n32297), .S(n32223));   // verilog/coms.v(126[12] 293[6])
    SB_DFFSS \FRAME_MATCHER.state_i25  (.Q(\FRAME_MATCHER.state [25]), .C(clk32MHz), 
            .D(n32299), .S(n32221));   // verilog/coms.v(126[12] 293[6])
    SB_DFFSS \FRAME_MATCHER.state_i26  (.Q(\FRAME_MATCHER.state [26]), .C(clk32MHz), 
            .D(n32301), .S(n32219));   // verilog/coms.v(126[12] 293[6])
    SB_DFFSS \FRAME_MATCHER.state_i27  (.Q(\FRAME_MATCHER.state [27]), .C(clk32MHz), 
            .D(n32171), .S(n29611));   // verilog/coms.v(126[12] 293[6])
    SB_DFFSS \FRAME_MATCHER.state_i28  (.Q(\FRAME_MATCHER.state [28]), .C(clk32MHz), 
            .D(n32273), .S(n32271));   // verilog/coms.v(126[12] 293[6])
    SB_DFFSS \FRAME_MATCHER.state_i29  (.Q(\FRAME_MATCHER.state [29]), .C(clk32MHz), 
            .D(n32173), .S(n29609));   // verilog/coms.v(126[12] 293[6])
    SB_DFFSS \FRAME_MATCHER.state_i30  (.Q(\FRAME_MATCHER.state [30]), .C(clk32MHz), 
            .D(n32175), .S(n29613));   // verilog/coms.v(126[12] 293[6])
    SB_DFFSS \FRAME_MATCHER.state_i31  (.Q(\FRAME_MATCHER.state [31]), .C(clk32MHz), 
            .D(n32179), .S(n29607));   // verilog/coms.v(126[12] 293[6])
    SB_LUT4 i14_3_lut (.I0(\data_out_frame[16] [7]), .I1(n28_adj_4554), 
            .I2(n30968), .I3(GND_net), .O(n32_adj_4558));
    defparam i14_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 i13355_3_lut_4_lut (.I0(n8), .I1(n32952), .I2(rx_data[6]), 
            .I3(\data_in_frame[21] [6]), .O(n18184));
    defparam i13355_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13354_3_lut_4_lut (.I0(n8), .I1(n32952), .I2(rx_data[5]), 
            .I3(\data_in_frame[21] [5]), .O(n18183));
    defparam i13354_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 equal_132_i8_2_lut_3_lut (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(\FRAME_MATCHER.i [0]), .I3(GND_net), .O(n8));   // verilog/coms.v(153[7:23])
    defparam equal_132_i8_2_lut_3_lut.LUT_INIT = 16'hbfbf;
    SB_LUT4 equal_133_i8_2_lut_3_lut (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(\FRAME_MATCHER.i [0]), .I3(GND_net), .O(n8_adj_4353));   // verilog/coms.v(153[7:23])
    defparam equal_133_i8_2_lut_3_lut.LUT_INIT = 16'hfbfb;
    SB_LUT4 i12_4_lut_adj_1152 (.I0(\data_out_frame[20] [4]), .I1(n33511), 
            .I2(n33570), .I3(n33442), .O(n30_adj_4559));
    defparam i12_4_lut_adj_1152.LUT_INIT = 16'h6996;
    SB_LUT4 i13_4_lut_adj_1153 (.I0(n33195), .I1(n34672), .I2(n33168), 
            .I3(\data_out_frame[14] [5]), .O(n31_adj_4560));
    defparam i13_4_lut_adj_1153.LUT_INIT = 16'h9669;
    SB_LUT4 i11_4_lut_adj_1154 (.I0(n33616), .I1(n33175), .I2(n33467), 
            .I3(\data_out_frame[18] [7]), .O(n29_adj_4561));
    defparam i11_4_lut_adj_1154.LUT_INIT = 16'h6996;
    SB_DFFESR driver_enable_3433 (.Q(PIN_11_c), .C(clk32MHz), .E(n33781), 
            .D(n5034), .R(n34073));   // verilog/coms.v(126[12] 293[6])
    SB_DFF data_in_0___i16 (.Q(\data_in[1] [7]), .C(clk32MHz), .D(n17805));   // verilog/coms.v(126[12] 293[6])
    SB_LUT4 i13309_3_lut_4_lut (.I0(n8_adj_4463), .I1(n32952), .I2(rx_data[0]), 
            .I3(\data_in_frame[16] [0]), .O(n18138));
    defparam i13309_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i17_4_lut_adj_1155 (.I0(n29_adj_4561), .I1(n31_adj_4560), .I2(n30_adj_4559), 
            .I3(n32_adj_4558), .O(n34726));
    defparam i17_4_lut_adj_1155.LUT_INIT = 16'h6996;
    SB_LUT4 i13310_3_lut_4_lut (.I0(n8_adj_4463), .I1(n32952), .I2(rx_data[1]), 
            .I3(\data_in_frame[16] [1]), .O(n18139));
    defparam i13310_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13311_3_lut_4_lut (.I0(n8_adj_4463), .I1(n32952), .I2(rx_data[2]), 
            .I3(\data_in_frame[16] [2]), .O(n18140));
    defparam i13311_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i3_4_lut_adj_1156 (.I0(n34726), .I1(n33198), .I2(n30192), 
            .I3(n16477), .O(n34130));
    defparam i3_4_lut_adj_1156.LUT_INIT = 16'h6996;
    SB_LUT4 i13312_3_lut_4_lut (.I0(n8_adj_4463), .I1(n32952), .I2(rx_data[3]), 
            .I3(\data_in_frame[16] [3]), .O(n18141));
    defparam i13312_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13200_3_lut_4_lut (.I0(n8_adj_4435), .I1(n32959), .I2(rx_data[3]), 
            .I3(\data_in_frame[2] [3]), .O(n18029));
    defparam i13200_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_2_lut_3_lut_4_lut (.I0(\data_in_frame[3] [7]), .I1(\data_in_frame[3] [6]), 
            .I2(\data_in_frame[4] [0]), .I3(\data_in_frame[6] [3]), .O(n10));   // verilog/coms.v(72[16:42])
    defparam i2_2_lut_3_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1157 (.I0(n33198), .I1(n33273), .I2(\data_out_frame[19] [3]), 
            .I3(GND_net), .O(n34502));
    defparam i2_3_lut_adj_1157.LUT_INIT = 16'h9696;
    SB_LUT4 i13313_3_lut_4_lut (.I0(n8_adj_4463), .I1(n32952), .I2(rx_data[4]), 
            .I3(\data_in_frame[16] [4]), .O(n18142));
    defparam i13313_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13201_3_lut_4_lut (.I0(n8_adj_4435), .I1(n32959), .I2(rx_data[4]), 
            .I3(\data_in_frame[2] [4]), .O(n18030));
    defparam i13201_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i9_4_lut_adj_1158 (.I0(n17_adj_4489), .I1(\data_in_frame[3] [0]), 
            .I2(n16_adj_4488), .I3(\data_in_frame[2] [6]), .O(Kp_23__N_996));   // verilog/coms.v(74[16:43])
    defparam i9_4_lut_adj_1158.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1159 (.I0(\data_out_frame[19] [1]), .I1(n30899), 
            .I2(GND_net), .I3(GND_net), .O(n33273));
    defparam i1_2_lut_adj_1159.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_4_lut_adj_1160 (.I0(\data_in_frame[2] [0]), .I1(\data_in_frame[2] [1]), 
            .I2(\data_in_frame[4] [2]), .I3(\data_in_frame[0] [0]), .O(n32982));   // verilog/coms.v(72[16:42])
    defparam i2_3_lut_4_lut_adj_1160.LUT_INIT = 16'h6996;
    SB_LUT4 i13202_3_lut_4_lut (.I0(n8_adj_4435), .I1(n32959), .I2(rx_data[5]), 
            .I3(\data_in_frame[2] [5]), .O(n18031));
    defparam i13202_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i8_4_lut_adj_1161 (.I0(n33081), .I1(n16855), .I2(\data_in_frame[7] [6]), 
            .I3(n33397), .O(n20_adj_4562));   // verilog/coms.v(84[17:28])
    defparam i8_4_lut_adj_1161.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1162 (.I0(\data_in_frame[5] [1]), .I1(Kp_23__N_996), 
            .I2(GND_net), .I3(GND_net), .O(n33259));   // verilog/coms.v(78[16:35])
    defparam i1_2_lut_adj_1162.LUT_INIT = 16'h6666;
    SB_LUT4 i7_4_lut_adj_1163 (.I0(\data_in_frame[19] [1]), .I1(n33464), 
            .I2(n33039), .I3(n16335), .O(n19));   // verilog/coms.v(84[17:28])
    defparam i7_4_lut_adj_1163.LUT_INIT = 16'h6996;
    SB_LUT4 i9_4_lut_adj_1164 (.I0(n33045), .I1(\data_in_frame[8] [1]), 
            .I2(\data_in_frame[17] [0]), .I3(\data_in_frame[18] [7]), .O(n21_adj_4563));   // verilog/coms.v(84[17:28])
    defparam i9_4_lut_adj_1164.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_1165 (.I0(n33552), .I1(n33148), .I2(n31287), 
            .I3(n33613), .O(n10_adj_4564));
    defparam i4_4_lut_adj_1165.LUT_INIT = 16'h6996;
    SB_LUT4 i13314_3_lut_4_lut (.I0(n8_adj_4463), .I1(n32952), .I2(rx_data[5]), 
            .I3(\data_in_frame[16] [5]), .O(n18143));
    defparam i13314_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13315_3_lut_4_lut (.I0(n8_adj_4463), .I1(n32952), .I2(rx_data[6]), 
            .I3(\data_in_frame[16] [6]), .O(n18144));
    defparam i13315_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_3_lut_adj_1166 (.I0(n33127), .I1(\data_in_frame[10] [4]), 
            .I2(Kp_23__N_1046), .I3(GND_net), .O(n6_adj_4565));   // verilog/coms.v(84[17:28])
    defparam i1_2_lut_3_lut_adj_1166.LUT_INIT = 16'h9696;
    SB_LUT4 i2_4_lut_adj_1167 (.I0(\data_out_frame[19] [2]), .I1(n33273), 
            .I2(n9_adj_4566), .I3(n10_adj_4564), .O(n34501));
    defparam i2_4_lut_adj_1167.LUT_INIT = 16'h9669;
    SB_LUT4 i2_3_lut_4_lut_adj_1168 (.I0(n30900), .I1(\data_in_frame[4] [7]), 
            .I2(\data_in_frame[7] [3]), .I3(\data_in_frame[7] [4]), .O(n33500));
    defparam i2_3_lut_4_lut_adj_1168.LUT_INIT = 16'h6996;
    SB_LUT4 i13316_3_lut_4_lut (.I0(n8_adj_4463), .I1(n32952), .I2(rx_data[7]), 
            .I3(\data_in_frame[16] [7]), .O(n18145));
    defparam i13316_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_1169 (.I0(n16570), .I1(\data_out_frame[18] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n33613));
    defparam i1_2_lut_adj_1169.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1170 (.I0(\data_out_frame[19] [1]), .I1(\data_out_frame[18] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n33183));
    defparam i1_2_lut_adj_1170.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_4_lut_adj_1171 (.I0(\data_out_frame[17] [2]), .I1(n14584), 
            .I2(n34236), .I3(n4_adj_4567), .O(n33198));
    defparam i1_2_lut_4_lut_adj_1171.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_4_lut_adj_1172 (.I0(\data_out_frame[17] [2]), .I1(n14584), 
            .I2(n34236), .I3(\data_out_frame[19] [4]), .O(n4));
    defparam i1_2_lut_4_lut_adj_1172.LUT_INIT = 16'h9669;
    SB_LUT4 i6_4_lut_adj_1173 (.I0(n33183), .I1(n31287), .I2(n33613), 
            .I3(n33567), .O(n16_adj_4569));
    defparam i6_4_lut_adj_1173.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_3_lut_adj_1174 (.I0(\data_in_frame[16] [3]), .I1(Kp_23__N_843), 
            .I2(n34730), .I3(GND_net), .O(n31235));
    defparam i1_2_lut_3_lut_adj_1174.LUT_INIT = 16'h6969;
    SB_CARRY add_41_30 (.CI(n27936), .I0(\FRAME_MATCHER.i [28]), .I1(GND_net), 
            .CO(n27937));
    SB_LUT4 add_41_29_lut (.I0(n2290), .I1(\FRAME_MATCHER.i [27]), .I2(GND_net), 
            .I3(n27935), .O(n2_adj_4545)) /* synthesis syn_instantiated=1 */ ;
    defparam add_41_29_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i2_3_lut_4_lut_adj_1175 (.I0(\data_in_frame[1] [3]), .I1(\data_in_frame[1] [5]), 
            .I2(\data_in_frame[3] [6]), .I3(\data_in_frame[3] [5]), .O(Kp_23__N_1046));   // verilog/coms.v(95[12:25])
    defparam i2_3_lut_4_lut_adj_1175.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_1176 (.I0(\data_in_frame[1] [3]), .I1(\data_in_frame[1] [5]), 
            .I2(\data_in_frame[1] [7]), .I3(n16347), .O(n33406));   // verilog/coms.v(95[12:25])
    defparam i2_3_lut_4_lut_adj_1176.LUT_INIT = 16'h6996;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_4_i16_3_lut (.I0(\data_out_frame[16] [4]), 
            .I1(\data_out_frame[17] [4]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n16_adj_4570));   // verilog/coms.v(105[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_4_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF data_in_0___i15 (.Q(\data_in[1] [6]), .C(clk32MHz), .D(n17804));   // verilog/coms.v(126[12] 293[6])
    SB_DFF data_in_0___i14 (.Q(\data_in[1] [5]), .C(clk32MHz), .D(n17803));   // verilog/coms.v(126[12] 293[6])
    SB_LUT4 i27193_2_lut_3_lut (.I0(\FRAME_MATCHER.state [2]), .I1(n25118), 
            .I2(\FRAME_MATCHER.state [0]), .I3(GND_net), .O(n33789));
    defparam i27193_2_lut_3_lut.LUT_INIT = 16'hfefe;
    SB_DFF data_in_0___i13 (.Q(\data_in[1] [4]), .C(clk32MHz), .D(n17802));   // verilog/coms.v(126[12] 293[6])
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_4_i17_3_lut (.I0(\data_out_frame[18] [4]), 
            .I1(\data_out_frame[19] [4]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n17_adj_4571));   // verilog/coms.v(105[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_4_i17_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF data_in_0___i12 (.Q(\data_in[1] [3]), .C(clk32MHz), .D(n17801));   // verilog/coms.v(126[12] 293[6])
    SB_DFF data_in_0___i11 (.Q(\data_in[1] [2]), .C(clk32MHz), .D(n17800));   // verilog/coms.v(126[12] 293[6])
    SB_DFF data_in_0___i10 (.Q(\data_in[1] [1]), .C(clk32MHz), .D(n17799));   // verilog/coms.v(126[12] 293[6])
    SB_DFF data_in_0___i9 (.Q(\data_in[1] [0]), .C(clk32MHz), .D(n17798));   // verilog/coms.v(126[12] 293[6])
    SB_DFF data_in_0___i8 (.Q(\data_in[0][7] ), .C(clk32MHz), .D(n17797));   // verilog/coms.v(126[12] 293[6])
    SB_DFF data_in_0___i7 (.Q(\data_in[0][6] ), .C(clk32MHz), .D(n17796));   // verilog/coms.v(126[12] 293[6])
    SB_DFF data_in_0___i6 (.Q(\data_in[0][5] ), .C(clk32MHz), .D(n17795));   // verilog/coms.v(126[12] 293[6])
    SB_DFF data_in_0___i5 (.Q(\data_in[0][4] ), .C(clk32MHz), .D(n17794));   // verilog/coms.v(126[12] 293[6])
    SB_LUT4 i3_3_lut_4_lut_adj_1177 (.I0(\FRAME_MATCHER.state [2]), .I1(n25118), 
            .I2(\FRAME_MATCHER.state [3]), .I3(n13554), .O(n17308));
    defparam i3_3_lut_4_lut_adj_1177.LUT_INIT = 16'h0010;
    SB_DFF data_in_0___i4 (.Q(\data_in[0][3] ), .C(clk32MHz), .D(n17793));   // verilog/coms.v(126[12] 293[6])
    SB_DFF data_in_0___i3 (.Q(\data_in[0] [2]), .C(clk32MHz), .D(n17792));   // verilog/coms.v(126[12] 293[6])
    SB_DFF data_in_0___i2 (.Q(\data_in[0][1] ), .C(clk32MHz), .D(n17791));   // verilog/coms.v(126[12] 293[6])
    SB_DFF IntegralLimit_i0_i23 (.Q(IntegralLimit[23]), .C(clk32MHz), .D(n17790));   // verilog/coms.v(126[12] 293[6])
    SB_DFF IntegralLimit_i0_i22 (.Q(IntegralLimit[22]), .C(clk32MHz), .D(n17789));   // verilog/coms.v(126[12] 293[6])
    SB_LUT4 i30858_2_lut (.I0(\data_out_frame[23] [4]), .I1(byte_transmit_counter[0]), 
            .I2(GND_net), .I3(GND_net), .O(n37274));
    defparam i30858_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i30840_2_lut (.I0(\data_out_frame[20] [4]), .I1(byte_transmit_counter[0]), 
            .I2(GND_net), .I3(GND_net), .O(n37273));
    defparam i30840_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i13325_3_lut_4_lut (.I0(n8_adj_4435), .I1(n32952), .I2(rx_data[0]), 
            .I3(\data_in_frame[18] [0]), .O(n18154));
    defparam i13325_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13326_3_lut_4_lut (.I0(n8_adj_4435), .I1(n32952), .I2(rx_data[1]), 
            .I3(\data_in_frame[18] [1]), .O(n18155));
    defparam i13326_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13327_3_lut_4_lut (.I0(n8_adj_4435), .I1(n32952), .I2(rx_data[2]), 
            .I3(\data_in_frame[18] [2]), .O(n18156));
    defparam i13327_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13328_3_lut_4_lut (.I0(n8_adj_4435), .I1(n32952), .I2(rx_data[3]), 
            .I3(\data_in_frame[18] [3]), .O(n18157));
    defparam i13328_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13236_3_lut_4_lut (.I0(n8_adj_4355), .I1(n32959), .I2(rx_data[7]), 
            .I3(\data_in_frame[6] [7]), .O(n18065));
    defparam i13236_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i7_4_lut_adj_1178 (.I0(n31295), .I1(n33580), .I2(n33616), 
            .I3(n33448), .O(n17_adj_4572));
    defparam i7_4_lut_adj_1178.LUT_INIT = 16'h9669;
    SB_LUT4 i9_4_lut_adj_1179 (.I0(n17_adj_4572), .I1(n33158), .I2(n16_adj_4569), 
            .I3(n31178), .O(n34374));
    defparam i9_4_lut_adj_1179.LUT_INIT = 16'h9669;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_2_i16_3_lut (.I0(\data_out_frame[16] [2]), 
            .I1(\data_out_frame[17] [2]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n16_adj_4573));   // verilog/coms.v(105[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_2_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2_3_lut_adj_1180 (.I0(n16647), .I1(n33244), .I2(\data_out_frame[19] [0]), 
            .I3(GND_net), .O(n34864));
    defparam i2_3_lut_adj_1180.LUT_INIT = 16'h6969;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_2_i17_3_lut (.I0(\data_out_frame[18] [2]), 
            .I1(\data_out_frame[19] [2]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n17_adj_4574));   // verilog/coms.v(105[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_2_i17_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i30867_2_lut (.I0(\data_out_frame[23] [2]), .I1(byte_transmit_counter[0]), 
            .I2(GND_net), .I3(GND_net), .O(n37268));
    defparam i30867_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i30958_2_lut (.I0(\data_out_frame[20] [2]), .I1(byte_transmit_counter[0]), 
            .I2(GND_net), .I3(GND_net), .O(n37267));
    defparam i30958_2_lut.LUT_INIT = 16'h2222;
    SB_DFF IntegralLimit_i0_i21 (.Q(IntegralLimit[21]), .C(clk32MHz), .D(n17788));   // verilog/coms.v(126[12] 293[6])
    SB_LUT4 i1_2_lut_adj_1181 (.I0(\data_out_frame[14] [5]), .I1(\data_out_frame[14] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n33451));
    defparam i1_2_lut_adj_1181.LUT_INIT = 16'h6666;
    SB_DFF IntegralLimit_i0_i20 (.Q(IntegralLimit[20]), .C(clk32MHz), .D(n17787));   // verilog/coms.v(126[12] 293[6])
    SB_DFF IntegralLimit_i0_i19 (.Q(IntegralLimit[19]), .C(clk32MHz), .D(n17786));   // verilog/coms.v(126[12] 293[6])
    SB_LUT4 i1_2_lut_4_lut_adj_1182 (.I0(n16954), .I1(n16679), .I2(n16661), 
            .I3(\data_out_frame[19] [7]), .O(n6_adj_4433));   // verilog/coms.v(77[16:27])
    defparam i1_2_lut_4_lut_adj_1182.LUT_INIT = 16'h6996;
    SB_DFF IntegralLimit_i0_i18 (.Q(IntegralLimit[18]), .C(clk32MHz), .D(n17785));   // verilog/coms.v(126[12] 293[6])
    SB_DFF data_in_frame_0__i91 (.Q(\data_in_frame[11] [2]), .C(clk32MHz), 
           .D(n18100));   // verilog/coms.v(126[12] 293[6])
    SB_DFF IntegralLimit_i0_i17 (.Q(IntegralLimit[17]), .C(clk32MHz), .D(n17784));   // verilog/coms.v(126[12] 293[6])
    SB_DFF IntegralLimit_i0_i16 (.Q(IntegralLimit[16]), .C(clk32MHz), .D(n17783));   // verilog/coms.v(126[12] 293[6])
    SB_LUT4 i5_2_lut_4_lut (.I0(n34691), .I1(\data_in_frame[18] [4]), .I2(n17081), 
            .I3(\data_in_frame[17] [6]), .O(n19_adj_4575));
    defparam i5_2_lut_4_lut.LUT_INIT = 16'h9669;
    SB_DFF IntegralLimit_i0_i15 (.Q(IntegralLimit[15]), .C(clk32MHz), .D(n17782));   // verilog/coms.v(126[12] 293[6])
    SB_DFF IntegralLimit_i0_i14 (.Q(IntegralLimit[14]), .C(clk32MHz), .D(n17781));   // verilog/coms.v(126[12] 293[6])
    SB_DFF IntegralLimit_i0_i13 (.Q(IntegralLimit[13]), .C(clk32MHz), .D(n17780));   // verilog/coms.v(126[12] 293[6])
    SB_LUT4 i11_3_lut (.I0(n21_adj_4563), .I1(n19), .I2(n20_adj_4562), 
            .I3(GND_net), .O(n33269));   // verilog/coms.v(84[17:28])
    defparam i11_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1183 (.I0(n16304), .I1(\data_out_frame[12] [6]), 
            .I2(\data_out_frame[15] [0]), .I3(GND_net), .O(n33374));
    defparam i1_2_lut_3_lut_adj_1183.LUT_INIT = 16'h9696;
    SB_DFF IntegralLimit_i0_i12 (.Q(IntegralLimit[12]), .C(clk32MHz), .D(n17779));   // verilog/coms.v(126[12] 293[6])
    SB_LUT4 i3_4_lut_adj_1184 (.I0(\data_in_frame[5] [5]), .I1(n33094), 
            .I2(\data_in_frame[1] [2]), .I3(\data_in_frame[3] [4]), .O(n16335));   // verilog/coms.v(95[12:25])
    defparam i3_4_lut_adj_1184.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_1185 (.I0(n7_adj_4460), .I1(n34691), .I2(n31257), 
            .I3(Kp_23__N_1662), .O(n33471));
    defparam i4_4_lut_adj_1185.LUT_INIT = 16'h6996;
    SB_DFF IntegralLimit_i0_i11 (.Q(IntegralLimit[11]), .C(clk32MHz), .D(n17778));   // verilog/coms.v(126[12] 293[6])
    SB_DFF data_in_frame_0__i90 (.Q(\data_in_frame[11] [1]), .C(clk32MHz), 
           .D(n18099));   // verilog/coms.v(126[12] 293[6])
    SB_LUT4 i4_4_lut_adj_1186 (.I0(n33595), .I1(n33503), .I2(\data_in_frame[13] [5]), 
            .I3(n33628), .O(n10_adj_4458));
    defparam i4_4_lut_adj_1186.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_1187 (.I0(\data_in_frame[1] [2]), .I1(\data_in_frame[1] [1]), 
            .I2(\data_in_frame[3] [3]), .I3(\data_in_frame[0] [7]), .O(n33354));   // verilog/coms.v(72[16:34])
    defparam i2_3_lut_4_lut_adj_1187.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1188 (.I0(n33063), .I1(\data_out_frame[12] [1]), 
            .I2(\data_out_frame[11] [7]), .I3(GND_net), .O(n33436));
    defparam i2_3_lut_adj_1188.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_4_lut_adj_1189 (.I0(\data_out_frame[11] [5]), .I1(n33576), 
            .I2(\data_out_frame[9] [5]), .I3(n33115), .O(n33394));
    defparam i2_3_lut_4_lut_adj_1189.LUT_INIT = 16'h6996;
    SB_LUT4 i13203_3_lut_4_lut (.I0(n8_adj_4435), .I1(n32959), .I2(rx_data[6]), 
            .I3(\data_in_frame[2] [6]), .O(n18032));
    defparam i13203_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1190 (.I0(\data_out_frame[5] [0]), .I1(\data_out_frame[6] [7]), 
            .I2(\data_out_frame[7] [1]), .I3(\data_out_frame[7] [2]), .O(n16880));   // verilog/coms.v(84[17:70])
    defparam i1_2_lut_3_lut_4_lut_adj_1190.LUT_INIT = 16'h6996;
    SB_LUT4 i13329_3_lut_4_lut (.I0(n8_adj_4435), .I1(n32952), .I2(rx_data[4]), 
            .I3(\data_in_frame[18] [4]), .O(n18158));
    defparam i13329_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13330_3_lut_4_lut (.I0(n8_adj_4435), .I1(n32952), .I2(rx_data[5]), 
            .I3(\data_in_frame[18] [5]), .O(n18159));
    defparam i13330_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_CARRY add_41_29 (.CI(n27935), .I0(\FRAME_MATCHER.i [27]), .I1(GND_net), 
            .CO(n27936));
    SB_LUT4 add_41_28_lut (.I0(n2290), .I1(\FRAME_MATCHER.i [26]), .I2(GND_net), 
            .I3(n27934), .O(n2_adj_4543)) /* synthesis syn_instantiated=1 */ ;
    defparam add_41_28_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i1_2_lut_3_lut_adj_1191 (.I0(\data_out_frame[11] [7]), .I1(n33066), 
            .I2(\data_out_frame[14] [1]), .I3(GND_net), .O(n33576));
    defparam i1_2_lut_3_lut_adj_1191.LUT_INIT = 16'h9696;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_31665 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[10] [0]), .I2(\data_out_frame[11] [0]), 
            .I3(byte_transmit_counter_c[1]), .O(n38351));
    defparam byte_transmit_counter_0__bdd_4_lut_31665.LUT_INIT = 16'he4aa;
    SB_CARRY add_41_28 (.CI(n27934), .I0(\FRAME_MATCHER.i [26]), .I1(GND_net), 
            .CO(n27935));
    SB_DFF data_in_frame_0__i89 (.Q(\data_in_frame[11] [0]), .C(clk32MHz), 
           .D(n18098));   // verilog/coms.v(126[12] 293[6])
    SB_DFF data_in_frame_0__i88 (.Q(\data_in_frame[10] [7]), .C(clk32MHz), 
           .D(n18097));   // verilog/coms.v(126[12] 293[6])
    SB_DFF data_in_frame_0__i87 (.Q(\data_in_frame[10] [6]), .C(clk32MHz), 
           .D(n18096));   // verilog/coms.v(126[12] 293[6])
    SB_DFF data_in_frame_0__i86 (.Q(\data_in_frame[10] [5]), .C(clk32MHz), 
           .D(n18095));   // verilog/coms.v(126[12] 293[6])
    SB_DFF data_in_frame_0__i85 (.Q(\data_in_frame[10] [4]), .C(clk32MHz), 
           .D(n18094));   // verilog/coms.v(126[12] 293[6])
    SB_DFF data_in_frame_0__i84 (.Q(\data_in_frame[10] [3]), .C(clk32MHz), 
           .D(n18093));   // verilog/coms.v(126[12] 293[6])
    SB_DFFESR LED_3432 (.Q(LED_c), .C(clk32MHz), .E(n33636), .D(n17449), 
            .R(n35075));   // verilog/coms.v(126[12] 293[6])
    SB_LUT4 n38351_bdd_4_lut (.I0(n38351), .I1(\data_out_frame[9] [0]), 
            .I2(\data_out_frame[8] [0]), .I3(byte_transmit_counter_c[1]), 
            .O(n38354));
    defparam n38351_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i20002_2_lut_3_lut_4_lut (.I0(n98), .I1(n1_c), .I2(n136), 
            .I3(\FRAME_MATCHER.state [4]), .O(n24819));
    defparam i20002_2_lut_3_lut_4_lut.LUT_INIT = 16'hfe00;
    SB_LUT4 add_41_27_lut (.I0(n2290), .I1(\FRAME_MATCHER.i [25]), .I2(GND_net), 
            .I3(n27933), .O(n2_adj_4541)) /* synthesis syn_instantiated=1 */ ;
    defparam add_41_27_lut.LUT_INIT = 16'h8228;
    SB_DFF data_in_frame_0__i83 (.Q(\data_in_frame[10] [2]), .C(clk32MHz), 
           .D(n18092));   // verilog/coms.v(126[12] 293[6])
    SB_LUT4 i13331_3_lut_4_lut (.I0(n8_adj_4435), .I1(n32952), .I2(rx_data[6]), 
            .I3(\data_in_frame[18] [6]), .O(n18160));
    defparam i13331_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_CARRY add_41_27 (.CI(n27933), .I0(\FRAME_MATCHER.i [25]), .I1(GND_net), 
            .CO(n27934));
    SB_LUT4 add_41_26_lut (.I0(n2290), .I1(\FRAME_MATCHER.i [24]), .I2(GND_net), 
            .I3(n27932), .O(n2_adj_4539)) /* synthesis syn_instantiated=1 */ ;
    defparam add_41_26_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_41_26 (.CI(n27932), .I0(\FRAME_MATCHER.i [24]), .I1(GND_net), 
            .CO(n27933));
    SB_LUT4 i13204_3_lut_4_lut (.I0(n8_adj_4435), .I1(n32959), .I2(rx_data[7]), 
            .I3(\data_in_frame[2] [7]), .O(n18033));
    defparam i13204_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13332_3_lut_4_lut (.I0(n8_adj_4435), .I1(n32952), .I2(rx_data[7]), 
            .I3(\data_in_frame[18] [7]), .O(n18161));
    defparam i13332_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF data_in_frame_0__i82 (.Q(\data_in_frame[10] [1]), .C(clk32MHz), 
           .D(n18091));   // verilog/coms.v(126[12] 293[6])
    SB_DFF data_in_frame_0__i149 (.Q(\data_in_frame[18] [4]), .C(clk32MHz), 
           .D(n18158));   // verilog/coms.v(126[12] 293[6])
    SB_DFF IntegralLimit_i0_i10 (.Q(IntegralLimit[10]), .C(clk32MHz), .D(n17777));   // verilog/coms.v(126[12] 293[6])
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1192 (.I0(n98), .I1(n1_c), .I2(n136), 
            .I3(\FRAME_MATCHER.state [7]), .O(n8_adj_4557));
    defparam i1_2_lut_3_lut_4_lut_adj_1192.LUT_INIT = 16'hfe00;
    SB_LUT4 i2_2_lut_3_lut (.I0(\data_out_frame[10] [7]), .I1(\data_out_frame[10] [6]), 
            .I2(n33265), .I3(GND_net), .O(n22));   // verilog/coms.v(70[16:27])
    defparam i2_2_lut_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 i4_4_lut_adj_1193 (.I0(\data_out_frame[12] [5]), .I1(n31249), 
            .I2(n33436), .I3(n6_adj_4576), .O(n33023));
    defparam i4_4_lut_adj_1193.LUT_INIT = 16'h9669;
    SB_LUT4 i3_4_lut_adj_1194 (.I0(\data_out_frame[18] [7]), .I1(n33374), 
            .I2(n33023), .I3(n16746), .O(n30899));
    defparam i3_4_lut_adj_1194.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1195 (.I0(n31178), .I1(n31295), .I2(GND_net), 
            .I3(GND_net), .O(n31204));
    defparam i1_2_lut_adj_1195.LUT_INIT = 16'h9999;
    SB_LUT4 i20003_2_lut_3_lut_4_lut (.I0(n98), .I1(n1_c), .I2(n136), 
            .I3(\FRAME_MATCHER.state [8]), .O(n24821));
    defparam i20003_2_lut_3_lut_4_lut.LUT_INIT = 16'hfe00;
    SB_LUT4 i1_2_lut_3_lut_adj_1196 (.I0(\data_out_frame[10] [7]), .I1(\data_out_frame[10] [6]), 
            .I2(n33344), .I3(GND_net), .O(n14531));   // verilog/coms.v(70[16:27])
    defparam i1_2_lut_3_lut_adj_1196.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1197 (.I0(n98), .I1(n1_c), .I2(n136), 
            .I3(\FRAME_MATCHER.state [9]), .O(n32113));
    defparam i1_2_lut_3_lut_4_lut_adj_1197.LUT_INIT = 16'hfe00;
    SB_LUT4 i1_2_lut_adj_1198 (.I0(\data_out_frame[16] [7]), .I1(n33439), 
            .I2(GND_net), .I3(GND_net), .O(n4_adj_4567));   // verilog/coms.v(70[16:27])
    defparam i1_2_lut_adj_1198.LUT_INIT = 16'h6666;
    SB_DFF IntegralLimit_i0_i9 (.Q(IntegralLimit[9]), .C(clk32MHz), .D(n17776));   // verilog/coms.v(126[12] 293[6])
    SB_LUT4 i1_2_lut_adj_1199 (.I0(n31168), .I1(n31235), .I2(GND_net), 
            .I3(GND_net), .O(n33186));
    defparam i1_2_lut_adj_1199.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1200 (.I0(n16292), .I1(\data_in_frame[8] [4]), 
            .I2(\data_in_frame[15] [2]), .I3(n33121), .O(n10_adj_4398));   // verilog/coms.v(73[16:43])
    defparam i4_4_lut_adj_1200.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1201 (.I0(n98), .I1(n1_c), .I2(n136), 
            .I3(\FRAME_MATCHER.state [10]), .O(n32117));
    defparam i1_2_lut_3_lut_4_lut_adj_1201.LUT_INIT = 16'hfe00;
    SB_LUT4 i1_2_lut_adj_1202 (.I0(\data_in_frame[10] [6]), .I1(\data_in_frame[13] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n16292));   // verilog/coms.v(75[16:43])
    defparam i1_2_lut_adj_1202.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_1203 (.I0(\data_in_frame[8] [1]), .I1(n16262), 
            .I2(n16292), .I3(\data_in_frame[12] [7]), .O(n33409));   // verilog/coms.v(84[17:28])
    defparam i3_4_lut_adj_1203.LUT_INIT = 16'h6996;
    SB_LUT4 i20004_2_lut_3_lut_4_lut (.I0(n98), .I1(n1_c), .I2(n136), 
            .I3(\FRAME_MATCHER.state [17]), .O(n24823));
    defparam i20004_2_lut_3_lut_4_lut.LUT_INIT = 16'hfe00;
    SB_LUT4 i6_4_lut_adj_1204 (.I0(n16521), .I1(\data_out_frame[7] [3]), 
            .I2(n33368), .I3(\data_out_frame[7] [0]), .O(n16_adj_4577));
    defparam i6_4_lut_adj_1204.LUT_INIT = 16'h6996;
    SB_LUT4 i8_4_lut_adj_1205 (.I0(\data_in_frame[12] [5]), .I1(n33409), 
            .I2(\data_in_frame[7] [7]), .I3(n16335), .O(n20_adj_4578));   // verilog/coms.v(84[17:28])
    defparam i8_4_lut_adj_1205.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut_adj_1206 (.I0(\data_in_frame[17] [3]), .I1(\data_in_frame[15] [3]), 
            .I2(n33000), .I3(n16447), .O(n19_adj_4579));   // verilog/coms.v(84[17:28])
    defparam i7_4_lut_adj_1206.LUT_INIT = 16'h6996;
    SB_LUT4 i9_4_lut_adj_1207 (.I0(n33555), .I1(\data_in_frame[5] [7]), 
            .I2(n33118), .I3(\data_in_frame[10] [3]), .O(n21_adj_4580));   // verilog/coms.v(84[17:28])
    defparam i9_4_lut_adj_1207.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut_adj_1208 (.I0(\data_out_frame[8] [5]), .I1(\data_out_frame[8] [4]), 
            .I2(n33537), .I3(\data_out_frame[5] [3]), .O(n17_adj_4581));
    defparam i7_4_lut_adj_1208.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1209 (.I0(\data_in_frame[19] [5]), .I1(n21_adj_4580), 
            .I2(n19_adj_4579), .I3(n20_adj_4578), .O(n33171));
    defparam i1_4_lut_adj_1209.LUT_INIT = 16'h6996;
    SB_LUT4 add_41_25_lut (.I0(n2290), .I1(\FRAME_MATCHER.i [23]), .I2(GND_net), 
            .I3(n27931), .O(n2_adj_4537)) /* synthesis syn_instantiated=1 */ ;
    defparam add_41_25_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_41_25 (.CI(n27931), .I0(\FRAME_MATCHER.i [23]), .I1(GND_net), 
            .CO(n27932));
    SB_LUT4 i9_4_lut_adj_1210 (.I0(n17_adj_4581), .I1(n1301), .I2(n16_adj_4577), 
            .I3(\data_out_frame[7] [4]), .O(n34934));
    defparam i9_4_lut_adj_1210.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1211 (.I0(\data_out_frame[10] [7]), .I1(n34934), 
            .I2(GND_net), .I3(GND_net), .O(n17072));
    defparam i1_2_lut_adj_1211.LUT_INIT = 16'h9999;
    SB_LUT4 i12703_2_lut_3_lut_4_lut (.I0(n63), .I1(\FRAME_MATCHER.state [2]), 
            .I2(\FRAME_MATCHER.state [0]), .I3(n16153), .O(n17527));   // verilog/coms.v(126[12] 293[6])
    defparam i12703_2_lut_3_lut_4_lut.LUT_INIT = 16'h5515;
    SB_DFF data_in_frame_0__i148 (.Q(\data_in_frame[18] [3]), .C(clk32MHz), 
           .D(n18157));   // verilog/coms.v(126[12] 293[6])
    SB_LUT4 i20005_2_lut_3_lut_4_lut (.I0(n98), .I1(n1_c), .I2(n136), 
            .I3(\FRAME_MATCHER.state [20]), .O(n24825));
    defparam i20005_2_lut_3_lut_4_lut.LUT_INIT = 16'hfe00;
    SB_LUT4 i4_4_lut_adj_1212 (.I0(\data_in_frame[19] [6]), .I1(n33357), 
            .I2(Kp_23__N_860), .I3(\data_in_frame[17] [5]), .O(n10_adj_4582));   // verilog/coms.v(75[16:43])
    defparam i4_4_lut_adj_1212.LUT_INIT = 16'h6996;
    SB_LUT4 i5_3_lut_adj_1213 (.I0(n33000), .I1(n10_adj_4582), .I2(n16466), 
            .I3(GND_net), .O(n33564));   // verilog/coms.v(75[16:43])
    defparam i5_3_lut_adj_1213.LUT_INIT = 16'h9696;
    SB_LUT4 i2_2_lut_3_lut_4_lut_adj_1214 (.I0(\data_out_frame[7] [7]), .I1(n16304), 
            .I2(\data_out_frame[12] [6]), .I3(\data_out_frame[15] [0]), 
            .O(n10_adj_4415));   // verilog/coms.v(84[17:28])
    defparam i2_2_lut_3_lut_4_lut_adj_1214.LUT_INIT = 16'h6996;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_31655 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[10] [2]), .I2(\data_out_frame[11] [2]), 
            .I3(byte_transmit_counter_c[1]), .O(n38345));
    defparam byte_transmit_counter_0__bdd_4_lut_31655.LUT_INIT = 16'he4aa;
    SB_LUT4 n38345_bdd_4_lut (.I0(n38345), .I1(\data_out_frame[9] [2]), 
            .I2(\data_out_frame[8] [2]), .I3(byte_transmit_counter_c[1]), 
            .O(n38348));
    defparam n38345_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_31650 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[10] [3]), .I2(\data_out_frame[11] [3]), 
            .I3(byte_transmit_counter_c[1]), .O(n38339));
    defparam byte_transmit_counter_0__bdd_4_lut_31650.LUT_INIT = 16'he4aa;
    SB_LUT4 n38339_bdd_4_lut (.I0(n38339), .I1(\data_out_frame[9] [3]), 
            .I2(\data_out_frame[8] [3]), .I3(byte_transmit_counter_c[1]), 
            .O(n38342));
    defparam n38339_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_31689 (.I0(byte_transmit_counter_c[1]), 
            .I1(n37258), .I2(n37259), .I3(byte_transmit_counter_c[2]), 
            .O(n38333));
    defparam byte_transmit_counter_1__bdd_4_lut_31689.LUT_INIT = 16'he4aa;
    SB_LUT4 n38333_bdd_4_lut (.I0(n38333), .I1(n17_adj_4583), .I2(n16_adj_4584), 
            .I3(byte_transmit_counter_c[2]), .O(n38336));
    defparam n38333_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_31645 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[10] [4]), .I2(\data_out_frame[11] [4]), 
            .I3(byte_transmit_counter_c[1]), .O(n38327));
    defparam byte_transmit_counter_0__bdd_4_lut_31645.LUT_INIT = 16'he4aa;
    SB_LUT4 n38327_bdd_4_lut (.I0(n38327), .I1(\data_out_frame[9] [4]), 
            .I2(\data_out_frame[8] [4]), .I3(byte_transmit_counter_c[1]), 
            .O(n38330));
    defparam n38327_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_31635 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[10] [5]), .I2(\data_out_frame[11] [5]), 
            .I3(byte_transmit_counter_c[1]), .O(n38321));
    defparam byte_transmit_counter_0__bdd_4_lut_31635.LUT_INIT = 16'he4aa;
    SB_LUT4 n38321_bdd_4_lut (.I0(n38321), .I1(\data_out_frame[9] [5]), 
            .I2(\data_out_frame[8] [5]), .I3(byte_transmit_counter_c[1]), 
            .O(n38324));
    defparam n38321_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_31630 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[14] [5]), .I2(\data_out_frame[15] [5]), 
            .I3(byte_transmit_counter_c[1]), .O(n38315));
    defparam byte_transmit_counter_0__bdd_4_lut_31630.LUT_INIT = 16'he4aa;
    SB_LUT4 n38315_bdd_4_lut (.I0(n38315), .I1(\data_out_frame[13] [5]), 
            .I2(\data_out_frame[12] [5]), .I3(byte_transmit_counter_c[1]), 
            .O(n38318));
    defparam n38315_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF data_in_frame_0__i147 (.Q(\data_in_frame[18] [2]), .C(clk32MHz), 
           .D(n18156));   // verilog/coms.v(126[12] 293[6])
    SB_DFF data_in_frame_0__i146 (.Q(\data_in_frame[18] [1]), .C(clk32MHz), 
           .D(n18155));   // verilog/coms.v(126[12] 293[6])
    SB_LUT4 i2_3_lut_4_lut_adj_1215 (.I0(\data_out_frame[9] [0]), .I1(\data_out_frame[8] [7]), 
            .I2(\data_out_frame[8] [6]), .I3(n16350), .O(n33517));
    defparam i2_3_lut_4_lut_adj_1215.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1216 (.I0(n16447), .I1(n16862), .I2(\data_in_frame[15] [4]), 
            .I3(GND_net), .O(n16740));   // verilog/coms.v(74[16:43])
    defparam i2_3_lut_adj_1216.LUT_INIT = 16'h9696;
    SB_LUT4 i7_4_lut_adj_1217 (.I0(n17072), .I1(n1251), .I2(n33110), .I3(\data_out_frame[7] [2]), 
            .O(n18_adj_4585));
    defparam i7_4_lut_adj_1217.LUT_INIT = 16'h6996;
    SB_LUT4 add_41_24_lut (.I0(n2290), .I1(\FRAME_MATCHER.i [22]), .I2(GND_net), 
            .I3(n27930), .O(n2_adj_4535)) /* synthesis syn_instantiated=1 */ ;
    defparam add_41_24_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_41_24 (.CI(n27930), .I0(\FRAME_MATCHER.i [22]), .I1(GND_net), 
            .CO(n27931));
    SB_LUT4 add_41_23_lut (.I0(n2290), .I1(\FRAME_MATCHER.i [21]), .I2(GND_net), 
            .I3(n27929), .O(n2_adj_4533)) /* synthesis syn_instantiated=1 */ ;
    defparam add_41_23_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i1_2_lut_3_lut_adj_1218 (.I0(\data_in_frame[13] [4]), .I1(\data_in_frame[13] [5]), 
            .I2(\data_in_frame[15] [6]), .I3(GND_net), .O(n16248));   // verilog/coms.v(73[16:43])
    defparam i1_2_lut_3_lut_adj_1218.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_4_lut_adj_1219 (.I0(\data_in_frame[7] [0]), .I1(\data_in_frame[4] [6]), 
            .I2(\data_in_frame[9] [1]), .I3(Kp_23__N_993), .O(n33054));   // verilog/coms.v(70[16:27])
    defparam i2_3_lut_4_lut_adj_1219.LUT_INIT = 16'h6996;
    SB_CARRY add_41_23 (.CI(n27929), .I0(\FRAME_MATCHER.i [21]), .I1(GND_net), 
            .CO(n27930));
    SB_LUT4 i2_3_lut_4_lut_adj_1220 (.I0(\data_in_frame[6] [6]), .I1(n16722), 
            .I2(\data_in_frame[6] [4]), .I3(\data_in_frame[11] [2]), .O(n33414));   // verilog/coms.v(73[16:43])
    defparam i2_3_lut_4_lut_adj_1220.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_adj_1221 (.I0(\data_in_frame[1] [6]), .I1(n16242), 
            .I2(\data_in_frame[4] [2]), .I3(\data_in_frame[0] [0]), .O(n16722));   // verilog/coms.v(72[16:42])
    defparam i1_2_lut_4_lut_adj_1221.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_1222 (.I0(n16746), .I1(n34982), .I2(\data_out_frame[18] [5]), 
            .I3(n33192), .O(n33020));
    defparam i2_3_lut_4_lut_adj_1222.LUT_INIT = 16'h9669;
    SB_LUT4 i9_4_lut_adj_1223 (.I0(n15783), .I1(n18_adj_4585), .I2(\data_out_frame[9] [1]), 
            .I3(n33341), .O(n20_adj_4586));
    defparam i9_4_lut_adj_1223.LUT_INIT = 16'h6996;
    SB_LUT4 add_41_22_lut (.I0(n2290), .I1(\FRAME_MATCHER.i [20]), .I2(GND_net), 
            .I3(n27928), .O(n2_adj_4531)) /* synthesis syn_instantiated=1 */ ;
    defparam add_41_22_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i1_2_lut_3_lut_adj_1224 (.I0(\data_out_frame[18] [4]), .I1(n34982), 
            .I2(n16711), .I3(GND_net), .O(n33371));
    defparam i1_2_lut_3_lut_adj_1224.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1225 (.I0(\data_out_frame[5] [6]), .I1(\data_out_frame[6] [0]), 
            .I2(\data_out_frame[5] [7]), .I3(\data_out_frame[8] [3]), .O(n33368));   // verilog/coms.v(84[17:28])
    defparam i1_2_lut_3_lut_4_lut_adj_1225.LUT_INIT = 16'h6996;
    SB_LUT4 i3_3_lut_4_lut_3_lut (.I0(\FRAME_MATCHER.state [0]), .I1(\FRAME_MATCHER.state [1]), 
            .I2(\FRAME_MATCHER.state [2]), .I3(GND_net), .O(n33634));   // verilog/coms.v(144[4] 292[11])
    defparam i3_3_lut_4_lut_3_lut.LUT_INIT = 16'habab;
    SB_LUT4 i1_2_lut_4_lut_adj_1226 (.I0(\data_in_frame[9] [0]), .I1(\data_in_frame[11] [1]), 
            .I2(n17169), .I3(n33151), .O(n6_adj_4587));   // verilog/coms.v(70[16:27])
    defparam i1_2_lut_4_lut_adj_1226.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1227 (.I0(n16722), .I1(\data_in_frame[6] [4]), 
            .I2(n16380), .I3(GND_net), .O(n16840));   // verilog/coms.v(75[16:43])
    defparam i1_2_lut_3_lut_adj_1227.LUT_INIT = 16'h9696;
    SB_LUT4 i10_4_lut_adj_1228 (.I0(n33115), .I1(n20_adj_4586), .I2(n16_adj_4588), 
            .I3(n33107), .O(n34996));
    defparam i10_4_lut_adj_1228.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1229 (.I0(Kp_23__N_993), .I1(Kp_23__N_996), 
            .I2(\data_in_frame[7] [1]), .I3(GND_net), .O(n33003));
    defparam i1_2_lut_3_lut_adj_1229.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_4_lut_adj_1230 (.I0(n16380), .I1(n16384), .I2(\data_in_frame[6] [5]), 
            .I3(n33388), .O(n6_adj_4589));   // verilog/coms.v(70[16:27])
    defparam i1_2_lut_4_lut_adj_1230.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1231 (.I0(\data_out_frame[7] [6]), .I1(\data_out_frame[9] [5]), 
            .I2(n33115), .I3(GND_net), .O(n6_adj_4590));   // verilog/coms.v(84[17:63])
    defparam i1_2_lut_3_lut_adj_1231.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1232 (.I0(\data_out_frame[16] [6]), .I1(\data_out_frame[18] [7]), 
            .I2(\data_out_frame[18] [6]), .I3(GND_net), .O(n6_adj_4591));
    defparam i1_2_lut_3_lut_adj_1232.LUT_INIT = 16'h9696;
    SB_LUT4 i19285_2_lut_3_lut (.I0(n24810), .I1(rx_data_ready), .I2(\FRAME_MATCHER.rx_data_ready_prev ), 
            .I3(GND_net), .O(n24089));
    defparam i19285_2_lut_3_lut.LUT_INIT = 16'h0404;
    SB_DFF data_in_frame_0__i145 (.Q(\data_in_frame[18] [0]), .C(clk32MHz), 
           .D(n18154));   // verilog/coms.v(126[12] 293[6])
    SB_DFF data_in_frame_0__i144 (.Q(\data_in_frame[17] [7]), .C(clk32MHz), 
           .D(n18153));   // verilog/coms.v(126[12] 293[6])
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_1_i16_3_lut (.I0(\data_out_frame[16] [1]), 
            .I1(\data_out_frame[17] [1]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n16_adj_4584));   // verilog/coms.v(105[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_1_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_1_i17_3_lut (.I0(\data_out_frame[18] [1]), 
            .I1(\data_out_frame[19] [1]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n17_adj_4583));   // verilog/coms.v(105[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_1_i17_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_3_lut_adj_1233 (.I0(\FRAME_MATCHER.state [2]), .I1(\FRAME_MATCHER.state [0]), 
            .I2(n16158), .I3(GND_net), .O(n16161));   // verilog/coms.v(218[5:21])
    defparam i1_2_lut_3_lut_adj_1233.LUT_INIT = 16'hf7f7;
    SB_LUT4 i30870_2_lut (.I0(\data_out_frame[23] [1]), .I1(byte_transmit_counter[0]), 
            .I2(GND_net), .I3(GND_net), .O(n37259));
    defparam i30870_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i3_4_lut_adj_1234 (.I0(\data_in_frame[17] [6]), .I1(n16248), 
            .I2(n30930), .I3(n17132), .O(n33323));
    defparam i3_4_lut_adj_1234.LUT_INIT = 16'h6996;
    SB_LUT4 i30959_2_lut (.I0(\data_out_frame[20] [1]), .I1(byte_transmit_counter[0]), 
            .I2(GND_net), .I3(GND_net), .O(n37258));
    defparam i30959_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i1_2_lut_4_lut_adj_1235 (.I0(\data_in_frame[6] [0]), .I1(\data_in_frame[10] [5]), 
            .I2(\data_in_frame[15] [1]), .I3(\data_in_frame[14] [7]), .O(n33118));   // verilog/coms.v(84[17:28])
    defparam i1_2_lut_4_lut_adj_1235.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1236 (.I0(\data_in_frame[13] [1]), .I1(n33151), 
            .I2(n33090), .I3(n16840), .O(n33421));   // verilog/coms.v(70[16:27])
    defparam i3_4_lut_adj_1236.LUT_INIT = 16'h6996;
    SB_CARRY add_41_22 (.CI(n27928), .I0(\FRAME_MATCHER.i [20]), .I1(GND_net), 
            .CO(n27929));
    SB_LUT4 i1_2_lut_adj_1237 (.I0(\data_in_frame[17] [5]), .I1(\data_in_frame[15] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n17042));
    defparam i1_2_lut_adj_1237.LUT_INIT = 16'h6666;
    SB_LUT4 i13261_3_lut_4_lut (.I0(n8_adj_4435), .I1(n32937), .I2(rx_data[0]), 
            .I3(\data_in_frame[10] [0]), .O(n18090));
    defparam i13261_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_3_lut_4_lut_adj_1238 (.I0(\data_out_frame[7] [0]), .I1(\data_out_frame[6] [7]), 
            .I2(n33537), .I3(n16536), .O(n33341));
    defparam i2_3_lut_4_lut_adj_1238.LUT_INIT = 16'h6996;
    SB_LUT4 i2_2_lut_4_lut_adj_1239 (.I0(n30900), .I1(\data_in_frame[5] [1]), 
            .I2(n17157), .I3(\data_in_frame[7] [1]), .O(n7_adj_4592));
    defparam i2_2_lut_4_lut_adj_1239.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1240 (.I0(\data_in_frame[18] [0]), .I1(n30438), 
            .I2(n31219), .I3(GND_net), .O(n17132));
    defparam i2_3_lut_adj_1240.LUT_INIT = 16'h9696;
    SB_LUT4 add_41_21_lut (.I0(n2290), .I1(\FRAME_MATCHER.i [19]), .I2(GND_net), 
            .I3(n27927), .O(n2_adj_4529)) /* synthesis syn_instantiated=1 */ ;
    defparam add_41_21_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i1_2_lut_4_lut_adj_1241 (.I0(n33505), .I1(n33598), .I2(n35345), 
            .I3(n16626), .O(Kp_23__N_843));
    defparam i1_2_lut_4_lut_adj_1241.LUT_INIT = 16'h9669;
    SB_LUT4 i2_3_lut_4_lut_adj_1242 (.I0(\data_out_frame[8] [7]), .I1(\data_out_frame[6] [5]), 
            .I2(\data_out_frame[7] [0]), .I3(\data_out_frame[6] [7]), .O(n1337));   // verilog/coms.v(70[16:27])
    defparam i2_3_lut_4_lut_adj_1242.LUT_INIT = 16'h6996;
    SB_LUT4 i5_2_lut_4_lut_adj_1243 (.I0(\data_out_frame[5] [0]), .I1(\data_out_frame[6] [7]), 
            .I2(n16521), .I3(\data_out_frame[11] [1]), .O(n16_adj_4588));
    defparam i5_2_lut_4_lut_adj_1243.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_adj_1244 (.I0(\data_in_frame[17] [4]), .I1(n16413), 
            .I2(n33421), .I3(\data_in_frame[12] [7]), .O(n33000));   // verilog/coms.v(75[16:43])
    defparam i1_2_lut_4_lut_adj_1244.LUT_INIT = 16'h6996;
    SB_CARRY add_41_21 (.CI(n27927), .I0(\FRAME_MATCHER.i [19]), .I1(GND_net), 
            .CO(n27928));
    SB_DFF data_in_frame_0__i143 (.Q(\data_in_frame[17] [6]), .C(clk32MHz), 
           .D(n18152));   // verilog/coms.v(126[12] 293[6])
    SB_DFF data_in_frame_0__i142 (.Q(\data_in_frame[17] [5]), .C(clk32MHz), 
           .D(n18151));   // verilog/coms.v(126[12] 293[6])
    SB_DFF data_in_frame_0__i141 (.Q(\data_in_frame[17] [4]), .C(clk32MHz), 
           .D(n18150));   // verilog/coms.v(126[12] 293[6])
    SB_DFF data_in_frame_0__i140 (.Q(\data_in_frame[17] [3]), .C(clk32MHz), 
           .D(n18149));   // verilog/coms.v(126[12] 293[6])
    SB_DFF data_in_frame_0__i81 (.Q(\data_in_frame[10] [0]), .C(clk32MHz), 
           .D(n18090));   // verilog/coms.v(126[12] 293[6])
    SB_DFF data_in_frame_0__i69 (.Q(\data_in_frame[8] [4]), .C(clk32MHz), 
           .D(n18078));   // verilog/coms.v(126[12] 293[6])
    SB_LUT4 i1_2_lut_3_lut_adj_1245 (.I0(\data_out_frame[16] [7]), .I1(n33439), 
            .I2(n33467), .I3(GND_net), .O(n33580));
    defparam i1_2_lut_3_lut_adj_1245.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_4_lut_adj_1246 (.I0(n31178), .I1(n31295), .I2(n30899), 
            .I3(\data_out_frame[20] [7]), .O(n33467));
    defparam i2_3_lut_4_lut_adj_1246.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1247 (.I0(\data_in_frame[1] [7]), .I1(\data_in_frame[1] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n33232));   // verilog/coms.v(71[16:41])
    defparam i1_2_lut_adj_1247.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_3_lut_adj_1248 (.I0(\data_out_frame[14] [7]), .I1(\data_out_frame[17] [1]), 
            .I2(n33567), .I3(GND_net), .O(n6_adj_4576));
    defparam i1_2_lut_3_lut_adj_1248.LUT_INIT = 16'h9696;
    SB_LUT4 i13262_3_lut_4_lut (.I0(n8_adj_4435), .I1(n32937), .I2(rx_data[1]), 
            .I3(\data_in_frame[10] [1]), .O(n18091));
    defparam i13262_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_1249 (.I0(\data_in_frame[11] [5]), .I1(\data_in_frame[9] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n33595));
    defparam i1_2_lut_adj_1249.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_4_lut_adj_1250 (.I0(\data_out_frame[14] [3]), .I1(\data_out_frame[16] [7]), 
            .I2(\data_out_frame[16] [6]), .I3(\data_out_frame[16] [5]), 
            .O(n33567));
    defparam i1_2_lut_4_lut_adj_1250.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1251 (.I0(n30900), .I1(\data_in_frame[5] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n31230));
    defparam i1_2_lut_adj_1251.LUT_INIT = 16'h6666;
    SB_DFF data_in_frame_0__i80 (.Q(\data_in_frame[9] [7]), .C(clk32MHz), 
           .D(n18089));   // verilog/coms.v(126[12] 293[6])
    SB_DFF IntegralLimit_i0_i8 (.Q(IntegralLimit[8]), .C(clk32MHz), .D(n17775));   // verilog/coms.v(126[12] 293[6])
    SB_LUT4 i4_4_lut_adj_1252 (.I0(n17126), .I1(n31230), .I2(n33320), 
            .I3(n6_adj_4409), .O(n31219));
    defparam i4_4_lut_adj_1252.LUT_INIT = 16'h9669;
    SB_LUT4 i4_4_lut_adj_1253 (.I0(n17072), .I1(\data_out_frame[15] [4]), 
            .I2(n31225), .I3(n6_adj_4432), .O(n33477));
    defparam i4_4_lut_adj_1253.LUT_INIT = 16'h6996;
    SB_LUT4 i3_2_lut_4_lut (.I0(\data_out_frame[16] [7]), .I1(\data_out_frame[16] [6]), 
            .I2(\data_out_frame[16] [5]), .I3(\data_out_frame[19] [0]), 
            .O(n9_adj_4566));
    defparam i3_2_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_adj_1254 (.I0(\data_out_frame[19] [1]), .I1(\data_out_frame[16] [4]), 
            .I2(\data_out_frame[14] [6]), .I3(\data_out_frame[17] [0]), 
            .O(n33148));
    defparam i1_2_lut_4_lut_adj_1254.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_adj_1255 (.I0(\data_in[1] [5]), .I1(n10_adj_4440), 
            .I2(\data_in[2] [2]), .I3(n158), .O(n22269));
    defparam i1_2_lut_4_lut_adj_1255.LUT_INIT = 16'hffdf;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_31625 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[14] [0]), .I2(\data_out_frame[15] [0]), 
            .I3(byte_transmit_counter_c[1]), .O(n38309));
    defparam byte_transmit_counter_0__bdd_4_lut_31625.LUT_INIT = 16'he4aa;
    SB_LUT4 i1_2_lut_4_lut_adj_1256 (.I0(\data_in[1] [5]), .I1(n10_adj_4440), 
            .I2(\data_in[2] [2]), .I3(n136_adj_4445), .O(n22275));
    defparam i1_2_lut_4_lut_adj_1256.LUT_INIT = 16'hffdf;
    SB_LUT4 i2_3_lut_adj_1257 (.I0(\data_in_frame[0] [2]), .I1(\data_in_frame[2] [4]), 
            .I2(\data_in_frame[0] [3]), .I3(GND_net), .O(n16816));   // verilog/coms.v(74[16:43])
    defparam i2_3_lut_adj_1257.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1258 (.I0(\data_out_frame[16] [4]), .I1(\data_out_frame[14] [6]), 
            .I2(\data_out_frame[17] [0]), .I3(GND_net), .O(n33424));
    defparam i1_2_lut_3_lut_adj_1258.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1259 (.I0(\data_in_frame[18] [7]), .I1(\data_in_frame[18] [6]), 
            .I2(n31196), .I3(GND_net), .O(n33445));
    defparam i1_2_lut_3_lut_adj_1259.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_adj_1260 (.I0(n33517), .I1(n33341), .I2(n33313), 
            .I3(GND_net), .O(n31225));
    defparam i2_3_lut_adj_1260.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1261 (.I0(\data_in_frame[0] [3]), .I1(\data_in_frame[0] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n33104));   // verilog/coms.v(75[16:43])
    defparam i1_2_lut_adj_1261.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1262 (.I0(n33595), .I1(\data_in_frame[9] [3]), 
            .I2(\data_in_frame[14] [1]), .I3(n33625), .O(n10_adj_4593));
    defparam i4_4_lut_adj_1262.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1263 (.I0(\data_in_frame[19] [4]), .I1(\data_in_frame[17] [2]), 
            .I2(\data_in_frame[17] [3]), .I3(GND_net), .O(n6_adj_4553));   // verilog/coms.v(70[16:27])
    defparam i1_2_lut_3_lut_adj_1263.LUT_INIT = 16'h9696;
    SB_LUT4 i5_4_lut_adj_1264 (.I0(n33505), .I1(n10_adj_4593), .I2(n7_adj_4592), 
            .I3(n8_adj_4408), .O(n16626));
    defparam i5_4_lut_adj_1264.LUT_INIT = 16'h9669;
    SB_LUT4 i2_3_lut_adj_1265 (.I0(n16626), .I1(n31219), .I2(\data_in_frame[11] [4]), 
            .I3(GND_net), .O(n33483));
    defparam i2_3_lut_adj_1265.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_adj_1266 (.I0(n33335), .I1(n33483), .I2(n33298), 
            .I3(GND_net), .O(n34691));
    defparam i2_3_lut_adj_1266.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1267 (.I0(\data_in_frame[17] [2]), .I1(\data_in_frame[17] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n16435));
    defparam i1_2_lut_adj_1267.LUT_INIT = 16'h6666;
    SB_DFF IntegralLimit_i0_i7 (.Q(IntegralLimit[7]), .C(clk32MHz), .D(n17774));   // verilog/coms.v(126[12] 293[6])
    SB_LUT4 i2_3_lut_adj_1268 (.I0(n33164), .I1(n33427), .I2(\data_out_frame[8] [6]), 
            .I3(GND_net), .O(n33057));   // verilog/coms.v(74[16:27])
    defparam i2_3_lut_adj_1268.LUT_INIT = 16'h9696;
    SB_DFF data_in_frame_0__i79 (.Q(\data_in_frame[9] [6]), .C(clk32MHz), 
           .D(n18088));   // verilog/coms.v(126[12] 293[6])
    SB_LUT4 i1_2_lut_adj_1269 (.I0(n30805), .I1(n31257), .I2(GND_net), 
            .I3(GND_net), .O(n16855));
    defparam i1_2_lut_adj_1269.LUT_INIT = 16'h6666;
    SB_LUT4 data_in_frame_18__7__I_0_3455_2_lut (.I0(\data_in_frame[18] [7]), 
            .I1(\data_in_frame[18] [6]), .I2(GND_net), .I3(GND_net), .O(Kp_23__N_1453));   // verilog/coms.v(77[16:27])
    defparam data_in_frame_18__7__I_0_3455_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i5_4_lut_adj_1270 (.I0(Kp_23__N_1046), .I1(\data_in_frame[12] [3]), 
            .I2(n33235), .I3(n16233), .O(n12_adj_4594));   // verilog/coms.v(84[17:28])
    defparam i5_4_lut_adj_1270.LUT_INIT = 16'h6996;
    SB_LUT4 i7_3_lut_4_lut (.I0(\data_out_frame[18] [0]), .I1(\data_out_frame[19] [1]), 
            .I2(\data_out_frame[18] [5]), .I3(n34236), .O(n20_adj_4552));
    defparam i7_3_lut_4_lut.LUT_INIT = 16'h9669;
    SB_LUT4 i3_3_lut_adj_1271 (.I0(n31228), .I1(n31196), .I2(n15781), 
            .I3(GND_net), .O(n11));
    defparam i3_3_lut_adj_1271.LUT_INIT = 16'h9696;
    SB_LUT4 i6_4_lut_adj_1272 (.I0(\data_in_frame[6] [0]), .I1(n12_adj_4594), 
            .I2(\data_in_frame[9] [7]), .I3(n16608), .O(n33036));   // verilog/coms.v(84[17:28])
    defparam i6_4_lut_adj_1272.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1273 (.I0(\data_in_frame[8] [6]), .I1(\data_in_frame[11] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n33090));   // verilog/coms.v(70[16:27])
    defparam i1_2_lut_adj_1273.LUT_INIT = 16'h6666;
    SB_LUT4 i5_4_lut_adj_1274 (.I0(\data_in_frame[8] [5]), .I1(n17036), 
            .I2(n16765), .I3(\data_in_frame[8] [4]), .O(n12_adj_4595));   // verilog/coms.v(70[16:27])
    defparam i5_4_lut_adj_1274.LUT_INIT = 16'h6996;
    SB_LUT4 add_41_20_lut (.I0(n2290), .I1(\FRAME_MATCHER.i [18]), .I2(GND_net), 
            .I3(n27926), .O(n2_adj_4527)) /* synthesis syn_instantiated=1 */ ;
    defparam add_41_20_lut.LUT_INIT = 16'h8228;
    SB_LUT4 add_3528_9_lut (.I0(byte_transmit_counter_c[7]), .I1(byte_transmit_counter_c[7]), 
            .I2(n25050), .I3(n28024), .O(n17656)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3528_9_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 i6_4_lut_adj_1275 (.I0(\data_in_frame[13] [2]), .I1(n12_adj_4595), 
            .I2(n33090), .I3(\data_in_frame[10] [6]), .O(n33010));   // verilog/coms.v(70[16:27])
    defparam i6_4_lut_adj_1275.LUT_INIT = 16'h6996;
    SB_LUT4 add_3528_8_lut (.I0(byte_transmit_counter_c[6]), .I1(byte_transmit_counter_c[6]), 
            .I2(n25050), .I3(n28023), .O(n17659)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3528_8_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 i2_2_lut_adj_1276 (.I0(\FRAME_MATCHER.state [2]), .I1(\FRAME_MATCHER.state [0]), 
            .I2(GND_net), .I3(GND_net), .O(n24786));   // verilog/coms.v(144[4] 292[11])
    defparam i2_2_lut_adj_1276.LUT_INIT = 16'h8888;
    SB_CARRY add_41_20 (.CI(n27926), .I0(\FRAME_MATCHER.i [18]), .I1(GND_net), 
            .CO(n27927));
    SB_LUT4 n38309_bdd_4_lut (.I0(n38309), .I1(\data_out_frame[13] [0]), 
            .I2(\data_out_frame[12] [0]), .I3(byte_transmit_counter_c[1]), 
            .O(n38312));
    defparam n38309_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i5_3_lut_adj_1277 (.I0(\FRAME_MATCHER.state [27]), .I1(\FRAME_MATCHER.state [23]), 
            .I2(\FRAME_MATCHER.state [14]), .I3(GND_net), .O(n14_adj_4596));   // verilog/coms.v(126[12] 293[6])
    defparam i5_3_lut_adj_1277.LUT_INIT = 16'hfefe;
    SB_LUT4 i6_4_lut_adj_1278 (.I0(\FRAME_MATCHER.state [17]), .I1(\FRAME_MATCHER.state [18]), 
            .I2(\FRAME_MATCHER.state [24]), .I3(\FRAME_MATCHER.state [13]), 
            .O(n15_adj_4597));   // verilog/coms.v(126[12] 293[6])
    defparam i6_4_lut_adj_1278.LUT_INIT = 16'hfffe;
    SB_CARRY add_3528_8 (.CI(n28023), .I0(byte_transmit_counter_c[6]), .I1(n25050), 
            .CO(n28024));
    SB_LUT4 i1_2_lut_adj_1279 (.I0(\data_in_frame[15] [3]), .I1(\data_in_frame[15] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n33491));
    defparam i1_2_lut_adj_1279.LUT_INIT = 16'h6666;
    SB_LUT4 i2_2_lut_adj_1280 (.I0(\FRAME_MATCHER.state [8]), .I1(\FRAME_MATCHER.state [29]), 
            .I2(GND_net), .I3(GND_net), .O(n22_adj_4598));   // verilog/coms.v(227[5:23])
    defparam i2_2_lut_adj_1280.LUT_INIT = 16'heeee;
    SB_LUT4 i12_4_lut_adj_1281 (.I0(\FRAME_MATCHER.state [5]), .I1(\FRAME_MATCHER.state [30]), 
            .I2(\FRAME_MATCHER.state [19]), .I3(\FRAME_MATCHER.state [26]), 
            .O(n32_adj_4599));   // verilog/coms.v(227[5:23])
    defparam i12_4_lut_adj_1281.LUT_INIT = 16'hfffe;
    SB_LUT4 i8_4_lut_adj_1282 (.I0(n15_adj_4597), .I1(\FRAME_MATCHER.state [20]), 
            .I2(n14_adj_4596), .I3(\FRAME_MATCHER.state [31]), .O(n35349));   // verilog/coms.v(126[12] 293[6])
    defparam i8_4_lut_adj_1282.LUT_INIT = 16'hfffe;
    SB_LUT4 i16_4_lut_adj_1283 (.I0(n35349), .I1(n32_adj_4599), .I2(n22_adj_4598), 
            .I3(\FRAME_MATCHER.state [22]), .O(n36_adj_4600));   // verilog/coms.v(227[5:23])
    defparam i16_4_lut_adj_1283.LUT_INIT = 16'hfffe;
    SB_LUT4 i14_4_lut_adj_1284 (.I0(\FRAME_MATCHER.state [16]), .I1(\FRAME_MATCHER.state [4]), 
            .I2(\FRAME_MATCHER.state [11]), .I3(\FRAME_MATCHER.state [6]), 
            .O(n34_adj_4601));   // verilog/coms.v(227[5:23])
    defparam i14_4_lut_adj_1284.LUT_INIT = 16'hfffe;
    SB_LUT4 i15_4_lut_adj_1285 (.I0(\FRAME_MATCHER.state [21]), .I1(\FRAME_MATCHER.state [9]), 
            .I2(\FRAME_MATCHER.state [28]), .I3(\FRAME_MATCHER.state [15]), 
            .O(n35_adj_4602));   // verilog/coms.v(227[5:23])
    defparam i15_4_lut_adj_1285.LUT_INIT = 16'hfffe;
    SB_LUT4 i13_4_lut_adj_1286 (.I0(\FRAME_MATCHER.state [10]), .I1(\FRAME_MATCHER.state [25]), 
            .I2(\FRAME_MATCHER.state [12]), .I3(\FRAME_MATCHER.state [7]), 
            .O(n33_adj_4603));   // verilog/coms.v(227[5:23])
    defparam i13_4_lut_adj_1286.LUT_INIT = 16'hfffe;
    SB_LUT4 i19_4_lut_adj_1287 (.I0(n33_adj_4603), .I1(n35_adj_4602), .I2(n34_adj_4601), 
            .I3(n36_adj_4600), .O(n25118));   // verilog/coms.v(227[5:23])
    defparam i19_4_lut_adj_1287.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_adj_1288 (.I0(\FRAME_MATCHER.state [2]), .I1(\FRAME_MATCHER.state [0]), 
            .I2(GND_net), .I3(GND_net), .O(n16080));   // verilog/coms.v(247[5:25])
    defparam i1_2_lut_adj_1288.LUT_INIT = 16'hbbbb;
    SB_LUT4 i14_2_lut (.I0(rx_data_ready), .I1(\FRAME_MATCHER.rx_data_ready_prev ), 
            .I2(GND_net), .I3(GND_net), .O(n161));   // verilog/coms.v(152[9:50])
    defparam i14_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i2_4_lut_adj_1289 (.I0(n16161), .I1(n16080), .I2(\FRAME_MATCHER.state [3]), 
            .I3(n25118), .O(n24810));
    defparam i2_4_lut_adj_1289.LUT_INIT = 16'haaa8;
    SB_LUT4 i1_2_lut_3_lut_adj_1290 (.I0(\data_out_frame[13] [4]), .I1(\data_out_frame[13] [3]), 
            .I2(\data_out_frame[15] [5]), .I3(GND_net), .O(n33210));
    defparam i1_2_lut_3_lut_adj_1290.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_4_lut_adj_1291 (.I0(\data_in_frame[1] [4]), .I1(\data_in_frame[1] [6]), 
            .I2(\data_in_frame[1] [0]), .I3(n33406), .O(n16319));   // verilog/coms.v(69[16:27])
    defparam i1_2_lut_4_lut_adj_1291.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1292 (.I0(\FRAME_MATCHER.state [2]), .I1(\FRAME_MATCHER.state [0]), 
            .I2(n16158), .I3(GND_net), .O(n16159));   // verilog/coms.v(150[5:27])
    defparam i1_2_lut_3_lut_adj_1292.LUT_INIT = 16'hfbfb;
    SB_LUT4 i1_2_lut_adj_1293 (.I0(\data_in_frame[14] [6]), .I1(\data_in_frame[8] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n33607));   // verilog/coms.v(84[17:28])
    defparam i1_2_lut_adj_1293.LUT_INIT = 16'h6666;
    SB_DFF data_in_frame_0__i78 (.Q(\data_in_frame[9] [5]), .C(clk32MHz), 
           .D(n18087));   // verilog/coms.v(126[12] 293[6])
    SB_DFF data_in_frame_0__i77 (.Q(\data_in_frame[9] [4]), .C(clk32MHz), 
           .D(n18086));   // verilog/coms.v(126[12] 293[6])
    SB_DFF data_in_frame_0__i118 (.Q(\data_in_frame[14] [5]), .C(clk32MHz), 
           .D(n18127));   // verilog/coms.v(126[12] 293[6])
    SB_DFF data_in_frame_0__i76 (.Q(\data_in_frame[9] [3]), .C(clk32MHz), 
           .D(n18085));   // verilog/coms.v(126[12] 293[6])
    SB_LUT4 i4_4_lut_adj_1294 (.I0(\data_in_frame[10] [2]), .I1(\data_in_frame[12] [5]), 
            .I2(\data_in_frame[15] [5]), .I3(n33607), .O(n10_adj_4604));   // verilog/coms.v(84[17:28])
    defparam i4_4_lut_adj_1294.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_1295 (.I0(n33549), .I1(\data_out_frame[6] [6]), 
            .I2(n33057), .I3(\data_out_frame[8] [7]), .O(n14_adj_4605));
    defparam i6_4_lut_adj_1295.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut_adj_1296 (.I0(\data_out_frame[15] [3]), .I1(n14_adj_4605), 
            .I2(n10_adj_4606), .I3(n34934), .O(n30769));
    defparam i7_4_lut_adj_1296.LUT_INIT = 16'h9669;
    SB_LUT4 i13263_3_lut_4_lut (.I0(n8_adj_4435), .I1(n32937), .I2(rx_data[2]), 
            .I3(\data_in_frame[10] [2]), .O(n18092));
    defparam i13263_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i3_4_lut_adj_1297 (.I0(n16676), .I1(n33477), .I2(n1337), .I3(n34996), 
            .O(n16661));
    defparam i3_4_lut_adj_1297.LUT_INIT = 16'h9669;
    SB_LUT4 add_41_19_lut (.I0(n2290), .I1(\FRAME_MATCHER.i [17]), .I2(GND_net), 
            .I3(n27925), .O(n2_adj_4525)) /* synthesis syn_instantiated=1 */ ;
    defparam add_41_19_lut.LUT_INIT = 16'h8228;
    SB_LUT4 add_3528_7_lut (.I0(byte_transmit_counter_c[5]), .I1(byte_transmit_counter_c[5]), 
            .I2(n25050), .I3(n28022), .O(n17662)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3528_7_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 i13301_3_lut_4_lut (.I0(n24185), .I1(n32937), .I2(rx_data[0]), 
            .I3(\data_in_frame[15] [0]), .O(n18130));
    defparam i13301_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i13302_3_lut_4_lut (.I0(n24185), .I1(n32937), .I2(rx_data[1]), 
            .I3(\data_in_frame[15] [1]), .O(n18131));
    defparam i13302_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1225_2_lut (.I0(\data_out_frame[18] [7]), .I1(\data_out_frame[18] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n1981));   // verilog/coms.v(70[16:27])
    defparam i1225_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_31640 (.I0(byte_transmit_counter_c[1]), 
            .I1(n37267), .I2(n37268), .I3(byte_transmit_counter_c[2]), 
            .O(n38303));
    defparam byte_transmit_counter_1__bdd_4_lut_31640.LUT_INIT = 16'he4aa;
    SB_LUT4 i4_4_lut_adj_1298 (.I0(n33520), .I1(n33204), .I2(\data_out_frame[16] [1]), 
            .I3(n33601), .O(n10_adj_4607));
    defparam i4_4_lut_adj_1298.LUT_INIT = 16'h6996;
    SB_LUT4 n38303_bdd_4_lut (.I0(n38303), .I1(n17_adj_4574), .I2(n16_adj_4573), 
            .I3(byte_transmit_counter_c[2]), .O(n38306));
    defparam n38303_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i5_3_lut_adj_1299 (.I0(n33344), .I1(n10_adj_4607), .I2(n16672), 
            .I3(GND_net), .O(n16726));
    defparam i5_3_lut_adj_1299.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_4_lut_adj_1300 (.I0(n4_adj_4462), .I1(n12_adj_4464), 
            .I2(n14531), .I3(\data_out_frame[17] [3]), .O(n31178));
    defparam i1_2_lut_4_lut_adj_1300.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1301 (.I0(\data_out_frame[18] [4]), .I1(n16726), 
            .I2(\data_out_frame[18] [3]), .I3(n34982), .O(n31163));
    defparam i3_4_lut_adj_1301.LUT_INIT = 16'h9669;
    SB_LUT4 i2_3_lut_4_lut_adj_1302 (.I0(\data_out_frame[17] [7]), .I1(n16726), 
            .I2(n16954), .I3(\data_out_frame[18] [1]), .O(n33087));
    defparam i2_3_lut_4_lut_adj_1302.LUT_INIT = 16'h6996;
    SB_LUT4 i5_4_lut_adj_1303 (.I0(\data_in_frame[18] [7]), .I1(n33220), 
            .I2(n31235), .I3(n31257), .O(n13));
    defparam i5_4_lut_adj_1303.LUT_INIT = 16'h6996;
    SB_CARRY add_41_19 (.CI(n27925), .I0(\FRAME_MATCHER.i [17]), .I1(GND_net), 
            .CO(n27926));
    SB_CARRY add_3528_7 (.CI(n28022), .I0(byte_transmit_counter_c[5]), .I1(n25050), 
            .CO(n28023));
    SB_LUT4 i4_4_lut_adj_1304 (.I0(n33451), .I1(n33192), .I2(n16570), 
            .I3(n6_adj_4591), .O(n33244));
    defparam i4_4_lut_adj_1304.LUT_INIT = 16'h6996;
    SB_LUT4 add_3528_6_lut (.I0(byte_transmit_counter_c[4]), .I1(byte_transmit_counter_c[4]), 
            .I2(n25050), .I3(n28021), .O(n17665)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3528_6_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 i5_4_lut_adj_1305 (.I0(n33020), .I1(n33244), .I2(n31295), 
            .I3(n31163), .O(n12_adj_4608));
    defparam i5_4_lut_adj_1305.LUT_INIT = 16'h6996;
    SB_DFF data_in_frame_0__i75 (.Q(\data_in_frame[9] [2]), .C(clk32MHz), 
           .D(n18084));   // verilog/coms.v(126[12] 293[6])
    SB_DFF data_in_frame_0__i74 (.Q(\data_in_frame[9] [1]), .C(clk32MHz), 
           .D(n18083));   // verilog/coms.v(126[12] 293[6])
    SB_LUT4 add_41_18_lut (.I0(n2290), .I1(\FRAME_MATCHER.i [16]), .I2(GND_net), 
            .I3(n27924), .O(n2_adj_4523)) /* synthesis syn_instantiated=1 */ ;
    defparam add_41_18_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i6_4_lut_adj_1306 (.I0(\data_out_frame[20] [5]), .I1(n12_adj_4608), 
            .I2(n33580), .I3(n31178), .O(n35248));
    defparam i6_4_lut_adj_1306.LUT_INIT = 16'h9669;
    SB_CARRY add_3528_6 (.CI(n28021), .I0(byte_transmit_counter_c[4]), .I1(n25050), 
            .CO(n28022));
    SB_DFF data_in_frame_0__i73 (.Q(\data_in_frame[9] [0]), .C(clk32MHz), 
           .D(n18082));   // verilog/coms.v(126[12] 293[6])
    SB_CARRY add_41_18 (.CI(n27924), .I0(\FRAME_MATCHER.i [16]), .I1(GND_net), 
            .CO(n27925));
    SB_LUT4 i1_2_lut_adj_1307 (.I0(\data_in_frame[0] [1]), .I1(\data_in_frame[2] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n32989));   // verilog/coms.v(232[9:81])
    defparam i1_2_lut_adj_1307.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_4_lut_adj_1308 (.I0(\data_out_frame[20] [2]), .I1(n33303), 
            .I2(n10_adj_4416), .I3(n16975), .O(n33168));
    defparam i1_2_lut_4_lut_adj_1308.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1309 (.I0(n33104), .I1(n16816), .I2(\data_in_frame[2] [5]), 
            .I3(GND_net), .O(Kp_23__N_993));   // verilog/coms.v(75[16:43])
    defparam i2_3_lut_adj_1309.LUT_INIT = 16'h9696;
    SB_LUT4 i4_4_lut_adj_1310 (.I0(n16795), .I1(n16951), .I2(\data_out_frame[10] [0]), 
            .I3(n6_adj_4590), .O(n33063));   // verilog/coms.v(84[17:63])
    defparam i4_4_lut_adj_1310.LUT_INIT = 16'h6996;
    SB_LUT4 i5_3_lut_adj_1311 (.I0(n16791), .I1(n10_adj_4604), .I2(\data_in_frame[10] [4]), 
            .I3(GND_net), .O(n33039));   // verilog/coms.v(84[17:28])
    defparam i5_3_lut_adj_1311.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1312 (.I0(\data_in_frame[7] [2]), .I1(\data_in_frame[9] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n33320));
    defparam i1_2_lut_adj_1312.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1313 (.I0(\data_in_frame[6] [7]), .I1(n16834), 
            .I2(GND_net), .I3(GND_net), .O(n17126));
    defparam i1_2_lut_adj_1313.LUT_INIT = 16'h6666;
    SB_LUT4 i2_4_lut_adj_1314 (.I0(n16740), .I1(n33564), .I2(n33171), 
            .I3(\data_in_frame[21] [7]), .O(n35077));
    defparam i2_4_lut_adj_1314.LUT_INIT = 16'h6996;
    SB_LUT4 i13303_3_lut_4_lut (.I0(n24185), .I1(n32937), .I2(rx_data[2]), 
            .I3(\data_in_frame[15] [2]), .O(n18132));
    defparam i13303_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4_4_lut_adj_1315 (.I0(\data_in_frame[11] [4]), .I1(n33054), 
            .I2(n17126), .I3(n6_adj_4589), .O(n30438));   // verilog/coms.v(70[16:27])
    defparam i4_4_lut_adj_1315.LUT_INIT = 16'h6996;
    SB_LUT4 i13304_3_lut_4_lut (.I0(n24185), .I1(n32937), .I2(rx_data[3]), 
            .I3(\data_in_frame[15] [3]), .O(n18133));
    defparam i13304_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i2_3_lut_adj_1316 (.I0(\data_in_frame[15] [7]), .I1(n30438), 
            .I2(\data_in_frame[14] [0]), .I3(GND_net), .O(n33628));
    defparam i2_3_lut_adj_1316.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_4_lut_adj_1317 (.I0(n16608), .I1(\data_in_frame[7] [5]), 
            .I2(\data_in_frame[12] [0]), .I3(n16791), .O(n33631));
    defparam i2_3_lut_4_lut_adj_1317.LUT_INIT = 16'h6996;
    SB_LUT4 add_3528_5_lut (.I0(byte_transmit_counter_c[3]), .I1(byte_transmit_counter_c[3]), 
            .I2(n25050), .I3(n28020), .O(n17668)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3528_5_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 i13305_3_lut_4_lut (.I0(n24185), .I1(n32937), .I2(rx_data[4]), 
            .I3(\data_in_frame[15] [4]), .O(n18134));
    defparam i13305_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i2_3_lut_4_lut_adj_1318 (.I0(\data_in_frame[21] [3]), .I1(\data_in_frame[19] [2]), 
            .I2(n33269), .I3(n31228), .O(n34664));
    defparam i2_3_lut_4_lut_adj_1318.LUT_INIT = 16'h6996;
    SB_LUT4 i13306_3_lut_4_lut (.I0(n24185), .I1(n32937), .I2(rx_data[5]), 
            .I3(\data_in_frame[15] [5]), .O(n18135));
    defparam i13306_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i13307_3_lut_4_lut (.I0(n24185), .I1(n32937), .I2(rx_data[6]), 
            .I3(\data_in_frame[15] [6]), .O(n18136));
    defparam i13307_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1_2_lut_adj_1319 (.I0(\data_in_frame[16] [4]), .I1(\data_in_frame[16] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n17081));
    defparam i1_2_lut_adj_1319.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1320 (.I0(n33394), .I1(\data_out_frame[11] [6]), 
            .I2(\data_out_frame[16] [3]), .I3(n33552), .O(n10_adj_4405));
    defparam i4_4_lut_adj_1320.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_adj_1321 (.I0(\data_out_frame[6] [4]), .I1(\data_out_frame[6] [2]), 
            .I2(\data_out_frame[8] [4]), .I3(\data_out_frame[6] [3]), .O(n16350));
    defparam i1_2_lut_4_lut_adj_1321.LUT_INIT = 16'h6996;
    SB_LUT4 i2_2_lut_3_lut_adj_1322 (.I0(\data_out_frame[6] [2]), .I1(\data_out_frame[8] [4]), 
            .I2(\data_out_frame[6] [3]), .I3(GND_net), .O(n33110));   // verilog/coms.v(73[16:27])
    defparam i2_2_lut_3_lut_adj_1322.LUT_INIT = 16'h9696;
    SB_LUT4 i13308_3_lut_4_lut (.I0(n24185), .I1(n32937), .I2(rx_data[7]), 
            .I3(\data_in_frame[15] [7]), .O(n18137));
    defparam i13308_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1_2_lut_4_lut_adj_1323 (.I0(\data_out_frame[6] [4]), .I1(\data_out_frame[6] [3]), 
            .I2(\data_out_frame[8] [5]), .I3(n33223), .O(n33457));   // verilog/coms.v(70[16:27])
    defparam i1_2_lut_4_lut_adj_1323.LUT_INIT = 16'h6996;
    SB_LUT4 i2205_3_lut_4_lut (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(\FRAME_MATCHER.i [3]), .I3(\FRAME_MATCHER.i [4]), .O(n10_adj_4417));
    defparam i2205_3_lut_4_lut.LUT_INIT = 16'hf800;
    SB_LUT4 i19353_3_lut_4_lut (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(n15982), .I3(\FRAME_MATCHER.i [31]), .O(n3007));
    defparam i19353_3_lut_4_lut.LUT_INIT = 16'h00f8;
    SB_LUT4 i1_2_lut_3_lut_adj_1324 (.I0(\data_out_frame[6] [4]), .I1(\data_out_frame[6] [3]), 
            .I2(\data_out_frame[8] [5]), .I3(GND_net), .O(n16545));
    defparam i1_2_lut_3_lut_adj_1324.LUT_INIT = 16'h9696;
    SB_LUT4 equal_131_i8_2_lut_3_lut (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(\FRAME_MATCHER.i [0]), .I3(GND_net), .O(n8_adj_4355));
    defparam equal_131_i8_2_lut_3_lut.LUT_INIT = 16'hf7f7;
    SB_LUT4 i19375_2_lut_3_lut (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(\FRAME_MATCHER.i [0]), .I3(GND_net), .O(n24185));
    defparam i19375_2_lut_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 select_365_Select_31_i3_2_lut_4_lut (.I0(n24810), .I1(n16090), 
            .I2(n16158), .I3(\FRAME_MATCHER.i [31]), .O(n3_adj_4550));
    defparam select_365_Select_31_i3_2_lut_4_lut.LUT_INIT = 16'ha800;
    SB_LUT4 select_365_Select_30_i3_2_lut_4_lut (.I0(n24810), .I1(n16090), 
            .I2(n16158), .I3(\FRAME_MATCHER.i [30]), .O(n3_adj_4549));
    defparam select_365_Select_30_i3_2_lut_4_lut.LUT_INIT = 16'ha800;
    SB_LUT4 select_365_Select_29_i3_2_lut_4_lut (.I0(n24810), .I1(n16090), 
            .I2(n16158), .I3(\FRAME_MATCHER.i [29]), .O(n3_adj_4548));
    defparam select_365_Select_29_i3_2_lut_4_lut.LUT_INIT = 16'ha800;
    SB_LUT4 i2_3_lut_adj_1325 (.I0(n16765), .I1(\data_in_frame[8] [5]), 
            .I2(n16380), .I3(GND_net), .O(n33142));   // verilog/coms.v(73[16:43])
    defparam i2_3_lut_adj_1325.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_adj_1326 (.I0(n16380), .I1(n16384), .I2(\data_in_frame[6] [5]), 
            .I3(GND_net), .O(n16399));   // verilog/coms.v(70[16:27])
    defparam i2_3_lut_adj_1326.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_adj_1327 (.I0(\data_in_frame[6] [3]), .I1(n33142), 
            .I2(\data_in_frame[6] [4]), .I3(GND_net), .O(n16262));   // verilog/coms.v(73[16:43])
    defparam i2_3_lut_adj_1327.LUT_INIT = 16'h9696;
    SB_LUT4 select_365_Select_28_i3_2_lut_4_lut (.I0(n24810), .I1(n16090), 
            .I2(n16158), .I3(\FRAME_MATCHER.i [28]), .O(n3_adj_4547));
    defparam select_365_Select_28_i3_2_lut_4_lut.LUT_INIT = 16'ha800;
    SB_LUT4 select_365_Select_27_i3_2_lut_4_lut (.I0(n24810), .I1(n16090), 
            .I2(n16158), .I3(\FRAME_MATCHER.i [27]), .O(n3_adj_4546));
    defparam select_365_Select_27_i3_2_lut_4_lut.LUT_INIT = 16'ha800;
    SB_LUT4 i1_2_lut_adj_1328 (.I0(\data_in_frame[2] [0]), .I1(\data_in_frame[2] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n16242));   // verilog/coms.v(69[16:27])
    defparam i1_2_lut_adj_1328.LUT_INIT = 16'h6666;
    SB_LUT4 add_41_17_lut (.I0(n2290), .I1(\FRAME_MATCHER.i [15]), .I2(GND_net), 
            .I3(n27923), .O(n2_adj_4521)) /* synthesis syn_instantiated=1 */ ;
    defparam add_41_17_lut.LUT_INIT = 16'h8228;
    SB_LUT4 select_365_Select_26_i3_2_lut_4_lut (.I0(n24810), .I1(n16090), 
            .I2(n16158), .I3(\FRAME_MATCHER.i [26]), .O(n3_adj_4544));
    defparam select_365_Select_26_i3_2_lut_4_lut.LUT_INIT = 16'ha800;
    SB_LUT4 i1_2_lut_3_lut_adj_1329 (.I0(\data_in[0][6] ), .I1(n22566), 
            .I2(n35535), .I3(GND_net), .O(n10599));   // verilog/coms.v(94[12:19])
    defparam i1_2_lut_3_lut_adj_1329.LUT_INIT = 16'h0d0d;
    SB_LUT4 select_365_Select_25_i3_2_lut_4_lut (.I0(n24810), .I1(n16090), 
            .I2(n16158), .I3(\FRAME_MATCHER.i [25]), .O(n3_adj_4542));
    defparam select_365_Select_25_i3_2_lut_4_lut.LUT_INIT = 16'ha800;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_31620 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[14] [7]), .I2(\data_out_frame[15] [7]), 
            .I3(byte_transmit_counter_c[1]), .O(n38291));
    defparam byte_transmit_counter_0__bdd_4_lut_31620.LUT_INIT = 16'he4aa;
    SB_LUT4 n38291_bdd_4_lut (.I0(n38291), .I1(\data_out_frame[13] [7]), 
            .I2(\data_out_frame[12] [7]), .I3(byte_transmit_counter_c[1]), 
            .O(n38294));
    defparam n38291_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 select_365_Select_24_i3_2_lut_4_lut (.I0(n24810), .I1(n16090), 
            .I2(n16158), .I3(\FRAME_MATCHER.i [24]), .O(n3_adj_4540));
    defparam select_365_Select_24_i3_2_lut_4_lut.LUT_INIT = 16'ha800;
    SB_LUT4 select_365_Select_23_i3_2_lut_4_lut (.I0(n24810), .I1(n16090), 
            .I2(n16158), .I3(\FRAME_MATCHER.i [23]), .O(n3_adj_4538));
    defparam select_365_Select_23_i3_2_lut_4_lut.LUT_INIT = 16'ha800;
    SB_LUT4 select_365_Select_22_i3_2_lut_4_lut (.I0(n24810), .I1(n16090), 
            .I2(n16158), .I3(\FRAME_MATCHER.i [22]), .O(n3_adj_4536));
    defparam select_365_Select_22_i3_2_lut_4_lut.LUT_INIT = 16'ha800;
    SB_LUT4 select_365_Select_21_i3_2_lut_4_lut (.I0(n24810), .I1(n16090), 
            .I2(n16158), .I3(\FRAME_MATCHER.i [21]), .O(n3_adj_4534));
    defparam select_365_Select_21_i3_2_lut_4_lut.LUT_INIT = 16'ha800;
    SB_LUT4 select_365_Select_20_i3_2_lut_4_lut (.I0(n24810), .I1(n16090), 
            .I2(n16158), .I3(\FRAME_MATCHER.i [20]), .O(n3_adj_4532));
    defparam select_365_Select_20_i3_2_lut_4_lut.LUT_INIT = 16'ha800;
    SB_LUT4 select_365_Select_19_i3_2_lut_4_lut (.I0(n24810), .I1(n16090), 
            .I2(n16158), .I3(\FRAME_MATCHER.i [19]), .O(n3_adj_4530));
    defparam select_365_Select_19_i3_2_lut_4_lut.LUT_INIT = 16'ha800;
    SB_LUT4 i1_2_lut_adj_1330 (.I0(\data_in_frame[3] [5]), .I1(\data_in_frame[3] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n33076));   // verilog/coms.v(75[16:43])
    defparam i1_2_lut_adj_1330.LUT_INIT = 16'h6666;
    SB_LUT4 select_365_Select_18_i3_2_lut_4_lut (.I0(n24810), .I1(n16090), 
            .I2(n16158), .I3(\FRAME_MATCHER.i [18]), .O(n3_adj_4528));
    defparam select_365_Select_18_i3_2_lut_4_lut.LUT_INIT = 16'ha800;
    SB_CARRY add_41_17 (.CI(n27923), .I0(\FRAME_MATCHER.i [15]), .I1(GND_net), 
            .CO(n27924));
    SB_LUT4 select_365_Select_17_i3_2_lut_4_lut (.I0(n24810), .I1(n16090), 
            .I2(n16158), .I3(\FRAME_MATCHER.i [17]), .O(n3_adj_4526));
    defparam select_365_Select_17_i3_2_lut_4_lut.LUT_INIT = 16'ha800;
    SB_LUT4 i1_2_lut_3_lut_adj_1331 (.I0(\data_out_frame[19] [5]), .I1(\data_out_frame[19] [2]), 
            .I2(n31178), .I3(GND_net), .O(n6_adj_4434));
    defparam i1_2_lut_3_lut_adj_1331.LUT_INIT = 16'h9696;
    SB_LUT4 select_365_Select_16_i3_2_lut_4_lut (.I0(n24810), .I1(n16090), 
            .I2(n16158), .I3(\FRAME_MATCHER.i [16]), .O(n3_adj_4524));
    defparam select_365_Select_16_i3_2_lut_4_lut.LUT_INIT = 16'ha800;
    SB_LUT4 i13264_3_lut_4_lut (.I0(n8_adj_4435), .I1(n32937), .I2(rx_data[3]), 
            .I3(\data_in_frame[10] [3]), .O(n18093));
    defparam i13264_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_3_lut_adj_1332 (.I0(n16262), .I1(n16399), .I2(\data_in_frame[10] [7]), 
            .I3(GND_net), .O(n33151));   // verilog/coms.v(70[16:27])
    defparam i2_3_lut_adj_1332.LUT_INIT = 16'h9696;
    SB_LUT4 select_365_Select_15_i3_2_lut_4_lut (.I0(n24810), .I1(n16090), 
            .I2(n16158), .I3(\FRAME_MATCHER.i [15]), .O(n3_adj_4522));
    defparam select_365_Select_15_i3_2_lut_4_lut.LUT_INIT = 16'ha800;
    SB_LUT4 i2_3_lut_adj_1333 (.I0(\data_in_frame[9] [0]), .I1(\data_in_frame[11] [1]), 
            .I2(n17169), .I3(GND_net), .O(n17036));   // verilog/coms.v(70[16:27])
    defparam i2_3_lut_adj_1333.LUT_INIT = 16'h9696;
    SB_LUT4 i3_4_lut_adj_1334 (.I0(\data_in_frame[4] [3]), .I1(n32989), 
            .I2(\data_in_frame[1] [7]), .I3(\data_in_frame[2] [1]), .O(n16380));   // verilog/coms.v(232[9:81])
    defparam i3_4_lut_adj_1334.LUT_INIT = 16'h6996;
    SB_CARRY add_3528_5 (.CI(n28020), .I0(byte_transmit_counter_c[3]), .I1(n25050), 
            .CO(n28021));
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_31606 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[14] [6]), .I2(\data_out_frame[15] [6]), 
            .I3(byte_transmit_counter_c[1]), .O(n38285));
    defparam byte_transmit_counter_0__bdd_4_lut_31606.LUT_INIT = 16'he4aa;
    SB_LUT4 add_41_16_lut (.I0(n2290), .I1(\FRAME_MATCHER.i [14]), .I2(GND_net), 
            .I3(n27922), .O(n2_adj_4519)) /* synthesis syn_instantiated=1 */ ;
    defparam add_41_16_lut.LUT_INIT = 16'h8228;
    SB_DFF data_in_frame_0__i139 (.Q(\data_in_frame[17] [2]), .C(clk32MHz), 
           .D(n18148));   // verilog/coms.v(126[12] 293[6])
    SB_LUT4 n38285_bdd_4_lut (.I0(n38285), .I1(\data_out_frame[13] [6]), 
            .I2(\data_out_frame[12] [6]), .I3(byte_transmit_counter_c[1]), 
            .O(n38288));
    defparam n38285_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i2_3_lut_adj_1335 (.I0(\data_in_frame[4] [5]), .I1(n16816), 
            .I2(n4_adj_4410), .I3(GND_net), .O(n16834));   // verilog/coms.v(232[9:81])
    defparam i2_3_lut_adj_1335.LUT_INIT = 16'h9696;
    SB_LUT4 i3_3_lut_4_lut_adj_1336 (.I0(\data_in_frame[16] [3]), .I1(Kp_23__N_843), 
            .I2(\data_in_frame[20] [5]), .I3(n33279), .O(n8_adj_4449));
    defparam i3_3_lut_4_lut_adj_1336.LUT_INIT = 16'h6996;
    SB_LUT4 i13265_3_lut_4_lut (.I0(n8_adj_4435), .I1(n32937), .I2(rx_data[4]), 
            .I3(\data_in_frame[10] [4]), .O(n18094));
    defparam i13265_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 select_365_Select_14_i3_2_lut_4_lut (.I0(n24810), .I1(n16090), 
            .I2(n16158), .I3(\FRAME_MATCHER.i [14]), .O(n3_adj_4520));
    defparam select_365_Select_14_i3_2_lut_4_lut.LUT_INIT = 16'ha800;
    SB_LUT4 select_365_Select_13_i3_2_lut_4_lut (.I0(n24810), .I1(n16090), 
            .I2(n16158), .I3(\FRAME_MATCHER.i [13]), .O(n3_adj_4518));
    defparam select_365_Select_13_i3_2_lut_4_lut.LUT_INIT = 16'ha800;
    SB_LUT4 i3_4_lut_adj_1337 (.I0(n30801), .I1(\data_out_frame[14] [2]), 
            .I2(\data_out_frame[16] [4]), .I3(\data_out_frame[14] [3]), 
            .O(n33192));
    defparam i3_4_lut_adj_1337.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1338 (.I0(n16384), .I1(n16834), .I2(\data_in_frame[6] [6]), 
            .I3(GND_net), .O(n17169));
    defparam i2_3_lut_adj_1338.LUT_INIT = 16'h9696;
    SB_DFF data_in_frame_0__i138 (.Q(\data_in_frame[17] [1]), .C(clk32MHz), 
           .D(n18147));   // verilog/coms.v(126[12] 293[6])
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_31615 (.I0(byte_transmit_counter_c[1]), 
            .I1(n37273), .I2(n37274), .I3(byte_transmit_counter_c[2]), 
            .O(n38279));
    defparam byte_transmit_counter_1__bdd_4_lut_31615.LUT_INIT = 16'he4aa;
    SB_LUT4 i3_4_lut_adj_1339 (.I0(n33503), .I1(\data_in_frame[11] [3]), 
            .I2(\data_in_frame[8] [7]), .I3(n33529), .O(n33388));
    defparam i3_4_lut_adj_1339.LUT_INIT = 16'h9669;
    SB_LUT4 select_365_Select_12_i3_2_lut_4_lut (.I0(n24810), .I1(n16090), 
            .I2(n16158), .I3(\FRAME_MATCHER.i [12]), .O(n3_adj_4516));
    defparam select_365_Select_12_i3_2_lut_4_lut.LUT_INIT = 16'ha800;
    SB_LUT4 i1_2_lut_3_lut_adj_1340 (.I0(\data_out_frame[5] [3]), .I1(\data_out_frame[5] [5]), 
            .I2(n33589), .I3(GND_net), .O(n33543));
    defparam i1_2_lut_3_lut_adj_1340.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1341 (.I0(n16746), .I1(n34982), .I2(GND_net), 
            .I3(GND_net), .O(n33448));
    defparam i1_2_lut_adj_1341.LUT_INIT = 16'h9999;
    SB_LUT4 i4_4_lut_adj_1342 (.I0(\data_in_frame[11] [2]), .I1(n17169), 
            .I2(n16840), .I3(n6_adj_4406), .O(n30930));   // verilog/coms.v(73[16:43])
    defparam i4_4_lut_adj_1342.LUT_INIT = 16'h6996;
    SB_LUT4 n38279_bdd_4_lut (.I0(n38279), .I1(n17_adj_4571), .I2(n16_adj_4570), 
            .I3(byte_transmit_counter_c[2]), .O(n38282));
    defparam n38279_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 select_365_Select_11_i3_2_lut_4_lut (.I0(n24810), .I1(n16090), 
            .I2(n16158), .I3(\FRAME_MATCHER.i [11]), .O(n3_adj_4514));
    defparam select_365_Select_11_i3_2_lut_4_lut.LUT_INIT = 16'ha800;
    SB_DFF IntegralLimit_i0_i0 (.Q(IntegralLimit[0]), .C(clk32MHz), .D(n17550));   // verilog/coms.v(126[12] 293[6])
    SB_DFF IntegralLimit_i0_i6 (.Q(IntegralLimit[6]), .C(clk32MHz), .D(n17773));   // verilog/coms.v(126[12] 293[6])
    SB_DFF IntegralLimit_i0_i5 (.Q(IntegralLimit[5]), .C(clk32MHz), .D(n17772));   // verilog/coms.v(126[12] 293[6])
    SB_DFF IntegralLimit_i0_i4 (.Q(IntegralLimit[4]), .C(clk32MHz), .D(n17771));   // verilog/coms.v(126[12] 293[6])
    SB_DFF IntegralLimit_i0_i3 (.Q(IntegralLimit[3]), .C(clk32MHz), .D(n17770));   // verilog/coms.v(126[12] 293[6])
    SB_DFF IntegralLimit_i0_i2 (.Q(IntegralLimit[2]), .C(clk32MHz), .D(n17769));   // verilog/coms.v(126[12] 293[6])
    SB_DFF IntegralLimit_i0_i1 (.Q(IntegralLimit[1]), .C(clk32MHz), .D(n17768));   // verilog/coms.v(126[12] 293[6])
    SB_LUT4 select_365_Select_10_i3_2_lut_4_lut (.I0(n24810), .I1(n16090), 
            .I2(n16158), .I3(\FRAME_MATCHER.i [10]), .O(n3_adj_4512));
    defparam select_365_Select_10_i3_2_lut_4_lut.LUT_INIT = 16'ha800;
    SB_LUT4 select_365_Select_9_i3_2_lut_4_lut (.I0(n24810), .I1(n16090), 
            .I2(n16158), .I3(\FRAME_MATCHER.i [9]), .O(n3_adj_4510));
    defparam select_365_Select_9_i3_2_lut_4_lut.LUT_INIT = 16'ha800;
    SB_LUT4 i13266_3_lut_4_lut (.I0(n8_adj_4435), .I1(n32937), .I2(rx_data[5]), 
            .I3(\data_in_frame[10] [5]), .O(n18095));
    defparam i13266_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 select_365_Select_8_i3_2_lut_4_lut (.I0(n24810), .I1(n16090), 
            .I2(n16158), .I3(\FRAME_MATCHER.i [8]), .O(n3_adj_4508));
    defparam select_365_Select_8_i3_2_lut_4_lut.LUT_INIT = 16'ha800;
    SB_DFF data_in_frame_0__i68 (.Q(\data_in_frame[8] [3]), .C(clk32MHz), 
           .D(n18077));   // verilog/coms.v(126[12] 293[6])
    SB_LUT4 i4_4_lut_adj_1343 (.I0(\data_in_frame[13] [3]), .I1(\data_in_frame[8] [7]), 
            .I2(n16418), .I3(n6_adj_4587), .O(n16862));   // verilog/coms.v(70[16:27])
    defparam i4_4_lut_adj_1343.LUT_INIT = 16'h6996;
    SB_LUT4 select_365_Select_7_i3_2_lut_4_lut (.I0(n24810), .I1(n16090), 
            .I2(n16158), .I3(\FRAME_MATCHER.i [7]), .O(n3_adj_4506));
    defparam select_365_Select_7_i3_2_lut_4_lut.LUT_INIT = 16'ha800;
    SB_LUT4 i2_3_lut_adj_1344 (.I0(\data_in_frame[13] [4]), .I1(n16862), 
            .I2(n30930), .I3(GND_net), .O(n35410));
    defparam i2_3_lut_adj_1344.LUT_INIT = 16'h9696;
    SB_LUT4 i3_4_lut_adj_1345 (.I0(\data_in_frame[16] [6]), .I1(\data_in_frame[16] [3]), 
            .I2(\data_in_frame[16] [1]), .I3(n17081), .O(n33081));   // verilog/coms.v(77[16:27])
    defparam i3_4_lut_adj_1345.LUT_INIT = 16'h6996;
    SB_LUT4 select_365_Select_6_i3_2_lut_4_lut (.I0(n24810), .I1(n16090), 
            .I2(n16158), .I3(\FRAME_MATCHER.i [6]), .O(n3_adj_4504));
    defparam select_365_Select_6_i3_2_lut_4_lut.LUT_INIT = 16'ha800;
    SB_LUT4 select_365_Select_5_i3_2_lut_4_lut (.I0(n24810), .I1(n16090), 
            .I2(n16158), .I3(\FRAME_MATCHER.i [5]), .O(n3_adj_4502));
    defparam select_365_Select_5_i3_2_lut_4_lut.LUT_INIT = 16'ha800;
    SB_LUT4 i1_2_lut_adj_1346 (.I0(\data_in_frame[3] [7]), .I1(\data_in_frame[3] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n16299));   // verilog/coms.v(84[17:28])
    defparam i1_2_lut_adj_1346.LUT_INIT = 16'h6666;
    SB_LUT4 add_3528_4_lut (.I0(byte_transmit_counter_c[2]), .I1(byte_transmit_counter_c[2]), 
            .I2(n25050), .I3(n28019), .O(n17671)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3528_4_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 i1_2_lut_adj_1347 (.I0(n34982), .I1(n16711), .I2(GND_net), 
            .I3(GND_net), .O(n31209));
    defparam i1_2_lut_adj_1347.LUT_INIT = 16'h9999;
    SB_LUT4 select_365_Select_4_i3_2_lut_4_lut (.I0(n24810), .I1(n16090), 
            .I2(n16158), .I3(\FRAME_MATCHER.i [4]), .O(n3_adj_4500));
    defparam select_365_Select_4_i3_2_lut_4_lut.LUT_INIT = 16'ha800;
    SB_LUT4 i13267_3_lut_4_lut (.I0(n8_adj_4435), .I1(n32937), .I2(rx_data[6]), 
            .I3(\data_in_frame[10] [6]), .O(n18096));
    defparam i13267_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_3_lut_adj_1348 (.I0(n14758), .I1(n35410), .I2(\data_in_frame[16] [0]), 
            .I3(GND_net), .O(n33045));
    defparam i2_3_lut_adj_1348.LUT_INIT = 16'h6969;
    SB_CARRY add_41_16 (.CI(n27922), .I0(\FRAME_MATCHER.i [14]), .I1(GND_net), 
            .CO(n27923));
    SB_LUT4 i2_3_lut_adj_1349 (.I0(\data_in_frame[16] [5]), .I1(n33081), 
            .I2(\data_in_frame[16] [7]), .I3(GND_net), .O(Kp_23__N_1662));   // verilog/coms.v(77[16:27])
    defparam i2_3_lut_adj_1349.LUT_INIT = 16'h9696;
    SB_LUT4 data_in_frame_12__7__I_0_3451_2_lut (.I0(\data_in_frame[12] [7]), 
            .I1(\data_in_frame[12] [6]), .I2(GND_net), .I3(GND_net), .O(Kp_23__N_860));   // verilog/coms.v(70[16:27])
    defparam data_in_frame_12__7__I_0_3451_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_1350 (.I0(\data_in_frame[5] [7]), .I1(\data_in_frame[8] [1]), 
            .I2(n33036), .I3(GND_net), .O(n16780));   // verilog/coms.v(84[17:28])
    defparam i2_3_lut_adj_1350.LUT_INIT = 16'h9696;
    SB_LUT4 i3_2_lut_4_lut_adj_1351 (.I0(\data_out_frame[10] [6]), .I1(\data_out_frame[13] [0]), 
            .I2(\data_out_frame[12] [7]), .I3(\data_out_frame[12] [4]), 
            .O(n16_adj_4426));
    defparam i3_2_lut_4_lut_adj_1351.LUT_INIT = 16'h6996;
    SB_LUT4 i13268_3_lut_4_lut (.I0(n8_adj_4435), .I1(n32937), .I2(rx_data[7]), 
            .I3(\data_in_frame[10] [7]), .O(n18097));
    defparam i13268_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i4_4_lut_adj_1352 (.I0(Kp_23__N_1662), .I1(\data_in_frame[15] [5]), 
            .I2(n33045), .I3(n6_adj_4609), .O(n30805));
    defparam i4_4_lut_adj_1352.LUT_INIT = 16'h6996;
    SB_LUT4 i17_3_lut (.I0(\data_in_frame[14] [4]), .I1(\data_in_frame[15] [0]), 
            .I2(\data_in_frame[6] [3]), .I3(GND_net), .O(n50));
    defparam i17_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 select_365_Select_3_i3_2_lut_4_lut (.I0(n24810), .I1(n16090), 
            .I2(n16158), .I3(\FRAME_MATCHER.i [3]), .O(n3_adj_4498));
    defparam select_365_Select_3_i3_2_lut_4_lut.LUT_INIT = 16'ha800;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_31597 (.I0(byte_transmit_counter_c[1]), 
            .I1(n37276), .I2(n37277), .I3(byte_transmit_counter_c[2]), 
            .O(n38273));
    defparam byte_transmit_counter_1__bdd_4_lut_31597.LUT_INIT = 16'he4aa;
    SB_LUT4 i2_3_lut_4_lut_adj_1353 (.I0(\FRAME_MATCHER.state [0]), .I1(\FRAME_MATCHER.state [1]), 
            .I2(\FRAME_MATCHER.state_31__N_2630 [3]), .I3(\FRAME_MATCHER.state [2]), 
            .O(n35045));   // verilog/coms.v(144[4] 292[11])
    defparam i2_3_lut_4_lut_adj_1353.LUT_INIT = 16'hfffb;
    SB_LUT4 select_365_Select_2_i3_2_lut_4_lut (.I0(n24810), .I1(n16090), 
            .I2(n16158), .I3(\FRAME_MATCHER.i [2]), .O(n3_adj_4496));
    defparam select_365_Select_2_i3_2_lut_4_lut.LUT_INIT = 16'ha800;
    SB_LUT4 i24_4_lut_adj_1354 (.I0(n17111), .I1(Kp_23__N_860), .I2(n17157), 
            .I3(\data_in_frame[13] [3]), .O(n57));
    defparam i24_4_lut_adj_1354.LUT_INIT = 16'h6996;
    SB_LUT4 select_365_Select_1_i3_2_lut_4_lut (.I0(n24810), .I1(n16090), 
            .I2(n16158), .I3(\FRAME_MATCHER.i [1]), .O(n3_adj_4485));
    defparam select_365_Select_1_i3_2_lut_4_lut.LUT_INIT = 16'ha800;
    SB_LUT4 i21_4_lut (.I0(\data_in_frame[13] [1]), .I1(\data_in_frame[15] [2]), 
            .I2(\data_in_frame[14] [1]), .I3(n33628), .O(n54));
    defparam i21_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 select_365_Select_0_i3_2_lut_4_lut (.I0(n24810), .I1(n16090), 
            .I2(n16158), .I3(\FRAME_MATCHER.i [0]), .O(n3));
    defparam select_365_Select_0_i3_2_lut_4_lut.LUT_INIT = 16'ha800;
    SB_LUT4 i19_4_lut_adj_1355 (.I0(\data_in_frame[6] [2]), .I1(n33631), 
            .I2(\data_in_frame[13] [7]), .I3(n33508), .O(n52));
    defparam i19_4_lut_adj_1355.LUT_INIT = 16'h6996;
    SB_LUT4 n38273_bdd_4_lut (.I0(n38273), .I1(n17_adj_4481), .I2(n16_adj_4480), 
            .I3(byte_transmit_counter_c[2]), .O(n38276));
    defparam n38273_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_CARRY add_3528_4 (.CI(n28019), .I0(byte_transmit_counter_c[2]), .I1(n25050), 
            .CO(n28020));
    SB_LUT4 add_3528_3_lut (.I0(byte_transmit_counter_c[1]), .I1(byte_transmit_counter_c[1]), 
            .I2(n25050), .I3(n28018), .O(n17674)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3528_3_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY add_3528_3 (.CI(n28018), .I0(byte_transmit_counter_c[1]), .I1(n25050), 
            .CO(n28019));
    SB_LUT4 i13297_3_lut_4_lut (.I0(n8_adj_4355), .I1(n32937), .I2(rx_data[4]), 
            .I3(\data_in_frame[14] [4]), .O(n18126));
    defparam i13297_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_31592 (.I0(byte_transmit_counter_c[1]), 
            .I1(n37279), .I2(n37280), .I3(byte_transmit_counter_c[2]), 
            .O(n38267));
    defparam byte_transmit_counter_1__bdd_4_lut_31592.LUT_INIT = 16'he4aa;
    SB_LUT4 i13298_3_lut_4_lut (.I0(n8_adj_4355), .I1(n32937), .I2(rx_data[5]), 
            .I3(\data_in_frame[14] [5]), .O(n18127));
    defparam i13298_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 n38267_bdd_4_lut (.I0(n38267), .I1(n17_adj_4479), .I2(n16_adj_4478), 
            .I3(byte_transmit_counter_c[2]), .O(n38270));
    defparam n38267_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i13299_3_lut_4_lut (.I0(n8_adj_4355), .I1(n32937), .I2(rx_data[6]), 
            .I3(\data_in_frame[14] [6]), .O(n18128));
    defparam i13299_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 add_3528_2_lut (.I0(GND_net), .I1(byte_transmit_counter[0]), 
            .I2(tx_transmit_N_3355), .I3(GND_net), .O(n8014)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3528_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i13300_3_lut_4_lut (.I0(n8_adj_4355), .I1(n32937), .I2(rx_data[7]), 
            .I3(\data_in_frame[14] [7]), .O(n18129));
    defparam i13300_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13296_3_lut_4_lut (.I0(n8_adj_4355), .I1(n32937), .I2(rx_data[3]), 
            .I3(\data_in_frame[14] [3]), .O(n18125));
    defparam i13296_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 add_41_15_lut (.I0(n2290), .I1(\FRAME_MATCHER.i [13]), .I2(GND_net), 
            .I3(n27921), .O(n2_adj_4517)) /* synthesis syn_instantiated=1 */ ;
    defparam add_41_15_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i13293_3_lut_4_lut (.I0(n8_adj_4355), .I1(n32937), .I2(rx_data[0]), 
            .I3(\data_in_frame[14] [0]), .O(n18122));
    defparam i13293_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_CARRY add_3528_2 (.CI(GND_net), .I0(byte_transmit_counter[0]), .I1(tx_transmit_N_3355), 
            .CO(n28018));
    SB_LUT4 i13294_3_lut_4_lut (.I0(n8_adj_4355), .I1(n32937), .I2(rx_data[1]), 
            .I3(\data_in_frame[14] [1]), .O(n18123));
    defparam i13294_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13295_3_lut_4_lut (.I0(n8_adj_4355), .I1(n32937), .I2(rx_data[2]), 
            .I3(\data_in_frame[14] [2]), .O(n18124));
    defparam i13295_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_2_lut_3_lut_adj_1356 (.I0(\data_out_frame[13] [1]), .I1(\data_out_frame[13] [2]), 
            .I2(n16687), .I3(GND_net), .O(n10_adj_4606));
    defparam i2_2_lut_3_lut_adj_1356.LUT_INIT = 16'h9696;
    SB_LUT4 i20_4_lut (.I0(n33320), .I1(\data_in_frame[10] [7]), .I2(n33039), 
            .I3(n30900), .O(n53_adj_4610));
    defparam i20_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i18_4_lut_adj_1357 (.I0(n33454), .I1(n33598), .I2(\data_in_frame[11] [5]), 
            .I3(n33155), .O(n51));
    defparam i18_4_lut_adj_1357.LUT_INIT = 16'h6996;
    SB_CARRY add_41_15 (.CI(n27921), .I0(\FRAME_MATCHER.i [13]), .I1(GND_net), 
            .CO(n27922));
    SB_LUT4 i1_2_lut_3_lut_adj_1358 (.I0(\data_out_frame[5] [6]), .I1(\data_out_frame[6] [0]), 
            .I2(\data_out_frame[6] [1]), .I3(GND_net), .O(n32985));   // verilog/coms.v(84[17:28])
    defparam i1_2_lut_3_lut_adj_1358.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1359 (.I0(n16404), .I1(n31204), .I2(n35262), 
            .I3(GND_net), .O(n32999));
    defparam i1_2_lut_3_lut_adj_1359.LUT_INIT = 16'h6969;
    SB_LUT4 i1_2_lut_3_lut_adj_1360 (.I0(\data_out_frame[13] [1]), .I1(\data_out_frame[13] [2]), 
            .I2(\data_out_frame[13] [3]), .I3(GND_net), .O(n33073));
    defparam i1_2_lut_3_lut_adj_1360.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_4_lut_adj_1361 (.I0(n16404), .I1(n31204), .I2(n30192), 
            .I3(n31190), .O(n34495));
    defparam i2_3_lut_4_lut_adj_1361.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1362 (.I0(\data_out_frame[8] [1]), .I1(\data_out_frame[8] [2]), 
            .I2(n30857), .I3(GND_net), .O(n33537));
    defparam i1_2_lut_3_lut_adj_1362.LUT_INIT = 16'h9696;
    SB_LUT4 i23_4_lut_adj_1363 (.I0(n33118), .I1(\data_in_frame[7] [3]), 
            .I2(n33010), .I3(Kp_23__N_1183), .O(n56));
    defparam i23_4_lut_adj_1363.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_1364 (.I0(\data_out_frame[8] [1]), .I1(\data_out_frame[8] [2]), 
            .I2(\data_out_frame[10] [3]), .I3(n32985), .O(n33287));
    defparam i2_3_lut_4_lut_adj_1364.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1365 (.I0(\data_out_frame[14] [6]), .I1(\data_out_frame[17] [0]), 
            .I2(n31287), .I3(GND_net), .O(n33570));
    defparam i1_2_lut_3_lut_adj_1365.LUT_INIT = 16'h9696;
    SB_LUT4 i29_4_lut (.I0(n57), .I1(\data_in_frame[13] [0]), .I2(n50), 
            .I3(\data_in_frame[14] [3]), .O(n62));
    defparam i29_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1366 (.I0(\data_out_frame[5] [2]), .I1(\data_out_frame[5] [1]), 
            .I2(n16163), .I3(\data_out_frame[7] [3]), .O(n33115));
    defparam i1_2_lut_3_lut_4_lut_adj_1366.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1367 (.I0(\data_out_frame[5] [2]), .I1(\data_out_frame[5] [1]), 
            .I2(\data_out_frame[5] [0]), .I3(GND_net), .O(n33381));
    defparam i1_2_lut_3_lut_adj_1367.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1368 (.I0(\data_out_frame[5] [2]), .I1(\data_out_frame[5] [1]), 
            .I2(n16687), .I3(\data_out_frame[7] [3]), .O(n33241));
    defparam i1_2_lut_3_lut_4_lut_adj_1368.LUT_INIT = 16'h6996;
    SB_LUT4 i22_4_lut (.I0(n33592), .I1(n33414), .I2(n33491), .I3(n16248), 
            .O(n55));
    defparam i22_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1369 (.I0(\FRAME_MATCHER.state [2]), .I1(\FRAME_MATCHER.state [0]), 
            .I2(n16153), .I3(GND_net), .O(n16154));   // verilog/coms.v(247[5:25])
    defparam i1_2_lut_3_lut_adj_1369.LUT_INIT = 16'hfbfb;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1370 (.I0(n118), .I1(n10599), .I2(n24786), 
            .I3(n3007), .O(n7_adj_4402));   // verilog/coms.v(94[12:19])
    defparam i1_2_lut_3_lut_4_lut_adj_1370.LUT_INIT = 16'h0080;
    SB_LUT4 i119_2_lut_3_lut_4_lut (.I0(n118), .I1(n10599), .I2(n16161), 
            .I3(n3007), .O(n98));   // verilog/coms.v(94[12:19])
    defparam i119_2_lut_3_lut_4_lut.LUT_INIT = 16'h0008;
    SB_LUT4 i1_2_lut_3_lut_adj_1371 (.I0(n118), .I1(n10599), .I2(n2958), 
            .I3(GND_net), .O(n1_c));   // verilog/coms.v(94[12:19])
    defparam i1_2_lut_3_lut_adj_1371.LUT_INIT = 16'h8080;
    SB_LUT4 i30_4_lut (.I0(n51), .I1(n53_adj_4610), .I2(n52), .I3(n54), 
            .O(n63_adj_4611));
    defparam i30_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 add_41_14_lut (.I0(n2290), .I1(\FRAME_MATCHER.i [12]), .I2(GND_net), 
            .I3(n27920), .O(n2_adj_4515)) /* synthesis syn_instantiated=1 */ ;
    defparam add_41_14_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i1_3_lut_4_lut (.I0(n118), .I1(n10599), .I2(n16154), .I3(n3893), 
            .O(n3_adj_4430));   // verilog/coms.v(94[12:19])
    defparam i1_3_lut_4_lut.LUT_INIT = 16'h0008;
    SB_LUT4 i1_3_lut_4_lut_adj_1372 (.I0(n118), .I1(n10599), .I2(n16157), 
            .I3(n1502), .O(n53));   // verilog/coms.v(94[12:19])
    defparam i1_3_lut_4_lut_adj_1372.LUT_INIT = 16'h0800;
    SB_LUT4 i32_4_lut (.I0(n63_adj_4611), .I1(n55), .I2(n62), .I3(n56), 
            .O(n14758));
    defparam i32_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1373 (.I0(n16722), .I1(\data_in_frame[6] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n33121));   // verilog/coms.v(73[16:43])
    defparam i1_2_lut_adj_1373.LUT_INIT = 16'h6666;
    SB_LUT4 i1_4_lut_adj_1374 (.I0(\data_in_frame[13] [7]), .I1(n33259), 
            .I2(n33500), .I3(n16608), .O(n33625));
    defparam i1_4_lut_adj_1374.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_adj_1375 (.I0(\data_out_frame[7] [0]), .I1(\data_out_frame[6] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n16392));   // verilog/coms.v(70[16:27])
    defparam i1_2_lut_adj_1375.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_1376 (.I0(n16299), .I1(n33076), .I2(n16242), 
            .I3(\data_in_frame[3] [2]), .O(n33558));   // verilog/coms.v(95[12:25])
    defparam i3_4_lut_adj_1376.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_1377 (.I0(n33505), .I1(\data_in_frame[11] [6]), 
            .I2(\data_in_frame[14] [2]), .I3(n35345), .O(n16620));
    defparam i2_3_lut_4_lut_adj_1377.LUT_INIT = 16'h9669;
    SB_LUT4 i2_3_lut_adj_1378 (.I0(\data_in_frame[9] [4]), .I1(\data_in_frame[13] [6]), 
            .I2(\data_in_frame[9] [5]), .I3(GND_net), .O(n33454));
    defparam i2_3_lut_adj_1378.LUT_INIT = 16'h9696;
    SB_LUT4 i31544_2_lut_3_lut (.I0(byte_transmit_counter_c[3]), .I1(byte_transmit_counter_c[4]), 
            .I2(n16000), .I3(GND_net), .O(tx_transmit_N_3355));
    defparam i31544_2_lut_3_lut.LUT_INIT = 16'h0707;
    SB_LUT4 i1_2_lut_adj_1379 (.I0(\data_in_frame[11] [6]), .I1(n33625), 
            .I2(GND_net), .I3(GND_net), .O(n33207));
    defparam i1_2_lut_adj_1379.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1380 (.I0(\data_out_frame[9] [2]), .I1(\data_out_frame[9] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n33069));   // verilog/coms.v(84[17:63])
    defparam i1_2_lut_adj_1380.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1381 (.I0(\data_in_frame[7] [0]), .I1(\data_in_frame[4] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n17111));   // verilog/coms.v(73[16:43])
    defparam i1_2_lut_adj_1381.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1382 (.I0(n118), .I1(n737), .I2(n16080), 
            .I3(n10599), .O(n4_adj_4401));   // verilog/coms.v(94[12:19])
    defparam i1_2_lut_3_lut_4_lut_adj_1382.LUT_INIT = 16'h0200;
    SB_LUT4 i1_2_lut_3_lut_adj_1383 (.I0(\FRAME_MATCHER.state [2]), .I1(\FRAME_MATCHER.state [0]), 
            .I2(n16153), .I3(GND_net), .O(n16157));   // verilog/coms.v(208[5:16])
    defparam i1_2_lut_3_lut_adj_1383.LUT_INIT = 16'hf7f7;
    SB_LUT4 i2_3_lut_4_lut_adj_1384 (.I0(n118), .I1(n737), .I2(n92[2]), 
            .I3(n16159), .O(n34531));   // verilog/coms.v(94[12:19])
    defparam i2_3_lut_4_lut_adj_1384.LUT_INIT = 16'h0020;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1385 (.I0(n118), .I1(n737), .I2(n16159), 
            .I3(n10599), .O(n136));   // verilog/coms.v(94[12:19])
    defparam i1_2_lut_3_lut_4_lut_adj_1385.LUT_INIT = 16'h0200;
    SB_LUT4 i2_3_lut_4_lut_adj_1386 (.I0(\data_out_frame[7] [7]), .I1(\data_out_frame[7] [6]), 
            .I2(\data_out_frame[8] [0]), .I3(\data_out_frame[5] [6]), .O(n33145));
    defparam i2_3_lut_4_lut_adj_1386.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_1387 (.I0(\data_in_frame[6] [5]), .I1(\data_in_frame[6] [7]), 
            .I2(n33414), .I3(n6_adj_4407), .O(n16418));   // verilog/coms.v(73[16:43])
    defparam i4_4_lut_adj_1387.LUT_INIT = 16'h6996;
    SB_LUT4 i1_3_lut_4_lut_adj_1388 (.I0(n35535), .I1(\data_in[0][6] ), 
            .I2(n22566), .I3(\FRAME_MATCHER.state [2]), .O(n92[2]));
    defparam i1_3_lut_4_lut_adj_1388.LUT_INIT = 16'h5d0c;
    SB_LUT4 i1_2_lut_3_lut_adj_1389 (.I0(\data_out_frame[9] [7]), .I1(\data_out_frame[7] [5]), 
            .I2(\data_out_frame[12] [3]), .I3(GND_net), .O(n33622));
    defparam i1_2_lut_3_lut_adj_1389.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_4_lut_adj_1390 (.I0(Kp_23__N_1453), .I1(n31196), .I2(n31228), 
            .I3(n15781), .O(n6_adj_4421));
    defparam i2_3_lut_4_lut_adj_1390.LUT_INIT = 16'h9669;
    SB_LUT4 i2_3_lut_4_lut_adj_1391 (.I0(\data_out_frame[12] [4]), .I1(n16951), 
            .I2(\data_out_frame[12] [3]), .I3(\data_out_frame[5] [4]), .O(n33540));   // verilog/coms.v(84[17:28])
    defparam i2_3_lut_4_lut_adj_1391.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1392 (.I0(\data_in_frame[14] [0]), .I1(n33207), 
            .I2(n33454), .I3(n15795), .O(n33298));
    defparam i1_4_lut_adj_1392.LUT_INIT = 16'h9669;
    SB_LUT4 i1_4_lut_adj_1393 (.I0(\data_out_frame[14] [0]), .I1(n33069), 
            .I2(n16163), .I3(\data_out_frame[9] [5]), .O(n6_adj_4612));
    defparam i1_4_lut_adj_1393.LUT_INIT = 16'h6996;
    SB_CARRY add_41_14 (.CI(n27920), .I0(\FRAME_MATCHER.i [12]), .I1(GND_net), 
            .CO(n27921));
    SB_LUT4 i1_2_lut_3_lut_adj_1394 (.I0(n53), .I1(n3_adj_4430), .I2(\FRAME_MATCHER.state [31]), 
            .I3(GND_net), .O(n32179));
    defparam i1_2_lut_3_lut_adj_1394.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_2_lut_3_lut_adj_1395 (.I0(n53), .I1(n3_adj_4430), .I2(\FRAME_MATCHER.state [30]), 
            .I3(GND_net), .O(n32175));
    defparam i1_2_lut_3_lut_adj_1395.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_2_lut_3_lut_adj_1396 (.I0(n53), .I1(n3_adj_4430), .I2(\FRAME_MATCHER.state [29]), 
            .I3(GND_net), .O(n32173));
    defparam i1_2_lut_3_lut_adj_1396.LUT_INIT = 16'he0e0;
    SB_LUT4 i4_4_lut_adj_1397 (.I0(n33060), .I1(n16392), .I2(\data_out_frame[9] [4]), 
            .I3(n6_adj_4612), .O(n33520));
    defparam i4_4_lut_adj_1397.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1398 (.I0(n53), .I1(n3_adj_4430), .I2(\FRAME_MATCHER.state [28]), 
            .I3(GND_net), .O(n32273));
    defparam i1_2_lut_3_lut_adj_1398.LUT_INIT = 16'he0e0;
    SB_LUT4 i2_3_lut_adj_1399 (.I0(n16418), .I1(n16248), .I2(\data_in_frame[16] [0]), 
            .I3(GND_net), .O(n33217));
    defparam i2_3_lut_adj_1399.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1400 (.I0(n53), .I1(n3_adj_4430), .I2(\FRAME_MATCHER.state [27]), 
            .I3(GND_net), .O(n32171));
    defparam i1_2_lut_3_lut_adj_1400.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_2_lut_3_lut_adj_1401 (.I0(n53), .I1(n3_adj_4430), .I2(\FRAME_MATCHER.state [26]), 
            .I3(GND_net), .O(n32301));
    defparam i1_2_lut_3_lut_adj_1401.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_2_lut_3_lut_adj_1402 (.I0(n53), .I1(n3_adj_4430), .I2(\FRAME_MATCHER.state [25]), 
            .I3(GND_net), .O(n32299));
    defparam i1_2_lut_3_lut_adj_1402.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_2_lut_3_lut_adj_1403 (.I0(n53), .I1(n3_adj_4430), .I2(\FRAME_MATCHER.state [24]), 
            .I3(GND_net), .O(n32297));
    defparam i1_2_lut_3_lut_adj_1403.LUT_INIT = 16'he0e0;
    SB_LUT4 add_41_13_lut (.I0(n2290), .I1(\FRAME_MATCHER.i [11]), .I2(GND_net), 
            .I3(n27919), .O(n2_adj_4513)) /* synthesis syn_instantiated=1 */ ;
    defparam add_41_13_lut.LUT_INIT = 16'h8228;
    SB_DFF data_in_frame_0__i137 (.Q(\data_in_frame[17] [0]), .C(clk32MHz), 
           .D(n18146));   // verilog/coms.v(126[12] 293[6])
    SB_LUT4 i23019_2_lut_3_lut (.I0(n53), .I1(n3_adj_4430), .I2(\FRAME_MATCHER.state [23]), 
            .I3(GND_net), .O(n29601));
    defparam i23019_2_lut_3_lut.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_2_lut_3_lut_adj_1404 (.I0(n53), .I1(n3_adj_4430), .I2(\FRAME_MATCHER.state [22]), 
            .I3(GND_net), .O(n32295));
    defparam i1_2_lut_3_lut_adj_1404.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_2_lut_3_lut_adj_1405 (.I0(n53), .I1(n3_adj_4430), .I2(\FRAME_MATCHER.state [21]), 
            .I3(GND_net), .O(n32293));
    defparam i1_2_lut_3_lut_adj_1405.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_2_lut_3_lut_adj_1406 (.I0(\data_out_frame[5] [0]), .I1(\data_out_frame[6] [7]), 
            .I2(\data_out_frame[7] [1]), .I3(GND_net), .O(n17182));   // verilog/coms.v(84[17:70])
    defparam i1_2_lut_3_lut_adj_1406.LUT_INIT = 16'h9696;
    SB_LUT4 i19302_2_lut_3_lut (.I0(n53), .I1(n3_adj_4430), .I2(\FRAME_MATCHER.state [20]), 
            .I3(GND_net), .O(n24112));
    defparam i19302_2_lut_3_lut.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_2_lut_4_lut_adj_1407 (.I0(n118), .I1(n35535), .I2(n42_adj_4411), 
            .I3(\FRAME_MATCHER.state [2]), .O(\FRAME_MATCHER.state_31__N_2566[2] ));   // verilog/coms.v(94[12:19])
    defparam i1_2_lut_4_lut_adj_1407.LUT_INIT = 16'ha2a0;
    SB_LUT4 i1_2_lut_3_lut_adj_1408 (.I0(n53), .I1(n3_adj_4430), .I2(\FRAME_MATCHER.state [19]), 
            .I3(GND_net), .O(n32185));
    defparam i1_2_lut_3_lut_adj_1408.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_2_lut_3_lut_adj_1409 (.I0(n53), .I1(n3_adj_4430), .I2(\FRAME_MATCHER.state [18]), 
            .I3(GND_net), .O(n32275));
    defparam i1_2_lut_3_lut_adj_1409.LUT_INIT = 16'he0e0;
    SB_LUT4 i19301_2_lut_3_lut (.I0(n53), .I1(n3_adj_4430), .I2(\FRAME_MATCHER.state [17]), 
            .I3(GND_net), .O(n24110));
    defparam i19301_2_lut_3_lut.LUT_INIT = 16'he0e0;
    SB_LUT4 i3_4_lut_adj_1410 (.I0(\data_in_frame[18] [1]), .I1(n14758), 
            .I2(n30805), .I3(n34514), .O(n33583));
    defparam i3_4_lut_adj_1410.LUT_INIT = 16'h9669;
    SB_LUT4 i2_3_lut_adj_1411 (.I0(n33217), .I1(n33298), .I2(\data_in_frame[16] [1]), 
            .I3(GND_net), .O(n34605));   // verilog/coms.v(73[16:43])
    defparam i2_3_lut_adj_1411.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_4_lut_adj_1412 (.I0(\data_out_frame[11] [6]), .I1(n17182), 
            .I2(\data_out_frame[9] [3]), .I3(n33517), .O(n33060));   // verilog/coms.v(84[17:63])
    defparam i2_3_lut_4_lut_adj_1412.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1413 (.I0(\data_in_frame[17] [7]), .I1(n33583), 
            .I2(\data_in_frame[18] [2]), .I3(n34605), .O(n33247));
    defparam i3_4_lut_adj_1413.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1414 (.I0(n53), .I1(n3_adj_4430), .I2(\FRAME_MATCHER.state [16]), 
            .I3(GND_net), .O(n32291));
    defparam i1_2_lut_3_lut_adj_1414.LUT_INIT = 16'he0e0;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_31587 (.I0(byte_transmit_counter_c[1]), 
            .I1(n37282), .I2(n37283), .I3(byte_transmit_counter_c[2]), 
            .O(n38261));
    defparam byte_transmit_counter_1__bdd_4_lut_31587.LUT_INIT = 16'he4aa;
    SB_CARRY add_41_13 (.CI(n27919), .I0(\FRAME_MATCHER.i [11]), .I1(GND_net), 
            .CO(n27920));
    SB_DFF data_in_frame_0__i136 (.Q(\data_in_frame[16] [7]), .C(clk32MHz), 
           .D(n18145));   // verilog/coms.v(126[12] 293[6])
    SB_DFF data_in_frame_0__i135 (.Q(\data_in_frame[16] [6]), .C(clk32MHz), 
           .D(n18144));   // verilog/coms.v(126[12] 293[6])
    SB_LUT4 i1_2_lut_adj_1415 (.I0(\data_in_frame[1] [2]), .I1(\data_in_frame[1] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n16347));   // verilog/coms.v(72[16:34])
    defparam i1_2_lut_adj_1415.LUT_INIT = 16'h6666;
    SB_DFF data_in_frame_0__i134 (.Q(\data_in_frame[16] [5]), .C(clk32MHz), 
           .D(n18143));   // verilog/coms.v(126[12] 293[6])
    SB_LUT4 i1_2_lut_3_lut_adj_1416 (.I0(n53), .I1(n3_adj_4430), .I2(\FRAME_MATCHER.state [15]), 
            .I3(GND_net), .O(n32289));
    defparam i1_2_lut_3_lut_adj_1416.LUT_INIT = 16'he0e0;
    SB_LUT4 add_41_12_lut (.I0(n2290), .I1(\FRAME_MATCHER.i [10]), .I2(GND_net), 
            .I3(n27918), .O(n2_adj_4511)) /* synthesis syn_instantiated=1 */ ;
    defparam add_41_12_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i1_2_lut_3_lut_adj_1417 (.I0(\data_out_frame[5] [3]), .I1(\data_out_frame[5] [5]), 
            .I2(\data_out_frame[8] [0]), .I3(GND_net), .O(n33546));   // verilog/coms.v(70[16:27])
    defparam i1_2_lut_3_lut_adj_1417.LUT_INIT = 16'h9696;
    SB_CARRY add_41_12 (.CI(n27918), .I0(\FRAME_MATCHER.i [10]), .I1(GND_net), 
            .CO(n27919));
    SB_LUT4 add_41_11_lut (.I0(n2290), .I1(\FRAME_MATCHER.i [9]), .I2(GND_net), 
            .I3(n27917), .O(n2_adj_4509)) /* synthesis syn_instantiated=1 */ ;
    defparam add_41_11_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_41_11 (.CI(n27917), .I0(\FRAME_MATCHER.i [9]), .I1(GND_net), 
            .CO(n27918));
    SB_LUT4 i1_2_lut_3_lut_adj_1418 (.I0(n53), .I1(n3_adj_4430), .I2(\FRAME_MATCHER.state [14]), 
            .I3(GND_net), .O(n32287));
    defparam i1_2_lut_3_lut_adj_1418.LUT_INIT = 16'he0e0;
    SB_DFF \FRAME_MATCHER.state_i0  (.Q(\FRAME_MATCHER.state [0]), .C(clk32MHz), 
           .D(n34351));   // verilog/coms.v(126[12] 293[6])
    SB_LUT4 i1_2_lut_3_lut_adj_1419 (.I0(n53), .I1(n3_adj_4430), .I2(\FRAME_MATCHER.state [13]), 
            .I3(GND_net), .O(n32285));
    defparam i1_2_lut_3_lut_adj_1419.LUT_INIT = 16'he0e0;
    SB_LUT4 i2_2_lut_4_lut_adj_1420 (.I0(\data_in_frame[7] [7]), .I1(\data_in_frame[7] [6]), 
            .I2(\data_in_frame[10] [2]), .I3(\data_in_frame[6] [0]), .O(n10_adj_4372));   // verilog/coms.v(84[17:28])
    defparam i2_2_lut_4_lut_adj_1420.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1421 (.I0(\data_in_frame[7] [7]), .I1(\data_in_frame[7] [6]), 
            .I2(\data_in_frame[10] [2]), .I3(GND_net), .O(n33235));   // verilog/coms.v(84[17:28])
    defparam i1_2_lut_3_lut_adj_1421.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1422 (.I0(n53), .I1(n3_adj_4430), .I2(\FRAME_MATCHER.state [12]), 
            .I3(GND_net), .O(n32283));
    defparam i1_2_lut_3_lut_adj_1422.LUT_INIT = 16'he0e0;
    SB_DFF PWMLimit_i0_i0 (.Q(PWMLimit[0]), .C(clk32MHz), .D(n17696));   // verilog/coms.v(126[12] 293[6])
    SB_DFF data_in_frame_0__i1 (.Q(\data_in_frame[0] [0]), .C(clk32MHz), 
           .D(n17695));   // verilog/coms.v(126[12] 293[6])
    SB_DFF control_mode_i0_i0 (.Q(control_mode[0]), .C(clk32MHz), .D(n17694));   // verilog/coms.v(126[12] 293[6])
    SB_LUT4 i1_2_lut_3_lut_adj_1423 (.I0(\data_out_frame[11] [6]), .I1(n17182), 
            .I2(\data_out_frame[9] [6]), .I3(GND_net), .O(n6));   // verilog/coms.v(84[17:63])
    defparam i1_2_lut_3_lut_adj_1423.LUT_INIT = 16'h9696;
    SB_DFF setpoint__i0 (.Q(setpoint[0]), .C(clk32MHz), .D(n17693));   // verilog/coms.v(126[12] 293[6])
    SB_DFF Ki_i0 (.Q(\Ki[0] ), .C(clk32MHz), .D(n17692));   // verilog/coms.v(126[12] 293[6])
    SB_DFF Kp_i0 (.Q(\Kp[0] ), .C(clk32MHz), .D(n17691));   // verilog/coms.v(126[12] 293[6])
    SB_DFF data_in_0___i1 (.Q(\data_in[0][0] ), .C(clk32MHz), .D(n17690));   // verilog/coms.v(126[12] 293[6])
    SB_LUT4 i1_2_lut_3_lut_adj_1424 (.I0(n53), .I1(n3_adj_4430), .I2(\FRAME_MATCHER.state [11]), 
            .I3(GND_net), .O(n32281));
    defparam i1_2_lut_3_lut_adj_1424.LUT_INIT = 16'he0e0;
    SB_LUT4 i19300_2_lut_3_lut (.I0(n53), .I1(n3_adj_4430), .I2(\FRAME_MATCHER.state [10]), 
            .I3(GND_net), .O(n24108));
    defparam i19300_2_lut_3_lut.LUT_INIT = 16'he0e0;
    SB_LUT4 add_41_10_lut (.I0(n2290), .I1(\FRAME_MATCHER.i [8]), .I2(GND_net), 
            .I3(n27916), .O(n2_adj_4507)) /* synthesis syn_instantiated=1 */ ;
    defparam add_41_10_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i19299_2_lut_3_lut (.I0(n53), .I1(n3_adj_4430), .I2(\FRAME_MATCHER.state [9]), 
            .I3(GND_net), .O(n24106));
    defparam i19299_2_lut_3_lut.LUT_INIT = 16'he0e0;
    SB_CARRY add_41_10 (.CI(n27916), .I0(\FRAME_MATCHER.i [8]), .I1(GND_net), 
            .CO(n27917));
    SB_LUT4 add_41_9_lut (.I0(n2290), .I1(\FRAME_MATCHER.i [7]), .I2(GND_net), 
            .I3(n27915), .O(n2_adj_4505)) /* synthesis syn_instantiated=1 */ ;
    defparam add_41_9_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i31547_2_lut_3_lut (.I0(\FRAME_MATCHER.state [1]), .I1(\FRAME_MATCHER.state [2]), 
            .I2(\FRAME_MATCHER.state [0]), .I3(GND_net), .O(n17449));
    defparam i31547_2_lut_3_lut.LUT_INIT = 16'h0e0e;
    SB_LUT4 i1_2_lut_4_lut_adj_1425 (.I0(n33020), .I1(n33371), .I2(\data_out_frame[20] [6]), 
            .I3(n33201), .O(n33202));
    defparam i1_2_lut_4_lut_adj_1425.LUT_INIT = 16'h9669;
    SB_LUT4 i19298_2_lut_3_lut (.I0(n53), .I1(n3_adj_4430), .I2(\FRAME_MATCHER.state [8]), 
            .I3(GND_net), .O(n24104));
    defparam i19298_2_lut_3_lut.LUT_INIT = 16'he0e0;
    SB_LUT4 i4_4_lut_4_lut (.I0(n16153), .I1(n16158), .I2(n63), .I3(n16090), 
            .O(n2958));
    defparam i4_4_lut_4_lut.LUT_INIT = 16'h80a0;
    SB_LUT4 i2_2_lut_4_lut_adj_1426 (.I0(\data_out_frame[11] [5]), .I1(n33576), 
            .I2(n16548), .I3(n17068), .O(n10_adj_4346));
    defparam i2_2_lut_4_lut_adj_1426.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1427 (.I0(n53), .I1(n3_adj_4430), .I2(\FRAME_MATCHER.state [7]), 
            .I3(GND_net), .O(n7_adj_4556));
    defparam i1_2_lut_3_lut_adj_1427.LUT_INIT = 16'he0e0;
    SB_LUT4 i2_3_lut_4_lut_adj_1428 (.I0(\FRAME_MATCHER.state [2]), .I1(\FRAME_MATCHER.state [1]), 
            .I2(\FRAME_MATCHER.state [0]), .I3(n25118), .O(n5069));
    defparam i2_3_lut_4_lut_adj_1428.LUT_INIT = 16'hfffe;
    SB_LUT4 i9_4_lut_adj_1429 (.I0(n33220), .I1(Kp_23__N_1453), .I2(n16855), 
            .I3(n33474), .O(n23));
    defparam i9_4_lut_adj_1429.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1430 (.I0(n53), .I1(n3_adj_4430), .I2(\FRAME_MATCHER.state [6]), 
            .I3(GND_net), .O(n32279));
    defparam i1_2_lut_3_lut_adj_1430.LUT_INIT = 16'he0e0;
    SB_LUT4 i8_4_lut_adj_1431 (.I0(n33247), .I1(\data_in_frame[16] [6]), 
            .I2(\data_in_frame[17] [4]), .I3(\data_in_frame[16] [7]), .O(n22_adj_4613));
    defparam i8_4_lut_adj_1431.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1432 (.I0(n53), .I1(n3_adj_4430), .I2(\FRAME_MATCHER.state [5]), 
            .I3(GND_net), .O(n32277));
    defparam i1_2_lut_3_lut_adj_1432.LUT_INIT = 16'he0e0;
    SB_LUT4 n38261_bdd_4_lut (.I0(n38261), .I1(n17_adj_4443), .I2(n16_adj_4442), 
            .I3(byte_transmit_counter_c[2]), .O(n38264));
    defparam n38261_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i19297_2_lut_3_lut (.I0(n53), .I1(n3_adj_4430), .I2(\FRAME_MATCHER.state [4]), 
            .I3(GND_net), .O(n24102));
    defparam i19297_2_lut_3_lut.LUT_INIT = 16'he0e0;
    SB_LUT4 i2_3_lut_4_lut_adj_1433 (.I0(\data_out_frame[13] [7]), .I1(n10_adj_4342), 
            .I2(\data_out_frame[15] [7]), .I3(GND_net), .O(n33601));
    defparam i2_3_lut_4_lut_adj_1433.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1434 (.I0(\data_in[3][7] ), .I1(\data_in[0][5] ), 
            .I2(n22269), .I3(GND_net), .O(n4_adj_4469));
    defparam i1_2_lut_3_lut_adj_1434.LUT_INIT = 16'hfbfb;
    SB_LUT4 i2_3_lut_4_lut_adj_1435 (.I0(\data_out_frame[7] [1]), .I1(\data_out_frame[7] [2]), 
            .I2(\data_out_frame[6] [7]), .I3(\data_out_frame[5] [1]), .O(n1251));   // verilog/coms.v(84[17:70])
    defparam i2_3_lut_4_lut_adj_1435.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1436 (.I0(\data_in_frame[1] [3]), .I1(n33354), 
            .I2(GND_net), .I3(GND_net), .O(n33094));   // verilog/coms.v(95[12:25])
    defparam i1_2_lut_adj_1436.LUT_INIT = 16'h6666;
    SB_LUT4 i12_4_lut_adj_1437 (.I0(n23), .I1(n19_adj_4575), .I2(n35410), 
            .I3(n17042), .O(n26_adj_4614));
    defparam i12_4_lut_adj_1437.LUT_INIT = 16'h9669;
    SB_LUT4 i2_3_lut_4_lut_adj_1438 (.I0(\data_in[3][7] ), .I1(\data_in[0][5] ), 
            .I2(n158), .I3(n22275), .O(n118));
    defparam i2_3_lut_4_lut_adj_1438.LUT_INIT = 16'hfffb;
    SB_LUT4 i30763_2_lut_4_lut (.I0(byte_transmit_counter[0]), .I1(byte_transmit_counter_c[2]), 
            .I2(byte_transmit_counter_c[1]), .I3(\data_out_frame[24] [1]), 
            .O(n37257));   // verilog/coms.v(105[34:55])
    defparam i30763_2_lut_4_lut.LUT_INIT = 16'h0100;
    SB_LUT4 i30752_2_lut_4_lut (.I0(byte_transmit_counter[0]), .I1(byte_transmit_counter_c[2]), 
            .I2(byte_transmit_counter_c[1]), .I3(\data_out_frame[24] [2]), 
            .O(n37266));   // verilog/coms.v(105[34:55])
    defparam i30752_2_lut_4_lut.LUT_INIT = 16'h0100;
    SB_LUT4 i1_2_lut_4_lut_adj_1439 (.I0(n1301), .I1(n33107), .I2(\data_out_frame[6] [4]), 
            .I3(n16672), .O(n33253));   // verilog/coms.v(75[16:27])
    defparam i1_2_lut_4_lut_adj_1439.LUT_INIT = 16'h6996;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_31582 (.I0(byte_transmit_counter_c[1]), 
            .I1(n37291), .I2(n37292), .I3(byte_transmit_counter_c[2]), 
            .O(n38255));
    defparam byte_transmit_counter_1__bdd_4_lut_31582.LUT_INIT = 16'he4aa;
    SB_LUT4 i13_4_lut_adj_1440 (.I0(n16435), .I1(n26_adj_4614), .I2(n22_adj_4613), 
            .I3(\data_in_frame[18] [3]), .O(n31168));
    defparam i13_4_lut_adj_1440.LUT_INIT = 16'h6996;
    SB_LUT4 i30868_2_lut_4_lut (.I0(byte_transmit_counter[0]), .I1(byte_transmit_counter_c[2]), 
            .I2(byte_transmit_counter_c[1]), .I3(\data_out_frame[24] [3]), 
            .O(n37269));   // verilog/coms.v(105[34:55])
    defparam i30868_2_lut_4_lut.LUT_INIT = 16'h0100;
    SB_LUT4 i30864_2_lut_4_lut (.I0(byte_transmit_counter[0]), .I1(byte_transmit_counter_c[2]), 
            .I2(byte_transmit_counter_c[1]), .I3(\data_out_frame[24] [4]), 
            .O(n37272));   // verilog/coms.v(105[34:55])
    defparam i30864_2_lut_4_lut.LUT_INIT = 16'h0100;
    SB_LUT4 i1_2_lut_4_lut_adj_1441 (.I0(n1301), .I1(n33107), .I2(\data_out_frame[6] [4]), 
            .I3(n33042), .O(n6_adj_4472));   // verilog/coms.v(75[16:27])
    defparam i1_2_lut_4_lut_adj_1441.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1442 (.I0(\data_in_frame[4] [7]), .I1(\data_in_frame[7] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n33316));
    defparam i1_2_lut_adj_1442.LUT_INIT = 16'h6666;
    SB_CARRY add_41_9 (.CI(n27915), .I0(\FRAME_MATCHER.i [7]), .I1(GND_net), 
            .CO(n27916));
    SB_LUT4 add_41_8_lut (.I0(n2290), .I1(\FRAME_MATCHER.i [6]), .I2(GND_net), 
            .I3(n27914), .O(n2_adj_4503)) /* synthesis syn_instantiated=1 */ ;
    defparam add_41_8_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i2_2_lut_adj_1443 (.I0(n33558), .I1(\data_in_frame[3] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n10_adj_4615));   // verilog/coms.v(95[12:25])
    defparam i2_2_lut_adj_1443.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1444 (.I0(n30241), .I1(\data_out_frame[13] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n31188));
    defparam i1_2_lut_adj_1444.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_4_lut_adj_1445 (.I0(\data_out_frame[13] [1]), .I1(\data_out_frame[13] [7]), 
            .I2(n10_adj_4342), .I3(\data_out_frame[15] [7]), .O(n6_adj_4343));
    defparam i1_2_lut_4_lut_adj_1445.LUT_INIT = 16'h6996;
    SB_CARRY add_41_8 (.CI(n27914), .I0(\FRAME_MATCHER.i [6]), .I1(GND_net), 
            .CO(n27915));
    SB_LUT4 add_41_7_lut (.I0(n2290), .I1(\FRAME_MATCHER.i [5]), .I2(GND_net), 
            .I3(n27913), .O(n2_adj_4501)) /* synthesis syn_instantiated=1 */ ;
    defparam add_41_7_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i30859_2_lut_4_lut (.I0(byte_transmit_counter[0]), .I1(byte_transmit_counter_c[2]), 
            .I2(byte_transmit_counter_c[1]), .I3(\data_out_frame[24] [5]), 
            .O(n37275));   // verilog/coms.v(105[34:55])
    defparam i30859_2_lut_4_lut.LUT_INIT = 16'h0100;
    SB_LUT4 i2_3_lut_4_lut_adj_1446 (.I0(\data_out_frame[7] [0]), .I1(\data_out_frame[6] [7]), 
            .I2(\data_out_frame[6] [6]), .I3(n17182), .O(n15783));
    defparam i2_3_lut_4_lut_adj_1446.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_adj_1447 (.I0(\data_out_frame[7] [2]), .I1(\data_out_frame[5] [2]), 
            .I2(\data_out_frame[5] [0]), .I3(\data_out_frame[7] [3]), .O(n1254));
    defparam i1_2_lut_4_lut_adj_1447.LUT_INIT = 16'h6996;
    SB_LUT4 i30857_2_lut_4_lut (.I0(byte_transmit_counter[0]), .I1(byte_transmit_counter_c[2]), 
            .I2(byte_transmit_counter_c[1]), .I3(\data_out_frame[24] [6]), 
            .O(n37278));   // verilog/coms.v(105[34:55])
    defparam i30857_2_lut_4_lut.LUT_INIT = 16'h0100;
    SB_LUT4 i1_2_lut_adj_1448 (.I0(\data_in_frame[13] [5]), .I1(\data_in_frame[15] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n33295));
    defparam i1_2_lut_adj_1448.LUT_INIT = 16'h6666;
    SB_LUT4 i30852_2_lut_4_lut (.I0(byte_transmit_counter[0]), .I1(byte_transmit_counter_c[2]), 
            .I2(byte_transmit_counter_c[1]), .I3(\data_out_frame[24] [7]), 
            .O(n37281));   // verilog/coms.v(105[34:55])
    defparam i30852_2_lut_4_lut.LUT_INIT = 16'h0100;
    SB_LUT4 i6_4_lut_adj_1449 (.I0(n33604), .I1(n33094), .I2(n33403), 
            .I3(\data_in_frame[0] [3]), .O(n14_adj_4616));   // verilog/coms.v(95[12:25])
    defparam i6_4_lut_adj_1449.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1450 (.I0(n16413), .I1(n33421), .I2(\data_in_frame[12] [7]), 
            .I3(GND_net), .O(n17004));   // verilog/coms.v(70[16:27])
    defparam i2_3_lut_adj_1450.LUT_INIT = 16'h9696;
    SB_LUT4 i30714_2_lut_4_lut (.I0(byte_transmit_counter[0]), .I1(byte_transmit_counter_c[2]), 
            .I2(byte_transmit_counter_c[1]), .I3(\data_out_frame[24] [0]), 
            .O(n37290));   // verilog/coms.v(105[34:55])
    defparam i30714_2_lut_4_lut.LUT_INIT = 16'h0100;
    SB_LUT4 i5_4_lut_adj_1451 (.I0(n17004), .I1(n33295), .I2(n16179), 
            .I3(n31168), .O(n12_adj_4617));
    defparam i5_4_lut_adj_1451.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut_adj_1452 (.I0(\data_in_frame[2] [6]), .I1(n14_adj_4616), 
            .I2(n10_adj_4615), .I3(n33232), .O(n30900));   // verilog/coms.v(95[12:25])
    defparam i7_4_lut_adj_1452.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_1453 (.I0(n17132), .I1(n12_adj_4617), .I2(n33491), 
            .I3(n17042), .O(n34730));
    defparam i6_4_lut_adj_1453.LUT_INIT = 16'h6996;
    SB_CARRY add_41_7 (.CI(n27913), .I0(\FRAME_MATCHER.i [5]), .I1(GND_net), 
            .CO(n27914));
    SB_LUT4 i23023_2_lut_4_lut (.I0(n16158), .I1(n4_adj_4403), .I2(n7_adj_4402), 
            .I3(\FRAME_MATCHER.state [31]), .O(n29607));   // verilog/coms.v(114[11:12])
    defparam i23023_2_lut_4_lut.LUT_INIT = 16'hdc00;
    SB_LUT4 add_41_6_lut (.I0(n2290), .I1(\FRAME_MATCHER.i [4]), .I2(GND_net), 
            .I3(n27912), .O(n2_adj_4499)) /* synthesis syn_instantiated=1 */ ;
    defparam add_41_6_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i23026_2_lut_4_lut (.I0(n16158), .I1(n4_adj_4403), .I2(n7_adj_4402), 
            .I3(\FRAME_MATCHER.state [30]), .O(n29613));   // verilog/coms.v(114[11:12])
    defparam i23026_2_lut_4_lut.LUT_INIT = 16'hdc00;
    SB_DFF byte_transmit_counter_i0_i7 (.Q(byte_transmit_counter_c[7]), .C(clk32MHz), 
           .D(n17658));   // verilog/coms.v(126[12] 293[6])
    SB_LUT4 i23024_2_lut_4_lut (.I0(n16158), .I1(n4_adj_4403), .I2(n7_adj_4402), 
            .I3(\FRAME_MATCHER.state [29]), .O(n29609));   // verilog/coms.v(114[11:12])
    defparam i23024_2_lut_4_lut.LUT_INIT = 16'hdc00;
    SB_DFF byte_transmit_counter_i0_i6 (.Q(byte_transmit_counter_c[6]), .C(clk32MHz), 
           .D(n17661));   // verilog/coms.v(126[12] 293[6])
    SB_LUT4 i23025_2_lut_4_lut (.I0(n16158), .I1(n4_adj_4403), .I2(n7_adj_4402), 
            .I3(\FRAME_MATCHER.state [27]), .O(n29611));   // verilog/coms.v(114[11:12])
    defparam i23025_2_lut_4_lut.LUT_INIT = 16'hdc00;
    SB_DFF byte_transmit_counter_i0_i5 (.Q(byte_transmit_counter_c[5]), .C(clk32MHz), 
           .D(n17664));   // verilog/coms.v(126[12] 293[6])
    SB_DFF byte_transmit_counter_i0_i4 (.Q(byte_transmit_counter_c[4]), .C(clk32MHz), 
           .D(n17667));   // verilog/coms.v(126[12] 293[6])
    SB_LUT4 i23022_2_lut_4_lut (.I0(n16158), .I1(n4_adj_4403), .I2(n7_adj_4402), 
            .I3(\FRAME_MATCHER.state [23]), .O(n29605));   // verilog/coms.v(114[11:12])
    defparam i23022_2_lut_4_lut.LUT_INIT = 16'hdc00;
    SB_DFF byte_transmit_counter_i0_i3 (.Q(byte_transmit_counter_c[3]), .C(clk32MHz), 
           .D(n17670));   // verilog/coms.v(126[12] 293[6])
    SB_LUT4 i13229_3_lut_4_lut (.I0(n8_adj_4355), .I1(n32959), .I2(rx_data[0]), 
            .I3(\data_in_frame[6] [0]), .O(n18058));
    defparam i13229_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13343_3_lut_4_lut (.I0(n8_adj_4353), .I1(n32952), .I2(rx_data[2]), 
            .I3(\data_in_frame[20] [2]), .O(n18172));
    defparam i13343_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF byte_transmit_counter_i0_i2 (.Q(byte_transmit_counter_c[2]), .C(clk32MHz), 
           .D(n17673));   // verilog/coms.v(126[12] 293[6])
    SB_DFF byte_transmit_counter_i0_i1 (.Q(byte_transmit_counter_c[1]), .C(clk32MHz), 
           .D(n17676));   // verilog/coms.v(126[12] 293[6])
    SB_DFF byte_transmit_counter_i0_i0 (.Q(byte_transmit_counter[0]), .C(clk32MHz), 
           .D(n17731));   // verilog/coms.v(126[12] 293[6])
    SB_LUT4 i13230_3_lut_4_lut (.I0(n8_adj_4355), .I1(n32959), .I2(rx_data[1]), 
            .I3(\data_in_frame[6] [1]), .O(n18059));
    defparam i13230_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_1454 (.I0(\data_in_frame[16] [3]), .I1(Kp_23__N_843), 
            .I2(GND_net), .I3(GND_net), .O(n16179));
    defparam i1_2_lut_adj_1454.LUT_INIT = 16'h6666;
    SB_LUT4 i13342_3_lut_4_lut (.I0(n8_adj_4353), .I1(n32952), .I2(rx_data[1]), 
            .I3(\data_in_frame[20] [1]), .O(n18171));
    defparam i13342_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF data_in_frame_0__i117 (.Q(\data_in_frame[14] [4]), .C(clk32MHz), 
           .D(n18126));   // verilog/coms.v(126[12] 293[6])
    SB_LUT4 n38255_bdd_4_lut (.I0(n38255), .I1(n17_adj_4379), .I2(n16_adj_4378), 
            .I3(byte_transmit_counter_c[2]), .O(n38258));
    defparam n38255_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_CARRY add_41_6 (.CI(n27912), .I0(\FRAME_MATCHER.i [4]), .I1(GND_net), 
            .CO(n27913));
    SB_DFF data_in_frame_0__i72 (.Q(\data_in_frame[8] [7]), .C(clk32MHz), 
           .D(n18081));   // verilog/coms.v(126[12] 293[6])
    SB_LUT4 add_41_5_lut (.I0(n2290), .I1(\FRAME_MATCHER.i [3]), .I2(GND_net), 
            .I3(n27911), .O(n2_adj_4497)) /* synthesis syn_instantiated=1 */ ;
    defparam add_41_5_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i13341_3_lut_4_lut (.I0(n8_adj_4353), .I1(n32952), .I2(rx_data[0]), 
            .I3(\data_in_frame[20] [0]), .O(n18170));
    defparam i13341_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_CARRY add_41_5 (.CI(n27911), .I0(\FRAME_MATCHER.i [3]), .I1(GND_net), 
            .CO(n27912));
    SB_LUT4 i13231_3_lut_4_lut (.I0(n8_adj_4355), .I1(n32959), .I2(rx_data[2]), 
            .I3(\data_in_frame[6] [2]), .O(n18060));
    defparam i13231_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13345_3_lut_4_lut (.I0(n8_adj_4353), .I1(n32952), .I2(rx_data[4]), 
            .I3(\data_in_frame[20] [4]), .O(n18174));
    defparam i13345_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13344_3_lut_4_lut (.I0(n8_adj_4353), .I1(n32952), .I2(rx_data[3]), 
            .I3(\data_in_frame[20] [3]), .O(n18173));
    defparam i13344_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_3_lut_adj_1455 (.I0(\data_out_frame[9] [3]), .I1(\data_out_frame[11] [5]), 
            .I2(\data_out_frame[9] [4]), .I3(GND_net), .O(n33256));   // verilog/coms.v(84[17:63])
    defparam i2_3_lut_adj_1455.LUT_INIT = 16'h9696;
    SB_LUT4 i13347_3_lut_4_lut (.I0(n8_adj_4353), .I1(n32952), .I2(rx_data[6]), 
            .I3(\data_in_frame[20] [6]), .O(n18176));
    defparam i13347_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i3_4_lut_adj_1456 (.I0(n16335), .I1(\data_in_frame[12] [1]), 
            .I2(\data_in_frame[11] [7]), .I3(n33259), .O(n33592));   // verilog/coms.v(78[16:35])
    defparam i3_4_lut_adj_1456.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1457 (.I0(\data_in_frame[18] [5]), .I1(\data_in_frame[16] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n33220));
    defparam i1_2_lut_adj_1457.LUT_INIT = 16'h6666;
    SB_LUT4 i13346_3_lut_4_lut (.I0(n8_adj_4353), .I1(n32952), .I2(rx_data[5]), 
            .I3(\data_in_frame[20] [5]), .O(n18175));
    defparam i13346_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i3_4_lut_adj_1458 (.I0(\data_in_frame[4] [1]), .I1(n33232), 
            .I2(\data_in_frame[2] [0]), .I3(\data_in_frame[3] [7]), .O(n16765));   // verilog/coms.v(71[16:41])
    defparam i3_4_lut_adj_1458.LUT_INIT = 16'h6996;
    SB_LUT4 i5_4_lut_adj_1459 (.I0(\data_in_frame[10] [0]), .I1(n33500), 
            .I2(\data_in_frame[9] [5]), .I3(\data_in_frame[7] [5]), .O(n12_adj_4618));
    defparam i5_4_lut_adj_1459.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1460 (.I0(\data_out_frame[7] [5]), .I1(\data_out_frame[5] [4]), 
            .I2(\data_out_frame[5] [3]), .I3(GND_net), .O(n16687));   // verilog/coms.v(75[16:43])
    defparam i1_2_lut_3_lut_adj_1460.LUT_INIT = 16'h9696;
    SB_LUT4 i13348_3_lut_4_lut (.I0(n8_adj_4353), .I1(n32952), .I2(rx_data[7]), 
            .I3(\data_in_frame[20] [7]), .O(n18177));
    defparam i13348_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_3_lut_adj_1461 (.I0(n16314), .I1(\data_in_frame[14] [5]), 
            .I2(n16780), .I3(GND_net), .O(n6_adj_4609));
    defparam i1_2_lut_3_lut_adj_1461.LUT_INIT = 16'h9696;
    SB_LUT4 i6_4_lut_adj_1462 (.I0(\data_in_frame[9] [7]), .I1(n12_adj_4618), 
            .I2(n33592), .I3(\data_in_frame[7] [6]), .O(n35345));
    defparam i6_4_lut_adj_1462.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_1463 (.I0(n16314), .I1(\data_in_frame[14] [5]), 
            .I2(n30694), .I3(\data_in_frame[14] [4]), .O(n34514));
    defparam i2_3_lut_4_lut_adj_1463.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1464 (.I0(\data_in_frame[10] [4]), .I1(Kp_23__N_1046), 
            .I2(GND_net), .I3(GND_net), .O(n33555));   // verilog/coms.v(84[17:28])
    defparam i1_2_lut_adj_1464.LUT_INIT = 16'h6666;
    SB_LUT4 add_41_4_lut (.I0(n2290), .I1(\FRAME_MATCHER.i [2]), .I2(GND_net), 
            .I3(n27910), .O(n2_adj_4495)) /* synthesis syn_instantiated=1 */ ;
    defparam add_41_4_lut.LUT_INIT = 16'h8228;
    SB_DFF data_in_frame_0__i71 (.Q(\data_in_frame[8] [6]), .C(clk32MHz), 
           .D(n18080));   // verilog/coms.v(126[12] 293[6])
    SB_LUT4 i2_3_lut_4_lut_adj_1465 (.I0(\data_in_frame[14] [3]), .I1(n35345), 
            .I2(\data_in_frame[14] [4]), .I3(n16780), .O(n31257));
    defparam i2_3_lut_4_lut_adj_1465.LUT_INIT = 16'h9669;
    SB_LUT4 i4_4_lut_adj_1466 (.I0(\data_in_frame[6] [0]), .I1(n33007), 
            .I2(n33397), .I3(n6_adj_4565), .O(n16466));   // verilog/coms.v(84[17:28])
    defparam i4_4_lut_adj_1466.LUT_INIT = 16'h6996;
    SB_DFF data_in_frame_0__i133 (.Q(\data_in_frame[16] [4]), .C(clk32MHz), 
           .D(n18142));   // verilog/coms.v(126[12] 293[6])
    SB_LUT4 i1_2_lut_adj_1467 (.I0(\data_in_frame[5] [7]), .I1(\data_in_frame[8] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n33007));   // verilog/coms.v(84[17:28])
    defparam i1_2_lut_adj_1467.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1468 (.I0(\data_in_frame[7] [5]), .I1(\data_in_frame[10] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n16233));
    defparam i1_2_lut_adj_1468.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1469 (.I0(\data_in_frame[17] [0]), .I1(\data_in_frame[17] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n33474));
    defparam i1_2_lut_adj_1469.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_4_lut_adj_1470 (.I0(\data_in_frame[14] [3]), .I1(n35345), 
            .I2(n30694), .I3(n16620), .O(n33335));
    defparam i2_3_lut_4_lut_adj_1470.LUT_INIT = 16'h9669;
    SB_DFF data_in_frame_0__i132 (.Q(\data_in_frame[16] [3]), .C(clk32MHz), 
           .D(n18141));   // verilog/coms.v(126[12] 293[6])
    SB_DFF data_in_frame_0__i131 (.Q(\data_in_frame[16] [2]), .C(clk32MHz), 
           .D(n18140));   // verilog/coms.v(126[12] 293[6])
    SB_DFF data_in_frame_0__i130 (.Q(\data_in_frame[16] [1]), .C(clk32MHz), 
           .D(n18139));   // verilog/coms.v(126[12] 293[6])
    SB_DFF data_in_frame_0__i129 (.Q(\data_in_frame[16] [0]), .C(clk32MHz), 
           .D(n18138));   // verilog/coms.v(126[12] 293[6])
    SB_LUT4 i1_2_lut_3_lut_adj_1471 (.I0(\data_out_frame[5] [3]), .I1(\data_out_frame[5] [2]), 
            .I2(\data_out_frame[7] [4]), .I3(GND_net), .O(n16163));   // verilog/coms.v(75[16:43])
    defparam i1_2_lut_3_lut_adj_1471.LUT_INIT = 16'h9696;
    SB_LUT4 i6_4_lut_adj_1472 (.I0(n33532), .I1(\data_in_frame[1] [4]), 
            .I2(n33007), .I3(\data_in_frame[8] [4]), .O(n14));   // verilog/coms.v(72[16:42])
    defparam i6_4_lut_adj_1472.LUT_INIT = 16'h6996;
    SB_LUT4 i13221_3_lut_4_lut (.I0(n8), .I1(n32959), .I2(rx_data[0]), 
            .I3(\data_in_frame[5] [0]), .O(n18050));
    defparam i13221_3_lut_4_lut.LUT_INIT = 16'hfe10;
    uart_tx tx (.clk32MHz(clk32MHz), .tx_data({tx_data}), .\r_SM_Main[2] (\r_SM_Main[2] ), 
            .GND_net(GND_net), .r_Bit_Index({r_Bit_Index}), .n17362(n17362), 
            .n17534(n17534), .n5600(n5600), .\r_Clock_Count[6] (\r_Clock_Count[6] ), 
            .\r_Clock_Count[7] (\r_Clock_Count[7] ), .\r_Clock_Count[8] (\r_Clock_Count[8] ), 
            .\r_Clock_Count[0] (\r_Clock_Count[0] ), .\r_Clock_Count[3] (\r_Clock_Count[3] ), 
            .n313(n313), .n314(n314), .n315(n315), .n316(n316), .\r_Clock_Count[5] (\r_Clock_Count[5] ), 
            .tx_active(tx_active), .\r_SM_Main_2__N_3458[0] (\r_SM_Main_2__N_3458[0] ), 
            .n5478(n5478), .n318(n318), .n321(n321), .VCC_net(VCC_net), 
            .tx_o(tx_o), .tx_enable(tx_enable), .n17559(n17559), .tx_transmit_N_3355(tx_transmit_N_3355), 
            .n1502(n1502), .n63(n63), .n16157(n16157), .n25050(n25050), 
            .\byte_transmit_counter[4] (byte_transmit_counter_c[4]), .\byte_transmit_counter[3] (byte_transmit_counter_c[3]), 
            .n7(n7), .n18278(n18278), .n17652(n17652), .n17655(n17655), 
            .n17708(n17708), .n17713(n17713), .n17728(n17728), .n17549(n17549), 
            .n17553(n17553)) /* synthesis lattice_noprune=1, syn_preserve=0, syn_module_defined=1, syn_noprune=0 */ ;   // verilog/coms.v(106[10:70])
    uart_rx rx (.n25112(n25112), .r_SM_Main({Open_7, \r_SM_Main[1] , Open_8}), 
            .clk32MHz(clk32MHz), .VCC_net(VCC_net), .rx_data_ready(rx_data_ready), 
            .n18260(n18260), .rx_data({rx_data}), .r_Rx_Data(r_Rx_Data), 
            .n37332(n37332), .GND_net(GND_net), .PIN_13_N_105(PIN_13_N_105), 
            .\r_SM_Main[2] (\r_SM_Main[2]_adj_3 ), .n33769(n33769), .n17681(n17681), 
            .r_Bit_Index({r_Bit_Index_adj_10}), .n5578(n5578), .n24193(n24193), 
            .n4(n4_adj_7), .n4_adj_1(n4_adj_8), .n16148(n16148), .n25070(n25070), 
            .n1(n1), .n37333(n37333), .n17701(n17701), .n17689(n17689), 
            .n17688(n17688), .n17687(n17687), .n17686(n17686), .n17685(n17685), 
            .n17684(n17684), .n17683(n17683), .n16143(n16143), .n17679(n17679), 
            .n17682(n17682), .n17735(n17735), .n4_adj_2(n4_adj_9)) /* synthesis lattice_noprune=1, syn_preserve=0, syn_module_defined=1, syn_noprune=0 */ ;   // verilog/coms.v(92[10:44])
    
endmodule
//
// Verilog Description of module uart_tx
//

module uart_tx (clk32MHz, tx_data, \r_SM_Main[2] , GND_net, r_Bit_Index, 
            n17362, n17534, n5600, \r_Clock_Count[6] , \r_Clock_Count[7] , 
            \r_Clock_Count[8] , \r_Clock_Count[0] , \r_Clock_Count[3] , 
            n313, n314, n315, n316, \r_Clock_Count[5] , tx_active, 
            \r_SM_Main_2__N_3458[0] , n5478, n318, n321, VCC_net, 
            tx_o, tx_enable, n17559, tx_transmit_N_3355, n1502, n63, 
            n16157, n25050, \byte_transmit_counter[4] , \byte_transmit_counter[3] , 
            n7, n18278, n17652, n17655, n17708, n17713, n17728, 
            n17549, n17553) /* synthesis lattice_noprune=1, syn_preserve=0, syn_module_defined=1, syn_noprune=0 */ ;
    input clk32MHz;
    input [7:0]tx_data;
    output \r_SM_Main[2] ;
    input GND_net;
    output [2:0]r_Bit_Index;
    output n17362;
    output n17534;
    output n5600;
    output \r_Clock_Count[6] ;
    output \r_Clock_Count[7] ;
    output \r_Clock_Count[8] ;
    output \r_Clock_Count[0] ;
    output \r_Clock_Count[3] ;
    output n313;
    output n314;
    output n315;
    output n316;
    output \r_Clock_Count[5] ;
    output tx_active;
    input \r_SM_Main_2__N_3458[0] ;
    output n5478;
    output n318;
    output n321;
    input VCC_net;
    output tx_o;
    output tx_enable;
    input n17559;
    input tx_transmit_N_3355;
    output n1502;
    input n63;
    input n16157;
    output n25050;
    input \byte_transmit_counter[4] ;
    input \byte_transmit_counter[3] ;
    output n7;
    input n18278;
    input n17652;
    input n17655;
    input n17708;
    input n17713;
    input n17728;
    input n17549;
    input n17553;
    
    wire clk32MHz /* synthesis SET_AS_NETWORK=clk32MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(34[6:14])
    
    wire n32645;
    wire [2:0]r_SM_Main;   // verilog/uart_tx.v(31[16:25])
    
    wire n13717;
    wire [7:0]r_Tx_Data;   // verilog/uart_tx.v(34[16:25])
    wire [8:0]r_Clock_Count;   // verilog/uart_tx.v(32[16:29])
    
    wire n37307, n32443, n18, n37331, n38360, n38300, n2, n33833, 
        n24692, n19424, n12;
    wire [2:0]r_SM_Main_2__N_3455;
    
    wire n24489, n10, n28039, n28038, n28037, n28036, n28035, 
        n79, n34119, n4, n17282, n17703, n19438;
    wire [2:0]r_SM_Main_2__N_3426;
    
    wire n37306, n32445;
    wire [8:0]n312;
    
    wire n17732, n38429, n38432, n38357, n28034, n28033, n28032, 
        n38297;
    
    SB_DFF r_SM_Main_i1 (.Q(r_SM_Main[1]), .C(clk32MHz), .D(n32645));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFE r_Tx_Data_i0 (.Q(r_Tx_Data[0]), .C(clk32MHz), .E(n13717), 
            .D(tx_data[0]));   // verilog/uart_tx.v(40[10] 143[8])
    SB_LUT4 i25_3_lut (.I0(r_Clock_Count[4]), .I1(n37307), .I2(\r_SM_Main[2] ), 
            .I3(GND_net), .O(n32443));
    defparam i25_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i19873_2_lut (.I0(r_SM_Main[0]), .I1(\r_SM_Main[2] ), .I2(GND_net), 
            .I3(GND_net), .O(n18));
    defparam i19873_2_lut.LUT_INIT = 16'h1111;
    SB_LUT4 i30839_2_lut (.I0(r_SM_Main[0]), .I1(\r_SM_Main[2] ), .I2(GND_net), 
            .I3(GND_net), .O(n37331));
    defparam i30839_2_lut.LUT_INIT = 16'hdddd;
    SB_LUT4 i19537_4_lut (.I0(n38360), .I1(r_SM_Main[0]), .I2(n38300), 
            .I3(r_Bit_Index[2]), .O(n2));   // verilog/uart_tx.v(43[7] 142[14])
    defparam i19537_4_lut.LUT_INIT = 16'hfcee;
    SB_LUT4 i27236_2_lut (.I0(r_SM_Main[1]), .I1(r_SM_Main[0]), .I2(GND_net), 
            .I3(GND_net), .O(n33833));
    defparam i27236_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i1_4_lut (.I0(\r_SM_Main[2] ), .I1(n24692), .I2(n19424), .I3(n33833), 
            .O(n12));
    defparam i1_4_lut.LUT_INIT = 16'habaa;
    SB_LUT4 i2_4_lut (.I0(r_SM_Main[0]), .I1(\r_SM_Main[2] ), .I2(r_SM_Main[1]), 
            .I3(r_SM_Main_2__N_3455[1]), .O(n17362));
    defparam i2_4_lut.LUT_INIT = 16'h1101;
    SB_LUT4 i12705_3_lut (.I0(n17362), .I1(r_SM_Main[1]), .I2(n24489), 
            .I3(GND_net), .O(n17534));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i12705_3_lut.LUT_INIT = 16'ha2a2;
    SB_LUT4 i1814_2_lut (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[0]), .I2(GND_net), 
            .I3(GND_net), .O(n5600));   // verilog/uart_tx.v(98[36:51])
    defparam i1814_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i2_3_lut (.I0(\r_Clock_Count[6] ), .I1(\r_Clock_Count[7] ), 
            .I2(\r_Clock_Count[8] ), .I3(GND_net), .O(n24692));
    defparam i2_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i5_3_lut (.I0(\r_Clock_Count[0] ), .I1(n10), .I2(\r_Clock_Count[3] ), 
            .I3(GND_net), .O(n19424));   // verilog/uart_tx.v(32[16:29])
    defparam i5_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 add_59_10_lut (.I0(GND_net), .I1(\r_Clock_Count[8] ), .I2(GND_net), 
            .I3(n28039), .O(n313)) /* synthesis syn_instantiated=1 */ ;
    defparam add_59_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_59_9_lut (.I0(GND_net), .I1(\r_Clock_Count[7] ), .I2(GND_net), 
            .I3(n28038), .O(n314)) /* synthesis syn_instantiated=1 */ ;
    defparam add_59_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_59_9 (.CI(n28038), .I0(\r_Clock_Count[7] ), .I1(GND_net), 
            .CO(n28039));
    SB_LUT4 add_59_8_lut (.I0(GND_net), .I1(\r_Clock_Count[6] ), .I2(GND_net), 
            .I3(n28037), .O(n315)) /* synthesis syn_instantiated=1 */ ;
    defparam add_59_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_59_8 (.CI(n28037), .I0(\r_Clock_Count[6] ), .I1(GND_net), 
            .CO(n28038));
    SB_LUT4 add_59_7_lut (.I0(GND_net), .I1(\r_Clock_Count[5] ), .I2(GND_net), 
            .I3(n28036), .O(n316)) /* synthesis syn_instantiated=1 */ ;
    defparam add_59_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_59_7 (.CI(n28036), .I0(\r_Clock_Count[5] ), .I1(GND_net), 
            .CO(n28037));
    SB_LUT4 add_59_6_lut (.I0(n12), .I1(r_Clock_Count[4]), .I2(GND_net), 
            .I3(n28035), .O(n37307)) /* synthesis syn_instantiated=1 */ ;
    defparam add_59_6_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_59_6 (.CI(n28035), .I0(r_Clock_Count[4]), .I1(GND_net), 
            .CO(n28036));
    SB_LUT4 i2_3_lut_adj_869 (.I0(n79), .I1(r_SM_Main[1]), .I2(\r_SM_Main[2] ), 
            .I3(GND_net), .O(n34119));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i2_3_lut_adj_869.LUT_INIT = 16'h0808;
    SB_LUT4 i2_4_lut_adj_870 (.I0(n4), .I1(\r_SM_Main[2] ), .I2(r_SM_Main[1]), 
            .I3(n79), .O(n17282));
    defparam i2_4_lut_adj_870.LUT_INIT = 16'h3202;
    SB_LUT4 i15244_3_lut (.I0(n17282), .I1(r_SM_Main[1]), .I2(tx_active), 
            .I3(GND_net), .O(n17703));   // verilog/uart_tx.v(31[16:25])
    defparam i15244_3_lut.LUT_INIT = 16'h7272;
    SB_LUT4 i2_3_lut_adj_871 (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[2]), 
            .I2(r_Bit_Index[0]), .I3(GND_net), .O(n24489));
    defparam i2_3_lut_adj_871.LUT_INIT = 16'h8080;
    SB_LUT4 i14610_4_lut (.I0(\r_SM_Main_2__N_3458[0] ), .I1(n24489), .I2(r_SM_Main[1]), 
            .I3(r_SM_Main_2__N_3455[1]), .O(n19438));   // verilog/uart_tx.v(31[16:25])
    defparam i14610_4_lut.LUT_INIT = 16'hca0a;
    SB_LUT4 i1_4_lut_adj_872 (.I0(\r_SM_Main[2] ), .I1(n19438), .I2(r_SM_Main_2__N_3455[1]), 
            .I3(r_SM_Main[0]), .O(r_SM_Main_2__N_3426[0]));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i1_4_lut_adj_872.LUT_INIT = 16'h0544;
    SB_LUT4 i25_3_lut_adj_873 (.I0(r_Clock_Count[1]), .I1(n37306), .I2(\r_SM_Main[2] ), 
            .I3(GND_net), .O(n32445));
    defparam i25_3_lut_adj_873.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_874 (.I0(n5478), .I1(r_Clock_Count[2]), .I2(n312[2]), 
            .I3(\r_SM_Main[2] ), .O(n17732));
    defparam i1_4_lut_adj_874.LUT_INIT = 16'h4450;
    SB_LUT4 n38429_bdd_4_lut (.I0(n38429), .I1(n37331), .I2(n18), .I3(r_SM_Main[1]), 
            .O(n38432));
    defparam n38429_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 r_Bit_Index_0__bdd_4_lut (.I0(r_Bit_Index[0]), .I1(r_Tx_Data[2]), 
            .I2(r_Tx_Data[3]), .I3(r_Bit_Index[1]), .O(n38357));
    defparam r_Bit_Index_0__bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_LUT4 add_59_5_lut (.I0(GND_net), .I1(\r_Clock_Count[3] ), .I2(GND_net), 
            .I3(n28034), .O(n318)) /* synthesis syn_instantiated=1 */ ;
    defparam add_59_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_59_5 (.CI(n28034), .I0(\r_Clock_Count[3] ), .I1(GND_net), 
            .CO(n28035));
    SB_LUT4 add_59_4_lut (.I0(GND_net), .I1(r_Clock_Count[2]), .I2(GND_net), 
            .I3(n28033), .O(n312[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_59_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_59_4 (.CI(n28033), .I0(r_Clock_Count[2]), .I1(GND_net), 
            .CO(n28034));
    SB_LUT4 add_59_3_lut (.I0(n12), .I1(r_Clock_Count[1]), .I2(GND_net), 
            .I3(n28032), .O(n37306)) /* synthesis syn_instantiated=1 */ ;
    defparam add_59_3_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_59_3 (.CI(n28032), .I0(r_Clock_Count[1]), .I1(GND_net), 
            .CO(n28033));
    SB_LUT4 add_59_2_lut (.I0(GND_net), .I1(\r_Clock_Count[0] ), .I2(GND_net), 
            .I3(VCC_net), .O(n321)) /* synthesis syn_instantiated=1 */ ;
    defparam add_59_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_59_2 (.CI(VCC_net), .I0(\r_Clock_Count[0] ), .I1(GND_net), 
            .CO(n28032));
    SB_LUT4 n38357_bdd_4_lut (.I0(n38357), .I1(r_Tx_Data[1]), .I2(r_Tx_Data[0]), 
            .I3(r_Bit_Index[1]), .O(n38360));
    defparam n38357_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i4_4_lut (.I0(r_Clock_Count[2]), .I1(r_Clock_Count[1]), .I2(r_Clock_Count[4]), 
            .I3(\r_Clock_Count[5] ), .O(n10));   // verilog/uart_tx.v(32[16:29])
    defparam i4_4_lut.LUT_INIT = 16'h8000;
    SB_DFFE r_Tx_Data_i1 (.Q(r_Tx_Data[1]), .C(clk32MHz), .E(n13717), 
            .D(tx_data[1]));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFE r_Tx_Data_i2 (.Q(r_Tx_Data[2]), .C(clk32MHz), .E(n13717), 
            .D(tx_data[2]));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFE r_Tx_Data_i3 (.Q(r_Tx_Data[3]), .C(clk32MHz), .E(n13717), 
            .D(tx_data[3]));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFE r_Tx_Data_i4 (.Q(r_Tx_Data[4]), .C(clk32MHz), .E(n13717), 
            .D(tx_data[4]));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFE r_Tx_Data_i5 (.Q(r_Tx_Data[5]), .C(clk32MHz), .E(n13717), 
            .D(tx_data[5]));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFE r_Tx_Data_i6 (.Q(r_Tx_Data[6]), .C(clk32MHz), .E(n13717), 
            .D(tx_data[6]));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFE r_Tx_Data_i7 (.Q(r_Tx_Data[7]), .C(clk32MHz), .E(n13717), 
            .D(tx_data[7]));   // verilog/uart_tx.v(40[10] 143[8])
    SB_LUT4 i1_3_lut (.I0(\r_SM_Main[2] ), .I1(n79), .I2(r_SM_Main[1]), 
            .I3(GND_net), .O(n32645));   // verilog/uart_tx.v(31[16:25])
    defparam i1_3_lut.LUT_INIT = 16'h1414;
    SB_LUT4 i2_3_lut_4_lut (.I0(r_SM_Main[1]), .I1(r_SM_Main[0]), .I2(\r_SM_Main_2__N_3458[0] ), 
            .I3(\r_SM_Main[2] ), .O(n13717));
    defparam i2_3_lut_4_lut.LUT_INIT = 16'h0010;
    SB_LUT4 i1_3_lut_4_lut (.I0(\r_SM_Main[2] ), .I1(r_SM_Main[1]), .I2(r_SM_Main[0]), 
            .I3(r_SM_Main_2__N_3455[1]), .O(n5478));   // verilog/uart_tx.v(31[16:25])
    defparam i1_3_lut_4_lut.LUT_INIT = 16'h5501;
    SB_LUT4 tx_o_bdd_4_lut_4_lut (.I0(tx_o), .I1(n2), .I2(\r_SM_Main[2] ), 
            .I3(r_SM_Main[1]), .O(n38429));
    defparam tx_o_bdd_4_lut_4_lut.LUT_INIT = 16'hacaa;
    SB_LUT4 o_Tx_Serial_I_0_1_lut (.I0(tx_o), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(tx_enable));   // verilog/uart_tx.v(38[24:36])
    defparam o_Tx_Serial_I_0_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 r_Bit_Index_0__bdd_4_lut_31660 (.I0(r_Bit_Index[0]), .I1(r_Tx_Data[6]), 
            .I2(r_Tx_Data[7]), .I3(r_Bit_Index[1]), .O(n38297));
    defparam r_Bit_Index_0__bdd_4_lut_31660.LUT_INIT = 16'he4aa;
    SB_LUT4 n38297_bdd_4_lut (.I0(n38297), .I1(r_Tx_Data[5]), .I2(r_Tx_Data[4]), 
            .I3(r_Bit_Index[1]), .O(n38300));
    defparam n38297_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF r_Clock_Count__i3 (.Q(\r_Clock_Count[3] ), .C(clk32MHz), .D(n17559));   // verilog/uart_tx.v(40[10] 143[8])
    SB_LUT4 i1_2_lut_3_lut (.I0(tx_active), .I1(\r_SM_Main_2__N_3458[0] ), 
            .I2(tx_transmit_N_3355), .I3(GND_net), .O(n1502));
    defparam i1_2_lut_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i20228_3_lut_4_lut (.I0(tx_active), .I1(\r_SM_Main_2__N_3458[0] ), 
            .I2(n63), .I3(n16157), .O(n25050));
    defparam i20228_3_lut_4_lut.LUT_INIT = 16'hf0e0;
    SB_LUT4 i2_2_lut_3_lut_4_lut (.I0(tx_active), .I1(\r_SM_Main_2__N_3458[0] ), 
            .I2(\byte_transmit_counter[4] ), .I3(\byte_transmit_counter[3] ), 
            .O(n7));
    defparam i2_2_lut_3_lut_4_lut.LUT_INIT = 16'hfeee;
    SB_LUT4 i1_2_lut_3_lut_adj_875 (.I0(r_SM_Main[0]), .I1(n24692), .I2(n19424), 
            .I3(GND_net), .O(n79));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i1_2_lut_3_lut_adj_875.LUT_INIT = 16'ha8a8;
    SB_LUT4 i1_2_lut (.I0(r_SM_Main[0]), .I1(\r_SM_Main_2__N_3458[0] ), 
            .I2(GND_net), .I3(GND_net), .O(n4));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i1_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i1_2_lut_adj_876 (.I0(n24692), .I1(n19424), .I2(GND_net), 
            .I3(GND_net), .O(r_SM_Main_2__N_3455[1]));   // verilog/uart_tx.v(31[16:25])
    defparam i1_2_lut_adj_876.LUT_INIT = 16'heeee;
    SB_DFF r_Clock_Count__i2 (.Q(r_Clock_Count[2]), .C(clk32MHz), .D(n17732));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFF r_Clock_Count__i1 (.Q(r_Clock_Count[1]), .C(clk32MHz), .D(n32445));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFF r_SM_Main_i0 (.Q(r_SM_Main[0]), .C(clk32MHz), .D(r_SM_Main_2__N_3426[0]));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFF r_Tx_Active_47 (.Q(tx_active), .C(clk32MHz), .D(n17703));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFF o_Tx_Serial_45 (.Q(tx_o), .C(clk32MHz), .D(n38432));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFF r_SM_Main_i2 (.Q(\r_SM_Main[2] ), .C(clk32MHz), .D(n34119));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFF r_Clock_Count__i0 (.Q(\r_Clock_Count[0] ), .C(clk32MHz), .D(n18278));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFF r_Bit_Index_i2 (.Q(r_Bit_Index[2]), .C(clk32MHz), .D(n17652));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFF r_Bit_Index_i1 (.Q(r_Bit_Index[1]), .C(clk32MHz), .D(n17655));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFF r_Clock_Count__i8 (.Q(\r_Clock_Count[8] ), .C(clk32MHz), .D(n17708));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFF r_Clock_Count__i7 (.Q(\r_Clock_Count[7] ), .C(clk32MHz), .D(n17713));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFF r_Bit_Index_i0 (.Q(r_Bit_Index[0]), .C(clk32MHz), .D(n17728));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFF r_Clock_Count__i6 (.Q(\r_Clock_Count[6] ), .C(clk32MHz), .D(n17549));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFF r_Clock_Count__i5 (.Q(\r_Clock_Count[5] ), .C(clk32MHz), .D(n17553));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFF r_Clock_Count__i4 (.Q(r_Clock_Count[4]), .C(clk32MHz), .D(n32443));   // verilog/uart_tx.v(40[10] 143[8])
    
endmodule
//
// Verilog Description of module uart_rx
//

module uart_rx (n25112, r_SM_Main, clk32MHz, VCC_net, rx_data_ready, 
            n18260, rx_data, r_Rx_Data, n37332, GND_net, PIN_13_N_105, 
            \r_SM_Main[2] , n33769, n17681, r_Bit_Index, n5578, n24193, 
            n4, n4_adj_1, n16148, n25070, n1, n37333, n17701, 
            n17689, n17688, n17687, n17686, n17685, n17684, n17683, 
            n16143, n17679, n17682, n17735, n4_adj_2) /* synthesis lattice_noprune=1, syn_preserve=0, syn_module_defined=1, syn_noprune=0 */ ;
    input n25112;
    output [2:0]r_SM_Main;
    input clk32MHz;
    input VCC_net;
    output rx_data_ready;
    input n18260;
    output [7:0]rx_data;
    output r_Rx_Data;
    output n37332;
    input GND_net;
    input PIN_13_N_105;
    output \r_SM_Main[2] ;
    output n33769;
    output n17681;
    output [2:0]r_Bit_Index;
    output n5578;
    output n24193;
    output n4;
    output n4_adj_1;
    output n16148;
    output n25070;
    output n1;
    output n37333;
    input n17701;
    input n17689;
    input n17688;
    input n17687;
    input n17686;
    input n17685;
    input n17684;
    input n17683;
    output n16143;
    input n17679;
    input n17682;
    input n17735;
    output n4_adj_2;
    
    wire clk32MHz /* synthesis SET_AS_NETWORK=clk32MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(34[6:14])
    
    wire n32355;
    wire [2:0]r_SM_Main_c;   // verilog/uart_rx.v(36[17:26])
    wire [2:0]r_SM_Main_2__N_3390;
    
    wire r_Rx_Data_R;
    wire [31:0]n194;
    
    wire n17340;
    wire [7:0]r_Clock_Count;   // verilog/uart_rx.v(32[17:30])
    
    wire n17511;
    wire [2:0]r_SM_Main_2__N_3384;
    
    wire n32933, n24495, n32858, n15964, n28031, n28030, n28029, 
        n28028, n28027, n28026, n6, n28025, n17268, n36424, n37296, 
        n6_adj_4337;
    
    SB_DFF r_SM_Main_i1 (.Q(r_SM_Main[1]), .C(clk32MHz), .D(n25112));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFFE r_Rx_DV_52 (.Q(rx_data_ready), .C(clk32MHz), .E(VCC_net), 
            .D(n32355));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_Byte_i0 (.Q(rx_data[0]), .C(clk32MHz), .D(n18260));   // verilog/uart_rx.v(49[10] 144[8])
    SB_LUT4 i30964_3_lut (.I0(r_SM_Main_c[0]), .I1(r_SM_Main_2__N_3390[0]), 
            .I2(r_Rx_Data), .I3(GND_net), .O(n37332));   // verilog/uart_rx.v(52[7] 143[14])
    defparam i30964_3_lut.LUT_INIT = 16'hfdfd;
    SB_DFF r_Rx_Data_50 (.Q(r_Rx_Data), .C(clk32MHz), .D(r_Rx_Data_R));   // verilog/uart_rx.v(41[10] 45[8])
    SB_DFFESR r_Clock_Count__i7 (.Q(r_Clock_Count[7]), .C(clk32MHz), .E(n17340), 
            .D(n194[7]), .R(n17511));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_Data_R_49 (.Q(r_Rx_Data_R), .C(clk32MHz), .D(PIN_13_N_105));   // verilog/uart_rx.v(41[10] 45[8])
    SB_DFFESR r_Clock_Count__i6 (.Q(r_Clock_Count[6]), .C(clk32MHz), .E(n17340), 
            .D(n194[6]), .R(n17511));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFFESR r_Clock_Count__i5 (.Q(r_Clock_Count[5]), .C(clk32MHz), .E(n17340), 
            .D(n194[5]), .R(n17511));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFFSR r_SM_Main_i2 (.Q(\r_SM_Main[2] ), .C(clk32MHz), .D(r_SM_Main_2__N_3384[2]), 
            .R(n32933));   // verilog/uart_rx.v(49[10] 144[8])
    SB_LUT4 i2_4_lut (.I0(\r_SM_Main[2] ), .I1(r_SM_Main_2__N_3384[2]), 
            .I2(r_SM_Main_c[0]), .I3(r_SM_Main[1]), .O(n33769));
    defparam i2_4_lut.LUT_INIT = 16'hfbfa;
    SB_LUT4 i27181_3_lut (.I0(n33769), .I1(n24495), .I2(r_SM_Main[1]), 
            .I3(GND_net), .O(n17681));
    defparam i27181_3_lut.LUT_INIT = 16'hbaba;
    SB_LUT4 i1792_2_lut (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[0]), .I2(GND_net), 
            .I3(GND_net), .O(n5578));   // verilog/uart_rx.v(102[36:51])
    defparam i1792_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i2_3_lut_4_lut (.I0(r_Clock_Count[6]), .I1(r_Clock_Count[7]), 
            .I2(n32858), .I3(r_Clock_Count[5]), .O(r_SM_Main_2__N_3384[2]));   // verilog/uart_rx.v(68[17:52])
    defparam i2_3_lut_4_lut.LUT_INIT = 16'hfeee;
    SB_LUT4 i2_3_lut_4_lut_adj_865 (.I0(r_Clock_Count[6]), .I1(r_Clock_Count[7]), 
            .I2(n32858), .I3(r_Clock_Count[5]), .O(r_SM_Main_2__N_3390[0]));   // verilog/uart_rx.v(68[17:52])
    defparam i2_3_lut_4_lut_adj_865.LUT_INIT = 16'hffef;
    SB_LUT4 i19383_2_lut (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[2]), .I2(GND_net), 
            .I3(GND_net), .O(n24193));
    defparam i19383_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 equal_148_i4_2_lut (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[2]), 
            .I2(GND_net), .I3(GND_net), .O(n4));   // verilog/uart_rx.v(97[17:39])
    defparam equal_148_i4_2_lut.LUT_INIT = 16'hbbbb;
    SB_LUT4 equal_150_i4_2_lut (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[2]), 
            .I2(GND_net), .I3(GND_net), .O(n4_adj_1));   // verilog/uart_rx.v(97[17:39])
    defparam equal_150_i4_2_lut.LUT_INIT = 16'hdddd;
    SB_LUT4 i1_2_lut (.I0(n15964), .I1(r_Bit_Index[0]), .I2(GND_net), 
            .I3(GND_net), .O(n16148));   // verilog/uart_rx.v(52[7] 143[14])
    defparam i1_2_lut.LUT_INIT = 16'hbbbb;
    SB_LUT4 i2_3_lut (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[2]), .I2(r_Bit_Index[0]), 
            .I3(GND_net), .O(n24495));
    defparam i2_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 r_SM_Main_2__I_0_56_Mux_0_i2_3_lut (.I0(n24495), .I1(r_SM_Main_2__N_3384[2]), 
            .I2(r_SM_Main_c[0]), .I3(GND_net), .O(n25070));   // verilog/uart_rx.v(52[7] 143[14])
    defparam r_SM_Main_2__I_0_56_Mux_0_i2_3_lut.LUT_INIT = 16'hc7c7;
    SB_LUT4 r_SM_Main_2__I_0_56_Mux_0_i1_3_lut (.I0(r_Rx_Data), .I1(r_SM_Main_2__N_3390[0]), 
            .I2(r_SM_Main_c[0]), .I3(GND_net), .O(n1));   // verilog/uart_rx.v(52[7] 143[14])
    defparam r_SM_Main_2__I_0_56_Mux_0_i1_3_lut.LUT_INIT = 16'hc5c5;
    SB_DFFESR r_Clock_Count__i0 (.Q(r_Clock_Count[0]), .C(clk32MHz), .E(n17340), 
            .D(n194[0]), .R(n17511));   // verilog/uart_rx.v(49[10] 144[8])
    SB_LUT4 add_62_9_lut (.I0(GND_net), .I1(r_Clock_Count[7]), .I2(GND_net), 
            .I3(n28031), .O(n194[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_62_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_62_8_lut (.I0(GND_net), .I1(r_Clock_Count[6]), .I2(GND_net), 
            .I3(n28030), .O(n194[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_62_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_62_8 (.CI(n28030), .I0(r_Clock_Count[6]), .I1(GND_net), 
            .CO(n28031));
    SB_LUT4 i30842_2_lut (.I0(r_SM_Main_2__N_3384[2]), .I1(r_SM_Main_c[0]), 
            .I2(GND_net), .I3(GND_net), .O(n37333));   // verilog/uart_rx.v(52[7] 143[14])
    defparam i30842_2_lut.LUT_INIT = 16'h8888;
    SB_DFFESR r_Clock_Count__i4 (.Q(r_Clock_Count[4]), .C(clk32MHz), .E(n17340), 
            .D(n194[4]), .R(n17511));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFFESR r_Clock_Count__i3 (.Q(r_Clock_Count[3]), .C(clk32MHz), .E(n17340), 
            .D(n194[3]), .R(n17511));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFFESR r_Clock_Count__i2 (.Q(r_Clock_Count[2]), .C(clk32MHz), .E(n17340), 
            .D(n194[2]), .R(n17511));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFFESR r_Clock_Count__i1 (.Q(r_Clock_Count[1]), .C(clk32MHz), .E(n17340), 
            .D(n194[1]), .R(n17511));   // verilog/uart_rx.v(49[10] 144[8])
    SB_LUT4 add_62_7_lut (.I0(GND_net), .I1(r_Clock_Count[5]), .I2(GND_net), 
            .I3(n28029), .O(n194[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_62_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_62_7 (.CI(n28029), .I0(r_Clock_Count[5]), .I1(GND_net), 
            .CO(n28030));
    SB_LUT4 add_62_6_lut (.I0(GND_net), .I1(r_Clock_Count[4]), .I2(GND_net), 
            .I3(n28028), .O(n194[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_62_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_62_6 (.CI(n28028), .I0(r_Clock_Count[4]), .I1(GND_net), 
            .CO(n28029));
    SB_LUT4 add_62_5_lut (.I0(GND_net), .I1(r_Clock_Count[3]), .I2(GND_net), 
            .I3(n28027), .O(n194[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_62_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_62_5 (.CI(n28027), .I0(r_Clock_Count[3]), .I1(GND_net), 
            .CO(n28028));
    SB_LUT4 add_62_4_lut (.I0(GND_net), .I1(r_Clock_Count[2]), .I2(GND_net), 
            .I3(n28026), .O(n194[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_62_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i4_4_lut (.I0(r_Clock_Count[1]), .I1(r_Clock_Count[3]), .I2(r_Clock_Count[4]), 
            .I3(n6), .O(n32858));
    defparam i4_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i1_2_lut_adj_866 (.I0(r_Clock_Count[0]), .I1(r_Clock_Count[2]), 
            .I2(GND_net), .I3(GND_net), .O(n6));
    defparam i1_2_lut_adj_866.LUT_INIT = 16'h8888;
    SB_CARRY add_62_4 (.CI(n28026), .I0(r_Clock_Count[2]), .I1(GND_net), 
            .CO(n28027));
    SB_LUT4 add_62_3_lut (.I0(GND_net), .I1(r_Clock_Count[1]), .I2(GND_net), 
            .I3(n28025), .O(n194[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_62_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_62_3 (.CI(n28025), .I0(r_Clock_Count[1]), .I1(GND_net), 
            .CO(n28026));
    SB_LUT4 add_62_2_lut (.I0(GND_net), .I1(r_Clock_Count[0]), .I2(GND_net), 
            .I3(VCC_net), .O(n194[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_62_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_62_2 (.CI(VCC_net), .I0(r_Clock_Count[0]), .I1(GND_net), 
            .CO(n28025));
    SB_LUT4 i2_4_lut_adj_867 (.I0(r_SM_Main[1]), .I1(r_SM_Main_2__N_3384[2]), 
            .I2(\r_SM_Main[2] ), .I3(r_SM_Main_c[0]), .O(n15964));
    defparam i2_4_lut_adj_867.LUT_INIT = 16'hfff7;
    SB_LUT4 i31538_2_lut_3_lut (.I0(r_SM_Main[1]), .I1(\r_SM_Main[2] ), 
            .I2(r_SM_Main_c[0]), .I3(GND_net), .O(n32933));
    defparam i31538_2_lut_3_lut.LUT_INIT = 16'hdfdf;
    SB_LUT4 i13_4_lut_4_lut (.I0(r_SM_Main[1]), .I1(\r_SM_Main[2] ), .I2(r_SM_Main_2__N_3384[2]), 
            .I3(r_SM_Main_c[0]), .O(n17268));
    defparam i13_4_lut_4_lut.LUT_INIT = 16'h2055;
    SB_LUT4 i12_3_lut_4_lut (.I0(r_SM_Main[1]), .I1(\r_SM_Main[2] ), .I2(n17268), 
            .I3(rx_data_ready), .O(n32355));
    defparam i12_3_lut_4_lut.LUT_INIT = 16'h2f20;
    SB_LUT4 i29821_4_lut (.I0(r_Clock_Count[5]), .I1(r_Rx_Data), .I2(r_Clock_Count[7]), 
            .I3(r_SM_Main_2__N_3390[0]), .O(n36424));
    defparam i29821_4_lut.LUT_INIT = 16'hfafe;
    SB_LUT4 i30810_4_lut (.I0(r_Clock_Count[6]), .I1(r_SM_Main_c[0]), .I2(n36424), 
            .I3(n32858), .O(n37296));
    defparam i30810_4_lut.LUT_INIT = 16'h3733;
    SB_LUT4 i1_4_lut (.I0(\r_SM_Main[2] ), .I1(n37296), .I2(r_SM_Main_2__N_3384[2]), 
            .I3(r_SM_Main[1]), .O(n17511));
    defparam i1_4_lut.LUT_INIT = 16'h5044;
    SB_LUT4 i2_2_lut (.I0(r_SM_Main_2__N_3390[0]), .I1(r_SM_Main_c[0]), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_4337));
    defparam i2_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i31481_4_lut (.I0(\r_SM_Main[2] ), .I1(r_SM_Main[1]), .I2(n6_adj_4337), 
            .I3(r_Rx_Data), .O(n17340));   // verilog/uart_rx.v(52[7] 143[14])
    defparam i31481_4_lut.LUT_INIT = 16'h4555;
    SB_DFF r_SM_Main_i0 (.Q(r_SM_Main_c[0]), .C(clk32MHz), .D(n17701));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_Byte_i1 (.Q(rx_data[1]), .C(clk32MHz), .D(n17689));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_Byte_i2 (.Q(rx_data[2]), .C(clk32MHz), .D(n17688));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_Byte_i3 (.Q(rx_data[3]), .C(clk32MHz), .D(n17687));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_Byte_i4 (.Q(rx_data[4]), .C(clk32MHz), .D(n17686));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_Byte_i5 (.Q(rx_data[5]), .C(clk32MHz), .D(n17685));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_Byte_i6 (.Q(rx_data[6]), .C(clk32MHz), .D(n17684));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_Byte_i7 (.Q(rx_data[7]), .C(clk32MHz), .D(n17683));   // verilog/uart_rx.v(49[10] 144[8])
    SB_LUT4 i1_2_lut_adj_868 (.I0(r_Bit_Index[0]), .I1(n15964), .I2(GND_net), 
            .I3(GND_net), .O(n16143));   // verilog/uart_rx.v(52[7] 143[14])
    defparam i1_2_lut_adj_868.LUT_INIT = 16'heeee;
    SB_DFF r_Bit_Index_i2 (.Q(r_Bit_Index[2]), .C(clk32MHz), .D(n17679));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Bit_Index_i1 (.Q(r_Bit_Index[1]), .C(clk32MHz), .D(n17682));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Bit_Index_i0 (.Q(r_Bit_Index[0]), .C(clk32MHz), .D(n17735));   // verilog/uart_rx.v(49[10] 144[8])
    SB_LUT4 equal_152_i4_2_lut (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[2]), 
            .I2(GND_net), .I3(GND_net), .O(n4_adj_2));   // verilog/uart_rx.v(97[17:39])
    defparam equal_152_i4_2_lut.LUT_INIT = 16'heeee;
    
endmodule
//
// Verilog Description of module \quad(DEBOUNCE_TICKS=100) 
//

module \quad(DEBOUNCE_TICKS=100)  (n18254, encoder1_position, clk32MHz, 
            n18255, n18256, n18252, n18253, n18250, n18251, n18248, 
            n18249, n18246, n18247, n18244, n18245, n18241, n18242, 
            n18243, n18239, n18240, n18235, n18236, n18237, n18238, 
            n18234, data_o, GND_net, n3158, count_enable, n17699, 
            PIN_9_c_1, n18264, reg_B, n34971, PIN_10_c_0, n17705) /* synthesis lattice_noprune=1, syn_preserve=0, syn_module_defined=1, syn_noprune=0 */ ;
    input n18254;
    output [23:0]encoder1_position;
    input clk32MHz;
    input n18255;
    input n18256;
    input n18252;
    input n18253;
    input n18250;
    input n18251;
    input n18248;
    input n18249;
    input n18246;
    input n18247;
    input n18244;
    input n18245;
    input n18241;
    input n18242;
    input n18243;
    input n18239;
    input n18240;
    input n18235;
    input n18236;
    input n18237;
    input n18238;
    input n18234;
    output [1:0]data_o;
    input GND_net;
    output [23:0]n3158;
    output count_enable;
    input n17699;
    input PIN_9_c_1;
    input n18264;
    output [1:0]reg_B;
    output n34971;
    input PIN_10_c_0;
    input n17705;
    
    wire clk32MHz /* synthesis SET_AS_NETWORK=clk32MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(34[6:14])
    
    wire B_delayed, A_delayed, count_direction, n3142, n28155, n28154, 
        n28153, n28152, n28151, n28150, n28149, n28148, n28147, 
        n28146, n28145, n28144, n28143, n28142, n28141, n28140, 
        n28139, n28138, n28137, n28136, n28135, n28134, n28133, 
        n28132;
    
    SB_DFF count_i0_i21 (.Q(encoder1_position[21]), .C(clk32MHz), .D(n18254));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i22 (.Q(encoder1_position[22]), .C(clk32MHz), .D(n18255));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i23 (.Q(encoder1_position[23]), .C(clk32MHz), .D(n18256));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i19 (.Q(encoder1_position[19]), .C(clk32MHz), .D(n18252));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i20 (.Q(encoder1_position[20]), .C(clk32MHz), .D(n18253));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i17 (.Q(encoder1_position[17]), .C(clk32MHz), .D(n18250));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i18 (.Q(encoder1_position[18]), .C(clk32MHz), .D(n18251));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i15 (.Q(encoder1_position[15]), .C(clk32MHz), .D(n18248));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i16 (.Q(encoder1_position[16]), .C(clk32MHz), .D(n18249));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i13 (.Q(encoder1_position[13]), .C(clk32MHz), .D(n18246));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i14 (.Q(encoder1_position[14]), .C(clk32MHz), .D(n18247));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i11 (.Q(encoder1_position[11]), .C(clk32MHz), .D(n18244));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i12 (.Q(encoder1_position[12]), .C(clk32MHz), .D(n18245));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i8 (.Q(encoder1_position[8]), .C(clk32MHz), .D(n18241));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i9 (.Q(encoder1_position[9]), .C(clk32MHz), .D(n18242));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i10 (.Q(encoder1_position[10]), .C(clk32MHz), .D(n18243));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i6 (.Q(encoder1_position[6]), .C(clk32MHz), .D(n18239));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i7 (.Q(encoder1_position[7]), .C(clk32MHz), .D(n18240));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i2 (.Q(encoder1_position[2]), .C(clk32MHz), .D(n18235));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i3 (.Q(encoder1_position[3]), .C(clk32MHz), .D(n18236));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i4 (.Q(encoder1_position[4]), .C(clk32MHz), .D(n18237));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i5 (.Q(encoder1_position[5]), .C(clk32MHz), .D(n18238));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i1 (.Q(encoder1_position[1]), .C(clk32MHz), .D(n18234));   // quad.v(35[10] 41[6])
    SB_DFF B_delayed_16 (.Q(B_delayed), .C(clk32MHz), .D(data_o[0]));   // quad.v(23[10:54])
    SB_DFF A_delayed_15 (.Q(A_delayed), .C(clk32MHz), .D(data_o[1]));   // quad.v(22[10:54])
    SB_LUT4 quadA_debounced_I_0_2_lut (.I0(data_o[1]), .I1(B_delayed), .I2(GND_net), 
            .I3(GND_net), .O(count_direction));   // quad.v(26[26:53])
    defparam quadA_debounced_I_0_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_633_25_lut (.I0(GND_net), .I1(encoder1_position[23]), .I2(n3142), 
            .I3(n28155), .O(n3158[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_633_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_633_24_lut (.I0(GND_net), .I1(encoder1_position[22]), .I2(n3142), 
            .I3(n28154), .O(n3158[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_633_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_633_24 (.CI(n28154), .I0(encoder1_position[22]), .I1(n3142), 
            .CO(n28155));
    SB_LUT4 add_633_23_lut (.I0(GND_net), .I1(encoder1_position[21]), .I2(n3142), 
            .I3(n28153), .O(n3158[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_633_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_633_23 (.CI(n28153), .I0(encoder1_position[21]), .I1(n3142), 
            .CO(n28154));
    SB_LUT4 add_633_22_lut (.I0(GND_net), .I1(encoder1_position[20]), .I2(n3142), 
            .I3(n28152), .O(n3158[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_633_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_633_22 (.CI(n28152), .I0(encoder1_position[20]), .I1(n3142), 
            .CO(n28153));
    SB_LUT4 add_633_21_lut (.I0(GND_net), .I1(encoder1_position[19]), .I2(n3142), 
            .I3(n28151), .O(n3158[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_633_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_633_21 (.CI(n28151), .I0(encoder1_position[19]), .I1(n3142), 
            .CO(n28152));
    SB_LUT4 add_633_20_lut (.I0(GND_net), .I1(encoder1_position[18]), .I2(n3142), 
            .I3(n28150), .O(n3158[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_633_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_633_20 (.CI(n28150), .I0(encoder1_position[18]), .I1(n3142), 
            .CO(n28151));
    SB_LUT4 i3_4_lut (.I0(data_o[1]), .I1(A_delayed), .I2(B_delayed), 
            .I3(data_o[0]), .O(count_enable));   // quad.v(25[23:80])
    defparam i3_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 add_633_19_lut (.I0(GND_net), .I1(encoder1_position[17]), .I2(n3142), 
            .I3(n28149), .O(n3158[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_633_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_633_19 (.CI(n28149), .I0(encoder1_position[17]), .I1(n3142), 
            .CO(n28150));
    SB_LUT4 add_633_18_lut (.I0(GND_net), .I1(encoder1_position[16]), .I2(n3142), 
            .I3(n28148), .O(n3158[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_633_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_633_18 (.CI(n28148), .I0(encoder1_position[16]), .I1(n3142), 
            .CO(n28149));
    SB_LUT4 add_633_17_lut (.I0(GND_net), .I1(encoder1_position[15]), .I2(n3142), 
            .I3(n28147), .O(n3158[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_633_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_633_17 (.CI(n28147), .I0(encoder1_position[15]), .I1(n3142), 
            .CO(n28148));
    SB_LUT4 add_633_16_lut (.I0(GND_net), .I1(encoder1_position[14]), .I2(n3142), 
            .I3(n28146), .O(n3158[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_633_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_633_16 (.CI(n28146), .I0(encoder1_position[14]), .I1(n3142), 
            .CO(n28147));
    SB_LUT4 add_633_15_lut (.I0(GND_net), .I1(encoder1_position[13]), .I2(n3142), 
            .I3(n28145), .O(n3158[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_633_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_633_15 (.CI(n28145), .I0(encoder1_position[13]), .I1(n3142), 
            .CO(n28146));
    SB_LUT4 add_633_14_lut (.I0(GND_net), .I1(encoder1_position[12]), .I2(n3142), 
            .I3(n28144), .O(n3158[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_633_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_633_14 (.CI(n28144), .I0(encoder1_position[12]), .I1(n3142), 
            .CO(n28145));
    SB_LUT4 add_633_13_lut (.I0(GND_net), .I1(encoder1_position[11]), .I2(n3142), 
            .I3(n28143), .O(n3158[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_633_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_633_13 (.CI(n28143), .I0(encoder1_position[11]), .I1(n3142), 
            .CO(n28144));
    SB_LUT4 add_633_12_lut (.I0(GND_net), .I1(encoder1_position[10]), .I2(n3142), 
            .I3(n28142), .O(n3158[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_633_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_633_12 (.CI(n28142), .I0(encoder1_position[10]), .I1(n3142), 
            .CO(n28143));
    SB_LUT4 add_633_11_lut (.I0(GND_net), .I1(encoder1_position[9]), .I2(n3142), 
            .I3(n28141), .O(n3158[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_633_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_633_11 (.CI(n28141), .I0(encoder1_position[9]), .I1(n3142), 
            .CO(n28142));
    SB_LUT4 add_633_10_lut (.I0(GND_net), .I1(encoder1_position[8]), .I2(n3142), 
            .I3(n28140), .O(n3158[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_633_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_633_10 (.CI(n28140), .I0(encoder1_position[8]), .I1(n3142), 
            .CO(n28141));
    SB_LUT4 add_633_9_lut (.I0(GND_net), .I1(encoder1_position[7]), .I2(n3142), 
            .I3(n28139), .O(n3158[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_633_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_633_9 (.CI(n28139), .I0(encoder1_position[7]), .I1(n3142), 
            .CO(n28140));
    SB_LUT4 add_633_8_lut (.I0(GND_net), .I1(encoder1_position[6]), .I2(n3142), 
            .I3(n28138), .O(n3158[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_633_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_633_8 (.CI(n28138), .I0(encoder1_position[6]), .I1(n3142), 
            .CO(n28139));
    SB_LUT4 add_633_7_lut (.I0(GND_net), .I1(encoder1_position[5]), .I2(n3142), 
            .I3(n28137), .O(n3158[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_633_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_633_7 (.CI(n28137), .I0(encoder1_position[5]), .I1(n3142), 
            .CO(n28138));
    SB_LUT4 add_633_6_lut (.I0(GND_net), .I1(encoder1_position[4]), .I2(n3142), 
            .I3(n28136), .O(n3158[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_633_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_633_6 (.CI(n28136), .I0(encoder1_position[4]), .I1(n3142), 
            .CO(n28137));
    SB_LUT4 add_633_5_lut (.I0(GND_net), .I1(encoder1_position[3]), .I2(n3142), 
            .I3(n28135), .O(n3158[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_633_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_633_5 (.CI(n28135), .I0(encoder1_position[3]), .I1(n3142), 
            .CO(n28136));
    SB_LUT4 add_633_4_lut (.I0(GND_net), .I1(encoder1_position[2]), .I2(n3142), 
            .I3(n28134), .O(n3158[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_633_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_633_4 (.CI(n28134), .I0(encoder1_position[2]), .I1(n3142), 
            .CO(n28135));
    SB_LUT4 add_633_3_lut (.I0(GND_net), .I1(encoder1_position[1]), .I2(n3142), 
            .I3(n28133), .O(n3158[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_633_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_633_3 (.CI(n28133), .I0(encoder1_position[1]), .I1(n3142), 
            .CO(n28134));
    SB_LUT4 add_633_2_lut (.I0(GND_net), .I1(encoder1_position[0]), .I2(count_direction), 
            .I3(n28132), .O(n3158[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_633_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_633_2 (.CI(n28132), .I0(encoder1_position[0]), .I1(count_direction), 
            .CO(n28133));
    SB_CARRY add_633_1 (.CI(GND_net), .I0(n3142), .I1(n3142), .CO(n28132));
    SB_LUT4 i1109_1_lut_2_lut (.I0(data_o[1]), .I1(B_delayed), .I2(GND_net), 
            .I3(GND_net), .O(n3142));   // quad.v(37[5] 40[8])
    defparam i1109_1_lut_2_lut.LUT_INIT = 16'h9999;
    SB_DFF count_i0_i0 (.Q(encoder1_position[0]), .C(clk32MHz), .D(n17699));   // quad.v(35[10] 41[6])
    \grp_debouncer(2,5)  debounce (.PIN_9_c_1(PIN_9_c_1), .clk32MHz(clk32MHz), 
            .n18264(n18264), .data_o({data_o}), .reg_B({reg_B}), .n34971(n34971), 
            .GND_net(GND_net), .PIN_10_c_0(PIN_10_c_0), .n17705(n17705)) /* synthesis lattice_noprune=1, syn_preserve=0, syn_noprune=0 */ ;   // quad.v(15[24] 19[4])
    
endmodule
//
// Verilog Description of module \grp_debouncer(2,5) 
//

module \grp_debouncer(2,5)  (PIN_9_c_1, clk32MHz, n18264, data_o, reg_B, 
            n34971, GND_net, PIN_10_c_0, n17705) /* synthesis lattice_noprune=1, syn_preserve=0, syn_noprune=0 */ ;
    input PIN_9_c_1;
    input clk32MHz;
    input n18264;
    output [1:0]data_o;
    output [1:0]reg_B;
    output n34971;
    input GND_net;
    input PIN_10_c_0;
    input n17705;
    
    wire clk32MHz /* synthesis SET_AS_NETWORK=clk32MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(34[6:14])
    wire [1:0]reg_A;   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(142[12:17])
    wire [2:0]cnt_reg;   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(149[12:19])
    wire [2:0]n17;
    
    wire cnt_next_2__N_3694, n2;
    
    SB_DFF reg_A_i1 (.Q(reg_A[1]), .C(clk32MHz), .D(PIN_9_c_1));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(178[9] 184[16])
    SB_DFF reg_out_i0_i1 (.Q(data_o[1]), .C(clk32MHz), .D(n18264));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(186[9] 190[16])
    SB_DFF reg_B_i0 (.Q(reg_B[0]), .C(clk32MHz), .D(reg_A[0]));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(178[9] 184[16])
    SB_LUT4 i2_3_lut (.I0(cnt_reg[0]), .I1(cnt_reg[2]), .I2(cnt_reg[1]), 
            .I3(GND_net), .O(n34971));
    defparam i2_3_lut.LUT_INIT = 16'hf7f7;
    SB_DFFSR cnt_reg_1528__i0 (.Q(cnt_reg[0]), .C(clk32MHz), .D(n17[0]), 
            .R(cnt_next_2__N_3694));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[78:85])
    SB_LUT4 i22716_3_lut (.I0(cnt_reg[2]), .I1(cnt_reg[1]), .I2(cnt_reg[0]), 
            .I3(GND_net), .O(n17[2]));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[78:85])
    defparam i22716_3_lut.LUT_INIT = 16'h6a6a;
    SB_LUT4 i22709_2_lut (.I0(cnt_reg[1]), .I1(cnt_reg[0]), .I2(GND_net), 
            .I3(GND_net), .O(n17[1]));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[78:85])
    defparam i22709_2_lut.LUT_INIT = 16'h6666;
    SB_DFF reg_B_i1 (.Q(reg_B[1]), .C(clk32MHz), .D(reg_A[1]));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(178[9] 184[16])
    SB_DFF reg_A_i0 (.Q(reg_A[0]), .C(clk32MHz), .D(PIN_10_c_0));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(178[9] 184[16])
    SB_LUT4 reg_B_1__I_0_i2_2_lut (.I0(reg_B[1]), .I1(reg_A[1]), .I2(GND_net), 
            .I3(GND_net), .O(n2));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(193[46:60])
    defparam reg_B_1__I_0_i2_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i2_4_lut (.I0(reg_B[0]), .I1(n34971), .I2(reg_A[0]), .I3(n2), 
            .O(cnt_next_2__N_3694));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[40:72])
    defparam i2_4_lut.LUT_INIT = 16'hff7b;
    SB_LUT4 i22707_1_lut (.I0(cnt_reg[0]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n17[0]));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[78:85])
    defparam i22707_1_lut.LUT_INIT = 16'h5555;
    SB_DFFSR cnt_reg_1528__i1 (.Q(cnt_reg[1]), .C(clk32MHz), .D(n17[1]), 
            .R(cnt_next_2__N_3694));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[78:85])
    SB_DFFSR cnt_reg_1528__i2 (.Q(cnt_reg[2]), .C(clk32MHz), .D(n17[2]), 
            .R(cnt_next_2__N_3694));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[78:85])
    SB_DFF reg_out_i0_i0 (.Q(data_o[0]), .C(clk32MHz), .D(n17705));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(186[9] 190[16])
    
endmodule
//
// Verilog Description of module \quad(DEBOUNCE_TICKS=100)_U1 
//

module \quad(DEBOUNCE_TICKS=100)_U1  (n3208, encoder0_position, GND_net, 
            n18226, clk32MHz, n18227, n18228, n18229, n18230, n18231, 
            n18222, n18223, n18224, n18225, n18220, n18221, n18218, 
            n18219, n18216, n18217, n18214, n18215, n18212, n18213, 
            n18209, n18210, n18211, data_o, count_enable, n17697, 
            n18261, reg_B, n34970, PIN_2_c_0, PIN_1_c_1, n17700) /* synthesis lattice_noprune=1, syn_preserve=0, syn_module_defined=1, syn_noprune=0 */ ;
    output [23:0]n3208;
    output [23:0]encoder0_position;
    input GND_net;
    input n18226;
    input clk32MHz;
    input n18227;
    input n18228;
    input n18229;
    input n18230;
    input n18231;
    input n18222;
    input n18223;
    input n18224;
    input n18225;
    input n18220;
    input n18221;
    input n18218;
    input n18219;
    input n18216;
    input n18217;
    input n18214;
    input n18215;
    input n18212;
    input n18213;
    input n18209;
    input n18210;
    input n18211;
    output [1:0]data_o;
    output count_enable;
    input n17697;
    input n18261;
    output [1:0]reg_B;
    output n34970;
    input PIN_2_c_0;
    input PIN_1_c_1;
    input n17700;
    
    wire clk32MHz /* synthesis SET_AS_NETWORK=clk32MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(34[6:14])
    
    wire n3204, n28000, n28001, n27999, n27998, n27997, n27996, 
        B_delayed, A_delayed, n27995, count_direction, n27994, n28017, 
        n28016, n28015, n28014, n28013, n28012, n28011, n28010, 
        n28009, n28008, n28007, n28006, n28005, n28004, n28003, 
        n28002;
    
    SB_LUT4 add_659_8_lut (.I0(GND_net), .I1(encoder0_position[6]), .I2(n3204), 
            .I3(n28000), .O(n3208[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_659_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_659_8 (.CI(n28000), .I0(encoder0_position[6]), .I1(n3204), 
            .CO(n28001));
    SB_LUT4 add_659_7_lut (.I0(GND_net), .I1(encoder0_position[5]), .I2(n3204), 
            .I3(n27999), .O(n3208[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_659_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_659_7 (.CI(n27999), .I0(encoder0_position[5]), .I1(n3204), 
            .CO(n28000));
    SB_LUT4 add_659_6_lut (.I0(GND_net), .I1(encoder0_position[4]), .I2(n3204), 
            .I3(n27998), .O(n3208[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_659_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_659_6 (.CI(n27998), .I0(encoder0_position[4]), .I1(n3204), 
            .CO(n27999));
    SB_DFF count_i0_i18 (.Q(encoder0_position[18]), .C(clk32MHz), .D(n18226));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i19 (.Q(encoder0_position[19]), .C(clk32MHz), .D(n18227));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i20 (.Q(encoder0_position[20]), .C(clk32MHz), .D(n18228));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i21 (.Q(encoder0_position[21]), .C(clk32MHz), .D(n18229));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i22 (.Q(encoder0_position[22]), .C(clk32MHz), .D(n18230));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i23 (.Q(encoder0_position[23]), .C(clk32MHz), .D(n18231));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i14 (.Q(encoder0_position[14]), .C(clk32MHz), .D(n18222));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i15 (.Q(encoder0_position[15]), .C(clk32MHz), .D(n18223));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i16 (.Q(encoder0_position[16]), .C(clk32MHz), .D(n18224));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i17 (.Q(encoder0_position[17]), .C(clk32MHz), .D(n18225));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i12 (.Q(encoder0_position[12]), .C(clk32MHz), .D(n18220));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i13 (.Q(encoder0_position[13]), .C(clk32MHz), .D(n18221));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i10 (.Q(encoder0_position[10]), .C(clk32MHz), .D(n18218));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i11 (.Q(encoder0_position[11]), .C(clk32MHz), .D(n18219));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i8 (.Q(encoder0_position[8]), .C(clk32MHz), .D(n18216));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i9 (.Q(encoder0_position[9]), .C(clk32MHz), .D(n18217));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i6 (.Q(encoder0_position[6]), .C(clk32MHz), .D(n18214));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i7 (.Q(encoder0_position[7]), .C(clk32MHz), .D(n18215));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i4 (.Q(encoder0_position[4]), .C(clk32MHz), .D(n18212));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i5 (.Q(encoder0_position[5]), .C(clk32MHz), .D(n18213));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i1 (.Q(encoder0_position[1]), .C(clk32MHz), .D(n18209));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i2 (.Q(encoder0_position[2]), .C(clk32MHz), .D(n18210));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i3 (.Q(encoder0_position[3]), .C(clk32MHz), .D(n18211));   // quad.v(35[10] 41[6])
    SB_LUT4 add_659_5_lut (.I0(GND_net), .I1(encoder0_position[3]), .I2(n3204), 
            .I3(n27997), .O(n3208[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_659_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_659_5 (.CI(n27997), .I0(encoder0_position[3]), .I1(n3204), 
            .CO(n27998));
    SB_LUT4 add_659_4_lut (.I0(GND_net), .I1(encoder0_position[2]), .I2(n3204), 
            .I3(n27996), .O(n3208[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_659_4_lut.LUT_INIT = 16'hC33C;
    SB_DFF B_delayed_16 (.Q(B_delayed), .C(clk32MHz), .D(data_o[0]));   // quad.v(23[10:54])
    SB_DFF A_delayed_15 (.Q(A_delayed), .C(clk32MHz), .D(data_o[1]));   // quad.v(22[10:54])
    SB_CARRY add_659_4 (.CI(n27996), .I0(encoder0_position[2]), .I1(n3204), 
            .CO(n27997));
    SB_LUT4 add_659_3_lut (.I0(GND_net), .I1(encoder0_position[1]), .I2(n3204), 
            .I3(n27995), .O(n3208[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_659_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_659_3 (.CI(n27995), .I0(encoder0_position[1]), .I1(n3204), 
            .CO(n27996));
    SB_LUT4 add_659_2_lut (.I0(GND_net), .I1(encoder0_position[0]), .I2(count_direction), 
            .I3(n27994), .O(n3208[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_659_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_659_2 (.CI(n27994), .I0(encoder0_position[0]), .I1(count_direction), 
            .CO(n27995));
    SB_CARRY add_659_1 (.CI(GND_net), .I0(n3204), .I1(n3204), .CO(n27994));
    SB_LUT4 quadA_debounced_I_0_2_lut (.I0(data_o[1]), .I1(B_delayed), .I2(GND_net), 
            .I3(GND_net), .O(count_direction));   // quad.v(26[26:53])
    defparam quadA_debounced_I_0_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut (.I0(data_o[1]), .I1(A_delayed), .I2(B_delayed), 
            .I3(data_o[0]), .O(count_enable));   // quad.v(25[23:80])
    defparam i3_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i1104_1_lut_2_lut (.I0(data_o[1]), .I1(B_delayed), .I2(GND_net), 
            .I3(GND_net), .O(n3204));   // quad.v(37[5] 40[8])
    defparam i1104_1_lut_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 add_659_25_lut (.I0(GND_net), .I1(encoder0_position[23]), .I2(n3204), 
            .I3(n28017), .O(n3208[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_659_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_659_24_lut (.I0(GND_net), .I1(encoder0_position[22]), .I2(n3204), 
            .I3(n28016), .O(n3208[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_659_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_659_24 (.CI(n28016), .I0(encoder0_position[22]), .I1(n3204), 
            .CO(n28017));
    SB_LUT4 add_659_23_lut (.I0(GND_net), .I1(encoder0_position[21]), .I2(n3204), 
            .I3(n28015), .O(n3208[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_659_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_659_23 (.CI(n28015), .I0(encoder0_position[21]), .I1(n3204), 
            .CO(n28016));
    SB_LUT4 add_659_22_lut (.I0(GND_net), .I1(encoder0_position[20]), .I2(n3204), 
            .I3(n28014), .O(n3208[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_659_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_659_22 (.CI(n28014), .I0(encoder0_position[20]), .I1(n3204), 
            .CO(n28015));
    SB_LUT4 add_659_21_lut (.I0(GND_net), .I1(encoder0_position[19]), .I2(n3204), 
            .I3(n28013), .O(n3208[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_659_21_lut.LUT_INIT = 16'hC33C;
    SB_DFF count_i0_i0 (.Q(encoder0_position[0]), .C(clk32MHz), .D(n17697));   // quad.v(35[10] 41[6])
    SB_CARRY add_659_21 (.CI(n28013), .I0(encoder0_position[19]), .I1(n3204), 
            .CO(n28014));
    SB_LUT4 add_659_20_lut (.I0(GND_net), .I1(encoder0_position[18]), .I2(n3204), 
            .I3(n28012), .O(n3208[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_659_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_659_20 (.CI(n28012), .I0(encoder0_position[18]), .I1(n3204), 
            .CO(n28013));
    SB_LUT4 add_659_19_lut (.I0(GND_net), .I1(encoder0_position[17]), .I2(n3204), 
            .I3(n28011), .O(n3208[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_659_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_659_19 (.CI(n28011), .I0(encoder0_position[17]), .I1(n3204), 
            .CO(n28012));
    SB_LUT4 add_659_18_lut (.I0(GND_net), .I1(encoder0_position[16]), .I2(n3204), 
            .I3(n28010), .O(n3208[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_659_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_659_18 (.CI(n28010), .I0(encoder0_position[16]), .I1(n3204), 
            .CO(n28011));
    SB_LUT4 add_659_17_lut (.I0(GND_net), .I1(encoder0_position[15]), .I2(n3204), 
            .I3(n28009), .O(n3208[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_659_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_659_17 (.CI(n28009), .I0(encoder0_position[15]), .I1(n3204), 
            .CO(n28010));
    SB_LUT4 add_659_16_lut (.I0(GND_net), .I1(encoder0_position[14]), .I2(n3204), 
            .I3(n28008), .O(n3208[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_659_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_659_16 (.CI(n28008), .I0(encoder0_position[14]), .I1(n3204), 
            .CO(n28009));
    SB_LUT4 add_659_15_lut (.I0(GND_net), .I1(encoder0_position[13]), .I2(n3204), 
            .I3(n28007), .O(n3208[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_659_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_659_15 (.CI(n28007), .I0(encoder0_position[13]), .I1(n3204), 
            .CO(n28008));
    SB_LUT4 add_659_14_lut (.I0(GND_net), .I1(encoder0_position[12]), .I2(n3204), 
            .I3(n28006), .O(n3208[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_659_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_659_14 (.CI(n28006), .I0(encoder0_position[12]), .I1(n3204), 
            .CO(n28007));
    SB_LUT4 add_659_13_lut (.I0(GND_net), .I1(encoder0_position[11]), .I2(n3204), 
            .I3(n28005), .O(n3208[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_659_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_659_13 (.CI(n28005), .I0(encoder0_position[11]), .I1(n3204), 
            .CO(n28006));
    SB_LUT4 add_659_12_lut (.I0(GND_net), .I1(encoder0_position[10]), .I2(n3204), 
            .I3(n28004), .O(n3208[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_659_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_659_12 (.CI(n28004), .I0(encoder0_position[10]), .I1(n3204), 
            .CO(n28005));
    SB_LUT4 add_659_11_lut (.I0(GND_net), .I1(encoder0_position[9]), .I2(n3204), 
            .I3(n28003), .O(n3208[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_659_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_659_11 (.CI(n28003), .I0(encoder0_position[9]), .I1(n3204), 
            .CO(n28004));
    SB_LUT4 add_659_10_lut (.I0(GND_net), .I1(encoder0_position[8]), .I2(n3204), 
            .I3(n28002), .O(n3208[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_659_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_659_10 (.CI(n28002), .I0(encoder0_position[8]), .I1(n3204), 
            .CO(n28003));
    SB_LUT4 add_659_9_lut (.I0(GND_net), .I1(encoder0_position[7]), .I2(n3204), 
            .I3(n28001), .O(n3208[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_659_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_659_9 (.CI(n28001), .I0(encoder0_position[7]), .I1(n3204), 
            .CO(n28002));
    \grp_debouncer(2,5)_U0  debounce (.n18261(n18261), .data_o({data_o}), 
            .clk32MHz(clk32MHz), .reg_B({reg_B}), .n34970(n34970), .GND_net(GND_net), 
            .PIN_2_c_0(PIN_2_c_0), .PIN_1_c_1(PIN_1_c_1), .n17700(n17700)) /* synthesis lattice_noprune=1, syn_preserve=0, syn_noprune=0 */ ;   // quad.v(15[24] 19[4])
    
endmodule
//
// Verilog Description of module \grp_debouncer(2,5)_U0 
//

module \grp_debouncer(2,5)_U0  (n18261, data_o, clk32MHz, reg_B, n34970, 
            GND_net, PIN_2_c_0, PIN_1_c_1, n17700) /* synthesis lattice_noprune=1, syn_preserve=0, syn_noprune=0 */ ;
    input n18261;
    output [1:0]data_o;
    input clk32MHz;
    output [1:0]reg_B;
    output n34970;
    input GND_net;
    input PIN_2_c_0;
    input PIN_1_c_1;
    input n17700;
    
    wire clk32MHz /* synthesis SET_AS_NETWORK=clk32MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(34[6:14])
    wire [1:0]reg_A;   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(142[12:17])
    wire [2:0]cnt_reg;   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(149[12:19])
    wire [2:0]n17;
    
    wire cnt_next_2__N_3694, n2;
    
    SB_DFF reg_out_i0_i1 (.Q(data_o[1]), .C(clk32MHz), .D(n18261));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(186[9] 190[16])
    SB_DFF reg_B_i0 (.Q(reg_B[0]), .C(clk32MHz), .D(reg_A[0]));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(178[9] 184[16])
    SB_LUT4 i2_3_lut (.I0(cnt_reg[0]), .I1(cnt_reg[2]), .I2(cnt_reg[1]), 
            .I3(GND_net), .O(n34970));
    defparam i2_3_lut.LUT_INIT = 16'hf7f7;
    SB_DFFSR cnt_reg_1527__i0 (.Q(cnt_reg[0]), .C(clk32MHz), .D(n17[0]), 
            .R(cnt_next_2__N_3694));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[78:85])
    SB_LUT4 i22694_3_lut (.I0(cnt_reg[2]), .I1(cnt_reg[1]), .I2(cnt_reg[0]), 
            .I3(GND_net), .O(n17[2]));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[78:85])
    defparam i22694_3_lut.LUT_INIT = 16'h6a6a;
    SB_LUT4 i22687_2_lut (.I0(cnt_reg[1]), .I1(cnt_reg[0]), .I2(GND_net), 
            .I3(GND_net), .O(n17[1]));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[78:85])
    defparam i22687_2_lut.LUT_INIT = 16'h6666;
    SB_DFF reg_B_i1 (.Q(reg_B[1]), .C(clk32MHz), .D(reg_A[1]));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(178[9] 184[16])
    SB_DFF reg_A_i0 (.Q(reg_A[0]), .C(clk32MHz), .D(PIN_2_c_0));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(178[9] 184[16])
    SB_LUT4 reg_B_1__I_0_i2_2_lut (.I0(reg_B[1]), .I1(reg_A[1]), .I2(GND_net), 
            .I3(GND_net), .O(n2));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(193[46:60])
    defparam reg_B_1__I_0_i2_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i2_4_lut (.I0(reg_B[0]), .I1(n34970), .I2(reg_A[0]), .I3(n2), 
            .O(cnt_next_2__N_3694));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[40:72])
    defparam i2_4_lut.LUT_INIT = 16'hff7b;
    SB_LUT4 i22685_1_lut (.I0(cnt_reg[0]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n17[0]));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[78:85])
    defparam i22685_1_lut.LUT_INIT = 16'h5555;
    SB_DFF reg_A_i1 (.Q(reg_A[1]), .C(clk32MHz), .D(PIN_1_c_1));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(178[9] 184[16])
    SB_DFFSR cnt_reg_1527__i1 (.Q(cnt_reg[1]), .C(clk32MHz), .D(n17[1]), 
            .R(cnt_next_2__N_3694));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[78:85])
    SB_DFFSR cnt_reg_1527__i2 (.Q(cnt_reg[2]), .C(clk32MHz), .D(n17[2]), 
            .R(cnt_next_2__N_3694));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[78:85])
    SB_DFF reg_out_i0_i0 (.Q(data_o[0]), .C(clk32MHz), .D(n17700));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(186[9] 190[16])
    
endmodule
//
// Verilog Description of module \pwm(32000000,20000,32000000,23,1) 
//

module \pwm(32000000,20000,32000000,23,1)  (pwm_setpoint, GND_net, \half_duty_new[0] , 
            CLK_c, n1466, n18268, \half_duty[0][4] , n18270, \half_duty[0][6] , 
            n18271, \half_duty[0][7] , n18267, \half_duty[0][3] , n18265, 
            \half_duty[0][1] , n18266, \half_duty[0][2] , \half_duty[0][0] , 
            PIN_19_c_0, VCC_net, \half_duty_new[1] , \half_duty_new[2] , 
            \half_duty_new[3] , \half_duty_new[4] , \half_duty_new[6] , 
            \half_duty_new[7] , n17710) /* synthesis lattice_noprune=1, syn_preserve=0, syn_noprune=0 */ ;
    input [22:0]pwm_setpoint;
    input GND_net;
    output \half_duty_new[0] ;
    input CLK_c;
    output n1466;
    input n18268;
    output \half_duty[0][4] ;
    input n18270;
    output \half_duty[0][6] ;
    input n18271;
    output \half_duty[0][7] ;
    input n18267;
    output \half_duty[0][3] ;
    input n18265;
    output \half_duty[0][1] ;
    input n18266;
    output \half_duty[0][2] ;
    output \half_duty[0][0] ;
    output PIN_19_c_0;
    input VCC_net;
    output \half_duty_new[1] ;
    output \half_duty_new[2] ;
    output \half_duty_new[3] ;
    output \half_duty_new[4] ;
    output \half_duty_new[6] ;
    output \half_duty_new[7] ;
    input n17710;
    
    wire CLK_c /* synthesis SET_AS_NETWORK=CLK_c, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(3[9:12])
    
    wire n28266, n28267;
    wire [22:0]n6168;
    
    wire n28265;
    wire [9:0]half_duty_new_9__N_764;
    
    wire n28264;
    wire [10:0]n49;
    
    wire pause_counter_0__N_712;
    wire [10:0]\count[0] ;   // vhdl/pwm.vhd(51[11:16])
    
    wire n28263, n28262, n28261, n22073;
    wire [9:0]\half_duty[0] ;   // vhdl/pwm.vhd(55[11:20])
    
    wire n28260, n28259, n28258;
    wire [10:0]pwm_out_0__N_687;
    
    wire n28257, n28256, n28255, n28254, n28253, n28252, n28251, 
        n28250, n28249, pwm_out_0__N_682, n17287, n33687, pause_counter_0, 
        n28248, n12, n27907, pwm_out_0__N_686, n27906, n14, n18, 
        n19, n10, n27905, n38151, n27904, n8, n27903, n38147, 
        n27902, n4, n20, n5, n13, n38149, n22, n2, n3, n1, 
        n36420, n14_adj_4334, n18_adj_4335, n16, n17, n15;
    wire [9:0]half_duty_new;   // vhdl/pwm.vhd(53[12:25])
    
    wire n27901, n27900, n27899, n27898, n27897, n28475, n28474, 
        n28473, n28472, n28471, n28470, n28469, n28468, n28467, 
        n28466, n28290, n28289, n28288, n28287, n28286, n28285, 
        n28284, n28283, n28282, n28281, n28280, n28279, n28278, 
        n28277, n28276, n28275, n28274, n28273, n28272, n28271, 
        n28270, n28269, n28268;
    
    SB_CARRY add_2208_21 (.CI(n28266), .I0(pwm_setpoint[19]), .I1(GND_net), 
            .CO(n28267));
    SB_LUT4 add_2208_20_lut (.I0(GND_net), .I1(pwm_setpoint[18]), .I2(pwm_setpoint[22]), 
            .I3(n28265), .O(n6168[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2208_20_lut.LUT_INIT = 16'hC33C;
    SB_DFF half_duty_new_i1 (.Q(\half_duty_new[0] ), .C(CLK_c), .D(half_duty_new_9__N_764[0]));   // vhdl/pwm.vhd(59[5] 95[12])
    SB_CARRY add_2208_20 (.CI(n28265), .I0(pwm_setpoint[18]), .I1(pwm_setpoint[22]), 
            .CO(n28266));
    SB_LUT4 add_2208_19_lut (.I0(GND_net), .I1(pwm_setpoint[17]), .I2(pwm_setpoint[21]), 
            .I3(n28264), .O(n6168[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2208_19_lut.LUT_INIT = 16'hC33C;
    SB_DFFESR count_0__1525__i10 (.Q(\count[0] [10]), .C(CLK_c), .E(pause_counter_0__N_712), 
            .D(n49[10]), .R(n1466));   // vhdl/pwm.vhd(77[18:26])
    SB_CARRY add_2208_19 (.CI(n28264), .I0(pwm_setpoint[17]), .I1(pwm_setpoint[21]), 
            .CO(n28265));
    SB_LUT4 add_2208_18_lut (.I0(GND_net), .I1(pwm_setpoint[16]), .I2(pwm_setpoint[20]), 
            .I3(n28263), .O(n6168[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2208_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2208_18 (.CI(n28263), .I0(pwm_setpoint[16]), .I1(pwm_setpoint[20]), 
            .CO(n28264));
    SB_LUT4 add_2208_17_lut (.I0(GND_net), .I1(pwm_setpoint[15]), .I2(pwm_setpoint[19]), 
            .I3(n28262), .O(n6168[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2208_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2208_17 (.CI(n28262), .I0(pwm_setpoint[15]), .I1(pwm_setpoint[19]), 
            .CO(n28263));
    SB_LUT4 add_2208_16_lut (.I0(GND_net), .I1(pwm_setpoint[14]), .I2(pwm_setpoint[18]), 
            .I3(n28261), .O(n6168[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2208_16_lut.LUT_INIT = 16'hC33C;
    SB_DFFESR count_0__1525__i9 (.Q(\count[0] [9]), .C(CLK_c), .E(pause_counter_0__N_712), 
            .D(n49[9]), .R(n1466));   // vhdl/pwm.vhd(77[18:26])
    SB_DFFESR count_0__1525__i8 (.Q(\count[0] [8]), .C(CLK_c), .E(pause_counter_0__N_712), 
            .D(n49[8]), .R(n1466));   // vhdl/pwm.vhd(77[18:26])
    SB_DFF half_duty_0___i5 (.Q(\half_duty[0][4] ), .C(CLK_c), .D(n18268));   // vhdl/pwm.vhd(59[5] 95[12])
    SB_DFF half_duty_0___i6 (.Q(\half_duty[0] [5]), .C(CLK_c), .D(n22073));   // vhdl/pwm.vhd(59[5] 95[12])
    SB_DFF half_duty_0___i7 (.Q(\half_duty[0][6] ), .C(CLK_c), .D(n18270));   // vhdl/pwm.vhd(59[5] 95[12])
    SB_DFF half_duty_0___i8 (.Q(\half_duty[0][7] ), .C(CLK_c), .D(n18271));   // vhdl/pwm.vhd(59[5] 95[12])
    SB_DFFESR count_0__1525__i7 (.Q(\count[0] [7]), .C(CLK_c), .E(pause_counter_0__N_712), 
            .D(n49[7]), .R(n1466));   // vhdl/pwm.vhd(77[18:26])
    SB_DFF half_duty_0___i4 (.Q(\half_duty[0][3] ), .C(CLK_c), .D(n18267));   // vhdl/pwm.vhd(59[5] 95[12])
    SB_DFFESR count_0__1525__i6 (.Q(\count[0] [6]), .C(CLK_c), .E(pause_counter_0__N_712), 
            .D(n49[6]), .R(n1466));   // vhdl/pwm.vhd(77[18:26])
    SB_DFF half_duty_0___i2 (.Q(\half_duty[0][1] ), .C(CLK_c), .D(n18265));   // vhdl/pwm.vhd(59[5] 95[12])
    SB_DFF half_duty_0___i3 (.Q(\half_duty[0][2] ), .C(CLK_c), .D(n18266));   // vhdl/pwm.vhd(59[5] 95[12])
    SB_DFFESR count_0__1525__i5 (.Q(\count[0] [5]), .C(CLK_c), .E(pause_counter_0__N_712), 
            .D(n49[5]), .R(n1466));   // vhdl/pwm.vhd(77[18:26])
    SB_DFFESR count_0__1525__i4 (.Q(\count[0] [4]), .C(CLK_c), .E(pause_counter_0__N_712), 
            .D(n49[4]), .R(n1466));   // vhdl/pwm.vhd(77[18:26])
    SB_DFFESR count_0__1525__i3 (.Q(\count[0] [3]), .C(CLK_c), .E(pause_counter_0__N_712), 
            .D(n49[3]), .R(n1466));   // vhdl/pwm.vhd(77[18:26])
    SB_DFFESR count_0__1525__i2 (.Q(\count[0] [2]), .C(CLK_c), .E(pause_counter_0__N_712), 
            .D(n49[2]), .R(n1466));   // vhdl/pwm.vhd(77[18:26])
    SB_CARRY add_2208_16 (.CI(n28261), .I0(pwm_setpoint[14]), .I1(pwm_setpoint[18]), 
            .CO(n28262));
    SB_LUT4 add_2208_15_lut (.I0(GND_net), .I1(pwm_setpoint[13]), .I2(pwm_setpoint[17]), 
            .I3(n28260), .O(n6168[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2208_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2208_15 (.CI(n28260), .I0(pwm_setpoint[13]), .I1(pwm_setpoint[17]), 
            .CO(n28261));
    SB_LUT4 add_2208_14_lut (.I0(GND_net), .I1(pwm_setpoint[12]), .I2(pwm_setpoint[16]), 
            .I3(n28259), .O(n6168[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2208_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2208_14 (.CI(n28259), .I0(pwm_setpoint[12]), .I1(pwm_setpoint[16]), 
            .CO(n28260));
    SB_LUT4 add_2208_13_lut (.I0(GND_net), .I1(pwm_setpoint[11]), .I2(pwm_setpoint[15]), 
            .I3(n28258), .O(n6168[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2208_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 half_duty_0__9__I_0_i1_1_lut (.I0(\half_duty[0][0] ), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(pwm_out_0__N_687[0]));   // vhdl/pwm.vhd(84[22:28])
    defparam half_duty_0__9__I_0_i1_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 half_duty_0__9__I_0_i2_1_lut (.I0(\half_duty[0][1] ), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(pwm_out_0__N_687[1]));   // vhdl/pwm.vhd(84[22:28])
    defparam half_duty_0__9__I_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 half_duty_0__9__I_0_i3_1_lut (.I0(\half_duty[0][2] ), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(pwm_out_0__N_687[2]));   // vhdl/pwm.vhd(84[22:28])
    defparam half_duty_0__9__I_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_DFFESR count_0__1525__i1 (.Q(\count[0] [1]), .C(CLK_c), .E(pause_counter_0__N_712), 
            .D(n49[1]), .R(n1466));   // vhdl/pwm.vhd(77[18:26])
    SB_CARRY add_2208_13 (.CI(n28258), .I0(pwm_setpoint[11]), .I1(pwm_setpoint[15]), 
            .CO(n28259));
    SB_LUT4 add_2208_12_lut (.I0(GND_net), .I1(pwm_setpoint[10]), .I2(pwm_setpoint[14]), 
            .I3(n28257), .O(n6168[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2208_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2208_12 (.CI(n28257), .I0(pwm_setpoint[10]), .I1(pwm_setpoint[14]), 
            .CO(n28258));
    SB_LUT4 add_2208_11_lut (.I0(GND_net), .I1(pwm_setpoint[9]), .I2(pwm_setpoint[13]), 
            .I3(n28256), .O(n6168[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2208_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 half_duty_0__9__I_0_i4_1_lut (.I0(\half_duty[0][3] ), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(pwm_out_0__N_687[3]));   // vhdl/pwm.vhd(84[22:28])
    defparam half_duty_0__9__I_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 half_duty_0__9__I_0_i5_1_lut (.I0(\half_duty[0][4] ), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(pwm_out_0__N_687[4]));   // vhdl/pwm.vhd(84[22:28])
    defparam half_duty_0__9__I_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 half_duty_0__9__I_0_i6_1_lut (.I0(\half_duty[0] [5]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(pwm_out_0__N_687[5]));   // vhdl/pwm.vhd(84[22:28])
    defparam half_duty_0__9__I_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_2208_11 (.CI(n28256), .I0(pwm_setpoint[9]), .I1(pwm_setpoint[13]), 
            .CO(n28257));
    SB_LUT4 add_2208_10_lut (.I0(GND_net), .I1(pwm_setpoint[8]), .I2(pwm_setpoint[12]), 
            .I3(n28255), .O(n6168[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2208_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2208_10 (.CI(n28255), .I0(pwm_setpoint[8]), .I1(pwm_setpoint[12]), 
            .CO(n28256));
    SB_LUT4 add_2208_9_lut (.I0(GND_net), .I1(pwm_setpoint[7]), .I2(pwm_setpoint[11]), 
            .I3(n28254), .O(n6168[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2208_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2208_9 (.CI(n28254), .I0(pwm_setpoint[7]), .I1(pwm_setpoint[11]), 
            .CO(n28255));
    SB_LUT4 add_2208_8_lut (.I0(GND_net), .I1(pwm_setpoint[6]), .I2(pwm_setpoint[10]), 
            .I3(n28253), .O(n6168[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2208_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2208_8 (.CI(n28253), .I0(pwm_setpoint[6]), .I1(pwm_setpoint[10]), 
            .CO(n28254));
    SB_LUT4 add_2208_7_lut (.I0(GND_net), .I1(pwm_setpoint[5]), .I2(pwm_setpoint[9]), 
            .I3(n28252), .O(n6168[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2208_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2208_7 (.CI(n28252), .I0(pwm_setpoint[5]), .I1(pwm_setpoint[9]), 
            .CO(n28253));
    SB_LUT4 add_2208_6_lut (.I0(GND_net), .I1(pwm_setpoint[4]), .I2(pwm_setpoint[8]), 
            .I3(n28251), .O(n6168[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2208_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2208_6 (.CI(n28251), .I0(pwm_setpoint[4]), .I1(pwm_setpoint[8]), 
            .CO(n28252));
    SB_LUT4 add_2208_5_lut (.I0(GND_net), .I1(pwm_setpoint[3]), .I2(pwm_setpoint[7]), 
            .I3(n28250), .O(n6168[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2208_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2208_5 (.CI(n28250), .I0(pwm_setpoint[3]), .I1(pwm_setpoint[7]), 
            .CO(n28251));
    SB_LUT4 add_2208_4_lut (.I0(GND_net), .I1(pwm_setpoint[2]), .I2(pwm_setpoint[6]), 
            .I3(n28249), .O(n6168[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2208_4_lut.LUT_INIT = 16'hC33C;
    SB_DFFE pwm_out_0__39 (.Q(PIN_19_c_0), .C(CLK_c), .E(n17287), .D(pwm_out_0__N_682));   // vhdl/pwm.vhd(59[5] 95[12])
    SB_DFF pause_counter_0__38 (.Q(pause_counter_0), .C(CLK_c), .D(n33687));   // vhdl/pwm.vhd(59[5] 95[12])
    SB_CARRY add_2208_4 (.CI(n28249), .I0(pwm_setpoint[2]), .I1(pwm_setpoint[6]), 
            .CO(n28250));
    SB_LUT4 add_2208_3_lut (.I0(GND_net), .I1(pwm_setpoint[1]), .I2(pwm_setpoint[5]), 
            .I3(n28248), .O(n6168[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2208_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_2_lut (.I0(\count[0] [4]), .I1(\count[0] [5]), .I2(GND_net), 
            .I3(GND_net), .O(n12));
    defparam i1_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_2208_3 (.CI(n28248), .I0(pwm_setpoint[1]), .I1(pwm_setpoint[5]), 
            .CO(n28249));
    SB_LUT4 add_2208_2_lut (.I0(GND_net), .I1(pwm_setpoint[0]), .I2(pwm_setpoint[4]), 
            .I3(GND_net), .O(n6168[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2208_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2208_2 (.CI(GND_net), .I0(pwm_setpoint[0]), .I1(pwm_setpoint[4]), 
            .CO(n28248));
    SB_CARRY pwm_out_0__I_21_13 (.CI(n27907), .I0(GND_net), .I1(VCC_net), 
            .CO(pwm_out_0__N_686));
    SB_CARRY pwm_out_0__I_21_12 (.CI(n27906), .I0(VCC_net), .I1(VCC_net), 
            .CO(n27907));
    SB_LUT4 i7_4_lut (.I0(\count[0] [8]), .I1(n14), .I2(\count[0] [10]), 
            .I3(\count[0] [6]), .O(n18));
    defparam i7_4_lut.LUT_INIT = 16'h0040;
    SB_LUT4 i8_4_lut (.I0(\count[0] [9]), .I1(\count[0] [0]), .I2(\count[0] [1]), 
            .I3(\count[0] [2]), .O(n19));
    defparam i8_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i10_4_lut (.I0(n19), .I1(\count[0] [7]), .I2(n18), .I3(n12), 
            .O(n1466));
    defparam i10_4_lut.LUT_INIT = 16'h2000;
    SB_LUT4 pause_counter_0__I_0_48_1_lut (.I0(pause_counter_0), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(pause_counter_0__N_712));   // vhdl/pwm.vhd(72[7:27])
    defparam pause_counter_0__I_0_48_1_lut.LUT_INIT = 16'h5555;
    SB_DFFESR count_0__1525__i0 (.Q(\count[0] [0]), .C(CLK_c), .E(pause_counter_0__N_712), 
            .D(n49[0]), .R(n1466));   // vhdl/pwm.vhd(77[18:26])
    SB_LUT4 pwm_out_0__I_21_11_lut (.I0(\count[0] [9]), .I1(VCC_net), .I2(VCC_net), 
            .I3(n27905), .O(n10)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_out_0__I_21_11_lut.LUT_INIT = 16'h6996;
    SB_CARRY pwm_out_0__I_21_11 (.CI(n27905), .I0(VCC_net), .I1(VCC_net), 
            .CO(n27906));
    SB_LUT4 i17260_1_lut (.I0(\half_duty[0][6] ), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(pwm_out_0__N_687[6]));   // vhdl/pwm.vhd(59[5] 95[12])
    defparam i17260_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 pwm_out_0__I_21_10_lut (.I0(\count[0] [8]), .I1(GND_net), .I2(VCC_net), 
            .I3(n27904), .O(n38151)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_out_0__I_21_10_lut.LUT_INIT = 16'h6996;
    SB_CARRY pwm_out_0__I_21_10 (.CI(n27904), .I0(GND_net), .I1(VCC_net), 
            .CO(n27905));
    SB_LUT4 pwm_out_0__I_21_9_lut (.I0(\count[0] [7]), .I1(GND_net), .I2(pwm_out_0__N_687[7]), 
            .I3(n27903), .O(n8)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_out_0__I_21_9_lut.LUT_INIT = 16'h6996;
    SB_CARRY pwm_out_0__I_21_9 (.CI(n27903), .I0(GND_net), .I1(pwm_out_0__N_687[7]), 
            .CO(n27904));
    SB_LUT4 pwm_out_0__I_21_8_lut (.I0(\count[0] [6]), .I1(VCC_net), .I2(pwm_out_0__N_687[6]), 
            .I3(n27902), .O(n38147)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_out_0__I_21_8_lut.LUT_INIT = 16'h6996;
    SB_CARRY pwm_out_0__I_21_8 (.CI(n27902), .I0(VCC_net), .I1(pwm_out_0__N_687[6]), 
            .CO(n27903));
    SB_DFF half_duty_new_i2 (.Q(\half_duty_new[1] ), .C(CLK_c), .D(half_duty_new_9__N_764[1]));   // vhdl/pwm.vhd(59[5] 95[12])
    SB_LUT4 i31525_2_lut (.I0(pause_counter_0), .I1(pwm_out_0__N_682), .I2(GND_net), 
            .I3(GND_net), .O(n33687));
    defparam i31525_2_lut.LUT_INIT = 16'h1111;
    SB_LUT4 i8_4_lut_adj_860 (.I0(n4), .I1(n38151), .I2(n38147), .I3(pwm_out_0__N_686), 
            .O(n20));
    defparam i8_4_lut_adj_860.LUT_INIT = 16'h0100;
    SB_LUT4 i1_2_lut_adj_861 (.I0(\count[0] [10]), .I1(n5), .I2(GND_net), 
            .I3(GND_net), .O(n13));
    defparam i1_2_lut_adj_861.LUT_INIT = 16'h2222;
    SB_LUT4 i10_4_lut_adj_862 (.I0(n13), .I1(n20), .I2(n8), .I3(n38149), 
            .O(n22));
    defparam i10_4_lut_adj_862.LUT_INIT = 16'h0008;
    SB_LUT4 i29817_4_lut (.I0(n2), .I1(n3), .I2(n10), .I3(n1), .O(n36420));
    defparam i29817_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut (.I0(n36420), .I1(pause_counter_0__N_712), .I2(pwm_out_0__N_682), 
            .I3(n22), .O(n17287));
    defparam i1_4_lut.LUT_INIT = 16'h4c0c;
    SB_LUT4 i3_4_lut (.I0(\half_duty[0][4] ), .I1(\half_duty[0][1] ), .I2(\count[0] [4]), 
            .I3(\count[0] [1]), .O(n14_adj_4334));   // vhdl/pwm.vhd(80[8:31])
    defparam i3_4_lut.LUT_INIT = 16'h7bde;
    SB_LUT4 i7_4_lut_adj_863 (.I0(\count[0] [0]), .I1(n14_adj_4334), .I2(\count[0] [10]), 
            .I3(\half_duty[0][0] ), .O(n18_adj_4335));   // vhdl/pwm.vhd(80[8:31])
    defparam i7_4_lut_adj_863.LUT_INIT = 16'hfdfe;
    SB_LUT4 i5_4_lut (.I0(\half_duty[0][3] ), .I1(\half_duty[0][2] ), .I2(\count[0] [3]), 
            .I3(\count[0] [2]), .O(n16));   // vhdl/pwm.vhd(80[8:31])
    defparam i5_4_lut.LUT_INIT = 16'h7bde;
    SB_LUT4 i6_4_lut (.I0(\count[0] [6]), .I1(\count[0] [9]), .I2(\half_duty[0][6] ), 
            .I3(\count[0] [8]), .O(n17));   // vhdl/pwm.vhd(80[8:31])
    defparam i6_4_lut.LUT_INIT = 16'hffde;
    SB_LUT4 i4_4_lut (.I0(\half_duty[0][7] ), .I1(\count[0] [5]), .I2(\count[0] [7]), 
            .I3(\half_duty[0] [5]), .O(n15));   // vhdl/pwm.vhd(80[8:31])
    defparam i4_4_lut.LUT_INIT = 16'h7bde;
    SB_LUT4 i10_4_lut_adj_864 (.I0(n15), .I1(n17), .I2(n16), .I3(n18_adj_4335), 
            .O(pwm_out_0__N_682));   // vhdl/pwm.vhd(80[8:31])
    defparam i10_4_lut_adj_864.LUT_INIT = 16'hfffe;
    SB_DFF half_duty_new_i3 (.Q(\half_duty_new[2] ), .C(CLK_c), .D(half_duty_new_9__N_764[2]));   // vhdl/pwm.vhd(59[5] 95[12])
    SB_DFF half_duty_new_i4 (.Q(\half_duty_new[3] ), .C(CLK_c), .D(half_duty_new_9__N_764[3]));   // vhdl/pwm.vhd(59[5] 95[12])
    SB_DFF half_duty_new_i5 (.Q(\half_duty_new[4] ), .C(CLK_c), .D(half_duty_new_9__N_764[4]));   // vhdl/pwm.vhd(59[5] 95[12])
    SB_DFF half_duty_new_i6 (.Q(half_duty_new[5]), .C(CLK_c), .D(half_duty_new_9__N_764[5]));   // vhdl/pwm.vhd(59[5] 95[12])
    SB_DFF half_duty_new_i7 (.Q(\half_duty_new[6] ), .C(CLK_c), .D(half_duty_new_9__N_764[6]));   // vhdl/pwm.vhd(59[5] 95[12])
    SB_DFF half_duty_new_i8 (.Q(\half_duty_new[7] ), .C(CLK_c), .D(half_duty_new_9__N_764[7]));   // vhdl/pwm.vhd(59[5] 95[12])
    SB_LUT4 pwm_out_0__I_21_7_lut (.I0(\count[0] [5]), .I1(GND_net), .I2(pwm_out_0__N_687[5]), 
            .I3(n27901), .O(n38149)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_out_0__I_21_7_lut.LUT_INIT = 16'h6996;
    SB_CARRY pwm_out_0__I_21_7 (.CI(n27901), .I0(GND_net), .I1(pwm_out_0__N_687[5]), 
            .CO(n27902));
    SB_LUT4 pwm_out_0__I_21_6_lut (.I0(\count[0] [4]), .I1(GND_net), .I2(pwm_out_0__N_687[4]), 
            .I3(n27900), .O(n5)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_out_0__I_21_6_lut.LUT_INIT = 16'h6996;
    SB_CARRY pwm_out_0__I_21_6 (.CI(n27900), .I0(GND_net), .I1(pwm_out_0__N_687[4]), 
            .CO(n27901));
    SB_LUT4 half_duty_0__9__I_0_i8_1_lut (.I0(\half_duty[0][7] ), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(pwm_out_0__N_687[7]));   // vhdl/pwm.vhd(84[22:28])
    defparam half_duty_0__9__I_0_i8_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 pwm_out_0__I_21_5_lut (.I0(\count[0] [3]), .I1(GND_net), .I2(pwm_out_0__N_687[3]), 
            .I3(n27899), .O(n4)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_out_0__I_21_5_lut.LUT_INIT = 16'h6996;
    SB_CARRY pwm_out_0__I_21_5 (.CI(n27899), .I0(GND_net), .I1(pwm_out_0__N_687[3]), 
            .CO(n27900));
    SB_LUT4 pwm_out_0__I_21_4_lut (.I0(\count[0] [2]), .I1(GND_net), .I2(pwm_out_0__N_687[2]), 
            .I3(n27898), .O(n3)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_out_0__I_21_4_lut.LUT_INIT = 16'h6996;
    SB_CARRY pwm_out_0__I_21_4 (.CI(n27898), .I0(GND_net), .I1(pwm_out_0__N_687[2]), 
            .CO(n27899));
    SB_LUT4 pwm_out_0__I_21_3_lut (.I0(\count[0] [1]), .I1(GND_net), .I2(pwm_out_0__N_687[1]), 
            .I3(n27897), .O(n2)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_out_0__I_21_3_lut.LUT_INIT = 16'h6996;
    SB_CARRY pwm_out_0__I_21_3 (.CI(n27897), .I0(GND_net), .I1(pwm_out_0__N_687[1]), 
            .CO(n27898));
    SB_LUT4 pwm_out_0__I_21_2_lut (.I0(\count[0] [0]), .I1(GND_net), .I2(pwm_out_0__N_687[0]), 
            .I3(VCC_net), .O(n1)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_out_0__I_21_2_lut.LUT_INIT = 16'h6996;
    SB_CARRY pwm_out_0__I_21_2 (.CI(VCC_net), .I0(GND_net), .I1(pwm_out_0__N_687[0]), 
            .CO(n27897));
    SB_LUT4 count_0__1525_add_4_12_lut (.I0(GND_net), .I1(GND_net), .I2(\count[0] [10]), 
            .I3(n28475), .O(n49[10])) /* synthesis syn_instantiated=1 */ ;
    defparam count_0__1525_add_4_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 count_0__1525_add_4_11_lut (.I0(GND_net), .I1(GND_net), .I2(\count[0] [9]), 
            .I3(n28474), .O(n49[9])) /* synthesis syn_instantiated=1 */ ;
    defparam count_0__1525_add_4_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY count_0__1525_add_4_11 (.CI(n28474), .I0(GND_net), .I1(\count[0] [9]), 
            .CO(n28475));
    SB_LUT4 count_0__1525_add_4_10_lut (.I0(GND_net), .I1(GND_net), .I2(\count[0] [8]), 
            .I3(n28473), .O(n49[8])) /* synthesis syn_instantiated=1 */ ;
    defparam count_0__1525_add_4_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY count_0__1525_add_4_10 (.CI(n28473), .I0(GND_net), .I1(\count[0] [8]), 
            .CO(n28474));
    SB_LUT4 count_0__1525_add_4_9_lut (.I0(GND_net), .I1(GND_net), .I2(\count[0] [7]), 
            .I3(n28472), .O(n49[7])) /* synthesis syn_instantiated=1 */ ;
    defparam count_0__1525_add_4_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY count_0__1525_add_4_9 (.CI(n28472), .I0(GND_net), .I1(\count[0] [7]), 
            .CO(n28473));
    SB_LUT4 count_0__1525_add_4_8_lut (.I0(GND_net), .I1(GND_net), .I2(\count[0] [6]), 
            .I3(n28471), .O(n49[6])) /* synthesis syn_instantiated=1 */ ;
    defparam count_0__1525_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY count_0__1525_add_4_8 (.CI(n28471), .I0(GND_net), .I1(\count[0] [6]), 
            .CO(n28472));
    SB_LUT4 count_0__1525_add_4_7_lut (.I0(GND_net), .I1(GND_net), .I2(\count[0] [5]), 
            .I3(n28470), .O(n49[5])) /* synthesis syn_instantiated=1 */ ;
    defparam count_0__1525_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY count_0__1525_add_4_7 (.CI(n28470), .I0(GND_net), .I1(\count[0] [5]), 
            .CO(n28471));
    SB_LUT4 i17252_3_lut (.I0(\half_duty[0] [5]), .I1(half_duty_new[5]), 
            .I2(n1466), .I3(GND_net), .O(n22073));
    defparam i17252_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 count_0__1525_add_4_6_lut (.I0(GND_net), .I1(GND_net), .I2(\count[0] [4]), 
            .I3(n28469), .O(n49[4])) /* synthesis syn_instantiated=1 */ ;
    defparam count_0__1525_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY count_0__1525_add_4_6 (.CI(n28469), .I0(GND_net), .I1(\count[0] [4]), 
            .CO(n28470));
    SB_LUT4 count_0__1525_add_4_5_lut (.I0(GND_net), .I1(GND_net), .I2(\count[0] [3]), 
            .I3(n28468), .O(n49[3])) /* synthesis syn_instantiated=1 */ ;
    defparam count_0__1525_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY count_0__1525_add_4_5 (.CI(n28468), .I0(GND_net), .I1(\count[0] [3]), 
            .CO(n28469));
    SB_LUT4 count_0__1525_add_4_4_lut (.I0(GND_net), .I1(GND_net), .I2(\count[0] [2]), 
            .I3(n28467), .O(n49[2])) /* synthesis syn_instantiated=1 */ ;
    defparam count_0__1525_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY count_0__1525_add_4_4 (.CI(n28467), .I0(GND_net), .I1(\count[0] [2]), 
            .CO(n28468));
    SB_LUT4 count_0__1525_add_4_3_lut (.I0(GND_net), .I1(GND_net), .I2(\count[0] [1]), 
            .I3(n28466), .O(n49[1])) /* synthesis syn_instantiated=1 */ ;
    defparam count_0__1525_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY count_0__1525_add_4_3 (.CI(n28466), .I0(GND_net), .I1(\count[0] [1]), 
            .CO(n28467));
    SB_LUT4 count_0__1525_add_4_2_lut (.I0(GND_net), .I1(GND_net), .I2(\count[0] [0]), 
            .I3(VCC_net), .O(n49[0])) /* synthesis syn_instantiated=1 */ ;
    defparam count_0__1525_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY count_0__1525_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(\count[0] [0]), 
            .CO(n28466));
    SB_DFF half_duty_0___i1 (.Q(\half_duty[0][0] ), .C(CLK_c), .D(n17710));   // vhdl/pwm.vhd(59[5] 95[12])
    SB_LUT4 i3_2_lut_2_lut (.I0(\count[0] [3]), .I1(pause_counter_0), .I2(GND_net), 
            .I3(GND_net), .O(n14));
    defparam i3_2_lut_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 add_2202_24_lut (.I0(GND_net), .I1(n6168[22]), .I2(pwm_setpoint[22]), 
            .I3(n28290), .O(half_duty_new_9__N_764[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2202_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2202_23_lut (.I0(GND_net), .I1(n6168[21]), .I2(pwm_setpoint[21]), 
            .I3(n28289), .O(half_duty_new_9__N_764[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2202_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2202_23 (.CI(n28289), .I0(n6168[21]), .I1(pwm_setpoint[21]), 
            .CO(n28290));
    SB_LUT4 add_2202_22_lut (.I0(GND_net), .I1(n6168[20]), .I2(pwm_setpoint[20]), 
            .I3(n28288), .O(half_duty_new_9__N_764[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2202_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2202_22 (.CI(n28288), .I0(n6168[20]), .I1(pwm_setpoint[20]), 
            .CO(n28289));
    SB_LUT4 add_2202_21_lut (.I0(GND_net), .I1(n6168[19]), .I2(pwm_setpoint[19]), 
            .I3(n28287), .O(half_duty_new_9__N_764[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2202_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2202_21 (.CI(n28287), .I0(n6168[19]), .I1(pwm_setpoint[19]), 
            .CO(n28288));
    SB_LUT4 add_2202_20_lut (.I0(GND_net), .I1(n6168[18]), .I2(pwm_setpoint[18]), 
            .I3(n28286), .O(half_duty_new_9__N_764[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2202_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2202_20 (.CI(n28286), .I0(n6168[18]), .I1(pwm_setpoint[18]), 
            .CO(n28287));
    SB_LUT4 add_2202_19_lut (.I0(GND_net), .I1(n6168[17]), .I2(pwm_setpoint[17]), 
            .I3(n28285), .O(half_duty_new_9__N_764[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2202_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2202_19 (.CI(n28285), .I0(n6168[17]), .I1(pwm_setpoint[17]), 
            .CO(n28286));
    SB_LUT4 add_2202_18_lut (.I0(GND_net), .I1(n6168[16]), .I2(pwm_setpoint[16]), 
            .I3(n28284), .O(half_duty_new_9__N_764[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2202_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2202_18 (.CI(n28284), .I0(n6168[16]), .I1(pwm_setpoint[16]), 
            .CO(n28285));
    SB_LUT4 add_2202_17_lut (.I0(GND_net), .I1(n6168[15]), .I2(pwm_setpoint[15]), 
            .I3(n28283), .O(half_duty_new_9__N_764[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2202_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2202_17 (.CI(n28283), .I0(n6168[15]), .I1(pwm_setpoint[15]), 
            .CO(n28284));
    SB_CARRY add_2202_16 (.CI(n28282), .I0(n6168[14]), .I1(pwm_setpoint[14]), 
            .CO(n28283));
    SB_CARRY add_2202_15 (.CI(n28281), .I0(n6168[13]), .I1(pwm_setpoint[13]), 
            .CO(n28282));
    SB_CARRY add_2202_14 (.CI(n28280), .I0(n6168[12]), .I1(pwm_setpoint[12]), 
            .CO(n28281));
    SB_CARRY add_2202_13 (.CI(n28279), .I0(n6168[11]), .I1(pwm_setpoint[11]), 
            .CO(n28280));
    SB_CARRY add_2202_12 (.CI(n28278), .I0(n6168[10]), .I1(pwm_setpoint[10]), 
            .CO(n28279));
    SB_CARRY add_2202_11 (.CI(n28277), .I0(n6168[9]), .I1(pwm_setpoint[9]), 
            .CO(n28278));
    SB_CARRY add_2202_10 (.CI(n28276), .I0(n6168[8]), .I1(pwm_setpoint[8]), 
            .CO(n28277));
    SB_CARRY add_2202_9 (.CI(n28275), .I0(n6168[7]), .I1(pwm_setpoint[7]), 
            .CO(n28276));
    SB_CARRY add_2202_8 (.CI(n28274), .I0(n6168[6]), .I1(pwm_setpoint[6]), 
            .CO(n28275));
    SB_CARRY add_2202_7 (.CI(n28273), .I0(n6168[5]), .I1(pwm_setpoint[5]), 
            .CO(n28274));
    SB_CARRY add_2202_6 (.CI(n28272), .I0(n6168[4]), .I1(pwm_setpoint[4]), 
            .CO(n28273));
    SB_CARRY add_2202_5 (.CI(n28271), .I0(n6168[3]), .I1(pwm_setpoint[3]), 
            .CO(n28272));
    SB_CARRY add_2202_4 (.CI(n28270), .I0(n6168[2]), .I1(pwm_setpoint[2]), 
            .CO(n28271));
    SB_CARRY add_2202_3 (.CI(n28269), .I0(n6168[1]), .I1(pwm_setpoint[1]), 
            .CO(n28270));
    SB_CARRY add_2202_2 (.CI(GND_net), .I0(pwm_setpoint[3]), .I1(pwm_setpoint[0]), 
            .CO(n28269));
    SB_LUT4 add_2208_23_lut (.I0(GND_net), .I1(pwm_setpoint[21]), .I2(GND_net), 
            .I3(n28268), .O(n6168[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2208_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2208_22_lut (.I0(GND_net), .I1(pwm_setpoint[20]), .I2(GND_net), 
            .I3(n28267), .O(n6168[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2208_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2208_22 (.CI(n28267), .I0(pwm_setpoint[20]), .I1(GND_net), 
            .CO(n28268));
    SB_LUT4 add_2208_21_lut (.I0(GND_net), .I1(pwm_setpoint[19]), .I2(GND_net), 
            .I3(n28266), .O(n6168[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2208_21_lut.LUT_INIT = 16'hC33C;
    
endmodule
//
// Verilog Description of module motorControl
//

module motorControl (PWMLimit, duty, GND_net, \Ki[11] , \Kp[15] , 
            \Kp[9] , \Ki[6] , \Ki[13] , \Ki[14] , \Ki[1] , \Ki[0] , 
            \Ki[15] , \Ki[2] , \Ki[3] , \Ki[4] , IntegralLimit, \Ki[5] , 
            \Kp[10] , \Ki[7] , \Kp[2] , \Kp[1] , \Ki[12] , \Kp[11] , 
            \Kp[0] , n38238, \Kp[3] , \Ki[8] , \Kp[5] , \Kp[6] , 
            \Kp[7] , \Kp[8] , \Ki[9] , \Kp[4] , \Kp[12] , \Kp[13] , 
            setpoint, \Kp[14] , \Ki[10] , VCC_net, n25, clk32MHz, 
            motor_state) /* synthesis lattice_noprune=1, syn_preserve=0, syn_module_defined=1, syn_noprune=0 */ ;
    input [23:0]PWMLimit;
    output [23:0]duty;
    input GND_net;
    input \Ki[11] ;
    input \Kp[15] ;
    input \Kp[9] ;
    input \Ki[6] ;
    input \Ki[13] ;
    input \Ki[14] ;
    input \Ki[1] ;
    input \Ki[0] ;
    input \Ki[15] ;
    input \Ki[2] ;
    input \Ki[3] ;
    input \Ki[4] ;
    input [23:0]IntegralLimit;
    input \Ki[5] ;
    input \Kp[10] ;
    input \Ki[7] ;
    input \Kp[2] ;
    input \Kp[1] ;
    input \Ki[12] ;
    input \Kp[11] ;
    input \Kp[0] ;
    output n38238;
    input \Kp[3] ;
    input \Ki[8] ;
    input \Kp[5] ;
    input \Kp[6] ;
    input \Kp[7] ;
    input \Kp[8] ;
    input \Ki[9] ;
    input \Kp[4] ;
    input \Kp[12] ;
    input \Kp[13] ;
    input [23:0]setpoint;
    input \Kp[14] ;
    input \Ki[10] ;
    input VCC_net;
    input n25;
    input clk32MHz;
    input [23:0]motor_state;
    
    wire clk32MHz /* synthesis SET_AS_NETWORK=clk32MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(34[6:14])
    
    wire n31, n29107;
    wire [21:0]n8273;
    
    wire n366, n29108;
    wire [9:0]n8495;
    wire [8:0]n8507;
    
    wire n770, n29299, n23, n25_c;
    wire [23:0]n257;
    wire [23:0]n1;
    
    wire n28113;
    wire [23:0]n3265;
    
    wire n293, n29106, n24379, n28114;
    wire [23:0]\PID_CONTROLLER.integral ;   // verilog/motorControl.v(31[23:31])
    
    wire n840;
    wire [23:0]\PID_CONTROLLER.err ;   // verilog/motorControl.v(29[23:26])
    
    wire n1114;
    wire [15:0]n8699;
    wire [14:0]n8717;
    
    wire n29473, n697, n29298, n220, n29105, n1117, n29472, n147, 
        n29104, n33, n694, n460, n624, n29297, n1044, n29471, 
        n5, n74, n35, n551, n29296, n971, n29470, n11, n898, 
        n29469, n478, n29295, n13, n825, n29468, n405, n29294, 
        n752, n29467, n332, n29293, n259, n29292, n28112, n679, 
        n29466, n186, n29291, n606, n29465, n44, n113;
    wire [10:0]n8482;
    
    wire n840_adj_3906, n29290, n15, n533, n29464, n767, n29289, 
        n28111, n28110, n956, n29463, n29288, n1029, n113_adj_3907, 
        n44_adj_3908, n1102, n186_adj_3909, n259_adj_3910, n27;
    wire [47:0]n155;
    
    wire n256;
    wire [23:0]n3290;
    
    wire n9, n17, n19, n332_adj_3911, n21_adj_3912, n37509;
    wire [23:0]n1_adj_4332;
    
    wire n37502, n387, n29462, n12, n30, n37558, n37839, n405_adj_3913, 
        n37827, n38073, n29, n37959, n37, n38103, n6, n38019, 
        n38020, n621, n29287, n16, n45, n24_adj_3914, n43, n37482, 
        n8, n37480, n37929, n37744, n4, n37957, n314, n29461, 
        n241, n29460, n37958, n37498, n10, n37494, n38067, n37746, 
        n38117, n38118, n39, n38106, n41, n37484, n38055, n37752, 
        n38101, duty_23__N_3637;
    wire [23:0]duty_23__N_3613;
    wire [23:0]duty_23__N_3490;
    
    wire n822, n183, n95, n895, n168, n29459, n548, n29286, 
        n26, n256_adj_3915, n26_adj_3916, n95_adj_3917, n9_adj_3918, 
        n11_adj_3919, n13_adj_3920, n15_adj_3921, n21_adj_3923, n19_adj_3924, 
        n17_adj_3925, n23_adj_3926, n393;
    wire [16:0]n8680;
    
    wire n29458, n439, n116, n28109, n475, n29285, n47, n512, 
        n98, n29_adj_3928, n585, n658, n189, n478_adj_3930, n731, 
        n402, n29284, n387_adj_3931, n968, n1041, n83, n14, n262, 
        n329, n1114_adj_3933, n804, n460_adj_3934, n156, n335, n533_adj_3935, 
        n524, n229, n877, n606_adj_3937, n335_adj_3938, n302, n442, 
        n950, n408, n171, n408_adj_3939;
    wire [23:0]n1_adj_4333;
    
    wire n515, n29457, n588, n597, n661, n679_adj_3942, n466, 
        n752_adj_3944, n375, n539, n734, n825_adj_3945, n448, n481, 
        n898_adj_3946, n521, n971_adj_3947, n594, n1023, n481_adj_3948, 
        n554, n244, n1096, n1044_adj_3951, n554_adj_3952, n317, 
        n1117_adj_3955, n29456, n98_adj_3956, n29_adj_3957, n667, 
        n29283, n627, n29455, n29454, n171_adj_3959, n244_adj_3960, 
        n740, n700, n317_adj_3961, n37256, n627_adj_3963, n813, 
        n390, n886, n119, n50, n390_adj_3964, n700_adj_3965, n551_adj_3966, 
        n624_adj_3967, n168_adj_3969, n119_adj_3970;
    wire [23:0]\PID_CONTROLLER.integral_23__N_3589 ;
    
    wire n28108, n697_adj_3971, n50_adj_3972, n807, n770_adj_3974, 
        n241_adj_3975, n116_adj_3976, n47_adj_3977, n612, n314_adj_3978, 
        n880, n953, n1026, n1099, n463, n192_adj_3979, n685, n29282, 
        n45_adj_3983, n28107, n29453, n265, n338, n29281, n536, 
        n29452, n670, n411;
    wire [23:0]\PID_CONTROLLER.err_23__N_3514 ;
    
    wire n758, n609, n41_adj_3989, n110, n749, n29451;
    wire [11:0]n8468;
    
    wire n910, n29280, n682, n80, n11_adj_3990, n484, n153, n755, 
        n743, n557, n630, n676, n29450, n837, n29279, n764, 
        n29278, n691, n29277, n226, n603, n29449, n530, n29448, 
        n122, n53, n457, n29447, n618, n29276, n828, n384, n29446, 
        n299, n195_adj_3992, n901, n311, n29445, n189_adj_3994, 
        n545, n29275, n372, n268, n831, n238, n29444, n816, 
        n889, n43_adj_3997, n28106, n904, n165, n29443, n962, 
        n23_adj_4000, n92, n472, n29274;
    wire [17:0]n8660;
    
    wire n29442, n29441, n29440, n399, n29273, n326, n29272, n253, 
        n29271, n180, n29270, n1035, n1111, n29439, n977, n37_adj_4002, 
        n35_adj_4003, n33_adj_4004, n37935, n38095, n1050, n43_adj_4005, 
        n16_adj_4006, n38, n107, n1108, n104, n445, n341, n35_adj_4007, 
        n89, n20_adj_4009, n177, n162, n37312, n250, n235, n308, 
        n381, n323, n454, n396, n41_adj_4011, n28105, n1038, n29438, 
        n527;
    wire [12:0]n8453;
    
    wire n980, n29269, n965, n29437, n518, n892, n29436;
    wire [20:0]n8297;
    
    wire n28735, n28734, n907, n29268, n28733, n834, n29267, n600, 
        n469, n819, n29435, n39_adj_4014, n28104, n746, n29434, 
        n28732, n761, n29266, n6_adj_4016, n37949, n673, n29433, 
        n463_adj_4017, n542, n615, n688, n29265, n29264, n29263, 
        n29262, n591, n29432, n29431, n29261, n29430, n29260, 
        n29429, n29428, n37950, n414, n29427, n29259, n27993, 
        n29426, n29258;
    wire [18:0]n8639;
    
    wire n29425, n974, n29424, n29423, n29422, n29421, n1047;
    wire [13:0]n8437;
    
    wire n29257, n29256, n29420, n37_adj_4020, n28103, n959, n29419, 
        n1120, n192_adj_4022, n487, n29255, n27992, n560, n29418, 
        n664, n35_adj_4023, n28102, n29417, n29254, n27991, n29416, 
        n28731, n33_adj_4025, n28101, n29253, n27990, n29415, n1032, 
        n31_adj_4026, n28100, n29252, n265_adj_4027, n28730, n28729, 
        n28728, n28727, n28726, n28725, n29251, n536_adj_4029, n338_adj_4030, 
        n411_adj_4031, n609_adj_4033, n28724, n28723, n125, n29250, 
        n29249, n8_adj_4036, n56, n45_adj_4038, n24_adj_4039, n27989, 
        n28722, n29414, n28721, n1105, n484_adj_4040, n28720, n28719, 
        n682_adj_4041, n755_adj_4042, n737, n29413, n29248, n810, 
        n4_adj_4045;
    wire [3:0]n8849;
    
    wire n6_adj_4046;
    wire [4:0]n8842;
    wire [23:0]n28;
    
    wire \PID_CONTROLLER.integral_23__N_3586 , n25_adj_4049, n37464, n37425, 
        n29_adj_4050, n28099;
    wire [5:0]n8834;
    
    wire n35470, n490, n29568, n37423, n37931, n27_adj_4052, n28098, 
        n198, n451, n29412, n37754, n369, n28718, n417, n29567, 
        n883, n4_adj_4054, n378, n29411, n320, n29247, n27988, 
        n101, n32, n25_adj_4055, n28097, n27987, n27_adj_4058, n37947, 
        n344, n29566, n557_adj_4059, n296, n28717, n630_adj_4060, 
        n27714, n223, n28716, n150, n28715, n247, n29246, n305, 
        n29410, n271_adj_4061, n271_adj_4062, n29565, n232, n29409, 
        n174, n29245, n32_adj_4063, n101_adj_4064, n956_adj_4065, 
        n198_adj_4067, n29564, n159, n29408, n17_adj_4068, n86, 
        n8_adj_4069, n77, n344_adj_4070, n29_adj_4071, n37948, n1029_adj_4072, 
        n31_adj_4073, n37456, n37452, n174_adj_4074, n30_adj_4075, 
        n10_adj_4076, n37446, n38111, n27757, n37756, n828_adj_4077, 
        n1102_adj_4080, n417_adj_4081, n6_adj_4082;
    wire [3:0]n8552;
    wire [4:0]n8545;
    
    wire n38143, n38144, n39_adj_4084, n38134, n23_adj_4085, n28096, 
        n56_adj_4087, n125_adj_4088, n27986;
    wire [14:0]n8420;
    
    wire n1120_adj_4089, n29244;
    wire [19:0]n8617;
    
    wire n29407, n1047_adj_4090, n29243;
    wire [6:0]n8825;
    
    wire n560_adj_4091, n29563, n487_adj_4092, n29562, n414_adj_4093, 
        n29561, n29406, n122_adj_4094;
    wire [2:0]n8855;
    
    wire n4_adj_4095, n27791;
    wire [1:0]n8860;
    
    wire n4_adj_4096, n204;
    wire [1:0]n8563;
    
    wire n29405, n341_adj_4097, n29560, n974_adj_4098, n29242, n268_adj_4099, 
        n29559, n29404, n21_adj_4100, n28095, n901_adj_4102, n29241, 
        n19_adj_4103, n28094, n17_adj_4105, n28093, n195_adj_4107, 
        n29558, n29403, n53_adj_4108, n131, n15_adj_4109, n28092, 
        n29240;
    wire [7:0]n8815;
    
    wire n29557, n29556, n62, n27985, n13_adj_4110, n28091, n29239, 
        n29238, n29555, n29402, n4_adj_4111;
    wire [2:0]n8558;
    
    wire n490_adj_4112, n12_adj_4113, n29237, n8_adj_4114, n11_adj_4115, 
        n29554, n29553, n29236, n29552, n29401, n6_adj_4116, n27646, 
        n18_adj_4117, n13_adj_4118, n4_adj_4119, n34771, n29551, n29400, 
        n27984, n29235, n77_adj_4120, n8_adj_4121, n247_adj_4122;
    wire [0:0]n7788;
    
    wire n150_adj_4125, n83_adj_4126, n14_adj_4127, n223_adj_4128, n320_adj_4129, 
        n156_adj_4131, n393_adj_4132, n296_adj_4133, n229_adj_4134, 
        n302_adj_4135, n369_adj_4136, n466_adj_4137, n41_adj_4139, n37427, 
        n375_adj_4140, n442_adj_4141, n515_adj_4142, n448_adj_4143, 
        n539_adj_4144, n521_adj_4146, n38059, n588_adj_4147, n594_adj_4148, 
        n612_adj_4149, n40, n667_adj_4150, n661_adj_4151, n740_adj_4152, 
        n734_adj_4153, n685_adj_4154, n813_adj_4155, n886_adj_4156, 
        n807_adj_4157, n959_adj_4158, n880_adj_4159, n758_adj_4160, 
        n1032_adj_4161, n953_adj_4162, n1105_adj_4163, n1026_adj_4164, 
        n831_adj_4165, n1099_adj_4166, n904_adj_4167, n86_adj_4169, 
        n17_adj_4170, n977_adj_4171, n159_adj_4172, n1050_adj_4173, 
        n232_adj_4174, n305_adj_4175, n378_adj_4176, n104_adj_4177, 
        n35_adj_4178, n451_adj_4179, n524_adj_4180, n177_adj_4181, n74_adj_4182, 
        n5_adj_4183, n11_adj_4184, n28090, n597_adj_4185, n147_adj_4186, 
        n670_adj_4187, n250_adj_4188, n220_adj_4189, n743_adj_4190, 
        n38061, n293_adj_4192, n323_adj_4193, n816_adj_4195, n889_adj_4196, 
        n366_adj_4197, n962_adj_4198, n396_adj_4199, n439_adj_4200, 
        n1035_adj_4201, n512_adj_4202, n1108_adj_4203, n469_adj_4204, 
        n542_adj_4205, n615_adj_4206, n585_adj_4207, n688_adj_4208, 
        n658_adj_4209, n761_adj_4210, n89_adj_4211, n20_adj_4212, n162_adj_4213, 
        n731_adj_4214, n235_adj_4215, n804_adj_4216, n834_adj_4217, 
        n308_adj_4218, n877_adj_4219, n907_adj_4220, n381_adj_4221, 
        n29399, n29234, n29398, n29233, n454_adj_4222;
    wire [8:0]n8804;
    
    wire n29550, n29397, n29232, n29231, n29549, n29396, n950_adj_4223, 
        n980_adj_4224, n1023_adj_4225, n527_adj_4226, n107_adj_4227, 
        n38_adj_4228;
    wire [15:0]n8402;
    
    wire n29230, n29229, n600_adj_4229, n29228, n27983, n29548, 
        n29395, n29227, n29394, n29226, n27982, n29547, n29393, 
        n29225, n29392, n29224, n29223, n27981, n673_adj_4230, n29546, 
        n29391, n29222, n9_adj_4231, n28089, n29390, n29221, n1096_adj_4232, 
        n29545, n29389, n29220, n7_adj_4233, n28088, n29219, n180_adj_4234, 
        n746_adj_4235, n47_adj_4236, n262_adj_4237, n29544, n29543;
    wire [20:0]n8594;
    
    wire n29388, n29218, n29387, n29386, n29217, n27980, n29385;
    wire [9:0]n8792;
    
    wire n29542, n29541, n29216, n29384, n29540, n253_adj_4238, 
        n29539, n819_adj_4239, n326_adj_4240, n892_adj_4241, n965_adj_4242, 
        n1038_adj_4243, n399_adj_4244, n472_adj_4245, n1111_adj_4246, 
        n545_adj_4247, n80_adj_4248, n11_adj_4249, n27979, n153_adj_4250, 
        n618_adj_4251, n29538, n92_adj_4252, n23_adj_4253, n5_adj_4254, 
        n28087, n226_adj_4255, n165_adj_4256, n299_adj_4257, n691_adj_4258, 
        n238_adj_4259, n311_adj_4260, n372_adj_4261, n384_adj_4262, 
        n457_adj_4264, n445_adj_4265, n764_adj_4266, n837_adj_4267, 
        n910_adj_4268, n110_adj_4269, n29537, n41_adj_4270, n518_adj_4271, 
        n530_adj_4272, n183_adj_4273, n603_adj_4274, n29383, n3_adj_4275, 
        n28086, n591_adj_4276, n29536, n27978;
    wire [16:0]n8383;
    
    wire n29215, n29535, n29534, n256_adj_4277, n29214, n29382, 
        n29381, n29380, n29213;
    wire [10:0]n8779;
    
    wire n29533, n27977, n767_adj_4278, n29532, n1041_adj_4279, n29212, 
        n883_adj_4280, n29379, n694_adj_4281, n29531, n968_adj_4282, 
        n29211, n4_adj_4284, n676_adj_4285, n27544, n621_adj_4286, 
        n29530, n329_adj_4287, n402_adj_4288, n749_adj_4290, n475_adj_4291, 
        n664_adj_4292, n822_adj_4293, n548_adj_4294, n737_adj_4295, 
        n27976, n810_adj_4296, n895_adj_4297, n29210, n29378, n8_adj_4298, 
        n29377, n29529, n29209, n29376, n27621, n29528, n29208, 
        n27975, n29527, n29526, n29207, n12_adj_4300, n8_adj_4301, 
        n29525, n11_adj_4302, n6_adj_4303, n27816, n18_adj_4304, n13_adj_4305, 
        n29375, n29206, n29524, n29205, n29374, n27974;
    wire [11:0]n8765;
    
    wire n29523, n29522, n29521, n29373, n29204, n29203, n29372, 
        n29202, n29201, n29520, n29371, n29200, n29370, n29519, 
        n29369;
    wire [17:0]n8363;
    
    wire n29199, n27973, n17_adj_4306, n9_adj_4307, n29198, n11_adj_4308, 
        n37397, n37393, n39123, n37899, n37683, n27972, n29197, 
        n39105, n37681, n37679, n39098, n37603, n37609, n16_adj_4309, 
        n37560, n8_adj_4310, n24_adj_4311, n37625, n29518, n12_adj_4312;
    wire [21:0]n8570;
    
    wire n29368, n29196, n29367, n29517, n37871, n37867, n38083, 
        n29516, n29366, n29195, n37975, n27971, n29365, n28498, 
        n28497, n28496, n28495, n28494, n28493, n29194, n28492, 
        n29364, n29193, n28491, n28490, n29515, n29363, n38107, 
        n28489, n29192, n37685, n28488, n29514, n29362, n28487, 
        n39092, n28486, n37891, n39087, n28485, n12_adj_4320, n29191, 
        n37653, n39110, n28484, n10_adj_4321, n30_adj_4322, n29513, 
        n29361, n37993, n28483, n28482, n29360, n29190, n28481, 
        n29189, n28480, n28479, n28478, n28477, n28476, n29188, 
        n29359;
    wire [12:0]n8750;
    
    wire n29512, n29358, n29187, n29186, n29511, n37673, n37478, 
        n37788, n39090, n29357, n29185, n29510, n29356, n29184, 
        n29355, n37991, n29183, n39116, n29509, n29354, n38087;
    wire [18:0]n8342;
    
    wire n29182, n39081, n29508, n29181, n29353, n38127, n29180, 
        n29507, n29506, n29179, n29505, n39078, n29178, n29352, 
        n29177, n29351, n29504, n16_adj_4323, n29176, n29350, n29175, 
        n29174, n37627, n28131, n29503, n29349, n28130, n29173, 
        n29348, n29502, n29172, n29347, n29171, n29501, n29170, 
        n29169, n29346, n29345, n29168, n24_adj_4324, n29167, n6_adj_4325, 
        n38047, n29344, n38048, n29166, n37632;
    wire [13:0]n8734;
    
    wire n29500, n29343, n29165, n39076, n37925, n29499, n29342, 
        n29341;
    wire [19:0]n8320;
    
    wire n29164, n38006, n4_adj_4326, n29163, n28129, n29498, n29340, 
        n29162, n29161, n29339, n37784, n29160, n38025, n38026, 
        n12_adj_4327, n37573, n29497, n29338, n29159, n29337, n10_adj_4328, 
        n29158, n30_adj_4329, n37575, n38091, n29496, n29336, n29157, 
        n29335, n29156, n37736, n38131, n29155, n38132, n38122, 
        n6_adj_4330, n38027, n38028, n37562, n29495, n29334, n29154, 
        n37927, n37734, n29333, n29153, n37564, n29494, n29152, 
        n38053, n37742, n29332, n29151, n28128, n29493, n38099, 
        n29150, n29331, n4_adj_4331, n29330, n29149, n28127, n38031, 
        n38032, n29492, n29329, n29148, n29147, n29328, n29491, 
        n29146, n28126, n29490, n29327, n29145, n29144, n37656, 
        n29326, n29143, n28125, n28124, n38089, n29142, n29489, 
        n29141, n29140;
    wire [5:0]n8537;
    
    wire n29325, n37726, n38129, n29324, n38065, n29139, n28123, 
        n29488, n38130, n38124, n29138, n37635, n29323, n28122, 
        n29137, n29322, n29136, n29321, n28121, n29135, n28120, 
        n29134, n38051, n28313, n28312, n37732, n28311, \PID_CONTROLLER.integral_23__N_3588 , 
        n28310, n38097, n28309, n29133;
    wire [6:0]n8528;
    
    wire n29320, n29319, n29487, n28119, n28308, n29486, n29485, 
        n29318, n29132, n29131, n28307, n28306, n29317, n29130, 
        n28305, n28304, n29316, n29129, n28118, n28303, n29484, 
        n29315, n29128, n29483, n28302, n29127;
    wire [7:0]n8518;
    
    wire n29314, n29313, n29482, n29126, n29312, n29481, n28301, 
        n29480, n28117, n29311, n29125, n29124, n29479, n28300, 
        n29310, n29309, n28299, n29123, n28116, n29308, n29122, 
        n29478, n29121, n28298, n29120, n28115, n29119, n29307, 
        n29477, n28297, n29306, n29118, n28296, n28295, n29476, 
        n28294, n29305, n29117, n29475, n28293, n29304, n29116, 
        n28292, n28291, n29474, n29303, n29115, n29302, n29114, 
        n29113, n29301, n29112, n29300, n29111, n29110, n29109;
    
    SB_LUT4 duty_23__I_0_i31_2_lut (.I0(PWMLimit[15]), .I1(duty[15]), .I2(GND_net), 
            .I3(GND_net), .O(n31));   // verilog/motorControl.v(44[10:25])
    defparam duty_23__I_0_i31_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY mult_10_add_1225_6 (.CI(n29107), .I0(n8273[3]), .I1(n366), 
            .CO(n29108));
    SB_LUT4 add_4122_11_lut (.I0(GND_net), .I1(n8507[8]), .I2(n770), .I3(n29299), 
            .O(n8495[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4122_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 duty_23__I_0_i23_2_lut (.I0(PWMLimit[11]), .I1(duty[11]), .I2(GND_net), 
            .I3(GND_net), .O(n23));   // verilog/motorControl.v(44[10:25])
    defparam duty_23__I_0_i23_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i25_2_lut (.I0(PWMLimit[12]), .I1(duty[12]), .I2(GND_net), 
            .I3(GND_net), .O(n25_c));   // verilog/motorControl.v(44[10:25])
    defparam duty_23__I_0_i25_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 unary_minus_16_add_3_7_lut (.I0(GND_net), .I1(GND_net), .I2(n1[5]), 
            .I3(n28113), .O(n257[5])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_add_1225_5_lut (.I0(n24379), .I1(n8273[2]), .I2(n293), 
            .I3(n29106), .O(n3265[4])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_5_lut.LUT_INIT = 16'h8228;
    SB_CARRY unary_minus_16_add_3_7 (.CI(n28113), .I0(GND_net), .I1(n1[5]), 
            .CO(n28114));
    SB_LUT4 mult_11_i565_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral [12]), 
            .I2(GND_net), .I3(GND_net), .O(n840));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i565_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i749_2_lut (.I0(\Kp[15] ), .I1(\PID_CONTROLLER.err [6]), 
            .I2(GND_net), .I3(GND_net), .O(n1114));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i749_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_4138_17_lut (.I0(GND_net), .I1(n8717[14]), .I2(GND_net), 
            .I3(n29473), .O(n8699[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4138_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4122_10_lut (.I0(GND_net), .I1(n8507[7]), .I2(n697), .I3(n29298), 
            .O(n8495[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4122_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_1225_5 (.CI(n29106), .I0(n8273[2]), .I1(n293), 
            .CO(n29107));
    SB_LUT4 mult_10_add_1225_4_lut (.I0(n24379), .I1(n8273[1]), .I2(n220), 
            .I3(n29105), .O(n3265[3])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_4_lut.LUT_INIT = 16'h8228;
    SB_LUT4 add_4138_16_lut (.I0(GND_net), .I1(n8717[13]), .I2(n1117), 
            .I3(n29472), .O(n8699[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4138_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4122_10 (.CI(n29298), .I0(n8507[7]), .I1(n697), .CO(n29299));
    SB_CARRY mult_10_add_1225_4 (.CI(n29105), .I0(n8273[1]), .I1(n220), 
            .CO(n29106));
    SB_LUT4 mult_10_add_1225_3_lut (.I0(n24379), .I1(n8273[0]), .I2(n147), 
            .I3(n29104), .O(n3265[2])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_3_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_4138_16 (.CI(n29472), .I0(n8717[13]), .I1(n1117), .CO(n29473));
    SB_LUT4 duty_23__I_0_i33_2_lut (.I0(PWMLimit[16]), .I1(duty[16]), .I2(GND_net), 
            .I3(GND_net), .O(n33));   // verilog/motorControl.v(44[10:25])
    defparam duty_23__I_0_i33_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_10_i467_2_lut (.I0(\Kp[9] ), .I1(\PID_CONTROLLER.err [12]), 
            .I2(GND_net), .I3(GND_net), .O(n694));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i467_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i310_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral [7]), 
            .I2(GND_net), .I3(GND_net), .O(n460));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i310_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_4122_9_lut (.I0(GND_net), .I1(n8507[6]), .I2(n624), .I3(n29297), 
            .O(n8495[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4122_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4122_9 (.CI(n29297), .I0(n8507[6]), .I1(n624), .CO(n29298));
    SB_LUT4 add_4138_15_lut (.I0(GND_net), .I1(n8717[12]), .I2(n1044), 
            .I3(n29471), .O(n8699[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4138_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_16_inv_0_i3_1_lut (.I0(PWMLimit[2]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[2]));   // verilog/motorControl.v(47[19:28])
    defparam unary_minus_16_inv_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY mult_10_add_1225_3 (.CI(n29104), .I0(n8273[0]), .I1(n147), 
            .CO(n29105));
    SB_LUT4 mult_10_add_1225_2_lut (.I0(n24379), .I1(n5), .I2(n74), .I3(GND_net), 
            .O(n3265[1])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_2_lut.LUT_INIT = 16'h8228;
    SB_LUT4 duty_23__I_0_i35_2_lut (.I0(PWMLimit[17]), .I1(duty[17]), .I2(GND_net), 
            .I3(GND_net), .O(n35));   // verilog/motorControl.v(44[10:25])
    defparam duty_23__I_0_i35_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_4138_15 (.CI(n29471), .I0(n8717[12]), .I1(n1044), .CO(n29472));
    SB_LUT4 add_4122_8_lut (.I0(GND_net), .I1(n8507[5]), .I2(n551), .I3(n29296), 
            .O(n8495[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4122_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_1225_2 (.CI(GND_net), .I0(n5), .I1(n74), .CO(n29104));
    SB_LUT4 add_4138_14_lut (.I0(GND_net), .I1(n8717[11]), .I2(n971), 
            .I3(n29470), .O(n8699[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4138_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4122_8 (.CI(n29296), .I0(n8507[5]), .I1(n551), .CO(n29297));
    SB_CARRY add_4138_14 (.CI(n29470), .I0(n8717[11]), .I1(n971), .CO(n29471));
    SB_LUT4 duty_23__I_0_i11_2_lut (.I0(PWMLimit[5]), .I1(duty[5]), .I2(GND_net), 
            .I3(GND_net), .O(n11));   // verilog/motorControl.v(44[10:25])
    defparam duty_23__I_0_i11_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_4138_13_lut (.I0(GND_net), .I1(n8717[10]), .I2(n898), 
            .I3(n29469), .O(n8699[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4138_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4122_7_lut (.I0(GND_net), .I1(n8507[4]), .I2(n478), .I3(n29295), 
            .O(n8495[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4122_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4138_13 (.CI(n29469), .I0(n8717[10]), .I1(n898), .CO(n29470));
    SB_CARRY add_4122_7 (.CI(n29295), .I0(n8507[4]), .I1(n478), .CO(n29296));
    SB_LUT4 duty_23__I_0_i13_2_lut (.I0(PWMLimit[6]), .I1(duty[6]), .I2(GND_net), 
            .I3(GND_net), .O(n13));   // verilog/motorControl.v(44[10:25])
    defparam duty_23__I_0_i13_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_4138_12_lut (.I0(GND_net), .I1(n8717[9]), .I2(n825), .I3(n29468), 
            .O(n8699[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4138_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4122_6_lut (.I0(GND_net), .I1(n8507[3]), .I2(n405), .I3(n29294), 
            .O(n8495[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4122_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4138_12 (.CI(n29468), .I0(n8717[9]), .I1(n825), .CO(n29469));
    SB_CARRY add_4122_6 (.CI(n29294), .I0(n8507[3]), .I1(n405), .CO(n29295));
    SB_LUT4 add_4138_11_lut (.I0(GND_net), .I1(n8717[8]), .I2(n752), .I3(n29467), 
            .O(n8699[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4138_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4122_5_lut (.I0(GND_net), .I1(n8507[2]), .I2(n332), .I3(n29293), 
            .O(n8495[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4122_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4122_5 (.CI(n29293), .I0(n8507[2]), .I1(n332), .CO(n29294));
    SB_CARRY add_4138_11 (.CI(n29467), .I0(n8717[8]), .I1(n752), .CO(n29468));
    SB_LUT4 add_4122_4_lut (.I0(GND_net), .I1(n8507[1]), .I2(n259), .I3(n29292), 
            .O(n8495[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4122_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4122_4 (.CI(n29292), .I0(n8507[1]), .I1(n259), .CO(n29293));
    SB_LUT4 unary_minus_16_add_3_6_lut (.I0(GND_net), .I1(GND_net), .I2(n1[4]), 
            .I3(n28112), .O(n257[4])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4138_10_lut (.I0(GND_net), .I1(n8717[7]), .I2(n679), .I3(n29466), 
            .O(n8699[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4138_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4122_3_lut (.I0(GND_net), .I1(n8507[0]), .I2(n186), .I3(n29291), 
            .O(n8495[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4122_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4138_10 (.CI(n29466), .I0(n8717[7]), .I1(n679), .CO(n29467));
    SB_CARRY add_4122_3 (.CI(n29291), .I0(n8507[0]), .I1(n186), .CO(n29292));
    SB_LUT4 add_4138_9_lut (.I0(GND_net), .I1(n8717[6]), .I2(n606), .I3(n29465), 
            .O(n8699[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4138_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4122_2_lut (.I0(GND_net), .I1(n44), .I2(n113), .I3(GND_net), 
            .O(n8495[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4122_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4122_2 (.CI(GND_net), .I0(n44), .I1(n113), .CO(n29291));
    SB_CARRY add_4138_9 (.CI(n29465), .I0(n8717[6]), .I1(n606), .CO(n29466));
    SB_LUT4 add_4121_12_lut (.I0(GND_net), .I1(n8495[9]), .I2(n840_adj_3906), 
            .I3(n29290), .O(n8482[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4121_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 duty_23__I_0_i15_2_lut (.I0(PWMLimit[7]), .I1(duty[7]), .I2(GND_net), 
            .I3(GND_net), .O(n15));   // verilog/motorControl.v(44[10:25])
    defparam duty_23__I_0_i15_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_4138_8_lut (.I0(GND_net), .I1(n8717[5]), .I2(n533), .I3(n29464), 
            .O(n8699[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4138_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4121_11_lut (.I0(GND_net), .I1(n8495[8]), .I2(n767), .I3(n29289), 
            .O(n8482[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4121_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_6 (.CI(n28112), .I0(GND_net), .I1(n1[4]), 
            .CO(n28113));
    SB_LUT4 unary_minus_16_add_3_5_lut (.I0(GND_net), .I1(GND_net), .I2(n1[3]), 
            .I3(n28111), .O(n257[3])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_5 (.CI(n28111), .I0(GND_net), .I1(n1[3]), 
            .CO(n28112));
    SB_CARRY add_4138_8 (.CI(n29464), .I0(n8717[5]), .I1(n533), .CO(n29465));
    SB_CARRY add_4121_11 (.CI(n29289), .I0(n8495[8]), .I1(n767), .CO(n29290));
    SB_LUT4 unary_minus_16_add_3_4_lut (.I0(GND_net), .I1(GND_net), .I2(n1[2]), 
            .I3(n28110), .O(n257[2])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i643_2_lut (.I0(\Ki[13] ), .I1(\PID_CONTROLLER.integral [2]), 
            .I2(GND_net), .I3(GND_net), .O(n956));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i643_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_4138_7_lut (.I0(GND_net), .I1(n8717[4]), .I2(n460), .I3(n29463), 
            .O(n8699[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4138_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4121_10_lut (.I0(GND_net), .I1(n8495[7]), .I2(n694), .I3(n29288), 
            .O(n8482[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4121_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i692_2_lut (.I0(\Ki[14] ), .I1(\PID_CONTROLLER.integral [2]), 
            .I2(GND_net), .I3(GND_net), .O(n1029));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i692_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i77_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral [13]), 
            .I2(GND_net), .I3(GND_net), .O(n113_adj_3907));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i77_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i30_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral [14]), 
            .I2(GND_net), .I3(GND_net), .O(n44_adj_3908));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i30_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i741_2_lut (.I0(\Ki[15] ), .I1(\PID_CONTROLLER.integral [2]), 
            .I2(GND_net), .I3(GND_net), .O(n1102));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i741_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i126_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral [13]), 
            .I2(GND_net), .I3(GND_net), .O(n186_adj_3909));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i126_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i175_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral [13]), 
            .I2(GND_net), .I3(GND_net), .O(n259_adj_3910));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i175_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 duty_23__I_0_i27_2_lut (.I0(PWMLimit[13]), .I1(duty[13]), .I2(GND_net), 
            .I3(GND_net), .O(n27));   // verilog/motorControl.v(44[10:25])
    defparam duty_23__I_0_i27_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mux_666_i9_3_lut (.I0(n155[8]), .I1(PWMLimit[8]), .I2(n256), 
            .I3(GND_net), .O(n3290[8]));   // verilog/motorControl.v(46[16] 48[10])
    defparam mux_666_i9_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 duty_23__I_0_i9_2_lut (.I0(PWMLimit[4]), .I1(duty[4]), .I2(GND_net), 
            .I3(GND_net), .O(n9));   // verilog/motorControl.v(44[10:25])
    defparam duty_23__I_0_i9_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i17_2_lut (.I0(PWMLimit[8]), .I1(duty[8]), .I2(GND_net), 
            .I3(GND_net), .O(n17));   // verilog/motorControl.v(44[10:25])
    defparam duty_23__I_0_i17_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i19_2_lut (.I0(PWMLimit[9]), .I1(duty[9]), .I2(GND_net), 
            .I3(GND_net), .O(n19));   // verilog/motorControl.v(44[10:25])
    defparam duty_23__I_0_i19_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_11_i224_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral [13]), 
            .I2(GND_net), .I3(GND_net), .O(n332_adj_3911));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i224_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 duty_23__I_0_i21_2_lut (.I0(PWMLimit[10]), .I1(duty[10]), .I2(GND_net), 
            .I3(GND_net), .O(n21_adj_3912));   // verilog/motorControl.v(44[10:25])
    defparam duty_23__I_0_i21_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i30828_4_lut (.I0(n21_adj_3912), .I1(n19), .I2(n17), .I3(n9), 
            .O(n37509));
    defparam i30828_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 unary_minus_5_inv_0_i2_1_lut (.I0(IntegralLimit[1]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4332[1]));   // verilog/motorControl.v(39[48:62])
    defparam unary_minus_5_inv_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i30821_4_lut (.I0(n27), .I1(n15), .I2(n13), .I3(n11), .O(n37502));
    defparam i30821_4_lut.LUT_INIT = 16'haaab;
    SB_CARRY add_4138_7 (.CI(n29463), .I0(n8717[4]), .I1(n460), .CO(n29464));
    SB_LUT4 add_4138_6_lut (.I0(GND_net), .I1(n8717[3]), .I2(n387), .I3(n29462), 
            .O(n8699[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4138_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 duty_23__I_0_i30_3_lut (.I0(n12), .I1(duty[17]), .I2(n35), 
            .I3(GND_net), .O(n30));   // verilog/motorControl.v(44[10:25])
    defparam duty_23__I_0_i30_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i31157_4_lut (.I0(n13), .I1(n11), .I2(n9), .I3(n37558), 
            .O(n37839));
    defparam i31157_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 mult_11_i273_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral [13]), 
            .I2(GND_net), .I3(GND_net), .O(n405_adj_3913));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i273_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_4138_6 (.CI(n29462), .I0(n8717[3]), .I1(n387), .CO(n29463));
    SB_LUT4 i31145_4_lut (.I0(n19), .I1(n17), .I2(n15), .I3(n37839), 
            .O(n37827));
    defparam i31145_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i31391_4_lut (.I0(n25_c), .I1(n23), .I2(n21_adj_3912), .I3(n37827), 
            .O(n38073));
    defparam i31391_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i31277_4_lut (.I0(n31), .I1(n29), .I2(n27), .I3(n38073), 
            .O(n37959));
    defparam i31277_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 unary_minus_16_inv_0_i4_1_lut (.I0(PWMLimit[3]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[3]));   // verilog/motorControl.v(47[19:28])
    defparam unary_minus_16_inv_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i31421_4_lut (.I0(n37), .I1(n35), .I2(n33), .I3(n37959), 
            .O(n38103));
    defparam i31421_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i31337_3_lut (.I0(n6), .I1(duty[10]), .I2(n21_adj_3912), .I3(GND_net), 
            .O(n38019));   // verilog/motorControl.v(44[10:25])
    defparam i31337_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i31338_3_lut (.I0(n38019), .I1(duty[11]), .I2(n23), .I3(GND_net), 
            .O(n38020));   // verilog/motorControl.v(44[10:25])
    defparam i31338_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_4121_10 (.CI(n29288), .I0(n8495[7]), .I1(n694), .CO(n29289));
    SB_LUT4 add_4121_9_lut (.I0(GND_net), .I1(n8495[6]), .I2(n621), .I3(n29287), 
            .O(n8482[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4121_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 duty_23__I_0_i24_3_lut (.I0(n16), .I1(duty[22]), .I2(n45), 
            .I3(GND_net), .O(n24_adj_3914));   // verilog/motorControl.v(44[10:25])
    defparam duty_23__I_0_i24_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i30801_4_lut (.I0(n43), .I1(n25_c), .I2(n23), .I3(n37509), 
            .O(n37482));
    defparam i30801_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i31247_4_lut (.I0(n24_adj_3914), .I1(n8), .I2(n45), .I3(n37480), 
            .O(n37929));   // verilog/motorControl.v(44[10:25])
    defparam i31247_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i31062_3_lut (.I0(n38020), .I1(duty[12]), .I2(n25_c), .I3(GND_net), 
            .O(n37744));   // verilog/motorControl.v(44[10:25])
    defparam i31062_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i31275_3_lut (.I0(n4), .I1(duty[13]), .I2(n27), .I3(GND_net), 
            .O(n37957));   // verilog/motorControl.v(44[10:25])
    defparam i31275_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_4138_5_lut (.I0(GND_net), .I1(n8717[2]), .I2(n314), .I3(n29461), 
            .O(n8699[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4138_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4138_5 (.CI(n29461), .I0(n8717[2]), .I1(n314), .CO(n29462));
    SB_LUT4 add_4138_4_lut (.I0(GND_net), .I1(n8717[1]), .I2(n241), .I3(n29460), 
            .O(n8699[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4138_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i31276_3_lut (.I0(n37957), .I1(duty[14]), .I2(n29), .I3(GND_net), 
            .O(n37958));   // verilog/motorControl.v(44[10:25])
    defparam i31276_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i30817_4_lut (.I0(n33), .I1(n31), .I2(n29), .I3(n37502), 
            .O(n37498));
    defparam i30817_4_lut.LUT_INIT = 16'haaab;
    SB_CARRY add_4138_4 (.CI(n29460), .I0(n8717[1]), .I1(n241), .CO(n29461));
    SB_LUT4 i31385_4_lut (.I0(n30), .I1(n10), .I2(n35), .I3(n37494), 
            .O(n38067));   // verilog/motorControl.v(44[10:25])
    defparam i31385_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i31064_3_lut (.I0(n37958), .I1(duty[15]), .I2(n31), .I3(GND_net), 
            .O(n37746));   // verilog/motorControl.v(44[10:25])
    defparam i31064_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i31435_4_lut (.I0(n37746), .I1(n38067), .I2(n35), .I3(n37498), 
            .O(n38117));   // verilog/motorControl.v(44[10:25])
    defparam i31435_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i31436_3_lut (.I0(n38117), .I1(duty[18]), .I2(n37), .I3(GND_net), 
            .O(n38118));   // verilog/motorControl.v(44[10:25])
    defparam i31436_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i31424_3_lut (.I0(n38118), .I1(duty[19]), .I2(n39), .I3(GND_net), 
            .O(n38106));   // verilog/motorControl.v(44[10:25])
    defparam i31424_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_10_i516_2_lut (.I0(\Kp[10] ), .I1(\PID_CONTROLLER.err [12]), 
            .I2(GND_net), .I3(GND_net), .O(n767));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i516_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_4121_9 (.CI(n29287), .I0(n8495[6]), .I1(n621), .CO(n29288));
    SB_LUT4 i30803_4_lut (.I0(n43), .I1(n41), .I2(n39), .I3(n38103), 
            .O(n37484));
    defparam i30803_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i31373_4_lut (.I0(n37744), .I1(n37929), .I2(n45), .I3(n37482), 
            .O(n38055));   // verilog/motorControl.v(44[10:25])
    defparam i31373_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i31070_3_lut (.I0(n38106), .I1(duty[20]), .I2(n41), .I3(GND_net), 
            .O(n37752));   // verilog/motorControl.v(44[10:25])
    defparam i31070_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i31419_4_lut (.I0(n37752), .I1(n38055), .I2(n45), .I3(n37484), 
            .O(n38101));   // verilog/motorControl.v(44[10:25])
    defparam i31419_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i31420_3_lut (.I0(n38101), .I1(PWMLimit[23]), .I2(duty[23]), 
            .I3(GND_net), .O(duty_23__N_3637));   // verilog/motorControl.v(44[10:25])
    defparam i31420_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 mult_11_i359_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral [7]), 
            .I2(GND_net), .I3(GND_net), .O(n533));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i359_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 duty_23__I_0_29_i1_3_lut (.I0(duty_23__N_3613[0]), .I1(PWMLimit[0]), 
            .I2(duty_23__N_3637), .I3(GND_net), .O(duty_23__N_3490[0]));   // verilog/motorControl.v(46[16] 48[10])
    defparam duty_23__I_0_29_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_11_i553_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral [6]), 
            .I2(GND_net), .I3(GND_net), .O(n822));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i553_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i124_2_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err [12]), 
            .I2(GND_net), .I3(GND_net), .O(n183));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i124_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i65_2_lut (.I0(\Kp[1] ), .I1(\PID_CONTROLLER.err [7]), 
            .I2(GND_net), .I3(GND_net), .O(n95));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i65_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i602_2_lut (.I0(\Ki[12] ), .I1(\PID_CONTROLLER.integral [6]), 
            .I2(GND_net), .I3(GND_net), .O(n895));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i602_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_inv_0_i23_1_lut (.I0(IntegralLimit[22]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4332[22]));   // verilog/motorControl.v(39[48:62])
    defparam unary_minus_5_inv_0_i23_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_4138_3_lut (.I0(GND_net), .I1(n8717[0]), .I2(n168), .I3(n29459), 
            .O(n8699[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4138_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4121_8_lut (.I0(GND_net), .I1(n8495[5]), .I2(n548), .I3(n29286), 
            .O(n8482[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4121_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i565_2_lut (.I0(\Kp[11] ), .I1(\PID_CONTROLLER.err [12]), 
            .I2(GND_net), .I3(GND_net), .O(n840_adj_3906));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i565_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_4121_8 (.CI(n29286), .I0(n8495[5]), .I1(n548), .CO(n29287));
    SB_LUT4 mult_10_i18_2_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err [8]), 
            .I2(GND_net), .I3(GND_net), .O(n26));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i18_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i77_2_lut (.I0(\Kp[1] ), .I1(\PID_CONTROLLER.err [13]), 
            .I2(GND_net), .I3(GND_net), .O(n113));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i77_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i31558_1_lut (.I0(duty[23]), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n38238));   // verilog/motorControl.v(37[14] 56[8])
    defparam i31558_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i173_2_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err [12]), 
            .I2(GND_net), .I3(GND_net), .O(n256_adj_3915));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i173_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i30_2_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err [14]), 
            .I2(GND_net), .I3(GND_net), .O(n44));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i30_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_4138_3 (.CI(n29459), .I0(n8717[0]), .I1(n168), .CO(n29460));
    SB_LUT4 add_4138_2_lut (.I0(GND_net), .I1(n26_adj_3916), .I2(n95_adj_3917), 
            .I3(GND_net), .O(n8699[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4138_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_15_i9_2_lut (.I0(duty[4]), .I1(n257[4]), .I2(GND_net), 
            .I3(GND_net), .O(n9_adj_3918));   // verilog/motorControl.v(46[19:35])
    defparam LessThan_15_i9_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_15_i11_2_lut (.I0(duty[5]), .I1(n257[5]), .I2(GND_net), 
            .I3(GND_net), .O(n11_adj_3919));   // verilog/motorControl.v(46[19:35])
    defparam LessThan_15_i11_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_11_i408_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral [7]), 
            .I2(GND_net), .I3(GND_net), .O(n606));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i408_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_15_i13_2_lut (.I0(duty[6]), .I1(n257[6]), .I2(GND_net), 
            .I3(GND_net), .O(n13_adj_3920));   // verilog/motorControl.v(46[19:35])
    defparam LessThan_15_i13_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_15_i15_2_lut (.I0(duty[7]), .I1(n257[7]), .I2(GND_net), 
            .I3(GND_net), .O(n15_adj_3921));   // verilog/motorControl.v(46[19:35])
    defparam LessThan_15_i15_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 unary_minus_5_inv_0_i3_1_lut (.I0(IntegralLimit[2]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4332[2]));   // verilog/motorControl.v(39[48:62])
    defparam unary_minus_5_inv_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 LessThan_15_i21_2_lut (.I0(duty[10]), .I1(n257[10]), .I2(GND_net), 
            .I3(GND_net), .O(n21_adj_3923));   // verilog/motorControl.v(46[19:35])
    defparam LessThan_15_i21_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_15_i19_2_lut (.I0(duty[9]), .I1(n257[9]), .I2(GND_net), 
            .I3(GND_net), .O(n19_adj_3924));   // verilog/motorControl.v(46[19:35])
    defparam LessThan_15_i19_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_4138_2 (.CI(GND_net), .I0(n26_adj_3916), .I1(n95_adj_3917), 
            .CO(n29459));
    SB_LUT4 LessThan_15_i17_2_lut (.I0(duty[8]), .I1(n257[8]), .I2(GND_net), 
            .I3(GND_net), .O(n17_adj_3925));   // verilog/motorControl.v(46[19:35])
    defparam LessThan_15_i17_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY unary_minus_16_add_3_4 (.CI(n28110), .I0(GND_net), .I1(n1[2]), 
            .CO(n28111));
    SB_LUT4 LessThan_15_i23_2_lut (.I0(duty[11]), .I1(n257[11]), .I2(GND_net), 
            .I3(GND_net), .O(n23_adj_3926));   // verilog/motorControl.v(46[19:35])
    defparam LessThan_15_i23_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_10_i265_2_lut (.I0(\Kp[5] ), .I1(\PID_CONTROLLER.err [9]), 
            .I2(GND_net), .I3(GND_net), .O(n393));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i265_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_4137_18_lut (.I0(GND_net), .I1(n8699[15]), .I2(GND_net), 
            .I3(n29458), .O(n8680[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4137_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_5_inv_0_i24_1_lut (.I0(IntegralLimit[23]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4332[23]));   // verilog/motorControl.v(39[48:62])
    defparam unary_minus_5_inv_0_i24_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i296_2_lut (.I0(\Kp[6] ), .I1(\PID_CONTROLLER.err [0]), 
            .I2(GND_net), .I3(GND_net), .O(n439));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i296_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i79_2_lut (.I0(\Kp[1] ), .I1(\PID_CONTROLLER.err [14]), 
            .I2(GND_net), .I3(GND_net), .O(n116));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i79_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_16_add_3_3_lut (.I0(GND_net), .I1(GND_net), .I2(n1[1]), 
            .I3(n28109), .O(n257[1])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4121_7_lut (.I0(GND_net), .I1(n8495[4]), .I2(n475), .I3(n29285), 
            .O(n8482[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4121_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i32_2_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err [15]), 
            .I2(GND_net), .I3(GND_net), .O(n47));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i32_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i345_2_lut (.I0(\Kp[7] ), .I1(\PID_CONTROLLER.err [0]), 
            .I2(GND_net), .I3(GND_net), .O(n512));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i345_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i67_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral [8]), 
            .I2(GND_net), .I3(GND_net), .O(n98));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i67_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i20_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral [9]), 
            .I2(GND_net), .I3(GND_net), .O(n29_adj_3928));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i20_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i394_2_lut (.I0(\Kp[8] ), .I1(\PID_CONTROLLER.err [0]), 
            .I2(GND_net), .I3(GND_net), .O(n585));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i394_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i443_2_lut (.I0(\Kp[9] ), .I1(\PID_CONTROLLER.err [0]), 
            .I2(GND_net), .I3(GND_net), .O(n658));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i443_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i128_2_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err [14]), 
            .I2(GND_net), .I3(GND_net), .O(n189));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i128_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_16_inv_0_i1_1_lut (.I0(PWMLimit[0]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[0]));   // verilog/motorControl.v(47[19:28])
    defparam unary_minus_16_inv_0_i1_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_11_i322_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral [13]), 
            .I2(GND_net), .I3(GND_net), .O(n478_adj_3930));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i322_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_4121_7 (.CI(n29285), .I0(n8495[4]), .I1(n475), .CO(n29286));
    SB_LUT4 mult_10_i492_2_lut (.I0(\Kp[10] ), .I1(\PID_CONTROLLER.err [0]), 
            .I2(GND_net), .I3(GND_net), .O(n731));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i492_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_4121_6_lut (.I0(GND_net), .I1(n8495[3]), .I2(n402), .I3(n29284), 
            .O(n8482[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4121_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i261_2_lut (.I0(\Kp[5] ), .I1(\PID_CONTROLLER.err [7]), 
            .I2(GND_net), .I3(GND_net), .O(n387_adj_3931));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i261_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i126_2_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err [13]), 
            .I2(GND_net), .I3(GND_net), .O(n186));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i126_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_666_i10_3_lut (.I0(n155[9]), .I1(PWMLimit[9]), .I2(n256), 
            .I3(GND_net), .O(n3290[9]));   // verilog/motorControl.v(46[16] 48[10])
    defparam mux_666_i10_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 mult_11_i457_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral [7]), 
            .I2(GND_net), .I3(GND_net), .O(n679));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i457_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_16_inv_0_i5_1_lut (.I0(PWMLimit[4]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[4]));   // verilog/motorControl.v(47[19:28])
    defparam unary_minus_16_inv_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_11_i651_2_lut (.I0(\Ki[13] ), .I1(\PID_CONTROLLER.integral [6]), 
            .I2(GND_net), .I3(GND_net), .O(n968));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i651_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i700_2_lut (.I0(\Ki[14] ), .I1(\PID_CONTROLLER.integral [6]), 
            .I2(GND_net), .I3(GND_net), .O(n1041));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i700_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i57_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral [3]), 
            .I2(GND_net), .I3(GND_net), .O(n83));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i57_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i10_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral [4]), 
            .I2(GND_net), .I3(GND_net), .O(n14));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i10_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_inv_0_i4_1_lut (.I0(IntegralLimit[3]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4332[3]));   // verilog/motorControl.v(39[48:62])
    defparam unary_minus_5_inv_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i177_2_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err [14]), 
            .I2(GND_net), .I3(GND_net), .O(n262));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i177_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i222_2_lut (.I0(\Kp[4] ), .I1(\PID_CONTROLLER.err [12]), 
            .I2(GND_net), .I3(GND_net), .O(n329));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i222_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i749_2_lut (.I0(\Ki[15] ), .I1(\PID_CONTROLLER.integral [6]), 
            .I2(GND_net), .I3(GND_net), .O(n1114_adj_3933));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i749_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i541_2_lut (.I0(\Kp[11] ), .I1(\PID_CONTROLLER.err [0]), 
            .I2(GND_net), .I3(GND_net), .O(n804));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i541_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 duty_23__I_0_29_i24_3_lut (.I0(duty_23__N_3613[23]), .I1(PWMLimit[23]), 
            .I2(duty_23__N_3637), .I3(GND_net), .O(duty_23__N_3490[23]));   // verilog/motorControl.v(46[16] 48[10])
    defparam duty_23__I_0_29_i24_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_29_i23_3_lut (.I0(duty_23__N_3613[22]), .I1(PWMLimit[22]), 
            .I2(duty_23__N_3637), .I3(GND_net), .O(duty_23__N_3490[22]));   // verilog/motorControl.v(46[16] 48[10])
    defparam duty_23__I_0_29_i23_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_29_i22_3_lut (.I0(duty_23__N_3613[21]), .I1(PWMLimit[21]), 
            .I2(duty_23__N_3637), .I3(GND_net), .O(duty_23__N_3490[21]));   // verilog/motorControl.v(46[16] 48[10])
    defparam duty_23__I_0_29_i22_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_10_i310_2_lut (.I0(\Kp[6] ), .I1(\PID_CONTROLLER.err [7]), 
            .I2(GND_net), .I3(GND_net), .O(n460_adj_3934));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i310_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i106_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral [3]), 
            .I2(GND_net), .I3(GND_net), .O(n156));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i106_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i226_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral [14]), 
            .I2(GND_net), .I3(GND_net), .O(n335));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i226_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i359_2_lut (.I0(\Kp[7] ), .I1(\PID_CONTROLLER.err [7]), 
            .I2(GND_net), .I3(GND_net), .O(n533_adj_3935));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i359_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i353_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral [4]), 
            .I2(GND_net), .I3(GND_net), .O(n524));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i353_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 duty_23__I_0_29_i21_3_lut (.I0(duty_23__N_3613[20]), .I1(PWMLimit[20]), 
            .I2(duty_23__N_3637), .I3(GND_net), .O(duty_23__N_3490[20]));   // verilog/motorControl.v(46[16] 48[10])
    defparam duty_23__I_0_29_i21_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_11_i155_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral [3]), 
            .I2(GND_net), .I3(GND_net), .O(n229));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i155_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i590_2_lut (.I0(\Kp[12] ), .I1(\PID_CONTROLLER.err [0]), 
            .I2(GND_net), .I3(GND_net), .O(n877));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i590_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_inv_0_i5_1_lut (.I0(IntegralLimit[4]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4332[4]));   // verilog/motorControl.v(39[48:62])
    defparam unary_minus_5_inv_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 duty_23__I_0_29_i20_3_lut (.I0(duty_23__N_3613[19]), .I1(PWMLimit[19]), 
            .I2(duty_23__N_3637), .I3(GND_net), .O(duty_23__N_3490[19]));   // verilog/motorControl.v(46[16] 48[10])
    defparam duty_23__I_0_29_i20_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_10_i408_2_lut (.I0(\Kp[8] ), .I1(\PID_CONTROLLER.err [7]), 
            .I2(GND_net), .I3(GND_net), .O(n606_adj_3937));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i408_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i226_2_lut (.I0(\Kp[4] ), .I1(\PID_CONTROLLER.err [14]), 
            .I2(GND_net), .I3(GND_net), .O(n335_adj_3938));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i226_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i204_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral [3]), 
            .I2(GND_net), .I3(GND_net), .O(n302));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i204_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i298_2_lut (.I0(\Kp[6] ), .I1(\PID_CONTROLLER.err [1]), 
            .I2(GND_net), .I3(GND_net), .O(n442));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i298_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i639_2_lut (.I0(\Kp[13] ), .I1(\PID_CONTROLLER.err [0]), 
            .I2(GND_net), .I3(GND_net), .O(n950));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i639_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i275_2_lut (.I0(\Kp[5] ), .I1(\PID_CONTROLLER.err [14]), 
            .I2(GND_net), .I3(GND_net), .O(n408));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i275_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 duty_23__I_0_29_i19_3_lut (.I0(duty_23__N_3613[18]), .I1(PWMLimit[18]), 
            .I2(duty_23__N_3637), .I3(GND_net), .O(duty_23__N_3490[18]));   // verilog/motorControl.v(46[16] 48[10])
    defparam duty_23__I_0_29_i19_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_29_i18_3_lut (.I0(duty_23__N_3613[17]), .I1(PWMLimit[17]), 
            .I2(duty_23__N_3637), .I3(GND_net), .O(duty_23__N_3490[17]));   // verilog/motorControl.v(46[16] 48[10])
    defparam duty_23__I_0_29_i18_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_11_i116_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral [8]), 
            .I2(GND_net), .I3(GND_net), .O(n171));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i116_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i275_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral [14]), 
            .I2(GND_net), .I3(GND_net), .O(n408_adj_3939));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i275_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 state_23__I_0_inv_0_i1_1_lut (.I0(setpoint[0]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4333[0]));   // verilog/motorControl.v(38[14:30])
    defparam state_23__I_0_inv_0_i1_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mux_666_i12_3_lut (.I0(n155[11]), .I1(PWMLimit[11]), .I2(n256), 
            .I3(GND_net), .O(n3290[11]));   // verilog/motorControl.v(46[16] 48[10])
    defparam mux_666_i12_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 mult_10_i347_2_lut (.I0(\Kp[7] ), .I1(\PID_CONTROLLER.err [1]), 
            .I2(GND_net), .I3(GND_net), .O(n515));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i347_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 duty_23__I_0_29_i17_3_lut (.I0(duty_23__N_3613[16]), .I1(PWMLimit[16]), 
            .I2(duty_23__N_3637), .I3(GND_net), .O(duty_23__N_3490[16]));   // verilog/motorControl.v(46[16] 48[10])
    defparam duty_23__I_0_29_i17_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_29_i16_3_lut (.I0(duty_23__N_3613[15]), .I1(PWMLimit[15]), 
            .I2(duty_23__N_3637), .I3(GND_net), .O(duty_23__N_3490[15]));   // verilog/motorControl.v(46[16] 48[10])
    defparam duty_23__I_0_29_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 state_23__I_0_inv_0_i2_1_lut (.I0(setpoint[1]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4333[1]));   // verilog/motorControl.v(38[14:30])
    defparam state_23__I_0_inv_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_4137_17_lut (.I0(GND_net), .I1(n8699[14]), .I2(GND_net), 
            .I3(n29457), .O(n8680[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4137_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4121_6 (.CI(n29284), .I0(n8495[3]), .I1(n402), .CO(n29285));
    SB_LUT4 mult_10_i396_2_lut (.I0(\Kp[8] ), .I1(\PID_CONTROLLER.err [1]), 
            .I2(GND_net), .I3(GND_net), .O(n588));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i396_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i402_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral [4]), 
            .I2(GND_net), .I3(GND_net), .O(n597));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i402_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 duty_23__I_0_29_i15_3_lut (.I0(duty_23__N_3613[14]), .I1(PWMLimit[14]), 
            .I2(duty_23__N_3637), .I3(GND_net), .O(duty_23__N_3490[14]));   // verilog/motorControl.v(46[16] 48[10])
    defparam duty_23__I_0_29_i15_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_29_i14_3_lut (.I0(duty_23__N_3613[13]), .I1(PWMLimit[13]), 
            .I2(duty_23__N_3637), .I3(GND_net), .O(duty_23__N_3490[13]));   // verilog/motorControl.v(46[16] 48[10])
    defparam duty_23__I_0_29_i14_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_10_i445_2_lut (.I0(\Kp[9] ), .I1(\PID_CONTROLLER.err [1]), 
            .I2(GND_net), .I3(GND_net), .O(n661));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i445_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 duty_23__I_0_29_i13_3_lut (.I0(duty_23__N_3613[12]), .I1(PWMLimit[12]), 
            .I2(duty_23__N_3637), .I3(GND_net), .O(duty_23__N_3490[12]));   // verilog/motorControl.v(46[16] 48[10])
    defparam duty_23__I_0_29_i13_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_10_i457_2_lut (.I0(\Kp[9] ), .I1(\PID_CONTROLLER.err [7]), 
            .I2(GND_net), .I3(GND_net), .O(n679_adj_3942));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i457_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 state_23__I_0_inv_0_i3_1_lut (.I0(setpoint[2]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4333[2]));   // verilog/motorControl.v(38[14:30])
    defparam state_23__I_0_inv_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mux_666_i20_3_lut (.I0(n155[19]), .I1(PWMLimit[19]), .I2(n256), 
            .I3(GND_net), .O(n3290[19]));   // verilog/motorControl.v(46[16] 48[10])
    defparam mux_666_i20_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 mult_10_i314_2_lut (.I0(\Kp[6] ), .I1(\PID_CONTROLLER.err [9]), 
            .I2(GND_net), .I3(GND_net), .O(n466));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i314_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 duty_23__I_0_29_i12_3_lut (.I0(duty_23__N_3613[11]), .I1(PWMLimit[11]), 
            .I2(duty_23__N_3637), .I3(GND_net), .O(duty_23__N_3490[11]));   // verilog/motorControl.v(46[16] 48[10])
    defparam duty_23__I_0_29_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_10_i506_2_lut (.I0(\Kp[10] ), .I1(\PID_CONTROLLER.err [7]), 
            .I2(GND_net), .I3(GND_net), .O(n752_adj_3944));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i506_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i253_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral [3]), 
            .I2(GND_net), .I3(GND_net), .O(n375));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i253_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_4137_17 (.CI(n29457), .I0(n8699[14]), .I1(GND_net), .CO(n29458));
    SB_LUT4 mult_10_i363_2_lut (.I0(\Kp[7] ), .I1(\PID_CONTROLLER.err [9]), 
            .I2(GND_net), .I3(GND_net), .O(n539));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i363_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i494_2_lut (.I0(\Kp[10] ), .I1(\PID_CONTROLLER.err [1]), 
            .I2(GND_net), .I3(GND_net), .O(n734));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i494_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 duty_23__I_0_29_i11_3_lut (.I0(duty_23__N_3613[10]), .I1(PWMLimit[10]), 
            .I2(duty_23__N_3637), .I3(GND_net), .O(duty_23__N_3490[10]));   // verilog/motorControl.v(46[16] 48[10])
    defparam duty_23__I_0_29_i11_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_29_i10_3_lut (.I0(duty_23__N_3613[9]), .I1(PWMLimit[9]), 
            .I2(duty_23__N_3637), .I3(GND_net), .O(duty_23__N_3490[9]));   // verilog/motorControl.v(46[16] 48[10])
    defparam duty_23__I_0_29_i10_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_10_i555_2_lut (.I0(\Kp[11] ), .I1(\PID_CONTROLLER.err [7]), 
            .I2(GND_net), .I3(GND_net), .O(n825_adj_3945));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i555_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 duty_23__I_0_29_i9_3_lut (.I0(duty_23__N_3613[8]), .I1(PWMLimit[8]), 
            .I2(duty_23__N_3637), .I3(GND_net), .O(duty_23__N_3490[8]));   // verilog/motorControl.v(46[16] 48[10])
    defparam duty_23__I_0_29_i9_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_11_i302_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral [3]), 
            .I2(GND_net), .I3(GND_net), .O(n448));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i302_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i324_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral [14]), 
            .I2(GND_net), .I3(GND_net), .O(n481));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i324_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 duty_23__I_0_29_i8_3_lut (.I0(duty_23__N_3613[7]), .I1(PWMLimit[7]), 
            .I2(duty_23__N_3637), .I3(GND_net), .O(duty_23__N_3490[7]));   // verilog/motorControl.v(46[16] 48[10])
    defparam duty_23__I_0_29_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_29_i7_3_lut (.I0(duty_23__N_3613[6]), .I1(PWMLimit[6]), 
            .I2(duty_23__N_3637), .I3(GND_net), .O(duty_23__N_3490[6]));   // verilog/motorControl.v(46[16] 48[10])
    defparam duty_23__I_0_29_i7_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_666_i13_3_lut (.I0(n155[12]), .I1(PWMLimit[12]), .I2(n256), 
            .I3(GND_net), .O(n3290[12]));   // verilog/motorControl.v(46[16] 48[10])
    defparam mux_666_i13_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 duty_23__I_0_29_i6_3_lut (.I0(duty_23__N_3613[5]), .I1(PWMLimit[5]), 
            .I2(duty_23__N_3637), .I3(GND_net), .O(duty_23__N_3490[5]));   // verilog/motorControl.v(46[16] 48[10])
    defparam duty_23__I_0_29_i6_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_29_i5_3_lut (.I0(duty_23__N_3613[4]), .I1(PWMLimit[4]), 
            .I2(duty_23__N_3637), .I3(GND_net), .O(duty_23__N_3490[4]));   // verilog/motorControl.v(46[16] 48[10])
    defparam duty_23__I_0_29_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_29_i4_3_lut (.I0(duty_23__N_3613[3]), .I1(PWMLimit[3]), 
            .I2(duty_23__N_3637), .I3(GND_net), .O(duty_23__N_3490[3]));   // verilog/motorControl.v(46[16] 48[10])
    defparam duty_23__I_0_29_i4_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_29_i3_3_lut (.I0(duty_23__N_3613[2]), .I1(PWMLimit[2]), 
            .I2(duty_23__N_3637), .I3(GND_net), .O(duty_23__N_3490[2]));   // verilog/motorControl.v(46[16] 48[10])
    defparam duty_23__I_0_29_i3_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_10_i604_2_lut (.I0(\Kp[12] ), .I1(\PID_CONTROLLER.err [7]), 
            .I2(GND_net), .I3(GND_net), .O(n898_adj_3946));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i604_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i351_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral [3]), 
            .I2(GND_net), .I3(GND_net), .O(n521));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i351_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i653_2_lut (.I0(\Kp[13] ), .I1(\PID_CONTROLLER.err [7]), 
            .I2(GND_net), .I3(GND_net), .O(n971_adj_3947));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i653_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i400_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral [3]), 
            .I2(GND_net), .I3(GND_net), .O(n594));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i400_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i688_2_lut (.I0(\Kp[14] ), .I1(\PID_CONTROLLER.err [0]), 
            .I2(GND_net), .I3(GND_net), .O(n1023));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i688_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i324_2_lut (.I0(\Kp[6] ), .I1(\PID_CONTROLLER.err [14]), 
            .I2(GND_net), .I3(GND_net), .O(n481_adj_3948));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i324_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 state_23__I_0_inv_0_i4_1_lut (.I0(setpoint[3]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4333[3]));   // verilog/motorControl.v(38[14:30])
    defparam state_23__I_0_inv_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_11_i373_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral [14]), 
            .I2(GND_net), .I3(GND_net), .O(n554));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i373_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i175_2_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err [13]), 
            .I2(GND_net), .I3(GND_net), .O(n259));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i175_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i165_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral [8]), 
            .I2(GND_net), .I3(GND_net), .O(n244));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i165_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_666_i14_3_lut (.I0(n155[13]), .I1(PWMLimit[13]), .I2(n256), 
            .I3(GND_net), .O(n3290[13]));   // verilog/motorControl.v(46[16] 48[10])
    defparam mux_666_i14_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 unary_minus_16_inv_0_i7_1_lut (.I0(PWMLimit[6]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[6]));   // verilog/motorControl.v(47[19:28])
    defparam unary_minus_16_inv_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY unary_minus_16_add_3_3 (.CI(n28109), .I0(GND_net), .I1(n1[1]), 
            .CO(n28110));
    SB_LUT4 mult_10_i271_2_lut (.I0(\Kp[5] ), .I1(\PID_CONTROLLER.err [12]), 
            .I2(GND_net), .I3(GND_net), .O(n402));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i271_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i737_2_lut (.I0(\Kp[15] ), .I1(\PID_CONTROLLER.err [0]), 
            .I2(GND_net), .I3(GND_net), .O(n1096));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i737_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i320_2_lut (.I0(\Kp[6] ), .I1(\PID_CONTROLLER.err [12]), 
            .I2(GND_net), .I3(GND_net), .O(n475));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i320_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_16_inv_0_i2_1_lut (.I0(PWMLimit[1]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[1]));   // verilog/motorControl.v(47[19:28])
    defparam unary_minus_16_inv_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i702_2_lut (.I0(\Kp[14] ), .I1(\PID_CONTROLLER.err [7]), 
            .I2(GND_net), .I3(GND_net), .O(n1044_adj_3951));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i702_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i373_2_lut (.I0(\Kp[7] ), .I1(\PID_CONTROLLER.err [14]), 
            .I2(GND_net), .I3(GND_net), .O(n554_adj_3952));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i373_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 state_23__I_0_inv_0_i5_1_lut (.I0(setpoint[4]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4333[4]));   // verilog/motorControl.v(38[14:30])
    defparam state_23__I_0_inv_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_11_i65_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral [7]), 
            .I2(GND_net), .I3(GND_net), .O(n95_adj_3917));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i65_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i18_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral [8]), 
            .I2(GND_net), .I3(GND_net), .O(n26_adj_3916));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i18_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i369_2_lut (.I0(\Kp[7] ), .I1(\PID_CONTROLLER.err [12]), 
            .I2(GND_net), .I3(GND_net), .O(n548));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i369_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i114_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral [7]), 
            .I2(GND_net), .I3(GND_net), .O(n168));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i114_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i163_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral [7]), 
            .I2(GND_net), .I3(GND_net), .O(n241));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i163_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i214_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral [8]), 
            .I2(GND_net), .I3(GND_net), .O(n317));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i214_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 state_23__I_0_inv_0_i6_1_lut (.I0(setpoint[5]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4333[5]));   // verilog/motorControl.v(38[14:30])
    defparam state_23__I_0_inv_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_11_i212_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral [7]), 
            .I2(GND_net), .I3(GND_net), .O(n314));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i212_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i751_2_lut (.I0(\Kp[15] ), .I1(\PID_CONTROLLER.err [7]), 
            .I2(GND_net), .I3(GND_net), .O(n1117_adj_3955));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i751_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_4137_16_lut (.I0(GND_net), .I1(n8699[13]), .I2(n1114_adj_3933), 
            .I3(n29456), .O(n8680[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4137_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4137_16 (.CI(n29456), .I0(n8699[13]), .I1(n1114_adj_3933), 
            .CO(n29457));
    SB_LUT4 mult_10_i67_2_lut (.I0(\Kp[1] ), .I1(\PID_CONTROLLER.err [8]), 
            .I2(GND_net), .I3(GND_net), .O(n98_adj_3956));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i67_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i20_2_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err [9]), 
            .I2(GND_net), .I3(GND_net), .O(n29_adj_3957));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i20_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 state_23__I_0_inv_0_i7_1_lut (.I0(setpoint[6]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4333[6]));   // verilog/motorControl.v(38[14:30])
    defparam state_23__I_0_inv_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_11_i449_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral [3]), 
            .I2(GND_net), .I3(GND_net), .O(n667));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i449_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_4121_5_lut (.I0(GND_net), .I1(n8495[2]), .I2(n329), .I3(n29283), 
            .O(n8482[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4121_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i422_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral [14]), 
            .I2(GND_net), .I3(GND_net), .O(n627));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i422_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i418_2_lut (.I0(\Kp[8] ), .I1(\PID_CONTROLLER.err [12]), 
            .I2(GND_net), .I3(GND_net), .O(n621));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i418_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i224_2_lut (.I0(\Kp[4] ), .I1(\PID_CONTROLLER.err [13]), 
            .I2(GND_net), .I3(GND_net), .O(n332));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i224_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_4137_15_lut (.I0(GND_net), .I1(n8699[12]), .I2(n1041), 
            .I3(n29455), .O(n8680[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4137_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4137_15 (.CI(n29455), .I0(n8699[12]), .I1(n1041), .CO(n29456));
    SB_LUT4 add_4137_14_lut (.I0(GND_net), .I1(n8699[11]), .I2(n968), 
            .I3(n29454), .O(n8680[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4137_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i116_2_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err [8]), 
            .I2(GND_net), .I3(GND_net), .O(n171_adj_3959));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i116_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i165_2_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err [8]), 
            .I2(GND_net), .I3(GND_net), .O(n244_adj_3960));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i165_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i498_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral [3]), 
            .I2(GND_net), .I3(GND_net), .O(n740));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i498_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i471_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral [14]), 
            .I2(GND_net), .I3(GND_net), .O(n700));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i471_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_4137_14 (.CI(n29454), .I0(n8699[11]), .I1(n968), .CO(n29455));
    SB_CARRY add_4121_5 (.CI(n29283), .I0(n8495[2]), .I1(n329), .CO(n29284));
    SB_LUT4 mult_10_i214_2_lut (.I0(\Kp[4] ), .I1(\PID_CONTROLLER.err [8]), 
            .I2(GND_net), .I3(GND_net), .O(n317_adj_3961));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i214_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_16_add_3_2_lut (.I0(n25), .I1(GND_net), .I2(n1[0]), 
            .I3(VCC_net), .O(n37256)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_2_lut.LUT_INIT = 16'h8228;
    SB_LUT4 mult_10_i422_2_lut (.I0(\Kp[8] ), .I1(\PID_CONTROLLER.err [14]), 
            .I2(GND_net), .I3(GND_net), .O(n627_adj_3963));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i422_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i547_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral [3]), 
            .I2(GND_net), .I3(GND_net), .O(n813));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i547_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i263_2_lut (.I0(\Kp[5] ), .I1(\PID_CONTROLLER.err [8]), 
            .I2(GND_net), .I3(GND_net), .O(n390));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i263_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 state_23__I_0_inv_0_i8_1_lut (.I0(setpoint[7]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4333[7]));   // verilog/motorControl.v(38[14:30])
    defparam state_23__I_0_inv_0_i8_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_11_i596_2_lut (.I0(\Ki[12] ), .I1(\PID_CONTROLLER.integral [3]), 
            .I2(GND_net), .I3(GND_net), .O(n886));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i596_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i81_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral [15]), 
            .I2(GND_net), .I3(GND_net), .O(n119));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i81_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i34_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral [16]), 
            .I2(GND_net), .I3(GND_net), .O(n50));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i34_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i263_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral [8]), 
            .I2(GND_net), .I3(GND_net), .O(n390_adj_3964));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i263_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i471_2_lut (.I0(\Kp[9] ), .I1(\PID_CONTROLLER.err [14]), 
            .I2(GND_net), .I3(GND_net), .O(n700_adj_3965));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i471_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i371_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral [13]), 
            .I2(GND_net), .I3(GND_net), .O(n551_adj_3966));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i371_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i420_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral [13]), 
            .I2(GND_net), .I3(GND_net), .O(n624_adj_3967));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i420_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_16_inv_0_i8_1_lut (.I0(PWMLimit[7]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[7]));   // verilog/motorControl.v(47[19:28])
    defparam unary_minus_16_inv_0_i8_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i114_2_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err [7]), 
            .I2(GND_net), .I3(GND_net), .O(n168_adj_3969));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i114_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i81_2_lut (.I0(\Kp[1] ), .I1(\PID_CONTROLLER.err [15]), 
            .I2(GND_net), .I3(GND_net), .O(n119_adj_3970));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i81_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY unary_minus_16_add_3_2 (.CI(VCC_net), .I0(GND_net), .I1(n1[0]), 
            .CO(n28109));
    SB_LUT4 unary_minus_5_add_3_25_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4332[23]), 
            .I3(n28108), .O(\PID_CONTROLLER.integral_23__N_3589 [23])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i469_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral [13]), 
            .I2(GND_net), .I3(GND_net), .O(n697_adj_3971));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i469_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i34_2_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err [16]), 
            .I2(GND_net), .I3(GND_net), .O(n50_adj_3972));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i34_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 state_23__I_0_inv_0_i9_1_lut (.I0(setpoint[8]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4333[8]));   // verilog/motorControl.v(38[14:30])
    defparam state_23__I_0_inv_0_i9_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i543_2_lut (.I0(\Kp[11] ), .I1(\PID_CONTROLLER.err [1]), 
            .I2(GND_net), .I3(GND_net), .O(n807));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i543_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i518_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral [13]), 
            .I2(GND_net), .I3(GND_net), .O(n770_adj_3974));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i518_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_666_i11_3_lut (.I0(n155[10]), .I1(PWMLimit[10]), .I2(n256), 
            .I3(GND_net), .O(n3290[10]));   // verilog/motorControl.v(46[16] 48[10])
    defparam mux_666_i11_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 mult_10_i163_2_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err [7]), 
            .I2(GND_net), .I3(GND_net), .O(n241_adj_3975));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i163_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i79_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral [14]), 
            .I2(GND_net), .I3(GND_net), .O(n116_adj_3976));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i79_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i32_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral [15]), 
            .I2(GND_net), .I3(GND_net), .O(n47_adj_3977));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i32_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i412_2_lut (.I0(\Kp[8] ), .I1(\PID_CONTROLLER.err [9]), 
            .I2(GND_net), .I3(GND_net), .O(n612));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i412_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i212_2_lut (.I0(\Kp[4] ), .I1(\PID_CONTROLLER.err [7]), 
            .I2(GND_net), .I3(GND_net), .O(n314_adj_3978));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i212_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i592_2_lut (.I0(\Kp[12] ), .I1(\PID_CONTROLLER.err [1]), 
            .I2(GND_net), .I3(GND_net), .O(n880));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i592_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i641_2_lut (.I0(\Kp[13] ), .I1(\PID_CONTROLLER.err [1]), 
            .I2(GND_net), .I3(GND_net), .O(n953));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i641_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i690_2_lut (.I0(\Kp[14] ), .I1(\PID_CONTROLLER.err [1]), 
            .I2(GND_net), .I3(GND_net), .O(n1026));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i690_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i739_2_lut (.I0(\Kp[15] ), .I1(\PID_CONTROLLER.err [1]), 
            .I2(GND_net), .I3(GND_net), .O(n1099));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i739_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i312_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral [8]), 
            .I2(GND_net), .I3(GND_net), .O(n463));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i312_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i130_2_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err [15]), 
            .I2(GND_net), .I3(GND_net), .O(n192_adj_3979));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i130_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_16_inv_0_i9_1_lut (.I0(PWMLimit[8]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[8]));   // verilog/motorControl.v(47[19:28])
    defparam unary_minus_16_inv_0_i9_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i461_2_lut (.I0(\Kp[9] ), .I1(\PID_CONTROLLER.err [9]), 
            .I2(GND_net), .I3(GND_net), .O(n685));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i461_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 state_23__I_0_inv_0_i10_1_lut (.I0(setpoint[9]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4333[9]));   // verilog/motorControl.v(38[14:30])
    defparam state_23__I_0_inv_0_i10_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_5_inv_0_i16_1_lut (.I0(IntegralLimit[15]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4332[15]));   // verilog/motorControl.v(39[48:62])
    defparam unary_minus_5_inv_0_i16_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_11_i506_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral [7]), 
            .I2(GND_net), .I3(GND_net), .O(n752));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i506_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_4121_4_lut (.I0(GND_net), .I1(n8495[1]), .I2(n256_adj_3915), 
            .I3(n29282), .O(n8482[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4121_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i273_2_lut (.I0(\Kp[5] ), .I1(\PID_CONTROLLER.err [13]), 
            .I2(GND_net), .I3(GND_net), .O(n405));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i273_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_add_3_24_lut (.I0(\PID_CONTROLLER.integral [22]), 
            .I1(GND_net), .I2(n1_adj_4332[22]), .I3(n28107), .O(n45_adj_3983)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_24_lut.LUT_INIT = 16'h6996;
    SB_CARRY unary_minus_5_add_3_24 (.CI(n28107), .I0(GND_net), .I1(n1_adj_4332[22]), 
            .CO(n28108));
    SB_CARRY add_4121_4 (.CI(n29282), .I0(n8495[1]), .I1(n256_adj_3915), 
            .CO(n29283));
    SB_LUT4 add_4137_13_lut (.I0(GND_net), .I1(n8699[10]), .I2(n895), 
            .I3(n29453), .O(n8680[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4137_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i179_2_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err [15]), 
            .I2(GND_net), .I3(GND_net), .O(n265));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i179_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i555_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral [7]), 
            .I2(GND_net), .I3(GND_net), .O(n825));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i555_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i228_2_lut (.I0(\Kp[4] ), .I1(\PID_CONTROLLER.err [15]), 
            .I2(GND_net), .I3(GND_net), .O(n338));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i228_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i322_2_lut (.I0(\Kp[6] ), .I1(\PID_CONTROLLER.err [13]), 
            .I2(GND_net), .I3(GND_net), .O(n478));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i322_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 state_23__I_0_inv_0_i11_1_lut (.I0(setpoint[10]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4333[10]));   // verilog/motorControl.v(38[14:30])
    defparam state_23__I_0_inv_0_i11_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_4121_3_lut (.I0(GND_net), .I1(n8495[0]), .I2(n183), .I3(n29281), 
            .O(n8482[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4121_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i361_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral [8]), 
            .I2(GND_net), .I3(GND_net), .O(n536));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i361_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_4137_13 (.CI(n29453), .I0(n8699[10]), .I1(n895), .CO(n29454));
    SB_CARRY add_4121_3 (.CI(n29281), .I0(n8495[0]), .I1(n183), .CO(n29282));
    SB_LUT4 add_4137_12_lut (.I0(GND_net), .I1(n8699[9]), .I2(n822), .I3(n29452), 
            .O(n8680[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4137_12_lut.LUT_INIT = 16'hC33C;
    SB_DFF result_i0 (.Q(duty[0]), .C(clk32MHz), .D(duty_23__N_3490[0]));   // verilog/motorControl.v(37[14] 56[8])
    SB_LUT4 mult_11_i451_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral [4]), 
            .I2(GND_net), .I3(GND_net), .O(n670));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i451_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_666_i21_3_lut (.I0(n155[20]), .I1(PWMLimit[20]), .I2(n256), 
            .I3(GND_net), .O(n3290[20]));   // verilog/motorControl.v(46[16] 48[10])
    defparam mux_666_i21_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 mult_10_i277_2_lut (.I0(\Kp[5] ), .I1(\PID_CONTROLLER.err [15]), 
            .I2(GND_net), .I3(GND_net), .O(n411));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i277_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_16_inv_0_i10_1_lut (.I0(PWMLimit[9]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[9]));   // verilog/motorControl.v(47[19:28])
    defparam unary_minus_16_inv_0_i10_1_lut.LUT_INIT = 16'h5555;
    SB_DFF \PID_CONTROLLER.err_i0  (.Q(\PID_CONTROLLER.err [0]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_23__N_3514 [0]));   // verilog/motorControl.v(37[14] 56[8])
    SB_LUT4 mult_10_i510_2_lut (.I0(\Kp[10] ), .I1(\PID_CONTROLLER.err [9]), 
            .I2(GND_net), .I3(GND_net), .O(n758));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i510_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i410_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral [8]), 
            .I2(GND_net), .I3(GND_net), .O(n609));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i410_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 state_23__I_0_inv_0_i12_1_lut (.I0(setpoint[11]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4333[11]));   // verilog/motorControl.v(38[14:30])
    defparam state_23__I_0_inv_0_i12_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_5_inv_0_i17_1_lut (.I0(IntegralLimit[16]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4332[16]));   // verilog/motorControl.v(39[48:62])
    defparam unary_minus_5_inv_0_i17_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_4121_2_lut (.I0(GND_net), .I1(n41_adj_3989), .I2(n110), 
            .I3(GND_net), .O(n8482[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4121_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4121_2 (.CI(GND_net), .I0(n41_adj_3989), .I1(n110), .CO(n29281));
    SB_CARRY add_4137_12 (.CI(n29452), .I0(n8699[9]), .I1(n822), .CO(n29453));
    SB_LUT4 add_4137_11_lut (.I0(GND_net), .I1(n8699[8]), .I2(n749), .I3(n29451), 
            .O(n8680[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4137_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4120_13_lut (.I0(GND_net), .I1(n8482[10]), .I2(n910), 
            .I3(n29280), .O(n8468[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4120_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i459_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral [8]), 
            .I2(GND_net), .I3(GND_net), .O(n682));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i459_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i55_2_lut (.I0(\Kp[1] ), .I1(\PID_CONTROLLER.err [2]), 
            .I2(GND_net), .I3(GND_net), .O(n80));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i55_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i8_2_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err [3]), 
            .I2(GND_net), .I3(GND_net), .O(n11_adj_3990));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i8_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i326_2_lut (.I0(\Kp[6] ), .I1(\PID_CONTROLLER.err [15]), 
            .I2(GND_net), .I3(GND_net), .O(n484));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i326_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i104_2_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err [2]), 
            .I2(GND_net), .I3(GND_net), .O(n153));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i104_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i508_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral [8]), 
            .I2(GND_net), .I3(GND_net), .O(n755));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i508_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i500_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral [4]), 
            .I2(GND_net), .I3(GND_net), .O(n743));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i500_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_4137_11 (.CI(n29451), .I0(n8699[8]), .I1(n749), .CO(n29452));
    SB_LUT4 mult_10_i375_2_lut (.I0(\Kp[7] ), .I1(\PID_CONTROLLER.err [15]), 
            .I2(GND_net), .I3(GND_net), .O(n557));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i375_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i424_2_lut (.I0(\Kp[8] ), .I1(\PID_CONTROLLER.err [15]), 
            .I2(GND_net), .I3(GND_net), .O(n630));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i424_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_4137_10_lut (.I0(GND_net), .I1(n8699[7]), .I2(n676), .I3(n29450), 
            .O(n8680[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4137_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4120_12_lut (.I0(GND_net), .I1(n8482[9]), .I2(n837), .I3(n29279), 
            .O(n8468[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4120_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4120_12 (.CI(n29279), .I0(n8482[9]), .I1(n837), .CO(n29280));
    SB_LUT4 mux_666_i22_3_lut (.I0(n155[21]), .I1(PWMLimit[21]), .I2(n256), 
            .I3(GND_net), .O(n3290[21]));   // verilog/motorControl.v(46[16] 48[10])
    defparam mux_666_i22_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 add_4120_11_lut (.I0(GND_net), .I1(n8482[8]), .I2(n764), .I3(n29278), 
            .O(n8468[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4120_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4120_11 (.CI(n29278), .I0(n8482[8]), .I1(n764), .CO(n29279));
    SB_LUT4 add_4120_10_lut (.I0(GND_net), .I1(n8482[7]), .I2(n691), .I3(n29277), 
            .O(n8468[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4120_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i153_2_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err [2]), 
            .I2(GND_net), .I3(GND_net), .O(n226));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i153_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 state_23__I_0_inv_0_i13_1_lut (.I0(setpoint[12]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4333[12]));   // verilog/motorControl.v(38[14:30])
    defparam state_23__I_0_inv_0_i13_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_4120_10 (.CI(n29277), .I0(n8482[7]), .I1(n691), .CO(n29278));
    SB_CARRY add_4137_10 (.CI(n29450), .I0(n8699[7]), .I1(n676), .CO(n29451));
    SB_LUT4 add_4137_9_lut (.I0(GND_net), .I1(n8699[6]), .I2(n603), .I3(n29449), 
            .O(n8680[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4137_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4137_9 (.CI(n29449), .I0(n8699[6]), .I1(n603), .CO(n29450));
    SB_LUT4 add_4137_8_lut (.I0(GND_net), .I1(n8699[5]), .I2(n530), .I3(n29448), 
            .O(n8680[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4137_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i83_2_lut (.I0(\Kp[1] ), .I1(\PID_CONTROLLER.err [16]), 
            .I2(GND_net), .I3(GND_net), .O(n122));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i83_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i36_2_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err [17]), 
            .I2(GND_net), .I3(GND_net), .O(n53));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i36_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_4137_8 (.CI(n29448), .I0(n8699[5]), .I1(n530), .CO(n29449));
    SB_LUT4 add_4137_7_lut (.I0(GND_net), .I1(n8699[4]), .I2(n457), .I3(n29447), 
            .O(n8680[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4137_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4120_9_lut (.I0(GND_net), .I1(n8482[6]), .I2(n618), .I3(n29276), 
            .O(n8468[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4120_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i557_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral [8]), 
            .I2(GND_net), .I3(GND_net), .O(n828));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i557_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_4137_7 (.CI(n29447), .I0(n8699[4]), .I1(n457), .CO(n29448));
    SB_LUT4 add_4137_6_lut (.I0(GND_net), .I1(n8699[3]), .I2(n384), .I3(n29446), 
            .O(n8680[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4137_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i202_2_lut (.I0(\Kp[4] ), .I1(\PID_CONTROLLER.err [2]), 
            .I2(GND_net), .I3(GND_net), .O(n299));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i202_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i132_2_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err [16]), 
            .I2(GND_net), .I3(GND_net), .O(n195_adj_3992));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i132_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i606_2_lut (.I0(\Ki[12] ), .I1(\PID_CONTROLLER.integral [8]), 
            .I2(GND_net), .I3(GND_net), .O(n901));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i606_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_4137_6 (.CI(n29446), .I0(n8699[3]), .I1(n384), .CO(n29447));
    SB_LUT4 add_4137_5_lut (.I0(GND_net), .I1(n8699[2]), .I2(n311), .I3(n29445), 
            .O(n8680[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4137_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 state_23__I_0_inv_0_i14_1_lut (.I0(setpoint[13]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4333[13]));   // verilog/motorControl.v(38[14:30])
    defparam state_23__I_0_inv_0_i14_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_4120_9 (.CI(n29276), .I0(n8482[6]), .I1(n618), .CO(n29277));
    SB_LUT4 mult_11_i128_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral [14]), 
            .I2(GND_net), .I3(GND_net), .O(n189_adj_3994));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i128_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_4137_5 (.CI(n29445), .I0(n8699[2]), .I1(n311), .CO(n29446));
    SB_LUT4 add_4120_8_lut (.I0(GND_net), .I1(n8482[5]), .I2(n545), .I3(n29275), 
            .O(n8468[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4120_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_16_inv_0_i11_1_lut (.I0(PWMLimit[10]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[10]));   // verilog/motorControl.v(47[19:28])
    defparam unary_minus_16_inv_0_i11_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 duty_23__I_0_29_i2_3_lut (.I0(duty_23__N_3613[1]), .I1(PWMLimit[1]), 
            .I2(duty_23__N_3637), .I3(GND_net), .O(duty_23__N_3490[1]));   // verilog/motorControl.v(46[16] 48[10])
    defparam duty_23__I_0_29_i2_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_11_i604_2_lut (.I0(\Ki[12] ), .I1(\PID_CONTROLLER.integral [7]), 
            .I2(GND_net), .I3(GND_net), .O(n898));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i604_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i251_2_lut (.I0(\Kp[5] ), .I1(\PID_CONTROLLER.err [2]), 
            .I2(GND_net), .I3(GND_net), .O(n372));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i251_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i181_2_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err [16]), 
            .I2(GND_net), .I3(GND_net), .O(n268));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i181_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i559_2_lut (.I0(\Kp[11] ), .I1(\PID_CONTROLLER.err [9]), 
            .I2(GND_net), .I3(GND_net), .O(n831));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i559_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_4137_4_lut (.I0(GND_net), .I1(n8699[1]), .I2(n238), .I3(n29444), 
            .O(n8680[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4137_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4120_8 (.CI(n29275), .I0(n8482[5]), .I1(n545), .CO(n29276));
    SB_LUT4 mult_11_i549_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral [4]), 
            .I2(GND_net), .I3(GND_net), .O(n816));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i549_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_inv_0_i18_1_lut (.I0(IntegralLimit[17]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4332[17]));   // verilog/motorControl.v(39[48:62])
    defparam unary_minus_5_inv_0_i18_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_11_i598_2_lut (.I0(\Ki[12] ), .I1(\PID_CONTROLLER.integral [4]), 
            .I2(GND_net), .I3(GND_net), .O(n889));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i598_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_666_i23_3_lut (.I0(n155[22]), .I1(PWMLimit[22]), .I2(n256), 
            .I3(GND_net), .O(n3290[22]));   // verilog/motorControl.v(46[16] 48[10])
    defparam mux_666_i23_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 unary_minus_5_add_3_23_lut (.I0(\PID_CONTROLLER.integral [21]), 
            .I1(GND_net), .I2(n1_adj_4332[21]), .I3(n28106), .O(n43_adj_3997)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_23_lut.LUT_INIT = 16'h6996;
    SB_CARRY add_4137_4 (.CI(n29444), .I0(n8699[1]), .I1(n238), .CO(n29445));
    SB_LUT4 state_23__I_0_inv_0_i15_1_lut (.I0(setpoint[14]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4333[14]));   // verilog/motorControl.v(38[14:30])
    defparam state_23__I_0_inv_0_i15_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i608_2_lut (.I0(\Kp[12] ), .I1(\PID_CONTROLLER.err [9]), 
            .I2(GND_net), .I3(GND_net), .O(n904));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i608_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_4137_3_lut (.I0(GND_net), .I1(n8699[0]), .I2(n165), .I3(n29443), 
            .O(n8680[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4137_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i647_2_lut (.I0(\Ki[13] ), .I1(\PID_CONTROLLER.integral [4]), 
            .I2(GND_net), .I3(GND_net), .O(n962));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i647_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_4137_3 (.CI(n29443), .I0(n8699[0]), .I1(n165), .CO(n29444));
    SB_LUT4 add_4137_2_lut (.I0(GND_net), .I1(n23_adj_4000), .I2(n92), 
            .I3(GND_net), .O(n8680[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4137_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_5_inv_0_i19_1_lut (.I0(IntegralLimit[18]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4332[18]));   // verilog/motorControl.v(39[48:62])
    defparam unary_minus_5_inv_0_i19_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_4120_7_lut (.I0(GND_net), .I1(n8482[4]), .I2(n472), .I3(n29274), 
            .O(n8468[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4120_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4137_2 (.CI(GND_net), .I0(n23_adj_4000), .I1(n92), .CO(n29443));
    SB_LUT4 add_4136_19_lut (.I0(GND_net), .I1(n8680[16]), .I2(GND_net), 
            .I3(n29442), .O(n8660[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4136_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 state_23__I_0_inv_0_i16_1_lut (.I0(setpoint[15]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4333[15]));   // verilog/motorControl.v(38[14:30])
    defparam state_23__I_0_inv_0_i16_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_4120_7 (.CI(n29274), .I0(n8482[4]), .I1(n472), .CO(n29275));
    SB_LUT4 add_4136_18_lut (.I0(GND_net), .I1(n8680[15]), .I2(GND_net), 
            .I3(n29441), .O(n8660[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4136_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4136_18 (.CI(n29441), .I0(n8680[15]), .I1(GND_net), .CO(n29442));
    SB_LUT4 add_4136_17_lut (.I0(GND_net), .I1(n8680[14]), .I2(GND_net), 
            .I3(n29440), .O(n8660[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4136_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4120_6_lut (.I0(GND_net), .I1(n8482[3]), .I2(n399), .I3(n29273), 
            .O(n8468[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4120_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4120_6 (.CI(n29273), .I0(n8482[3]), .I1(n399), .CO(n29274));
    SB_LUT4 add_4120_5_lut (.I0(GND_net), .I1(n8482[2]), .I2(n326), .I3(n29272), 
            .O(n8468[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4120_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4120_5 (.CI(n29272), .I0(n8482[2]), .I1(n326), .CO(n29273));
    SB_LUT4 add_4120_4_lut (.I0(GND_net), .I1(n8482[1]), .I2(n253), .I3(n29271), 
            .O(n8468[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4120_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4120_4 (.CI(n29271), .I0(n8482[1]), .I1(n253), .CO(n29272));
    SB_LUT4 add_4120_3_lut (.I0(GND_net), .I1(n8482[0]), .I2(n180), .I3(n29270), 
            .O(n8468[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4120_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4136_17 (.CI(n29440), .I0(n8680[14]), .I1(GND_net), .CO(n29441));
    SB_CARRY unary_minus_5_add_3_23 (.CI(n28106), .I0(GND_net), .I1(n1_adj_4332[21]), 
            .CO(n28107));
    SB_LUT4 mult_11_i696_2_lut (.I0(\Ki[14] ), .I1(\PID_CONTROLLER.integral [4]), 
            .I2(GND_net), .I3(GND_net), .O(n1035));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i696_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_4136_16_lut (.I0(GND_net), .I1(n8680[13]), .I2(n1111), 
            .I3(n29439), .O(n8660[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4136_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i657_2_lut (.I0(\Kp[13] ), .I1(\PID_CONTROLLER.err [9]), 
            .I2(GND_net), .I3(GND_net), .O(n977));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i657_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i31413_4_lut (.I0(n37_adj_4002), .I1(n35_adj_4003), .I2(n33_adj_4004), 
            .I3(n37935), .O(n38095));
    defparam i31413_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 mult_10_i706_2_lut (.I0(\Kp[14] ), .I1(\PID_CONTROLLER.err [9]), 
            .I2(GND_net), .I3(GND_net), .O(n1050));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i706_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_15_i16_3_lut (.I0(n257[9]), .I1(n257[21]), .I2(n43_adj_4005), 
            .I3(GND_net), .O(n16_adj_4006));   // verilog/motorControl.v(46[19:35])
    defparam LessThan_15_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_4120_3 (.CI(n29270), .I0(n8482[0]), .I1(n180), .CO(n29271));
    SB_LUT4 add_4120_2_lut (.I0(GND_net), .I1(n38), .I2(n107), .I3(GND_net), 
            .O(n8468[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4120_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4136_16 (.CI(n29439), .I0(n8680[13]), .I1(n1111), .CO(n29440));
    SB_LUT4 mult_11_i745_2_lut (.I0(\Ki[15] ), .I1(\PID_CONTROLLER.integral [4]), 
            .I2(GND_net), .I3(GND_net), .O(n1108));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i745_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i71_2_lut (.I0(\Kp[1] ), .I1(\PID_CONTROLLER.err [10]), 
            .I2(GND_net), .I3(GND_net), .O(n104));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i71_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i751_2_lut (.I0(\Ki[15] ), .I1(\PID_CONTROLLER.integral [7]), 
            .I2(GND_net), .I3(GND_net), .O(n1117));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i751_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i300_2_lut (.I0(\Kp[6] ), .I1(\PID_CONTROLLER.err [2]), 
            .I2(GND_net), .I3(GND_net), .O(n445));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i300_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i230_2_lut (.I0(\Kp[4] ), .I1(\PID_CONTROLLER.err [16]), 
            .I2(GND_net), .I3(GND_net), .O(n341));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i230_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i24_2_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err [11]), 
            .I2(GND_net), .I3(GND_net), .O(n35_adj_4007));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i24_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i61_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral [5]), 
            .I2(GND_net), .I3(GND_net), .O(n89));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i61_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 state_23__I_0_inv_0_i17_1_lut (.I0(setpoint[16]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4333[16]));   // verilog/motorControl.v(38[14:30])
    defparam state_23__I_0_inv_0_i17_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_11_i14_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral [6]), 
            .I2(GND_net), .I3(GND_net), .O(n20_adj_4009));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i14_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i120_2_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err [10]), 
            .I2(GND_net), .I3(GND_net), .O(n177));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i120_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i110_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral [5]), 
            .I2(GND_net), .I3(GND_net), .O(n162));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i110_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_666_i24_3_lut (.I0(n37312), .I1(PWMLimit[23]), .I2(n256), 
            .I3(GND_net), .O(n3290[23]));   // verilog/motorControl.v(46[16] 48[10])
    defparam mux_666_i24_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 mult_10_i149_2_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err [0]), 
            .I2(GND_net), .I3(GND_net), .O(n220));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i149_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 state_23__I_0_inv_0_i18_1_lut (.I0(setpoint[17]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4333[17]));   // verilog/motorControl.v(38[14:30])
    defparam state_23__I_0_inv_0_i18_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i169_2_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err [10]), 
            .I2(GND_net), .I3(GND_net), .O(n250));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i169_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i159_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral [5]), 
            .I2(GND_net), .I3(GND_net), .O(n235));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i159_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i208_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral [5]), 
            .I2(GND_net), .I3(GND_net), .O(n308));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i208_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i257_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral [5]), 
            .I2(GND_net), .I3(GND_net), .O(n381));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i257_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i218_2_lut (.I0(\Kp[4] ), .I1(\PID_CONTROLLER.err [10]), 
            .I2(GND_net), .I3(GND_net), .O(n323));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i218_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i306_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral [5]), 
            .I2(GND_net), .I3(GND_net), .O(n454));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i306_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i267_2_lut (.I0(\Kp[5] ), .I1(\PID_CONTROLLER.err [10]), 
            .I2(GND_net), .I3(GND_net), .O(n396));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i267_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i261_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral [7]), 
            .I2(GND_net), .I3(GND_net), .O(n387));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i261_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_4120_2 (.CI(GND_net), .I0(n38), .I1(n107), .CO(n29270));
    SB_LUT4 unary_minus_5_add_3_22_lut (.I0(\PID_CONTROLLER.integral [20]), 
            .I1(GND_net), .I2(n1_adj_4332[20]), .I3(n28105), .O(n41_adj_4011)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_22_lut.LUT_INIT = 16'h6996;
    SB_LUT4 add_4136_15_lut (.I0(GND_net), .I1(n8680[12]), .I2(n1038), 
            .I3(n29438), .O(n8660[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4136_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i355_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral [5]), 
            .I2(GND_net), .I3(GND_net), .O(n527));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i355_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_4119_14_lut (.I0(GND_net), .I1(n8468[11]), .I2(n980), 
            .I3(n29269), .O(n8453[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4119_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4136_15 (.CI(n29438), .I0(n8680[12]), .I1(n1038), .CO(n29439));
    SB_LUT4 add_4136_14_lut (.I0(GND_net), .I1(n8680[11]), .I2(n965), 
            .I3(n29437), .O(n8660[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4136_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4136_14 (.CI(n29437), .I0(n8680[11]), .I1(n965), .CO(n29438));
    SB_LUT4 mult_10_i349_2_lut (.I0(\Kp[7] ), .I1(\PID_CONTROLLER.err [2]), 
            .I2(GND_net), .I3(GND_net), .O(n518));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i349_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_4136_13_lut (.I0(GND_net), .I1(n8680[10]), .I2(n892), 
            .I3(n29436), .O(n8660[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4136_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4110_23_lut (.I0(GND_net), .I1(n8297[20]), .I2(GND_net), 
            .I3(n28735), .O(n8273[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4110_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4110_22_lut (.I0(GND_net), .I1(n8297[19]), .I2(GND_net), 
            .I3(n28734), .O(n8273[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4110_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4119_13_lut (.I0(GND_net), .I1(n8468[10]), .I2(n907), 
            .I3(n29268), .O(n8453[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4119_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4136_13 (.CI(n29436), .I0(n8680[10]), .I1(n892), .CO(n29437));
    SB_CARRY add_4110_22 (.CI(n28734), .I0(n8297[19]), .I1(GND_net), .CO(n28735));
    SB_LUT4 add_4110_21_lut (.I0(GND_net), .I1(n8297[18]), .I2(GND_net), 
            .I3(n28733), .O(n8273[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4110_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4119_13 (.CI(n29268), .I0(n8468[10]), .I1(n907), .CO(n29269));
    SB_LUT4 add_4119_12_lut (.I0(GND_net), .I1(n8468[9]), .I2(n834), .I3(n29267), 
            .O(n8453[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4119_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i404_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral [5]), 
            .I2(GND_net), .I3(GND_net), .O(n600));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i404_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_inv_0_i6_1_lut (.I0(IntegralLimit[5]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4332[5]));   // verilog/motorControl.v(39[48:62])
    defparam unary_minus_5_inv_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY unary_minus_5_add_3_22 (.CI(n28105), .I0(GND_net), .I1(n1_adj_4332[20]), 
            .CO(n28106));
    SB_CARRY add_4119_12 (.CI(n29267), .I0(n8468[9]), .I1(n834), .CO(n29268));
    SB_LUT4 mult_10_i316_2_lut (.I0(\Kp[6] ), .I1(\PID_CONTROLLER.err [10]), 
            .I2(GND_net), .I3(GND_net), .O(n469));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i316_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_4136_12_lut (.I0(GND_net), .I1(n8680[9]), .I2(n819), .I3(n29435), 
            .O(n8660[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4136_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_5_add_3_21_lut (.I0(\PID_CONTROLLER.integral [19]), 
            .I1(GND_net), .I2(n1_adj_4332[19]), .I3(n28104), .O(n39_adj_4014)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_21_lut.LUT_INIT = 16'h6996;
    SB_CARRY add_4136_12 (.CI(n29435), .I0(n8680[9]), .I1(n819), .CO(n29436));
    SB_LUT4 add_4136_11_lut (.I0(GND_net), .I1(n8680[8]), .I2(n746), .I3(n29434), 
            .O(n8660[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4136_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4110_21 (.CI(n28733), .I0(n8297[18]), .I1(GND_net), .CO(n28734));
    SB_LUT4 add_4110_20_lut (.I0(GND_net), .I1(n8297[17]), .I2(GND_net), 
            .I3(n28732), .O(n8273[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4110_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4119_11_lut (.I0(GND_net), .I1(n8468[8]), .I2(n761), .I3(n29266), 
            .O(n8453[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4119_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i31267_3_lut (.I0(n6_adj_4016), .I1(n257[10]), .I2(n21_adj_3923), 
            .I3(GND_net), .O(n37949));   // verilog/motorControl.v(46[19:35])
    defparam i31267_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_4119_11 (.CI(n29266), .I0(n8468[8]), .I1(n761), .CO(n29267));
    SB_CARRY add_4136_11 (.CI(n29434), .I0(n8680[8]), .I1(n746), .CO(n29435));
    SB_LUT4 add_4136_10_lut (.I0(GND_net), .I1(n8680[7]), .I2(n673), .I3(n29433), 
            .O(n8660[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4136_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i312_2_lut (.I0(\Kp[6] ), .I1(\PID_CONTROLLER.err [8]), 
            .I2(GND_net), .I3(GND_net), .O(n463_adj_4017));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i312_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_666_i15_3_lut (.I0(n155[14]), .I1(PWMLimit[14]), .I2(n256), 
            .I3(GND_net), .O(n3290[14]));   // verilog/motorControl.v(46[16] 48[10])
    defparam mux_666_i15_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 mult_10_i365_2_lut (.I0(\Kp[7] ), .I1(\PID_CONTROLLER.err [10]), 
            .I2(GND_net), .I3(GND_net), .O(n542));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i365_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i414_2_lut (.I0(\Kp[8] ), .I1(\PID_CONTROLLER.err [10]), 
            .I2(GND_net), .I3(GND_net), .O(n615));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i414_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_4136_10 (.CI(n29433), .I0(n8680[7]), .I1(n673), .CO(n29434));
    SB_LUT4 add_4119_10_lut (.I0(GND_net), .I1(n8468[7]), .I2(n688), .I3(n29265), 
            .O(n8453[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4119_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4119_10 (.CI(n29265), .I0(n8468[7]), .I1(n688), .CO(n29266));
    SB_LUT4 add_4119_9_lut (.I0(GND_net), .I1(n8468[6]), .I2(n615), .I3(n29264), 
            .O(n8453[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4119_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i463_2_lut (.I0(\Kp[9] ), .I1(\PID_CONTROLLER.err [10]), 
            .I2(GND_net), .I3(GND_net), .O(n688));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i463_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_4119_9 (.CI(n29264), .I0(n8468[6]), .I1(n615), .CO(n29265));
    SB_LUT4 add_4119_8_lut (.I0(GND_net), .I1(n8468[5]), .I2(n542), .I3(n29263), 
            .O(n8453[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4119_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i453_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral [5]), 
            .I2(GND_net), .I3(GND_net), .O(n673));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i453_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_4119_8 (.CI(n29263), .I0(n8468[5]), .I1(n542), .CO(n29264));
    SB_LUT4 mult_10_i512_2_lut (.I0(\Kp[10] ), .I1(\PID_CONTROLLER.err [10]), 
            .I2(GND_net), .I3(GND_net), .O(n761));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i512_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_4119_7_lut (.I0(GND_net), .I1(n8468[4]), .I2(n469), .I3(n29262), 
            .O(n8453[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4119_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i398_2_lut (.I0(\Kp[8] ), .I1(\PID_CONTROLLER.err [2]), 
            .I2(GND_net), .I3(GND_net), .O(n591));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i398_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_4119_7 (.CI(n29262), .I0(n8468[4]), .I1(n469), .CO(n29263));
    SB_LUT4 add_4136_9_lut (.I0(GND_net), .I1(n8680[6]), .I2(n600), .I3(n29432), 
            .O(n8660[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4136_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4136_9 (.CI(n29432), .I0(n8680[6]), .I1(n600), .CO(n29433));
    SB_LUT4 add_4136_8_lut (.I0(GND_net), .I1(n8680[5]), .I2(n527), .I3(n29431), 
            .O(n8660[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4136_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4119_6_lut (.I0(GND_net), .I1(n8468[3]), .I2(n396), .I3(n29261), 
            .O(n8453[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4119_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4136_8 (.CI(n29431), .I0(n8680[5]), .I1(n527), .CO(n29432));
    SB_LUT4 add_4136_7_lut (.I0(GND_net), .I1(n8680[4]), .I2(n454), .I3(n29430), 
            .O(n8660[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4136_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4136_7 (.CI(n29430), .I0(n8680[4]), .I1(n454), .CO(n29431));
    SB_CARRY add_4119_6 (.CI(n29261), .I0(n8468[3]), .I1(n396), .CO(n29262));
    SB_LUT4 add_4119_5_lut (.I0(GND_net), .I1(n8468[2]), .I2(n323), .I3(n29260), 
            .O(n8453[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4119_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4136_6_lut (.I0(GND_net), .I1(n8680[3]), .I2(n381), .I3(n29429), 
            .O(n8660[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4136_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4136_6 (.CI(n29429), .I0(n8680[3]), .I1(n381), .CO(n29430));
    SB_LUT4 add_4136_5_lut (.I0(GND_net), .I1(n8680[2]), .I2(n308), .I3(n29428), 
            .O(n8660[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4136_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4136_5 (.CI(n29428), .I0(n8680[2]), .I1(n308), .CO(n29429));
    SB_LUT4 i31268_3_lut (.I0(n37949), .I1(n257[11]), .I2(n23_adj_3926), 
            .I3(GND_net), .O(n37950));   // verilog/motorControl.v(46[19:35])
    defparam i31268_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_10_i279_2_lut (.I0(\Kp[5] ), .I1(\PID_CONTROLLER.err [16]), 
            .I2(GND_net), .I3(GND_net), .O(n414));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i279_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY unary_minus_5_add_3_21 (.CI(n28104), .I0(GND_net), .I1(n1_adj_4332[19]), 
            .CO(n28105));
    SB_LUT4 add_4136_4_lut (.I0(GND_net), .I1(n8680[1]), .I2(n235), .I3(n29427), 
            .O(n8660[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4136_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4119_5 (.CI(n29260), .I0(n8468[2]), .I1(n323), .CO(n29261));
    SB_CARRY add_4136_4 (.CI(n29427), .I0(n8680[1]), .I1(n235), .CO(n29428));
    SB_LUT4 add_4119_4_lut (.I0(GND_net), .I1(n8468[1]), .I2(n250), .I3(n29259), 
            .O(n8453[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4119_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_668_25_lut (.I0(GND_net), .I1(n3265[23]), .I2(n3290[23]), 
            .I3(n27993), .O(duty_23__N_3613[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_668_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4119_4 (.CI(n29259), .I0(n8468[1]), .I1(n250), .CO(n29260));
    SB_LUT4 add_4136_3_lut (.I0(GND_net), .I1(n8680[0]), .I2(n162), .I3(n29426), 
            .O(n8660[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4136_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4119_3_lut (.I0(GND_net), .I1(n8468[0]), .I2(n177), .I3(n29258), 
            .O(n8453[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4119_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4119_3 (.CI(n29258), .I0(n8468[0]), .I1(n177), .CO(n29259));
    SB_CARRY add_4136_3 (.CI(n29426), .I0(n8680[0]), .I1(n162), .CO(n29427));
    SB_LUT4 add_4136_2_lut (.I0(GND_net), .I1(n20_adj_4009), .I2(n89), 
            .I3(GND_net), .O(n8660[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4136_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4136_2 (.CI(GND_net), .I0(n20_adj_4009), .I1(n89), .CO(n29426));
    SB_LUT4 add_4135_20_lut (.I0(GND_net), .I1(n8660[17]), .I2(GND_net), 
            .I3(n29425), .O(n8639[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4135_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i655_2_lut (.I0(\Ki[13] ), .I1(\PID_CONTROLLER.integral [8]), 
            .I2(GND_net), .I3(GND_net), .O(n974));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i655_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_4135_19_lut (.I0(GND_net), .I1(n8660[16]), .I2(GND_net), 
            .I3(n29424), .O(n8639[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4135_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4135_19 (.CI(n29424), .I0(n8660[16]), .I1(GND_net), .CO(n29425));
    SB_LUT4 add_4119_2_lut (.I0(GND_net), .I1(n35_adj_4007), .I2(n104), 
            .I3(GND_net), .O(n8453[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4119_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4135_18_lut (.I0(GND_net), .I1(n8660[15]), .I2(GND_net), 
            .I3(n29423), .O(n8639[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4135_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4135_18 (.CI(n29423), .I0(n8660[15]), .I1(GND_net), .CO(n29424));
    SB_LUT4 add_4135_17_lut (.I0(GND_net), .I1(n8660[14]), .I2(GND_net), 
            .I3(n29422), .O(n8639[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4135_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4119_2 (.CI(GND_net), .I0(n35_adj_4007), .I1(n104), .CO(n29258));
    SB_CARRY add_4135_17 (.CI(n29422), .I0(n8660[14]), .I1(GND_net), .CO(n29423));
    SB_LUT4 add_4135_16_lut (.I0(GND_net), .I1(n8660[13]), .I2(n1108), 
            .I3(n29421), .O(n8639[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4135_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4135_16 (.CI(n29421), .I0(n8660[13]), .I1(n1108), .CO(n29422));
    SB_LUT4 mult_11_i502_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral [5]), 
            .I2(GND_net), .I3(GND_net), .O(n746));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i502_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_inv_0_i20_1_lut (.I0(IntegralLimit[19]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4332[19]));   // verilog/motorControl.v(39[48:62])
    defparam unary_minus_5_inv_0_i20_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_11_i704_2_lut (.I0(\Ki[14] ), .I1(\PID_CONTROLLER.integral [8]), 
            .I2(GND_net), .I3(GND_net), .O(n1047));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i704_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_4118_15_lut (.I0(GND_net), .I1(n8453[12]), .I2(n1050), 
            .I3(n29257), .O(n8437[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4118_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4118_14_lut (.I0(GND_net), .I1(n8453[11]), .I2(n977), 
            .I3(n29256), .O(n8437[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4118_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 state_23__I_0_inv_0_i19_1_lut (.I0(setpoint[18]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4333[18]));   // verilog/motorControl.v(38[14:30])
    defparam state_23__I_0_inv_0_i19_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_11_i551_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral [5]), 
            .I2(GND_net), .I3(GND_net), .O(n819));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i551_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_4135_15_lut (.I0(GND_net), .I1(n8660[12]), .I2(n1035), 
            .I3(n29420), .O(n8639[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4135_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4135_15 (.CI(n29420), .I0(n8660[12]), .I1(n1035), .CO(n29421));
    SB_LUT4 unary_minus_5_add_3_20_lut (.I0(\PID_CONTROLLER.integral [18]), 
            .I1(GND_net), .I2(n1_adj_4332[18]), .I3(n28103), .O(n37_adj_4020)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_20_lut.LUT_INIT = 16'h6996;
    SB_CARRY add_4118_14 (.CI(n29256), .I0(n8453[11]), .I1(n977), .CO(n29257));
    SB_LUT4 mult_11_i645_2_lut (.I0(\Ki[13] ), .I1(\PID_CONTROLLER.integral [3]), 
            .I2(GND_net), .I3(GND_net), .O(n959));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i645_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_4135_14_lut (.I0(GND_net), .I1(n8660[11]), .I2(n962), 
            .I3(n29419), .O(n8639[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4135_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_16_inv_0_i12_1_lut (.I0(PWMLimit[11]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[11]));   // verilog/motorControl.v(47[19:28])
    defparam unary_minus_16_inv_0_i12_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_11_i753_2_lut (.I0(\Ki[15] ), .I1(\PID_CONTROLLER.integral [8]), 
            .I2(GND_net), .I3(GND_net), .O(n1120));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i753_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i130_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral [15]), 
            .I2(GND_net), .I3(GND_net), .O(n192_adj_4022));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i130_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i328_2_lut (.I0(\Kp[6] ), .I1(\PID_CONTROLLER.err [16]), 
            .I2(GND_net), .I3(GND_net), .O(n487));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i328_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_4118_13_lut (.I0(GND_net), .I1(n8453[10]), .I2(n904), 
            .I3(n29255), .O(n8437[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4118_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_668_24_lut (.I0(GND_net), .I1(n3265[22]), .I2(n3290[22]), 
            .I3(n27992), .O(duty_23__N_3613[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_668_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4135_14 (.CI(n29419), .I0(n8660[11]), .I1(n962), .CO(n29420));
    SB_LUT4 mult_10_i377_2_lut (.I0(\Kp[7] ), .I1(\PID_CONTROLLER.err [16]), 
            .I2(GND_net), .I3(GND_net), .O(n560));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i377_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_4135_13_lut (.I0(GND_net), .I1(n8660[10]), .I2(n889), 
            .I3(n29418), .O(n8639[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4135_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4135_13 (.CI(n29418), .I0(n8660[10]), .I1(n889), .CO(n29419));
    SB_LUT4 mult_10_i447_2_lut (.I0(\Kp[9] ), .I1(\PID_CONTROLLER.err [2]), 
            .I2(GND_net), .I3(GND_net), .O(n664));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i447_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY unary_minus_5_add_3_20 (.CI(n28103), .I0(GND_net), .I1(n1_adj_4332[18]), 
            .CO(n28104));
    SB_LUT4 unary_minus_5_add_3_19_lut (.I0(\PID_CONTROLLER.integral [17]), 
            .I1(GND_net), .I2(n1_adj_4332[17]), .I3(n28102), .O(n35_adj_4023)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_19_lut.LUT_INIT = 16'h6996;
    SB_LUT4 add_4135_12_lut (.I0(GND_net), .I1(n8660[9]), .I2(n816), .I3(n29417), 
            .O(n8639[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4135_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4135_12 (.CI(n29417), .I0(n8660[9]), .I1(n816), .CO(n29418));
    SB_CARRY add_4110_20 (.CI(n28732), .I0(n8297[17]), .I1(GND_net), .CO(n28733));
    SB_CARRY add_4118_13 (.CI(n29255), .I0(n8453[10]), .I1(n904), .CO(n29256));
    SB_LUT4 add_4118_12_lut (.I0(GND_net), .I1(n8453[9]), .I2(n831), .I3(n29254), 
            .O(n8437[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4118_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 state_23__I_0_inv_0_i20_1_lut (.I0(setpoint[19]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4333[19]));   // verilog/motorControl.v(38[14:30])
    defparam state_23__I_0_inv_0_i20_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY unary_minus_5_add_3_19 (.CI(n28102), .I0(GND_net), .I1(n1_adj_4332[17]), 
            .CO(n28103));
    SB_CARRY add_668_24 (.CI(n27992), .I0(n3265[22]), .I1(n3290[22]), 
            .CO(n27993));
    SB_LUT4 add_668_23_lut (.I0(GND_net), .I1(n3265[21]), .I2(n3290[21]), 
            .I3(n27991), .O(duty_23__N_3613[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_668_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4135_11_lut (.I0(GND_net), .I1(n8660[8]), .I2(n743), .I3(n29416), 
            .O(n8639[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4135_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4118_12 (.CI(n29254), .I0(n8453[9]), .I1(n831), .CO(n29255));
    SB_LUT4 add_4110_19_lut (.I0(GND_net), .I1(n8297[16]), .I2(GND_net), 
            .I3(n28731), .O(n8273[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4110_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_5_add_3_18_lut (.I0(\PID_CONTROLLER.integral [16]), 
            .I1(GND_net), .I2(n1_adj_4332[16]), .I3(n28101), .O(n33_adj_4025)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_18_lut.LUT_INIT = 16'h6996;
    SB_CARRY add_4135_11 (.CI(n29416), .I0(n8660[8]), .I1(n743), .CO(n29417));
    SB_CARRY add_668_23 (.CI(n27991), .I0(n3265[21]), .I1(n3290[21]), 
            .CO(n27992));
    SB_CARRY unary_minus_5_add_3_18 (.CI(n28101), .I0(GND_net), .I1(n1_adj_4332[16]), 
            .CO(n28102));
    SB_LUT4 add_4118_11_lut (.I0(GND_net), .I1(n8453[8]), .I2(n758), .I3(n29253), 
            .O(n8437[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4118_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_668_22_lut (.I0(GND_net), .I1(n3265[20]), .I2(n3290[20]), 
            .I3(n27990), .O(duty_23__N_3613[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_668_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4118_11 (.CI(n29253), .I0(n8453[8]), .I1(n758), .CO(n29254));
    SB_LUT4 add_4135_10_lut (.I0(GND_net), .I1(n8660[7]), .I2(n670), .I3(n29415), 
            .O(n8639[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4135_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_668_22 (.CI(n27990), .I0(n3265[20]), .I1(n3290[20]), 
            .CO(n27991));
    SB_LUT4 mult_11_i694_2_lut (.I0(\Ki[14] ), .I1(\PID_CONTROLLER.integral [3]), 
            .I2(GND_net), .I3(GND_net), .O(n1032));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i694_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_add_3_17_lut (.I0(\PID_CONTROLLER.integral [15]), 
            .I1(GND_net), .I2(n1_adj_4332[15]), .I3(n28100), .O(n31_adj_4026)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_17_lut.LUT_INIT = 16'h6996;
    SB_CARRY add_4110_19 (.CI(n28731), .I0(n8297[16]), .I1(GND_net), .CO(n28732));
    SB_LUT4 add_4118_10_lut (.I0(GND_net), .I1(n8453[7]), .I2(n685), .I3(n29252), 
            .O(n8437[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4118_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i179_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral [15]), 
            .I2(GND_net), .I3(GND_net), .O(n265_adj_4027));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i179_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_4110_18_lut (.I0(GND_net), .I1(n8297[15]), .I2(GND_net), 
            .I3(n28730), .O(n8273[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4110_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4110_18 (.CI(n28730), .I0(n8297[15]), .I1(GND_net), .CO(n28731));
    SB_LUT4 add_4110_17_lut (.I0(GND_net), .I1(n8297[14]), .I2(GND_net), 
            .I3(n28729), .O(n8273[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4110_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4110_17 (.CI(n28729), .I0(n8297[14]), .I1(GND_net), .CO(n28730));
    SB_LUT4 add_4110_16_lut (.I0(GND_net), .I1(n8297[13]), .I2(n1099), 
            .I3(n28728), .O(n8273[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4110_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4110_16 (.CI(n28728), .I0(n8297[13]), .I1(n1099), .CO(n28729));
    SB_LUT4 add_4110_15_lut (.I0(GND_net), .I1(n8297[12]), .I2(n1026), 
            .I3(n28727), .O(n8273[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4110_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4110_15 (.CI(n28727), .I0(n8297[12]), .I1(n1026), .CO(n28728));
    SB_LUT4 add_4110_14_lut (.I0(GND_net), .I1(n8297[11]), .I2(n953), 
            .I3(n28726), .O(n8273[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4110_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4110_14 (.CI(n28726), .I0(n8297[11]), .I1(n953), .CO(n28727));
    SB_LUT4 add_4110_13_lut (.I0(GND_net), .I1(n8297[10]), .I2(n880), 
            .I3(n28725), .O(n8273[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4110_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4118_10 (.CI(n29252), .I0(n8453[7]), .I1(n685), .CO(n29253));
    SB_LUT4 add_4118_9_lut (.I0(GND_net), .I1(n8453[6]), .I2(n612), .I3(n29251), 
            .O(n8437[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4118_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 state_23__I_0_inv_0_i21_1_lut (.I0(setpoint[20]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4333[20]));   // verilog/motorControl.v(38[14:30])
    defparam state_23__I_0_inv_0_i21_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_4110_13 (.CI(n28725), .I0(n8297[10]), .I1(n880), .CO(n28726));
    SB_CARRY add_4118_9 (.CI(n29251), .I0(n8453[6]), .I1(n612), .CO(n29252));
    SB_LUT4 mult_10_i361_2_lut (.I0(\Kp[7] ), .I1(\PID_CONTROLLER.err [8]), 
            .I2(GND_net), .I3(GND_net), .O(n536_adj_4029));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i361_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i228_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral [15]), 
            .I2(GND_net), .I3(GND_net), .O(n338_adj_4030));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i228_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i277_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral [15]), 
            .I2(GND_net), .I3(GND_net), .O(n411_adj_4031));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i277_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 state_23__I_0_inv_0_i22_1_lut (.I0(setpoint[21]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4333[21]));   // verilog/motorControl.v(38[14:30])
    defparam state_23__I_0_inv_0_i22_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i410_2_lut (.I0(\Kp[8] ), .I1(\PID_CONTROLLER.err [8]), 
            .I2(GND_net), .I3(GND_net), .O(n609_adj_4033));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i410_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 state_23__I_0_inv_0_i23_1_lut (.I0(setpoint[22]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4333[22]));   // verilog/motorControl.v(38[14:30])
    defparam state_23__I_0_inv_0_i23_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_4110_12_lut (.I0(GND_net), .I1(n8297[9]), .I2(n807), .I3(n28724), 
            .O(n8273[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4110_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4110_12 (.CI(n28724), .I0(n8297[9]), .I1(n807), .CO(n28725));
    SB_CARRY add_4135_10 (.CI(n29415), .I0(n8660[7]), .I1(n670), .CO(n29416));
    SB_LUT4 state_23__I_0_inv_0_i24_1_lut (.I0(setpoint[23]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4333[23]));   // verilog/motorControl.v(38[14:30])
    defparam state_23__I_0_inv_0_i24_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_4110_11_lut (.I0(GND_net), .I1(n8297[8]), .I2(n734), .I3(n28723), 
            .O(n8273[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4110_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i85_2_lut (.I0(\Kp[1] ), .I1(\PID_CONTROLLER.err [17]), 
            .I2(GND_net), .I3(GND_net), .O(n125));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i85_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_4118_8_lut (.I0(GND_net), .I1(n8453[5]), .I2(n539), .I3(n29250), 
            .O(n8437[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4118_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4118_8 (.CI(n29250), .I0(n8453[5]), .I1(n539), .CO(n29251));
    SB_CARRY add_4110_11 (.CI(n28723), .I0(n8297[8]), .I1(n734), .CO(n28724));
    SB_LUT4 add_4118_7_lut (.I0(GND_net), .I1(n8453[4]), .I2(n466), .I3(n29249), 
            .O(n8437[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4118_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_15_i8_3_lut (.I0(n257[4]), .I1(n257[8]), .I2(n17_adj_3925), 
            .I3(GND_net), .O(n8_adj_4036));   // verilog/motorControl.v(46[19:35])
    defparam LessThan_15_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_10_i38_2_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err [18]), 
            .I2(GND_net), .I3(GND_net), .O(n56));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i38_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY unary_minus_5_add_3_17 (.CI(n28100), .I0(GND_net), .I1(n1_adj_4332[15]), 
            .CO(n28101));
    SB_LUT4 LessThan_15_i24_3_lut (.I0(n16_adj_4006), .I1(n257[22]), .I2(n45_adj_4038), 
            .I3(GND_net), .O(n24_adj_4039));   // verilog/motorControl.v(46[19:35])
    defparam LessThan_15_i24_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_668_21_lut (.I0(GND_net), .I1(n3265[19]), .I2(n3290[19]), 
            .I3(n27989), .O(duty_23__N_3613[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_668_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4110_10_lut (.I0(GND_net), .I1(n8297[7]), .I2(n661), .I3(n28722), 
            .O(n8273[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4110_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4135_9_lut (.I0(GND_net), .I1(n8660[6]), .I2(n597), .I3(n29414), 
            .O(n8639[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4135_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4110_10 (.CI(n28722), .I0(n8297[7]), .I1(n661), .CO(n28723));
    SB_LUT4 add_4110_9_lut (.I0(GND_net), .I1(n8297[6]), .I2(n588), .I3(n28721), 
            .O(n8273[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4110_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4118_7 (.CI(n29249), .I0(n8453[4]), .I1(n466), .CO(n29250));
    SB_CARRY add_4110_9 (.CI(n28721), .I0(n8297[6]), .I1(n588), .CO(n28722));
    SB_LUT4 mult_11_i743_2_lut (.I0(\Ki[15] ), .I1(\PID_CONTROLLER.integral [3]), 
            .I2(GND_net), .I3(GND_net), .O(n1105));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i743_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i326_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral [15]), 
            .I2(GND_net), .I3(GND_net), .O(n484_adj_4040));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i326_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_4110_8_lut (.I0(GND_net), .I1(n8297[5]), .I2(n515), .I3(n28720), 
            .O(n8273[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4110_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4110_8 (.CI(n28720), .I0(n8297[5]), .I1(n515), .CO(n28721));
    SB_LUT4 add_4110_7_lut (.I0(GND_net), .I1(n8297[4]), .I2(n442), .I3(n28719), 
            .O(n8273[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4110_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i653_2_lut (.I0(\Ki[13] ), .I1(\PID_CONTROLLER.integral [7]), 
            .I2(GND_net), .I3(GND_net), .O(n971));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i653_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_4110_7 (.CI(n28719), .I0(n8297[4]), .I1(n442), .CO(n28720));
    SB_LUT4 mult_10_i459_2_lut (.I0(\Kp[9] ), .I1(\PID_CONTROLLER.err [8]), 
            .I2(GND_net), .I3(GND_net), .O(n682_adj_4041));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i459_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i508_2_lut (.I0(\Kp[10] ), .I1(\PID_CONTROLLER.err [8]), 
            .I2(GND_net), .I3(GND_net), .O(n755_adj_4042));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i508_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i496_2_lut (.I0(\Kp[10] ), .I1(\PID_CONTROLLER.err [2]), 
            .I2(GND_net), .I3(GND_net), .O(n737));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i496_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_inv_0_i7_1_lut (.I0(IntegralLimit[6]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4332[6]));   // verilog/motorControl.v(39[48:62])
    defparam unary_minus_5_inv_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mux_666_i16_3_lut (.I0(n155[15]), .I1(PWMLimit[15]), .I2(n256), 
            .I3(GND_net), .O(n3290[15]));   // verilog/motorControl.v(46[16] 48[10])
    defparam mux_666_i16_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 unary_minus_16_inv_0_i13_1_lut (.I0(PWMLimit[12]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[12]));   // verilog/motorControl.v(47[19:28])
    defparam unary_minus_16_inv_0_i13_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_4135_9 (.CI(n29414), .I0(n8660[6]), .I1(n597), .CO(n29415));
    SB_LUT4 add_4135_8_lut (.I0(GND_net), .I1(n8660[5]), .I2(n524), .I3(n29413), 
            .O(n8639[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4135_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i371_2_lut (.I0(\Kp[7] ), .I1(\PID_CONTROLLER.err [13]), 
            .I2(GND_net), .I3(GND_net), .O(n551));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i371_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i51_2_lut (.I0(\Kp[1] ), .I1(\PID_CONTROLLER.err [0]), 
            .I2(GND_net), .I3(GND_net), .O(n74));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i51_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i4_2_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err [1]), 
            .I2(GND_net), .I3(GND_net), .O(n5));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i4_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i702_2_lut (.I0(\Ki[14] ), .I1(\PID_CONTROLLER.integral [7]), 
            .I2(GND_net), .I3(GND_net), .O(n1044));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i702_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_4118_6_lut (.I0(GND_net), .I1(n8453[3]), .I2(n393), .I3(n29248), 
            .O(n8437[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4118_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i420_2_lut (.I0(\Kp[8] ), .I1(\PID_CONTROLLER.err [13]), 
            .I2(GND_net), .I3(GND_net), .O(n624));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i420_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i545_2_lut (.I0(\Kp[11] ), .I1(\PID_CONTROLLER.err [2]), 
            .I2(GND_net), .I3(GND_net), .O(n810));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i545_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_668_21 (.CI(n27989), .I0(n3265[19]), .I1(n3290[19]), 
            .CO(n27990));
    SB_LUT4 i22918_3_lut_4_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral [18]), 
            .I2(n4_adj_4045), .I3(n8849[1]), .O(n6_adj_4046));   // verilog/motorControl.v(42[26:37])
    defparam i22918_3_lut_4_lut.LUT_INIT = 16'hf880;
    SB_LUT4 i2_3_lut_4_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral [18]), 
            .I2(n8849[1]), .I3(n4_adj_4045), .O(n8842[2]));   // verilog/motorControl.v(42[26:37])
    defparam i2_3_lut_4_lut.LUT_INIT = 16'h8778;
    SB_LUT4 unary_minus_16_inv_0_i14_1_lut (.I0(PWMLimit[13]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[13]));   // verilog/motorControl.v(47[19:28])
    defparam unary_minus_16_inv_0_i14_1_lut.LUT_INIT = 16'h5555;
    SB_DFFE \PID_CONTROLLER.integral_1526__i0  (.Q(\PID_CONTROLLER.integral [0]), 
            .C(clk32MHz), .E(\PID_CONTROLLER.integral_23__N_3586 ), .D(n28[0]));   // verilog/motorControl.v(40[21:33])
    SB_LUT4 i30744_4_lut (.I0(n43_adj_4005), .I1(n25_adj_4049), .I2(n23_adj_3926), 
            .I3(n37464), .O(n37425));
    defparam i30744_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 unary_minus_5_add_3_16_lut (.I0(\PID_CONTROLLER.integral [14]), 
            .I1(GND_net), .I2(n1_adj_4332[14]), .I3(n28099), .O(n29_adj_4050)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_16_lut.LUT_INIT = 16'h6996;
    SB_LUT4 add_4148_7_lut (.I0(GND_net), .I1(n35470), .I2(n490), .I3(n29568), 
            .O(n8834[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4148_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i31249_4_lut (.I0(n24_adj_4039), .I1(n8_adj_4036), .I2(n45_adj_4038), 
            .I3(n37423), .O(n37931));   // verilog/motorControl.v(46[19:35])
    defparam i31249_4_lut.LUT_INIT = 16'haaac;
    SB_CARRY unary_minus_5_add_3_16 (.CI(n28099), .I0(GND_net), .I1(n1_adj_4332[14]), 
            .CO(n28100));
    SB_CARRY add_4135_8 (.CI(n29413), .I0(n8660[5]), .I1(n524), .CO(n29414));
    SB_LUT4 unary_minus_5_add_3_15_lut (.I0(\PID_CONTROLLER.integral [13]), 
            .I1(GND_net), .I2(n1_adj_4332[13]), .I3(n28098), .O(n27_adj_4052)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_15_lut.LUT_INIT = 16'h6996;
    SB_CARRY add_4118_6 (.CI(n29248), .I0(n8453[3]), .I1(n393), .CO(n29249));
    SB_CARRY unary_minus_5_add_3_15 (.CI(n28098), .I0(GND_net), .I1(n1_adj_4332[13]), 
            .CO(n28099));
    SB_LUT4 mult_10_i134_2_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err [17]), 
            .I2(GND_net), .I3(GND_net), .O(n198));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i134_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_4135_7_lut (.I0(GND_net), .I1(n8660[4]), .I2(n451), .I3(n29412), 
            .O(n8639[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4135_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i31072_3_lut (.I0(n37950), .I1(n257[12]), .I2(n25_adj_4049), 
            .I3(GND_net), .O(n37754));   // verilog/motorControl.v(46[19:35])
    defparam i31072_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_4135_7 (.CI(n29412), .I0(n8660[4]), .I1(n451), .CO(n29413));
    SB_LUT4 add_4110_6_lut (.I0(GND_net), .I1(n8297[3]), .I2(n369), .I3(n28718), 
            .O(n8273[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4110_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4148_6_lut (.I0(GND_net), .I1(n8842[3]), .I2(n417), .I3(n29567), 
            .O(n8834[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4148_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4148_6 (.CI(n29567), .I0(n8842[3]), .I1(n417), .CO(n29568));
    SB_LUT4 mult_10_i594_2_lut (.I0(\Kp[12] ), .I1(\PID_CONTROLLER.err [2]), 
            .I2(GND_net), .I3(GND_net), .O(n883));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i594_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_15_i4_3_lut (.I0(n37256), .I1(n257[1]), .I2(duty[1]), 
            .I3(GND_net), .O(n4_adj_4054));   // verilog/motorControl.v(46[19:35])
    defparam LessThan_15_i4_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 add_4135_6_lut (.I0(GND_net), .I1(n8660[3]), .I2(n378), .I3(n29411), 
            .O(n8639[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4135_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4118_5_lut (.I0(GND_net), .I1(n8453[2]), .I2(n320), .I3(n29247), 
            .O(n8437[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4118_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_668_20_lut (.I0(GND_net), .I1(n3265[18]), .I2(n3290[18]), 
            .I3(n27988), .O(duty_23__N_3613[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_668_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i69_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral [9]), 
            .I2(GND_net), .I3(GND_net), .O(n101));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i69_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_668_20 (.CI(n27988), .I0(n3265[18]), .I1(n3290[18]), 
            .CO(n27989));
    SB_LUT4 mult_11_i22_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral [10]), 
            .I2(GND_net), .I3(GND_net), .O(n32));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i22_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_add_3_14_lut (.I0(\PID_CONTROLLER.integral [12]), 
            .I1(GND_net), .I2(n1_adj_4332[12]), .I3(n28097), .O(n25_adj_4055)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_14_lut.LUT_INIT = 16'h6996;
    SB_LUT4 add_668_19_lut (.I0(GND_net), .I1(n3265[17]), .I2(n3290[17]), 
            .I3(n27987), .O(duty_23__N_3613[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_668_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4110_6 (.CI(n28718), .I0(n8297[3]), .I1(n369), .CO(n28719));
    SB_LUT4 i31265_3_lut (.I0(n4_adj_4054), .I1(n257[13]), .I2(n27_adj_4058), 
            .I3(GND_net), .O(n37947));   // verilog/motorControl.v(46[19:35])
    defparam i31265_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_4148_5_lut (.I0(GND_net), .I1(n8842[2]), .I2(n344), .I3(n29566), 
            .O(n8834[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4148_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i375_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral [15]), 
            .I2(GND_net), .I3(GND_net), .O(n557_adj_4059));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i375_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_4110_5_lut (.I0(GND_net), .I1(n8297[2]), .I2(n296), .I3(n28717), 
            .O(n8273[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4110_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i424_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral [15]), 
            .I2(GND_net), .I3(GND_net), .O(n630_adj_4060));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i424_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_4110_5 (.CI(n28717), .I0(n8297[2]), .I1(n296), .CO(n28718));
    SB_CARRY add_4118_5 (.CI(n29247), .I0(n8453[2]), .I1(n320), .CO(n29248));
    SB_LUT4 i2_3_lut_4_lut_adj_844 (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral [18]), 
            .I2(n8849[0]), .I3(n27714), .O(n8842[1]));   // verilog/motorControl.v(42[26:37])
    defparam i2_3_lut_4_lut_adj_844.LUT_INIT = 16'h8778;
    SB_LUT4 add_4110_4_lut (.I0(GND_net), .I1(n8297[1]), .I2(n223), .I3(n28716), 
            .O(n8273[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4110_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4148_5 (.CI(n29566), .I0(n8842[2]), .I1(n344), .CO(n29567));
    SB_CARRY add_4110_4 (.CI(n28716), .I0(n8297[1]), .I1(n223), .CO(n28717));
    SB_LUT4 add_4110_3_lut (.I0(GND_net), .I1(n8297[0]), .I2(n150), .I3(n28715), 
            .O(n8273[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4110_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4118_4_lut (.I0(GND_net), .I1(n8453[1]), .I2(n247), .I3(n29246), 
            .O(n8437[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4118_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4135_6 (.CI(n29411), .I0(n8660[3]), .I1(n378), .CO(n29412));
    SB_LUT4 add_4135_5_lut (.I0(GND_net), .I1(n8660[2]), .I2(n305), .I3(n29410), 
            .O(n8639[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4135_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i22910_3_lut_4_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral [18]), 
            .I2(n27714), .I3(n8849[0]), .O(n4_adj_4045));   // verilog/motorControl.v(42[26:37])
    defparam i22910_3_lut_4_lut.LUT_INIT = 16'hf880;
    SB_CARRY add_4118_4 (.CI(n29246), .I0(n8453[1]), .I1(n247), .CO(n29247));
    SB_LUT4 mult_10_i183_2_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err [17]), 
            .I2(GND_net), .I3(GND_net), .O(n271_adj_4061));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i183_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_4135_5 (.CI(n29410), .I0(n8660[2]), .I1(n305), .CO(n29411));
    SB_CARRY add_4110_3 (.CI(n28715), .I0(n8297[0]), .I1(n150), .CO(n28716));
    SB_LUT4 add_4148_4_lut (.I0(GND_net), .I1(n8842[1]), .I2(n271_adj_4062), 
            .I3(n29565), .O(n8834[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4148_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4148_4 (.CI(n29565), .I0(n8842[1]), .I1(n271_adj_4062), 
            .CO(n29566));
    SB_LUT4 add_4135_4_lut (.I0(GND_net), .I1(n8660[1]), .I2(n232), .I3(n29409), 
            .O(n8639[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4135_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4118_3_lut (.I0(GND_net), .I1(n8453[0]), .I2(n174), .I3(n29245), 
            .O(n8437[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4118_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i22897_2_lut_3_lut_4_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral [19]), 
            .I2(\PID_CONTROLLER.integral [18]), .I3(\Ki[1] ), .O(n8842[0]));   // verilog/motorControl.v(42[26:37])
    defparam i22897_2_lut_3_lut_4_lut.LUT_INIT = 16'h7888;
    SB_CARRY add_4118_3 (.CI(n29245), .I0(n8453[0]), .I1(n174), .CO(n29246));
    SB_LUT4 add_4118_2_lut (.I0(GND_net), .I1(n32_adj_4063), .I2(n101_adj_4064), 
            .I3(GND_net), .O(n8437[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4118_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i643_2_lut (.I0(\Kp[13] ), .I1(\PID_CONTROLLER.err [2]), 
            .I2(GND_net), .I3(GND_net), .O(n956_adj_4065));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i643_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_4118_2 (.CI(GND_net), .I0(n32_adj_4063), .I1(n101_adj_4064), 
            .CO(n29245));
    SB_CARRY add_4135_4 (.CI(n29409), .I0(n8660[1]), .I1(n232), .CO(n29410));
    SB_LUT4 unary_minus_16_inv_0_i15_1_lut (.I0(PWMLimit[14]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[14]));   // verilog/motorControl.v(47[19:28])
    defparam unary_minus_16_inv_0_i15_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_4148_3_lut (.I0(GND_net), .I1(n8842[0]), .I2(n198_adj_4067), 
            .I3(n29564), .O(n8834[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4148_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4135_3_lut (.I0(GND_net), .I1(n8660[0]), .I2(n159), .I3(n29408), 
            .O(n8639[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4135_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4135_3 (.CI(n29408), .I0(n8660[0]), .I1(n159), .CO(n29409));
    SB_LUT4 add_4135_2_lut (.I0(GND_net), .I1(n17_adj_4068), .I2(n86), 
            .I3(GND_net), .O(n8639[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4135_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4135_2 (.CI(GND_net), .I0(n17_adj_4068), .I1(n86), .CO(n29408));
    SB_LUT4 i22899_2_lut_3_lut_4_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral [19]), 
            .I2(\PID_CONTROLLER.integral [18]), .I3(\Ki[1] ), .O(n27714));   // verilog/motorControl.v(42[26:37])
    defparam i22899_2_lut_3_lut_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 add_4110_2_lut (.I0(GND_net), .I1(n8_adj_4069), .I2(n77), 
            .I3(GND_net), .O(n8273[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4110_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i232_2_lut (.I0(\Kp[4] ), .I1(\PID_CONTROLLER.err [17]), 
            .I2(GND_net), .I3(GND_net), .O(n344_adj_4070));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i232_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i31266_3_lut (.I0(n37947), .I1(n257[14]), .I2(n29_adj_4071), 
            .I3(GND_net), .O(n37948));   // verilog/motorControl.v(46[19:35])
    defparam i31266_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_10_i692_2_lut (.I0(\Kp[14] ), .I1(\PID_CONTROLLER.err [2]), 
            .I2(GND_net), .I3(GND_net), .O(n1029_adj_4072));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i692_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i30771_4_lut (.I0(n33_adj_4004), .I1(n31_adj_4073), .I2(n29_adj_4071), 
            .I3(n37456), .O(n37452));
    defparam i30771_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 mult_11_i118_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral [9]), 
            .I2(GND_net), .I3(GND_net), .O(n174_adj_4074));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i118_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i31429_4_lut (.I0(n30_adj_4075), .I1(n10_adj_4076), .I2(n35_adj_4003), 
            .I3(n37446), .O(n38111));   // verilog/motorControl.v(46[19:35])
    defparam i31429_4_lut.LUT_INIT = 16'haaac;
    SB_CARRY unary_minus_5_add_3_14 (.CI(n28097), .I0(GND_net), .I1(n1_adj_4332[12]), 
            .CO(n28098));
    SB_LUT4 i22938_2_lut_3_lut_4_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral [20]), 
            .I2(\PID_CONTROLLER.integral [19]), .I3(\Ki[1] ), .O(n27757));   // verilog/motorControl.v(42[26:37])
    defparam i22938_2_lut_3_lut_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i31074_3_lut (.I0(n37948), .I1(n257[15]), .I2(n31_adj_4073), 
            .I3(GND_net), .O(n37756));   // verilog/motorControl.v(46[19:35])
    defparam i31074_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_10_i557_2_lut (.I0(\Kp[11] ), .I1(\PID_CONTROLLER.err [8]), 
            .I2(GND_net), .I3(GND_net), .O(n828_adj_4077));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i557_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_inv_0_i8_1_lut (.I0(IntegralLimit[7]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4332[7]));   // verilog/motorControl.v(39[48:62])
    defparam unary_minus_5_inv_0_i8_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_16_inv_0_i16_1_lut (.I0(PWMLimit[15]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[15]));   // verilog/motorControl.v(47[19:28])
    defparam unary_minus_16_inv_0_i16_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i22936_2_lut_3_lut_4_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral [20]), 
            .I2(\PID_CONTROLLER.integral [19]), .I3(\Ki[1] ), .O(n8849[0]));   // verilog/motorControl.v(42[26:37])
    defparam i22936_2_lut_3_lut_4_lut.LUT_INIT = 16'h7888;
    SB_LUT4 mult_10_i741_2_lut (.I0(\Kp[15] ), .I1(\PID_CONTROLLER.err [2]), 
            .I2(GND_net), .I3(GND_net), .O(n1102_adj_4080));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i741_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i281_2_lut (.I0(\Kp[5] ), .I1(\PID_CONTROLLER.err [17]), 
            .I2(GND_net), .I3(GND_net), .O(n417_adj_4081));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i281_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i2_4_lut (.I0(n6_adj_4082), .I1(\Kp[4] ), .I2(n8552[2]), .I3(\PID_CONTROLLER.err [18]), 
            .O(n8545[3]));   // verilog/motorControl.v(42[17:23])
    defparam i2_4_lut.LUT_INIT = 16'h965a;
    SB_LUT4 i31461_4_lut (.I0(n37756), .I1(n38111), .I2(n35_adj_4003), 
            .I3(n37452), .O(n38143));   // verilog/motorControl.v(46[19:35])
    defparam i31461_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i31462_3_lut (.I0(n38143), .I1(n257[18]), .I2(n37_adj_4002), 
            .I3(GND_net), .O(n38144));   // verilog/motorControl.v(46[19:35])
    defparam i31462_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i31452_3_lut (.I0(n38144), .I1(n257[19]), .I2(n39_adj_4084), 
            .I3(GND_net), .O(n38134));   // verilog/motorControl.v(46[19:35])
    defparam i31452_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_4110_2 (.CI(GND_net), .I0(n8_adj_4069), .I1(n77), .CO(n28715));
    SB_CARRY add_4148_3 (.CI(n29564), .I0(n8842[0]), .I1(n198_adj_4067), 
            .CO(n29565));
    SB_LUT4 unary_minus_5_add_3_13_lut (.I0(\PID_CONTROLLER.integral [11]), 
            .I1(GND_net), .I2(n1_adj_4332[11]), .I3(n28096), .O(n23_adj_4085)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_13_lut.LUT_INIT = 16'h6996;
    SB_LUT4 add_4148_2_lut (.I0(GND_net), .I1(n56_adj_4087), .I2(n125_adj_4088), 
            .I3(GND_net), .O(n8834[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4148_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_668_19 (.CI(n27987), .I0(n3265[17]), .I1(n3290[17]), 
            .CO(n27988));
    SB_CARRY add_4148_2 (.CI(GND_net), .I0(n56_adj_4087), .I1(n125_adj_4088), 
            .CO(n29564));
    SB_LUT4 add_668_18_lut (.I0(GND_net), .I1(n3265[16]), .I2(n3290[16]), 
            .I3(n27986), .O(duty_23__N_3613[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_668_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4117_16_lut (.I0(GND_net), .I1(n8437[13]), .I2(n1120_adj_4089), 
            .I3(n29244), .O(n8420[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4117_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4134_21_lut (.I0(GND_net), .I1(n8639[18]), .I2(GND_net), 
            .I3(n29407), .O(n8617[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4134_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4117_15_lut (.I0(GND_net), .I1(n8437[12]), .I2(n1047_adj_4090), 
            .I3(n29243), .O(n8420[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4117_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4147_8_lut (.I0(GND_net), .I1(n8834[5]), .I2(n560_adj_4091), 
            .I3(n29563), .O(n8825[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4147_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_668_18 (.CI(n27986), .I0(n3265[16]), .I1(n3290[16]), 
            .CO(n27987));
    SB_LUT4 add_4147_7_lut (.I0(GND_net), .I1(n8834[4]), .I2(n487_adj_4092), 
            .I3(n29562), .O(n8825[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4147_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4147_7 (.CI(n29562), .I0(n8834[4]), .I1(n487_adj_4092), 
            .CO(n29563));
    SB_LUT4 add_4147_6_lut (.I0(GND_net), .I1(n8834[3]), .I2(n414_adj_4093), 
            .I3(n29561), .O(n8825[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4147_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4134_20_lut (.I0(GND_net), .I1(n8639[17]), .I2(GND_net), 
            .I3(n29406), .O(n8617[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4134_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i83_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral [16]), 
            .I2(GND_net), .I3(GND_net), .O(n122_adj_4094));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i83_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i2_3_lut_4_lut_adj_845 (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral [19]), 
            .I2(n8855[0]), .I3(n27757), .O(n8849[1]));   // verilog/motorControl.v(42[26:37])
    defparam i2_3_lut_4_lut_adj_845.LUT_INIT = 16'h8778;
    SB_LUT4 i22949_3_lut_4_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral [19]), 
            .I2(n27757), .I3(n8855[0]), .O(n4_adj_4095));   // verilog/motorControl.v(42[26:37])
    defparam i22949_3_lut_4_lut.LUT_INIT = 16'hf880;
    SB_LUT4 i22967_2_lut_3_lut_4_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral [21]), 
            .I2(\PID_CONTROLLER.integral [20]), .I3(\Ki[1] ), .O(n8855[0]));   // verilog/motorControl.v(42[26:37])
    defparam i22967_2_lut_3_lut_4_lut.LUT_INIT = 16'h7888;
    SB_LUT4 i22969_2_lut_3_lut_4_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral [21]), 
            .I2(\PID_CONTROLLER.integral [20]), .I3(\Ki[1] ), .O(n27791));   // verilog/motorControl.v(42[26:37])
    defparam i22969_2_lut_3_lut_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i22980_3_lut_4_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral [20]), 
            .I2(n27791), .I3(n8860[0]), .O(n4_adj_4096));   // verilog/motorControl.v(42[26:37])
    defparam i22980_3_lut_4_lut.LUT_INIT = 16'hf880;
    SB_CARRY add_4117_15 (.CI(n29243), .I0(n8437[12]), .I1(n1047_adj_4090), 
            .CO(n29244));
    SB_LUT4 mult_10_i138_2_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err [19]), 
            .I2(GND_net), .I3(GND_net), .O(n204));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i138_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i2_3_lut_4_lut_adj_846 (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral [20]), 
            .I2(n8860[0]), .I3(n27791), .O(n8855[1]));   // verilog/motorControl.v(42[26:37])
    defparam i2_3_lut_4_lut_adj_846.LUT_INIT = 16'h8778;
    SB_CARRY add_4134_20 (.CI(n29406), .I0(n8639[17]), .I1(GND_net), .CO(n29407));
    SB_LUT4 i22830_4_lut (.I0(\Kp[0] ), .I1(\Kp[1] ), .I2(\PID_CONTROLLER.err [22]), 
            .I3(\PID_CONTROLLER.err [21]), .O(n8563[0]));   // verilog/motorControl.v(42[17:23])
    defparam i22830_4_lut.LUT_INIT = 16'h6ca0;
    SB_LUT4 add_4134_19_lut (.I0(GND_net), .I1(n8639[16]), .I2(GND_net), 
            .I3(n29405), .O(n8617[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4134_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4147_6 (.CI(n29561), .I0(n8834[3]), .I1(n414_adj_4093), 
            .CO(n29562));
    SB_LUT4 add_4147_5_lut (.I0(GND_net), .I1(n8834[2]), .I2(n341_adj_4097), 
            .I3(n29560), .O(n8825[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4147_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_5_add_3_13 (.CI(n28096), .I0(GND_net), .I1(n1_adj_4332[11]), 
            .CO(n28097));
    SB_LUT4 add_4117_14_lut (.I0(GND_net), .I1(n8437[11]), .I2(n974_adj_4098), 
            .I3(n29242), .O(n8420[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4117_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4147_5 (.CI(n29560), .I0(n8834[2]), .I1(n341_adj_4097), 
            .CO(n29561));
    SB_CARRY add_4134_19 (.CI(n29405), .I0(n8639[16]), .I1(GND_net), .CO(n29406));
    SB_LUT4 add_4147_4_lut (.I0(GND_net), .I1(n8834[1]), .I2(n268_adj_4099), 
            .I3(n29559), .O(n8825[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4147_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4134_18_lut (.I0(GND_net), .I1(n8639[15]), .I2(GND_net), 
            .I3(n29404), .O(n8617[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4134_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4117_14 (.CI(n29242), .I0(n8437[11]), .I1(n974_adj_4098), 
            .CO(n29243));
    SB_CARRY add_4147_4 (.CI(n29559), .I0(n8834[1]), .I1(n268_adj_4099), 
            .CO(n29560));
    SB_LUT4 unary_minus_5_add_3_12_lut (.I0(\PID_CONTROLLER.integral [10]), 
            .I1(GND_net), .I2(n1_adj_4332[10]), .I3(n28095), .O(n21_adj_4100)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_12_lut.LUT_INIT = 16'h6996;
    SB_CARRY add_4134_18 (.CI(n29404), .I0(n8639[15]), .I1(GND_net), .CO(n29405));
    SB_CARRY unary_minus_5_add_3_12 (.CI(n28095), .I0(GND_net), .I1(n1_adj_4332[10]), 
            .CO(n28096));
    SB_LUT4 add_4117_13_lut (.I0(GND_net), .I1(n8437[10]), .I2(n901_adj_4102), 
            .I3(n29241), .O(n8420[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4117_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_5_add_3_11_lut (.I0(\PID_CONTROLLER.integral [9]), 
            .I1(GND_net), .I2(n1_adj_4332[9]), .I3(n28094), .O(n19_adj_4103)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_11_lut.LUT_INIT = 16'h6996;
    SB_CARRY unary_minus_5_add_3_11 (.CI(n28094), .I0(GND_net), .I1(n1_adj_4332[9]), 
            .CO(n28095));
    SB_LUT4 unary_minus_5_add_3_10_lut (.I0(\PID_CONTROLLER.integral [8]), 
            .I1(GND_net), .I2(n1_adj_4332[8]), .I3(n28093), .O(n17_adj_4105)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_10_lut.LUT_INIT = 16'h6996;
    SB_LUT4 add_4147_3_lut (.I0(GND_net), .I1(n8834[0]), .I2(n195_adj_4107), 
            .I3(n29558), .O(n8825[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4147_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4134_17_lut (.I0(GND_net), .I1(n8639[14]), .I2(GND_net), 
            .I3(n29403), .O(n8617[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4134_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4117_13 (.CI(n29241), .I0(n8437[10]), .I1(n901_adj_4102), 
            .CO(n29242));
    SB_CARRY unary_minus_5_add_3_10 (.CI(n28093), .I0(GND_net), .I1(n1_adj_4332[8]), 
            .CO(n28094));
    SB_CARRY add_4147_3 (.CI(n29558), .I0(n8834[0]), .I1(n195_adj_4107), 
            .CO(n29559));
    SB_LUT4 add_4147_2_lut (.I0(GND_net), .I1(n53_adj_4108), .I2(n122_adj_4094), 
            .I3(GND_net), .O(n8825[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4147_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i89_2_lut (.I0(\Kp[1] ), .I1(\PID_CONTROLLER.err [19]), 
            .I2(GND_net), .I3(GND_net), .O(n131));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i89_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_add_3_9_lut (.I0(\PID_CONTROLLER.integral [7]), 
            .I1(GND_net), .I2(n1_adj_4332[7]), .I3(n28092), .O(n15_adj_4109)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_9_lut.LUT_INIT = 16'h6996;
    SB_CARRY add_4134_17 (.CI(n29403), .I0(n8639[14]), .I1(GND_net), .CO(n29404));
    SB_LUT4 add_4117_12_lut (.I0(GND_net), .I1(n8437[9]), .I2(n828_adj_4077), 
            .I3(n29240), .O(n8420[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4117_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4147_2 (.CI(GND_net), .I0(n53_adj_4108), .I1(n122_adj_4094), 
            .CO(n29558));
    SB_LUT4 add_4146_9_lut (.I0(GND_net), .I1(n8825[6]), .I2(n630_adj_4060), 
            .I3(n29557), .O(n8815[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4146_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4146_8_lut (.I0(GND_net), .I1(n8825[5]), .I2(n557_adj_4059), 
            .I3(n29556), .O(n8815[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4146_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4117_12 (.CI(n29240), .I0(n8437[9]), .I1(n828_adj_4077), 
            .CO(n29241));
    SB_LUT4 mult_10_i42_2_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err [20]), 
            .I2(GND_net), .I3(GND_net), .O(n62));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i42_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_668_17_lut (.I0(GND_net), .I1(n3265[15]), .I2(n3290[15]), 
            .I3(n27985), .O(duty_23__N_3613[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_668_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4146_8 (.CI(n29556), .I0(n8825[5]), .I1(n557_adj_4059), 
            .CO(n29557));
    SB_CARRY unary_minus_5_add_3_9 (.CI(n28092), .I0(GND_net), .I1(n1_adj_4332[7]), 
            .CO(n28093));
    SB_LUT4 unary_minus_5_add_3_8_lut (.I0(\PID_CONTROLLER.integral [6]), 
            .I1(GND_net), .I2(n1_adj_4332[6]), .I3(n28091), .O(n13_adj_4110)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_8_lut.LUT_INIT = 16'h6996;
    SB_LUT4 add_4117_11_lut (.I0(GND_net), .I1(n8437[8]), .I2(n755_adj_4042), 
            .I3(n29239), .O(n8420[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4117_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4117_11 (.CI(n29239), .I0(n8437[8]), .I1(n755_adj_4042), 
            .CO(n29240));
    SB_LUT4 mult_11_i36_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral [17]), 
            .I2(GND_net), .I3(GND_net), .O(n53_adj_4108));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i36_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_4117_10_lut (.I0(GND_net), .I1(n8437[7]), .I2(n682_adj_4041), 
            .I3(n29238), .O(n8420[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4117_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4146_7_lut (.I0(GND_net), .I1(n8825[4]), .I2(n484_adj_4040), 
            .I3(n29555), .O(n8815[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4146_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4134_16_lut (.I0(GND_net), .I1(n8639[13]), .I2(n1105), 
            .I3(n29402), .O(n8617[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4134_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4117_10 (.CI(n29238), .I0(n8437[7]), .I1(n682_adj_4041), 
            .CO(n29239));
    SB_LUT4 i2_4_lut_adj_847 (.I0(n4_adj_4111), .I1(\Kp[3] ), .I2(n8558[1]), 
            .I3(\PID_CONTROLLER.err [19]), .O(n8552[2]));   // verilog/motorControl.v(42[17:23])
    defparam i2_4_lut_adj_847.LUT_INIT = 16'h965a;
    SB_LUT4 mult_10_i330_2_lut (.I0(\Kp[6] ), .I1(\PID_CONTROLLER.err [17]), 
            .I2(GND_net), .I3(GND_net), .O(n490_adj_4112));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i330_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i2_4_lut_adj_848 (.I0(\Kp[0] ), .I1(\Kp[3] ), .I2(\PID_CONTROLLER.err [23]), 
            .I3(\PID_CONTROLLER.err [20]), .O(n12_adj_4113));   // verilog/motorControl.v(42[17:23])
    defparam i2_4_lut_adj_848.LUT_INIT = 16'h9c50;
    SB_LUT4 add_4117_9_lut (.I0(GND_net), .I1(n8437[6]), .I2(n609_adj_4033), 
            .I3(n29237), .O(n8420[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4117_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_668_17 (.CI(n27985), .I0(n3265[15]), .I1(n3290[15]), 
            .CO(n27986));
    SB_LUT4 i22766_4_lut (.I0(n8552[2]), .I1(\Kp[4] ), .I2(n6_adj_4082), 
            .I3(\PID_CONTROLLER.err [18]), .O(n8_adj_4114));   // verilog/motorControl.v(42[17:23])
    defparam i22766_4_lut.LUT_INIT = 16'he8a0;
    SB_CARRY add_4146_7 (.CI(n29555), .I0(n8825[4]), .I1(n484_adj_4040), 
            .CO(n29556));
    SB_LUT4 i1_4_lut (.I0(\Kp[4] ), .I1(\Kp[2] ), .I2(\PID_CONTROLLER.err [19]), 
            .I3(\PID_CONTROLLER.err [21]), .O(n11_adj_4115));   // verilog/motorControl.v(42[17:23])
    defparam i1_4_lut.LUT_INIT = 16'h6ca0;
    SB_LUT4 add_4146_6_lut (.I0(GND_net), .I1(n8825[3]), .I2(n411_adj_4031), 
            .I3(n29554), .O(n8815[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4146_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4146_6 (.CI(n29554), .I0(n8825[3]), .I1(n411_adj_4031), 
            .CO(n29555));
    SB_CARRY add_4134_16 (.CI(n29402), .I0(n8639[13]), .I1(n1105), .CO(n29403));
    SB_CARRY add_4117_9 (.CI(n29237), .I0(n8437[6]), .I1(n609_adj_4033), 
            .CO(n29238));
    SB_LUT4 add_4146_5_lut (.I0(GND_net), .I1(n8825[2]), .I2(n338_adj_4030), 
            .I3(n29553), .O(n8815[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4146_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4117_8_lut (.I0(GND_net), .I1(n8437[5]), .I2(n536_adj_4029), 
            .I3(n29236), .O(n8420[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4117_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4146_5 (.CI(n29553), .I0(n8825[2]), .I1(n338_adj_4030), 
            .CO(n29554));
    SB_LUT4 add_4146_4_lut (.I0(GND_net), .I1(n8825[1]), .I2(n265_adj_4027), 
            .I3(n29552), .O(n8815[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4146_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4134_15_lut (.I0(GND_net), .I1(n8639[12]), .I2(n1032), 
            .I3(n29401), .O(n8617[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4134_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i22797_4_lut (.I0(n8558[1]), .I1(\Kp[3] ), .I2(n4_adj_4111), 
            .I3(\PID_CONTROLLER.err [19]), .O(n6_adj_4116));   // verilog/motorControl.v(42[17:23])
    defparam i22797_4_lut.LUT_INIT = 16'he8a0;
    SB_CARRY add_4146_4 (.CI(n29552), .I0(n8825[1]), .I1(n265_adj_4027), 
            .CO(n29553));
    SB_LUT4 i22832_4_lut (.I0(\Kp[0] ), .I1(\Kp[1] ), .I2(\PID_CONTROLLER.err [22]), 
            .I3(\PID_CONTROLLER.err [21]), .O(n27646));   // verilog/motorControl.v(42[17:23])
    defparam i22832_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 mult_11_i132_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral [16]), 
            .I2(GND_net), .I3(GND_net), .O(n195_adj_4107));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i132_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i8_4_lut (.I0(n6_adj_4116), .I1(n11_adj_4115), .I2(n8_adj_4114), 
            .I3(n12_adj_4113), .O(n18_adj_4117));   // verilog/motorControl.v(42[17:23])
    defparam i8_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 unary_minus_5_inv_0_i9_1_lut (.I0(IntegralLimit[8]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4332[8]));   // verilog/motorControl.v(39[48:62])
    defparam unary_minus_5_inv_0_i9_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i3_4_lut (.I0(\Kp[5] ), .I1(\Kp[1] ), .I2(\PID_CONTROLLER.err [18]), 
            .I3(\PID_CONTROLLER.err [22]), .O(n13_adj_4118));   // verilog/motorControl.v(42[17:23])
    defparam i3_4_lut.LUT_INIT = 16'h6ca0;
    SB_LUT4 i9_4_lut (.I0(n13_adj_4118), .I1(n18_adj_4117), .I2(n27646), 
            .I3(n4_adj_4119), .O(n34771));   // verilog/motorControl.v(42[17:23])
    defparam i9_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 add_4146_3_lut (.I0(GND_net), .I1(n8825[0]), .I2(n192_adj_4022), 
            .I3(n29551), .O(n8815[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4146_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4134_15 (.CI(n29401), .I0(n8639[12]), .I1(n1032), .CO(n29402));
    SB_CARRY add_4117_8 (.CI(n29236), .I0(n8437[5]), .I1(n536_adj_4029), 
            .CO(n29237));
    SB_LUT4 add_4134_14_lut (.I0(GND_net), .I1(n8639[11]), .I2(n959), 
            .I3(n29400), .O(n8617[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4134_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_5_inv_0_i10_1_lut (.I0(IntegralLimit[9]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4332[9]));   // verilog/motorControl.v(39[48:62])
    defparam unary_minus_5_inv_0_i10_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_668_16_lut (.I0(GND_net), .I1(n3265[14]), .I2(n3290[14]), 
            .I3(n27984), .O(duty_23__N_3613[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_668_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_668_16 (.CI(n27984), .I0(n3265[14]), .I1(n3290[14]), 
            .CO(n27985));
    SB_CARRY add_4134_14 (.CI(n29400), .I0(n8639[11]), .I1(n959), .CO(n29401));
    SB_LUT4 add_4117_7_lut (.I0(GND_net), .I1(n8437[4]), .I2(n463_adj_4017), 
            .I3(n29235), .O(n8420[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4117_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i606_2_lut (.I0(\Kp[12] ), .I1(\PID_CONTROLLER.err [8]), 
            .I2(GND_net), .I3(GND_net), .O(n901_adj_4102));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i606_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_inv_0_i11_1_lut (.I0(IntegralLimit[10]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4332[10]));   // verilog/motorControl.v(39[48:62])
    defparam unary_minus_5_inv_0_i11_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_11_i181_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral [16]), 
            .I2(GND_net), .I3(GND_net), .O(n268_adj_4099));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i181_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i53_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral [1]), 
            .I2(GND_net), .I3(GND_net), .O(n77_adj_4120));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i53_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i6_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral [2]), 
            .I2(GND_net), .I3(GND_net), .O(n8_adj_4121));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i6_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_4146_3 (.CI(n29551), .I0(n8825[0]), .I1(n192_adj_4022), 
            .CO(n29552));
    SB_LUT4 mult_11_i167_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral [9]), 
            .I2(GND_net), .I3(GND_net), .O(n247_adj_4122));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i167_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_16_inv_0_i17_1_lut (.I0(PWMLimit[16]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[16]));   // verilog/motorControl.v(47[19:28])
    defparam unary_minus_16_inv_0_i17_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i19586_2_lut_2_lut (.I0(n256), .I1(n7788[0]), .I2(GND_net), 
            .I3(GND_net), .O(n3265[23]));   // verilog/motorControl.v(46[19:35])
    defparam i19586_2_lut_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 unary_minus_16_inv_0_i18_1_lut (.I0(PWMLimit[17]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[17]));   // verilog/motorControl.v(47[19:28])
    defparam unary_minus_16_inv_0_i18_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_11_i102_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral [1]), 
            .I2(GND_net), .I3(GND_net), .O(n150_adj_4125));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i102_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i57_2_lut (.I0(\Kp[1] ), .I1(\PID_CONTROLLER.err [3]), 
            .I2(GND_net), .I3(GND_net), .O(n83_adj_4126));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i57_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i10_2_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err [4]), 
            .I2(GND_net), .I3(GND_net), .O(n14_adj_4127));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i10_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i151_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral [1]), 
            .I2(GND_net), .I3(GND_net), .O(n223_adj_4128));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i151_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i216_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral [9]), 
            .I2(GND_net), .I3(GND_net), .O(n320_adj_4129));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i216_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_16_inv_0_i19_1_lut (.I0(PWMLimit[18]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[18]));   // verilog/motorControl.v(47[19:28])
    defparam unary_minus_16_inv_0_i19_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i106_2_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err [3]), 
            .I2(GND_net), .I3(GND_net), .O(n156_adj_4131));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i106_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i265_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral [9]), 
            .I2(GND_net), .I3(GND_net), .O(n393_adj_4132));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i265_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i655_2_lut (.I0(\Kp[13] ), .I1(\PID_CONTROLLER.err [8]), 
            .I2(GND_net), .I3(GND_net), .O(n974_adj_4098));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i655_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i230_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral [16]), 
            .I2(GND_net), .I3(GND_net), .O(n341_adj_4097));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i230_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i200_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral [1]), 
            .I2(GND_net), .I3(GND_net), .O(n296_adj_4133));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i200_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i561_2_lut (.I0(\Kp[11] ), .I1(\PID_CONTROLLER.err [10]), 
            .I2(GND_net), .I3(GND_net), .O(n834));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i561_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i610_2_lut (.I0(\Kp[12] ), .I1(\PID_CONTROLLER.err [10]), 
            .I2(GND_net), .I3(GND_net), .O(n907));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i610_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i155_2_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err [3]), 
            .I2(GND_net), .I3(GND_net), .O(n229_adj_4134));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i155_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i600_2_lut (.I0(\Ki[12] ), .I1(\PID_CONTROLLER.integral [5]), 
            .I2(GND_net), .I3(GND_net), .O(n892));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i600_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i204_2_lut (.I0(\Kp[4] ), .I1(\PID_CONTROLLER.err [3]), 
            .I2(GND_net), .I3(GND_net), .O(n302_adj_4135));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i204_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i249_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral [1]), 
            .I2(GND_net), .I3(GND_net), .O(n369_adj_4136));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i249_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i314_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral [9]), 
            .I2(GND_net), .I3(GND_net), .O(n466_adj_4137));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i314_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_16_inv_0_i20_1_lut (.I0(PWMLimit[19]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[19]));   // verilog/motorControl.v(47[19:28])
    defparam unary_minus_16_inv_0_i20_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i30746_4_lut (.I0(n43_adj_4005), .I1(n41_adj_4139), .I2(n39_adj_4084), 
            .I3(n38095), .O(n37427));
    defparam i30746_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 mult_11_i649_2_lut (.I0(\Ki[13] ), .I1(\PID_CONTROLLER.integral [5]), 
            .I2(GND_net), .I3(GND_net), .O(n965));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i649_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i253_2_lut (.I0(\Kp[5] ), .I1(\PID_CONTROLLER.err [3]), 
            .I2(GND_net), .I3(GND_net), .O(n375_adj_4140));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i253_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i298_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral [1]), 
            .I2(GND_net), .I3(GND_net), .O(n442_adj_4141));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i298_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i347_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral [1]), 
            .I2(GND_net), .I3(GND_net), .O(n515_adj_4142));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i347_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i302_2_lut (.I0(\Kp[6] ), .I1(\PID_CONTROLLER.err [3]), 
            .I2(GND_net), .I3(GND_net), .O(n448_adj_4143));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i302_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i363_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral [9]), 
            .I2(GND_net), .I3(GND_net), .O(n539_adj_4144));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i363_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_16_inv_0_i21_1_lut (.I0(PWMLimit[20]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[20]));   // verilog/motorControl.v(47[19:28])
    defparam unary_minus_16_inv_0_i21_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i351_2_lut (.I0(\Kp[7] ), .I1(\PID_CONTROLLER.err [3]), 
            .I2(GND_net), .I3(GND_net), .O(n521_adj_4146));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i351_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i31377_4_lut (.I0(n37754), .I1(n37931), .I2(n45_adj_4038), 
            .I3(n37425), .O(n38059));   // verilog/motorControl.v(46[19:35])
    defparam i31377_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 mult_11_i396_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral [1]), 
            .I2(GND_net), .I3(GND_net), .O(n588_adj_4147));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i396_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i400_2_lut (.I0(\Kp[8] ), .I1(\PID_CONTROLLER.err [3]), 
            .I2(GND_net), .I3(GND_net), .O(n594_adj_4148));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i400_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i412_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral [9]), 
            .I2(GND_net), .I3(GND_net), .O(n612_adj_4149));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i412_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i31434_3_lut (.I0(n38134), .I1(n257[20]), .I2(n41_adj_4139), 
            .I3(GND_net), .O(n40));   // verilog/motorControl.v(46[19:35])
    defparam i31434_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_10_i449_2_lut (.I0(\Kp[9] ), .I1(\PID_CONTROLLER.err [3]), 
            .I2(GND_net), .I3(GND_net), .O(n667_adj_4150));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i449_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i445_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral [1]), 
            .I2(GND_net), .I3(GND_net), .O(n661_adj_4151));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i445_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i498_2_lut (.I0(\Kp[10] ), .I1(\PID_CONTROLLER.err [3]), 
            .I2(GND_net), .I3(GND_net), .O(n740_adj_4152));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i498_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i494_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral [1]), 
            .I2(GND_net), .I3(GND_net), .O(n734_adj_4153));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i494_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i659_2_lut (.I0(\Kp[13] ), .I1(\PID_CONTROLLER.err [10]), 
            .I2(GND_net), .I3(GND_net), .O(n980));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i659_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i461_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral [9]), 
            .I2(GND_net), .I3(GND_net), .O(n685_adj_4154));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i461_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i698_2_lut (.I0(\Ki[14] ), .I1(\PID_CONTROLLER.integral [5]), 
            .I2(GND_net), .I3(GND_net), .O(n1038));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i698_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i547_2_lut (.I0(\Kp[11] ), .I1(\PID_CONTROLLER.err [3]), 
            .I2(GND_net), .I3(GND_net), .O(n813_adj_4155));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i547_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_inv_0_i21_1_lut (.I0(IntegralLimit[20]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4332[20]));   // verilog/motorControl.v(39[48:62])
    defparam unary_minus_5_inv_0_i21_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i596_2_lut (.I0(\Kp[12] ), .I1(\PID_CONTROLLER.err [3]), 
            .I2(GND_net), .I3(GND_net), .O(n886_adj_4156));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i596_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i543_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral [1]), 
            .I2(GND_net), .I3(GND_net), .O(n807_adj_4157));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i543_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i100_2_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err [0]), 
            .I2(GND_net), .I3(GND_net), .O(n147));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i100_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i645_2_lut (.I0(\Kp[13] ), .I1(\PID_CONTROLLER.err [3]), 
            .I2(GND_net), .I3(GND_net), .O(n959_adj_4158));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i645_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i592_2_lut (.I0(\Ki[12] ), .I1(\PID_CONTROLLER.integral [1]), 
            .I2(GND_net), .I3(GND_net), .O(n880_adj_4159));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i592_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY unary_minus_5_add_3_8 (.CI(n28091), .I0(GND_net), .I1(n1_adj_4332[6]), 
            .CO(n28092));
    SB_LUT4 mult_11_i510_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral [9]), 
            .I2(GND_net), .I3(GND_net), .O(n758_adj_4160));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i510_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i694_2_lut (.I0(\Kp[14] ), .I1(\PID_CONTROLLER.err [3]), 
            .I2(GND_net), .I3(GND_net), .O(n1032_adj_4161));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i694_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i641_2_lut (.I0(\Ki[13] ), .I1(\PID_CONTROLLER.integral [1]), 
            .I2(GND_net), .I3(GND_net), .O(n953_adj_4162));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i641_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i743_2_lut (.I0(\Kp[15] ), .I1(\PID_CONTROLLER.err [3]), 
            .I2(GND_net), .I3(GND_net), .O(n1105_adj_4163));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i743_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i690_2_lut (.I0(\Ki[14] ), .I1(\PID_CONTROLLER.integral [1]), 
            .I2(GND_net), .I3(GND_net), .O(n1026_adj_4164));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i690_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i559_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral [9]), 
            .I2(GND_net), .I3(GND_net), .O(n831_adj_4165));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i559_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i739_2_lut (.I0(\Ki[15] ), .I1(\PID_CONTROLLER.integral [1]), 
            .I2(GND_net), .I3(GND_net), .O(n1099_adj_4166));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i739_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i608_2_lut (.I0(\Ki[12] ), .I1(\PID_CONTROLLER.integral [9]), 
            .I2(GND_net), .I3(GND_net), .O(n904_adj_4167));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i608_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_16_inv_0_i22_1_lut (.I0(PWMLimit[21]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[21]));   // verilog/motorControl.v(47[19:28])
    defparam unary_minus_16_inv_0_i22_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i59_2_lut (.I0(\Kp[1] ), .I1(\PID_CONTROLLER.err [4]), 
            .I2(GND_net), .I3(GND_net), .O(n86_adj_4169));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i59_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i12_2_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err [5]), 
            .I2(GND_net), .I3(GND_net), .O(n17_adj_4170));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i12_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i657_2_lut (.I0(\Ki[13] ), .I1(\PID_CONTROLLER.integral [9]), 
            .I2(GND_net), .I3(GND_net), .O(n977_adj_4171));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i657_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i279_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral [16]), 
            .I2(GND_net), .I3(GND_net), .O(n414_adj_4093));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i279_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i108_2_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err [4]), 
            .I2(GND_net), .I3(GND_net), .O(n159_adj_4172));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i108_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i706_2_lut (.I0(\Ki[14] ), .I1(\PID_CONTROLLER.integral [9]), 
            .I2(GND_net), .I3(GND_net), .O(n1050_adj_4173));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i706_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i157_2_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err [4]), 
            .I2(GND_net), .I3(GND_net), .O(n232_adj_4174));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i157_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i328_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral [16]), 
            .I2(GND_net), .I3(GND_net), .O(n487_adj_4092));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i328_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i206_2_lut (.I0(\Kp[4] ), .I1(\PID_CONTROLLER.err [4]), 
            .I2(GND_net), .I3(GND_net), .O(n305_adj_4175));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i206_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i255_2_lut (.I0(\Kp[5] ), .I1(\PID_CONTROLLER.err [4]), 
            .I2(GND_net), .I3(GND_net), .O(n378_adj_4176));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i255_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i73_2_lut (.I0(\Kp[1] ), .I1(\PID_CONTROLLER.err [11]), 
            .I2(GND_net), .I3(GND_net), .O(n107));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i73_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i26_2_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err [12]), 
            .I2(GND_net), .I3(GND_net), .O(n38));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i26_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i71_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral [10]), 
            .I2(GND_net), .I3(GND_net), .O(n104_adj_4177));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i71_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i24_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral [11]), 
            .I2(GND_net), .I3(GND_net), .O(n35_adj_4178));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i24_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i304_2_lut (.I0(\Kp[6] ), .I1(\PID_CONTROLLER.err [4]), 
            .I2(GND_net), .I3(GND_net), .O(n451_adj_4179));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i304_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i353_2_lut (.I0(\Kp[7] ), .I1(\PID_CONTROLLER.err [4]), 
            .I2(GND_net), .I3(GND_net), .O(n524_adj_4180));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i353_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i120_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral [10]), 
            .I2(GND_net), .I3(GND_net), .O(n177_adj_4181));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i120_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i747_2_lut (.I0(\Ki[15] ), .I1(\PID_CONTROLLER.integral [5]), 
            .I2(GND_net), .I3(GND_net), .O(n1111));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i747_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i51_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral [0]), 
            .I2(GND_net), .I3(GND_net), .O(n74_adj_4182));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i51_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i4_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral [1]), 
            .I2(GND_net), .I3(GND_net), .O(n5_adj_4183));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i4_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i122_2_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err [11]), 
            .I2(GND_net), .I3(GND_net), .O(n180));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i122_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_add_3_7_lut (.I0(\PID_CONTROLLER.integral [5]), 
            .I1(GND_net), .I2(n1_adj_4332[5]), .I3(n28090), .O(n11_adj_4184)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_7_lut.LUT_INIT = 16'h6996;
    SB_LUT4 mult_10_i171_2_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err [11]), 
            .I2(GND_net), .I3(GND_net), .O(n253));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i171_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i220_2_lut (.I0(\Kp[4] ), .I1(\PID_CONTROLLER.err [11]), 
            .I2(GND_net), .I3(GND_net), .O(n326));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i220_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i402_2_lut (.I0(\Kp[8] ), .I1(\PID_CONTROLLER.err [4]), 
            .I2(GND_net), .I3(GND_net), .O(n597_adj_4185));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i402_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i100_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral [0]), 
            .I2(GND_net), .I3(GND_net), .O(n147_adj_4186));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i100_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i451_2_lut (.I0(\Kp[9] ), .I1(\PID_CONTROLLER.err [4]), 
            .I2(GND_net), .I3(GND_net), .O(n670_adj_4187));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i451_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i169_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral [10]), 
            .I2(GND_net), .I3(GND_net), .O(n250_adj_4188));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i169_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i269_2_lut (.I0(\Kp[5] ), .I1(\PID_CONTROLLER.err [11]), 
            .I2(GND_net), .I3(GND_net), .O(n399));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i269_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i149_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral [0]), 
            .I2(GND_net), .I3(GND_net), .O(n220_adj_4189));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i149_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i500_2_lut (.I0(\Kp[10] ), .I1(\PID_CONTROLLER.err [4]), 
            .I2(GND_net), .I3(GND_net), .O(n743_adj_4190));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i500_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i31379_4_lut (.I0(n40), .I1(n38059), .I2(n45_adj_4038), .I3(n37427), 
            .O(n38061));   // verilog/motorControl.v(46[19:35])
    defparam i31379_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 unary_minus_16_inv_0_i23_1_lut (.I0(PWMLimit[22]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[22]));   // verilog/motorControl.v(47[19:28])
    defparam unary_minus_16_inv_0_i23_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_11_i198_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral [0]), 
            .I2(GND_net), .I3(GND_net), .O(n293_adj_4192));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i198_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i218_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral [10]), 
            .I2(GND_net), .I3(GND_net), .O(n323_adj_4193));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i218_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_16_inv_0_i24_1_lut (.I0(PWMLimit[23]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[23]));   // verilog/motorControl.v(47[19:28])
    defparam unary_minus_16_inv_0_i24_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i549_2_lut (.I0(\Kp[11] ), .I1(\PID_CONTROLLER.err [4]), 
            .I2(GND_net), .I3(GND_net), .O(n816_adj_4195));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i549_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i598_2_lut (.I0(\Kp[12] ), .I1(\PID_CONTROLLER.err [4]), 
            .I2(GND_net), .I3(GND_net), .O(n889_adj_4196));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i598_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i247_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral [0]), 
            .I2(GND_net), .I3(GND_net), .O(n366_adj_4197));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i247_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i647_2_lut (.I0(\Kp[13] ), .I1(\PID_CONTROLLER.err [4]), 
            .I2(GND_net), .I3(GND_net), .O(n962_adj_4198));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i647_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i267_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral [10]), 
            .I2(GND_net), .I3(GND_net), .O(n396_adj_4199));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i267_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i296_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral [0]), 
            .I2(GND_net), .I3(GND_net), .O(n439_adj_4200));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i296_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i696_2_lut (.I0(\Kp[14] ), .I1(\PID_CONTROLLER.err [4]), 
            .I2(GND_net), .I3(GND_net), .O(n1035_adj_4201));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i696_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i345_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral [0]), 
            .I2(GND_net), .I3(GND_net), .O(n512_adj_4202));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i345_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i745_2_lut (.I0(\Kp[15] ), .I1(\PID_CONTROLLER.err [4]), 
            .I2(GND_net), .I3(GND_net), .O(n1108_adj_4203));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i745_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i316_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral [10]), 
            .I2(GND_net), .I3(GND_net), .O(n469_adj_4204));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i316_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i365_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral [10]), 
            .I2(GND_net), .I3(GND_net), .O(n542_adj_4205));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i365_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i414_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral [10]), 
            .I2(GND_net), .I3(GND_net), .O(n615_adj_4206));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i414_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i394_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral [0]), 
            .I2(GND_net), .I3(GND_net), .O(n585_adj_4207));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i394_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i463_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral [10]), 
            .I2(GND_net), .I3(GND_net), .O(n688_adj_4208));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i463_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i443_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral [0]), 
            .I2(GND_net), .I3(GND_net), .O(n658_adj_4209));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i443_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i512_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral [10]), 
            .I2(GND_net), .I3(GND_net), .O(n761_adj_4210));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i512_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i61_2_lut (.I0(\Kp[1] ), .I1(\PID_CONTROLLER.err [5]), 
            .I2(GND_net), .I3(GND_net), .O(n89_adj_4211));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i61_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i14_2_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err [6]), 
            .I2(GND_net), .I3(GND_net), .O(n20_adj_4212));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i14_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i110_2_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err [5]), 
            .I2(GND_net), .I3(GND_net), .O(n162_adj_4213));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i110_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i492_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral [0]), 
            .I2(GND_net), .I3(GND_net), .O(n731_adj_4214));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i492_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i159_2_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err [5]), 
            .I2(GND_net), .I3(GND_net), .O(n235_adj_4215));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i159_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i541_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral [0]), 
            .I2(GND_net), .I3(GND_net), .O(n804_adj_4216));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i541_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i469_2_lut (.I0(\Kp[9] ), .I1(\PID_CONTROLLER.err [13]), 
            .I2(GND_net), .I3(GND_net), .O(n697));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i469_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i561_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral [10]), 
            .I2(GND_net), .I3(GND_net), .O(n834_adj_4217));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i561_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i208_2_lut (.I0(\Kp[4] ), .I1(\PID_CONTROLLER.err [5]), 
            .I2(GND_net), .I3(GND_net), .O(n308_adj_4218));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i208_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i590_2_lut (.I0(\Ki[12] ), .I1(\PID_CONTROLLER.integral [0]), 
            .I2(GND_net), .I3(GND_net), .O(n877_adj_4219));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i590_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i610_2_lut (.I0(\Ki[12] ), .I1(\PID_CONTROLLER.integral [10]), 
            .I2(GND_net), .I3(GND_net), .O(n907_adj_4220));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i610_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i257_2_lut (.I0(\Kp[5] ), .I1(\PID_CONTROLLER.err [5]), 
            .I2(GND_net), .I3(GND_net), .O(n381_adj_4221));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i257_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i318_2_lut (.I0(\Kp[6] ), .I1(\PID_CONTROLLER.err [11]), 
            .I2(GND_net), .I3(GND_net), .O(n472));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i318_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_4146_2_lut (.I0(GND_net), .I1(n50), .I2(n119), .I3(GND_net), 
            .O(n8815[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4146_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4134_13_lut (.I0(GND_net), .I1(n8639[10]), .I2(n886), 
            .I3(n29399), .O(n8617[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4134_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4117_7 (.CI(n29235), .I0(n8437[4]), .I1(n463_adj_4017), 
            .CO(n29236));
    SB_CARRY add_4134_13 (.CI(n29399), .I0(n8639[10]), .I1(n886), .CO(n29400));
    SB_LUT4 add_4117_6_lut (.I0(GND_net), .I1(n8437[3]), .I2(n390), .I3(n29234), 
            .O(n8420[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4117_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4146_2 (.CI(GND_net), .I0(n50), .I1(n119), .CO(n29551));
    SB_LUT4 add_4134_12_lut (.I0(GND_net), .I1(n8639[9]), .I2(n813), .I3(n29398), 
            .O(n8617[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4134_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4117_6 (.CI(n29234), .I0(n8437[3]), .I1(n390), .CO(n29235));
    SB_CARRY add_4134_12 (.CI(n29398), .I0(n8639[9]), .I1(n813), .CO(n29399));
    SB_LUT4 add_4117_5_lut (.I0(GND_net), .I1(n8437[2]), .I2(n317_adj_3961), 
            .I3(n29233), .O(n8420[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4117_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i19344_3_lut (.I0(\Kp[0] ), .I1(n256), .I2(\PID_CONTROLLER.err [0]), 
            .I3(GND_net), .O(n3265[0]));   // verilog/motorControl.v(46[16] 48[10])
    defparam i19344_3_lut.LUT_INIT = 16'hecec;
    SB_CARRY add_4117_5 (.CI(n29233), .I0(n8437[2]), .I1(n317_adj_3961), 
            .CO(n29234));
    SB_LUT4 mult_10_i306_2_lut (.I0(\Kp[6] ), .I1(\PID_CONTROLLER.err [5]), 
            .I2(GND_net), .I3(GND_net), .O(n454_adj_4222));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i306_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_4145_10_lut (.I0(GND_net), .I1(n8815[7]), .I2(n700), .I3(n29550), 
            .O(n8804[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4145_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4134_11_lut (.I0(GND_net), .I1(n8639[8]), .I2(n740), .I3(n29397), 
            .O(n8617[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4134_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4117_4_lut (.I0(GND_net), .I1(n8437[1]), .I2(n244_adj_3960), 
            .I3(n29232), .O(n8420[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4117_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4117_4 (.CI(n29232), .I0(n8437[1]), .I1(n244_adj_3960), 
            .CO(n29233));
    SB_CARRY add_4134_11 (.CI(n29397), .I0(n8639[8]), .I1(n740), .CO(n29398));
    SB_LUT4 add_4117_3_lut (.I0(GND_net), .I1(n8437[0]), .I2(n171_adj_3959), 
            .I3(n29231), .O(n8420[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4117_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4117_3 (.CI(n29231), .I0(n8437[0]), .I1(n171_adj_3959), 
            .CO(n29232));
    SB_LUT4 add_4145_9_lut (.I0(GND_net), .I1(n8815[6]), .I2(n627), .I3(n29549), 
            .O(n8804[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4145_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4134_10_lut (.I0(GND_net), .I1(n8639[7]), .I2(n667), .I3(n29396), 
            .O(n8617[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4134_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4117_2_lut (.I0(GND_net), .I1(n29_adj_3957), .I2(n98_adj_3956), 
            .I3(GND_net), .O(n8420[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4117_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4134_10 (.CI(n29396), .I0(n8639[7]), .I1(n667), .CO(n29397));
    SB_CARRY add_4117_2 (.CI(GND_net), .I0(n29_adj_3957), .I1(n98_adj_3956), 
            .CO(n29231));
    SB_LUT4 mult_11_i639_2_lut (.I0(\Ki[13] ), .I1(\PID_CONTROLLER.integral [0]), 
            .I2(GND_net), .I3(GND_net), .O(n950_adj_4223));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i639_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i659_2_lut (.I0(\Ki[13] ), .I1(\PID_CONTROLLER.integral [10]), 
            .I2(GND_net), .I3(GND_net), .O(n980_adj_4224));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i659_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i688_2_lut (.I0(\Ki[14] ), .I1(\PID_CONTROLLER.integral [0]), 
            .I2(GND_net), .I3(GND_net), .O(n1023_adj_4225));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i688_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i355_2_lut (.I0(\Kp[7] ), .I1(\PID_CONTROLLER.err [5]), 
            .I2(GND_net), .I3(GND_net), .O(n527_adj_4226));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i355_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i63_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral [6]), 
            .I2(GND_net), .I3(GND_net), .O(n92));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i63_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i16_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral [7]), 
            .I2(GND_net), .I3(GND_net), .O(n23_adj_4000));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i16_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i73_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral [11]), 
            .I2(GND_net), .I3(GND_net), .O(n107_adj_4227));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i73_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i26_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral [12]), 
            .I2(GND_net), .I3(GND_net), .O(n38_adj_4228));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i26_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_4116_17_lut (.I0(GND_net), .I1(n8420[14]), .I2(GND_net), 
            .I3(n29230), .O(n8402[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4116_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4116_16_lut (.I0(GND_net), .I1(n8420[13]), .I2(n1117_adj_3955), 
            .I3(n29229), .O(n8402[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4116_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4145_9 (.CI(n29549), .I0(n8815[6]), .I1(n627), .CO(n29550));
    SB_CARRY add_4116_16 (.CI(n29229), .I0(n8420[13]), .I1(n1117_adj_3955), 
            .CO(n29230));
    SB_LUT4 mult_10_i404_2_lut (.I0(\Kp[8] ), .I1(\PID_CONTROLLER.err [5]), 
            .I2(GND_net), .I3(GND_net), .O(n600_adj_4229));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i404_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_4116_15_lut (.I0(GND_net), .I1(n8420[12]), .I2(n1044_adj_3951), 
            .I3(n29228), .O(n8402[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4116_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_668_15_lut (.I0(GND_net), .I1(n3265[13]), .I2(n3290[13]), 
            .I3(n27983), .O(duty_23__N_3613[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_668_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4145_8_lut (.I0(GND_net), .I1(n8815[5]), .I2(n554), .I3(n29548), 
            .O(n8804[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4145_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4134_9_lut (.I0(GND_net), .I1(n8639[6]), .I2(n594), .I3(n29395), 
            .O(n8617[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4134_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4116_15 (.CI(n29228), .I0(n8420[12]), .I1(n1044_adj_3951), 
            .CO(n29229));
    SB_CARRY add_4134_9 (.CI(n29395), .I0(n8639[6]), .I1(n594), .CO(n29396));
    SB_LUT4 add_4116_14_lut (.I0(GND_net), .I1(n8420[11]), .I2(n971_adj_3947), 
            .I3(n29227), .O(n8402[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4116_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4145_8 (.CI(n29548), .I0(n8815[5]), .I1(n554), .CO(n29549));
    SB_LUT4 add_4134_8_lut (.I0(GND_net), .I1(n8639[5]), .I2(n521), .I3(n29394), 
            .O(n8617[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4134_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4116_14 (.CI(n29227), .I0(n8420[11]), .I1(n971_adj_3947), 
            .CO(n29228));
    SB_CARRY add_4134_8 (.CI(n29394), .I0(n8639[5]), .I1(n521), .CO(n29395));
    SB_LUT4 add_4116_13_lut (.I0(GND_net), .I1(n8420[10]), .I2(n898_adj_3946), 
            .I3(n29226), .O(n8402[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4116_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_668_15 (.CI(n27983), .I0(n3265[13]), .I1(n3290[13]), 
            .CO(n27984));
    SB_LUT4 add_668_14_lut (.I0(GND_net), .I1(n3265[12]), .I2(n3290[12]), 
            .I3(n27982), .O(duty_23__N_3613[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_668_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4145_7_lut (.I0(GND_net), .I1(n8815[4]), .I2(n481), .I3(n29547), 
            .O(n8804[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4145_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4134_7_lut (.I0(GND_net), .I1(n8639[4]), .I2(n448), .I3(n29393), 
            .O(n8617[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4134_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4116_13 (.CI(n29226), .I0(n8420[10]), .I1(n898_adj_3946), 
            .CO(n29227));
    SB_CARRY add_4134_7 (.CI(n29393), .I0(n8639[4]), .I1(n448), .CO(n29394));
    SB_LUT4 add_4116_12_lut (.I0(GND_net), .I1(n8420[9]), .I2(n825_adj_3945), 
            .I3(n29225), .O(n8402[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4116_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_668_14 (.CI(n27982), .I0(n3265[12]), .I1(n3290[12]), 
            .CO(n27983));
    SB_CARRY add_4145_7 (.CI(n29547), .I0(n8815[4]), .I1(n481), .CO(n29548));
    SB_LUT4 add_4134_6_lut (.I0(GND_net), .I1(n8639[3]), .I2(n375), .I3(n29392), 
            .O(n8617[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4134_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4116_12 (.CI(n29225), .I0(n8420[9]), .I1(n825_adj_3945), 
            .CO(n29226));
    SB_LUT4 add_4116_11_lut (.I0(GND_net), .I1(n8420[8]), .I2(n752_adj_3944), 
            .I3(n29224), .O(n8402[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4116_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_5_add_3_7 (.CI(n28090), .I0(GND_net), .I1(n1_adj_4332[5]), 
            .CO(n28091));
    SB_CARRY add_4134_6 (.CI(n29392), .I0(n8639[3]), .I1(n375), .CO(n29393));
    SB_CARRY add_4116_11 (.CI(n29224), .I0(n8420[8]), .I1(n752_adj_3944), 
            .CO(n29225));
    SB_LUT4 add_4116_10_lut (.I0(GND_net), .I1(n8420[7]), .I2(n679_adj_3942), 
            .I3(n29223), .O(n8402[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4116_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_668_13_lut (.I0(GND_net), .I1(n3265[11]), .I2(n3290[11]), 
            .I3(n27981), .O(duty_23__N_3613[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_668_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i453_2_lut (.I0(\Kp[9] ), .I1(\PID_CONTROLLER.err [5]), 
            .I2(GND_net), .I3(GND_net), .O(n673_adj_4230));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i453_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_4145_6_lut (.I0(GND_net), .I1(n8815[3]), .I2(n408_adj_3939), 
            .I3(n29546), .O(n8804[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4145_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4134_5_lut (.I0(GND_net), .I1(n8639[2]), .I2(n302), .I3(n29391), 
            .O(n8617[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4134_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4116_10 (.CI(n29223), .I0(n8420[7]), .I1(n679_adj_3942), 
            .CO(n29224));
    SB_CARRY add_4134_5 (.CI(n29391), .I0(n8639[2]), .I1(n302), .CO(n29392));
    SB_LUT4 add_4116_9_lut (.I0(GND_net), .I1(n8420[6]), .I2(n606_adj_3937), 
            .I3(n29222), .O(n8402[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4116_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_5_add_3_6_lut (.I0(\PID_CONTROLLER.integral [4]), 
            .I1(GND_net), .I2(n1_adj_4332[4]), .I3(n28089), .O(n9_adj_4231)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_6_lut.LUT_INIT = 16'h6996;
    SB_CARRY add_4145_6 (.CI(n29546), .I0(n8815[3]), .I1(n408_adj_3939), 
            .CO(n29547));
    SB_LUT4 add_4134_4_lut (.I0(GND_net), .I1(n8639[1]), .I2(n229), .I3(n29390), 
            .O(n8617[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4134_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4116_9 (.CI(n29222), .I0(n8420[6]), .I1(n606_adj_3937), 
            .CO(n29223));
    SB_LUT4 add_4116_8_lut (.I0(GND_net), .I1(n8420[5]), .I2(n533_adj_3935), 
            .I3(n29221), .O(n8402[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4116_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4134_4 (.CI(n29390), .I0(n8639[1]), .I1(n229), .CO(n29391));
    SB_CARRY add_4116_8 (.CI(n29221), .I0(n8420[5]), .I1(n533_adj_3935), 
            .CO(n29222));
    SB_LUT4 mult_11_i737_2_lut (.I0(\Ki[15] ), .I1(\PID_CONTROLLER.integral [0]), 
            .I2(GND_net), .I3(GND_net), .O(n1096_adj_4232));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i737_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_4145_5_lut (.I0(GND_net), .I1(n8815[2]), .I2(n335), .I3(n29545), 
            .O(n8804[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4145_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4134_3_lut (.I0(GND_net), .I1(n8639[0]), .I2(n156), .I3(n29389), 
            .O(n8617[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4134_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4116_7_lut (.I0(GND_net), .I1(n8420[4]), .I2(n460_adj_3934), 
            .I3(n29220), .O(n8402[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4116_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4134_3 (.CI(n29389), .I0(n8639[0]), .I1(n156), .CO(n29390));
    SB_CARRY add_4116_7 (.CI(n29220), .I0(n8420[4]), .I1(n460_adj_3934), 
            .CO(n29221));
    SB_CARRY unary_minus_5_add_3_6 (.CI(n28089), .I0(GND_net), .I1(n1_adj_4332[4]), 
            .CO(n28090));
    SB_LUT4 unary_minus_5_add_3_5_lut (.I0(\PID_CONTROLLER.integral [3]), 
            .I1(GND_net), .I2(n1_adj_4332[3]), .I3(n28088), .O(n7_adj_4233)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_5_lut.LUT_INIT = 16'h6996;
    SB_CARRY add_4145_5 (.CI(n29545), .I0(n8815[2]), .I1(n335), .CO(n29546));
    SB_LUT4 add_4134_2_lut (.I0(GND_net), .I1(n14), .I2(n83), .I3(GND_net), 
            .O(n8617[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4134_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4116_6_lut (.I0(GND_net), .I1(n8420[3]), .I2(n387_adj_3931), 
            .I3(n29219), .O(n8402[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4116_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i112_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral [6]), 
            .I2(GND_net), .I3(GND_net), .O(n165));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i112_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i122_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral [11]), 
            .I2(GND_net), .I3(GND_net), .O(n180_adj_4234));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i122_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i502_2_lut (.I0(\Kp[10] ), .I1(\PID_CONTROLLER.err [5]), 
            .I2(GND_net), .I3(GND_net), .O(n746_adj_4235));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i502_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i31380_3_lut (.I0(n38061), .I1(duty[23]), .I2(n47_adj_4236), 
            .I3(GND_net), .O(n256));   // verilog/motorControl.v(46[19:35])
    defparam i31380_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i19563_1_lut (.I0(n256), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n24379));   // verilog/motorControl.v(46[19:35])
    defparam i19563_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_5_inv_0_i22_1_lut (.I0(IntegralLimit[21]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4332[21]));   // verilog/motorControl.v(39[48:62])
    defparam unary_minus_5_inv_0_i22_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_11_i161_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral [6]), 
            .I2(GND_net), .I3(GND_net), .O(n238));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i161_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i367_2_lut (.I0(\Kp[7] ), .I1(\PID_CONTROLLER.err [11]), 
            .I2(GND_net), .I3(GND_net), .O(n545));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i367_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_4145_4_lut (.I0(GND_net), .I1(n8815[1]), .I2(n262_adj_4237), 
            .I3(n29544), .O(n8804[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4145_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i210_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral [6]), 
            .I2(GND_net), .I3(GND_net), .O(n311));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i210_2_lut.LUT_INIT = 16'h8888;
    SB_DFF result_i1 (.Q(duty[1]), .C(clk32MHz), .D(duty_23__N_3490[1]));   // verilog/motorControl.v(37[14] 56[8])
    SB_LUT4 mult_11_i377_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral [16]), 
            .I2(GND_net), .I3(GND_net), .O(n560_adj_4091));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i377_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_4145_4 (.CI(n29544), .I0(n8815[1]), .I1(n262_adj_4237), 
            .CO(n29545));
    SB_LUT4 mult_10_i704_2_lut (.I0(\Kp[14] ), .I1(\PID_CONTROLLER.err [8]), 
            .I2(GND_net), .I3(GND_net), .O(n1047_adj_4090));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i704_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i753_2_lut (.I0(\Kp[15] ), .I1(\PID_CONTROLLER.err [8]), 
            .I2(GND_net), .I3(GND_net), .O(n1120_adj_4089));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i753_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i259_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral [6]), 
            .I2(GND_net), .I3(GND_net), .O(n384));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i259_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_666_i17_3_lut (.I0(n155[16]), .I1(PWMLimit[16]), .I2(n256), 
            .I3(GND_net), .O(n3290[16]));   // verilog/motorControl.v(46[16] 48[10])
    defparam mux_666_i17_3_lut.LUT_INIT = 16'h3a3a;
    SB_CARRY add_4134_2 (.CI(GND_net), .I0(n14), .I1(n83), .CO(n29389));
    SB_LUT4 add_4145_3_lut (.I0(GND_net), .I1(n8815[0]), .I2(n189_adj_3994), 
            .I3(n29543), .O(n8804[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4145_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_668_13 (.CI(n27981), .I0(n3265[11]), .I1(n3290[11]), 
            .CO(n27982));
    SB_LUT4 mult_11_i85_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral [17]), 
            .I2(GND_net), .I3(GND_net), .O(n125_adj_4088));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i85_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_4116_6 (.CI(n29219), .I0(n8420[3]), .I1(n387_adj_3931), 
            .CO(n29220));
    SB_LUT4 mult_11_i38_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral [18]), 
            .I2(GND_net), .I3(GND_net), .O(n56_adj_4087));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i38_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_inv_0_i12_1_lut (.I0(IntegralLimit[11]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4332[11]));   // verilog/motorControl.v(39[48:62])
    defparam unary_minus_5_inv_0_i12_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i53_2_lut (.I0(\Kp[1] ), .I1(\PID_CONTROLLER.err [1]), 
            .I2(GND_net), .I3(GND_net), .O(n77));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i53_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i6_2_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err [2]), 
            .I2(GND_net), .I3(GND_net), .O(n8_adj_4069));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i6_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i59_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral [4]), 
            .I2(GND_net), .I3(GND_net), .O(n86));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i59_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i12_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral [5]), 
            .I2(GND_net), .I3(GND_net), .O(n17_adj_4068));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i12_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i108_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral [4]), 
            .I2(GND_net), .I3(GND_net), .O(n159));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i108_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i134_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral [17]), 
            .I2(GND_net), .I3(GND_net), .O(n198_adj_4067));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i134_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i69_2_lut (.I0(\Kp[1] ), .I1(\PID_CONTROLLER.err [9]), 
            .I2(GND_net), .I3(GND_net), .O(n101_adj_4064));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i69_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i22_2_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err [10]), 
            .I2(GND_net), .I3(GND_net), .O(n32_adj_4063));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i22_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i118_2_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err [9]), 
            .I2(GND_net), .I3(GND_net), .O(n174));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i118_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i198_2_lut (.I0(\Kp[4] ), .I1(\PID_CONTROLLER.err [0]), 
            .I2(GND_net), .I3(GND_net), .O(n293));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i198_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_4133_22_lut (.I0(GND_net), .I1(n8617[19]), .I2(GND_net), 
            .I3(n29388), .O(n8594[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4133_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i157_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral [4]), 
            .I2(GND_net), .I3(GND_net), .O(n232));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i157_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i183_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral [17]), 
            .I2(GND_net), .I3(GND_net), .O(n271_adj_4062));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i183_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_4116_5_lut (.I0(GND_net), .I1(n8420[2]), .I2(n314_adj_3978), 
            .I3(n29218), .O(n8402[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4116_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4145_3 (.CI(n29543), .I0(n8815[0]), .I1(n189_adj_3994), 
            .CO(n29544));
    SB_LUT4 mult_11_i206_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral [4]), 
            .I2(GND_net), .I3(GND_net), .O(n305));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i206_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_4133_21_lut (.I0(GND_net), .I1(n8617[18]), .I2(GND_net), 
            .I3(n29387), .O(n8594[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4133_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4145_2_lut (.I0(GND_net), .I1(n47_adj_3977), .I2(n116_adj_3976), 
            .I3(GND_net), .O(n8804[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4145_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4133_21 (.CI(n29387), .I0(n8617[18]), .I1(GND_net), .CO(n29388));
    SB_LUT4 mult_10_i167_2_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err [9]), 
            .I2(GND_net), .I3(GND_net), .O(n247));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i167_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_4145_2 (.CI(GND_net), .I0(n47_adj_3977), .I1(n116_adj_3976), 
            .CO(n29543));
    SB_LUT4 add_4133_20_lut (.I0(GND_net), .I1(n8617[17]), .I2(GND_net), 
            .I3(n29386), .O(n8594[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4133_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4116_5 (.CI(n29218), .I0(n8420[2]), .I1(n314_adj_3978), 
            .CO(n29219));
    SB_CARRY add_4133_20 (.CI(n29386), .I0(n8617[17]), .I1(GND_net), .CO(n29387));
    SB_LUT4 add_4116_4_lut (.I0(GND_net), .I1(n8420[1]), .I2(n241_adj_3975), 
            .I3(n29217), .O(n8402[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4116_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_668_12_lut (.I0(GND_net), .I1(n3265[10]), .I2(n3290[10]), 
            .I3(n27980), .O(duty_23__N_3613[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_668_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4133_19_lut (.I0(GND_net), .I1(n8617[16]), .I2(GND_net), 
            .I3(n29385), .O(n8594[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4133_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4133_19 (.CI(n29385), .I0(n8617[16]), .I1(GND_net), .CO(n29386));
    SB_LUT4 add_4144_11_lut (.I0(GND_net), .I1(n8804[8]), .I2(n770_adj_3974), 
            .I3(n29542), .O(n8792[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4144_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4116_4 (.CI(n29217), .I0(n8420[1]), .I1(n241_adj_3975), 
            .CO(n29218));
    SB_LUT4 add_4144_10_lut (.I0(GND_net), .I1(n8804[7]), .I2(n697_adj_3971), 
            .I3(n29541), .O(n8792[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4144_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4116_3_lut (.I0(GND_net), .I1(n8420[0]), .I2(n168_adj_3969), 
            .I3(n29216), .O(n8402[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4116_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4133_18_lut (.I0(GND_net), .I1(n8617[15]), .I2(GND_net), 
            .I3(n29384), .O(n8594[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4133_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4116_3 (.CI(n29216), .I0(n8420[0]), .I1(n168_adj_3969), 
            .CO(n29217));
    SB_CARRY add_4144_10 (.CI(n29541), .I0(n8804[7]), .I1(n697_adj_3971), 
            .CO(n29542));
    SB_LUT4 add_4144_9_lut (.I0(GND_net), .I1(n8804[6]), .I2(n624_adj_3967), 
            .I3(n29540), .O(n8792[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4144_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i171_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral [11]), 
            .I2(GND_net), .I3(GND_net), .O(n253_adj_4238));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i171_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_4144_9 (.CI(n29540), .I0(n8804[6]), .I1(n624_adj_3967), 
            .CO(n29541));
    SB_LUT4 add_4144_8_lut (.I0(GND_net), .I1(n8804[5]), .I2(n551_adj_3966), 
            .I3(n29539), .O(n8792[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4144_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i551_2_lut (.I0(\Kp[11] ), .I1(\PID_CONTROLLER.err [5]), 
            .I2(GND_net), .I3(GND_net), .O(n819_adj_4239));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i551_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i102_2_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err [1]), 
            .I2(GND_net), .I3(GND_net), .O(n150));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i102_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i220_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral [11]), 
            .I2(GND_net), .I3(GND_net), .O(n326_adj_4240));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i220_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i600_2_lut (.I0(\Kp[12] ), .I1(\PID_CONTROLLER.err [5]), 
            .I2(GND_net), .I3(GND_net), .O(n892_adj_4241));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i600_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i649_2_lut (.I0(\Kp[13] ), .I1(\PID_CONTROLLER.err [5]), 
            .I2(GND_net), .I3(GND_net), .O(n965_adj_4242));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i649_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_666_i2_3_lut (.I0(n155[1]), .I1(n1[1]), .I2(n256), .I3(GND_net), 
            .O(n3290[1]));   // verilog/motorControl.v(46[16] 48[10])
    defparam mux_666_i2_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_10_i698_2_lut (.I0(\Kp[14] ), .I1(\PID_CONTROLLER.err [5]), 
            .I2(GND_net), .I3(GND_net), .O(n1038_adj_4243));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i698_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i269_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral [11]), 
            .I2(GND_net), .I3(GND_net), .O(n399_adj_4244));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i269_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i318_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral [11]), 
            .I2(GND_net), .I3(GND_net), .O(n472_adj_4245));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i318_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i747_2_lut (.I0(\Kp[15] ), .I1(\PID_CONTROLLER.err [5]), 
            .I2(GND_net), .I3(GND_net), .O(n1111_adj_4246));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i747_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i367_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral [11]), 
            .I2(GND_net), .I3(GND_net), .O(n545_adj_4247));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i367_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i55_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral [2]), 
            .I2(GND_net), .I3(GND_net), .O(n80_adj_4248));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i55_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i8_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral [3]), 
            .I2(GND_net), .I3(GND_net), .O(n11_adj_4249));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i8_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_666_i3_3_lut (.I0(n155[2]), .I1(n1[2]), .I2(n256), .I3(GND_net), 
            .O(n3290[2]));   // verilog/motorControl.v(46[16] 48[10])
    defparam mux_666_i3_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_10_i151_2_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err [1]), 
            .I2(GND_net), .I3(GND_net), .O(n223));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i151_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i200_2_lut (.I0(\Kp[4] ), .I1(\PID_CONTROLLER.err [1]), 
            .I2(GND_net), .I3(GND_net), .O(n296));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i200_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i177_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral [14]), 
            .I2(GND_net), .I3(GND_net), .O(n262_adj_4237));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i177_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_666_i4_3_lut (.I0(n155[3]), .I1(n1[3]), .I2(n256), .I3(GND_net), 
            .O(n3290[3]));   // verilog/motorControl.v(46[16] 48[10])
    defparam mux_666_i4_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_11_i232_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral [17]), 
            .I2(GND_net), .I3(GND_net), .O(n344));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i232_2_lut.LUT_INIT = 16'h8888;
    SB_DFF result_i2 (.Q(duty[2]), .C(clk32MHz), .D(duty_23__N_3490[2]));   // verilog/motorControl.v(37[14] 56[8])
    SB_CARRY unary_minus_5_add_3_5 (.CI(n28088), .I0(GND_net), .I1(n1_adj_4332[3]), 
            .CO(n28089));
    SB_DFF result_i3 (.Q(duty[3]), .C(clk32MHz), .D(duty_23__N_3490[3]));   // verilog/motorControl.v(37[14] 56[8])
    SB_DFF result_i4 (.Q(duty[4]), .C(clk32MHz), .D(duty_23__N_3490[4]));   // verilog/motorControl.v(37[14] 56[8])
    SB_DFF result_i5 (.Q(duty[5]), .C(clk32MHz), .D(duty_23__N_3490[5]));   // verilog/motorControl.v(37[14] 56[8])
    SB_DFF result_i6 (.Q(duty[6]), .C(clk32MHz), .D(duty_23__N_3490[6]));   // verilog/motorControl.v(37[14] 56[8])
    SB_DFF result_i7 (.Q(duty[7]), .C(clk32MHz), .D(duty_23__N_3490[7]));   // verilog/motorControl.v(37[14] 56[8])
    SB_DFF result_i8 (.Q(duty[8]), .C(clk32MHz), .D(duty_23__N_3490[8]));   // verilog/motorControl.v(37[14] 56[8])
    SB_DFF result_i9 (.Q(duty[9]), .C(clk32MHz), .D(duty_23__N_3490[9]));   // verilog/motorControl.v(37[14] 56[8])
    SB_DFF result_i10 (.Q(duty[10]), .C(clk32MHz), .D(duty_23__N_3490[10]));   // verilog/motorControl.v(37[14] 56[8])
    SB_DFF result_i11 (.Q(duty[11]), .C(clk32MHz), .D(duty_23__N_3490[11]));   // verilog/motorControl.v(37[14] 56[8])
    SB_DFF result_i12 (.Q(duty[12]), .C(clk32MHz), .D(duty_23__N_3490[12]));   // verilog/motorControl.v(37[14] 56[8])
    SB_DFF result_i13 (.Q(duty[13]), .C(clk32MHz), .D(duty_23__N_3490[13]));   // verilog/motorControl.v(37[14] 56[8])
    SB_DFF result_i14 (.Q(duty[14]), .C(clk32MHz), .D(duty_23__N_3490[14]));   // verilog/motorControl.v(37[14] 56[8])
    SB_DFF result_i15 (.Q(duty[15]), .C(clk32MHz), .D(duty_23__N_3490[15]));   // verilog/motorControl.v(37[14] 56[8])
    SB_DFF result_i16 (.Q(duty[16]), .C(clk32MHz), .D(duty_23__N_3490[16]));   // verilog/motorControl.v(37[14] 56[8])
    SB_DFF result_i17 (.Q(duty[17]), .C(clk32MHz), .D(duty_23__N_3490[17]));   // verilog/motorControl.v(37[14] 56[8])
    SB_DFF result_i18 (.Q(duty[18]), .C(clk32MHz), .D(duty_23__N_3490[18]));   // verilog/motorControl.v(37[14] 56[8])
    SB_DFF result_i19 (.Q(duty[19]), .C(clk32MHz), .D(duty_23__N_3490[19]));   // verilog/motorControl.v(37[14] 56[8])
    SB_DFF result_i20 (.Q(duty[20]), .C(clk32MHz), .D(duty_23__N_3490[20]));   // verilog/motorControl.v(37[14] 56[8])
    SB_DFF result_i21 (.Q(duty[21]), .C(clk32MHz), .D(duty_23__N_3490[21]));   // verilog/motorControl.v(37[14] 56[8])
    SB_DFF result_i22 (.Q(duty[22]), .C(clk32MHz), .D(duty_23__N_3490[22]));   // verilog/motorControl.v(37[14] 56[8])
    SB_DFF result_i23 (.Q(duty[23]), .C(clk32MHz), .D(duty_23__N_3490[23]));   // verilog/motorControl.v(37[14] 56[8])
    SB_DFF \PID_CONTROLLER.err_i1  (.Q(\PID_CONTROLLER.err [1]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_23__N_3514 [1]));   // verilog/motorControl.v(37[14] 56[8])
    SB_DFF \PID_CONTROLLER.err_i2  (.Q(\PID_CONTROLLER.err [2]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_23__N_3514 [2]));   // verilog/motorControl.v(37[14] 56[8])
    SB_DFF \PID_CONTROLLER.err_i3  (.Q(\PID_CONTROLLER.err [3]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_23__N_3514 [3]));   // verilog/motorControl.v(37[14] 56[8])
    SB_DFF \PID_CONTROLLER.err_i4  (.Q(\PID_CONTROLLER.err [4]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_23__N_3514 [4]));   // verilog/motorControl.v(37[14] 56[8])
    SB_DFF \PID_CONTROLLER.err_i5  (.Q(\PID_CONTROLLER.err [5]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_23__N_3514 [5]));   // verilog/motorControl.v(37[14] 56[8])
    SB_DFF \PID_CONTROLLER.err_i6  (.Q(\PID_CONTROLLER.err [6]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_23__N_3514 [6]));   // verilog/motorControl.v(37[14] 56[8])
    SB_DFF \PID_CONTROLLER.err_i7  (.Q(\PID_CONTROLLER.err [7]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_23__N_3514 [7]));   // verilog/motorControl.v(37[14] 56[8])
    SB_DFF \PID_CONTROLLER.err_i8  (.Q(\PID_CONTROLLER.err [8]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_23__N_3514 [8]));   // verilog/motorControl.v(37[14] 56[8])
    SB_DFF \PID_CONTROLLER.err_i9  (.Q(\PID_CONTROLLER.err [9]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_23__N_3514 [9]));   // verilog/motorControl.v(37[14] 56[8])
    SB_DFF \PID_CONTROLLER.err_i10  (.Q(\PID_CONTROLLER.err [10]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_23__N_3514 [10]));   // verilog/motorControl.v(37[14] 56[8])
    SB_DFF \PID_CONTROLLER.err_i11  (.Q(\PID_CONTROLLER.err [11]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_23__N_3514 [11]));   // verilog/motorControl.v(37[14] 56[8])
    SB_DFF \PID_CONTROLLER.err_i12  (.Q(\PID_CONTROLLER.err [12]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_23__N_3514 [12]));   // verilog/motorControl.v(37[14] 56[8])
    SB_DFF \PID_CONTROLLER.err_i13  (.Q(\PID_CONTROLLER.err [13]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_23__N_3514 [13]));   // verilog/motorControl.v(37[14] 56[8])
    SB_DFF \PID_CONTROLLER.err_i14  (.Q(\PID_CONTROLLER.err [14]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_23__N_3514 [14]));   // verilog/motorControl.v(37[14] 56[8])
    SB_DFF \PID_CONTROLLER.err_i15  (.Q(\PID_CONTROLLER.err [15]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_23__N_3514 [15]));   // verilog/motorControl.v(37[14] 56[8])
    SB_DFF \PID_CONTROLLER.err_i16  (.Q(\PID_CONTROLLER.err [16]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_23__N_3514 [16]));   // verilog/motorControl.v(37[14] 56[8])
    SB_DFF \PID_CONTROLLER.err_i17  (.Q(\PID_CONTROLLER.err [17]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_23__N_3514 [17]));   // verilog/motorControl.v(37[14] 56[8])
    SB_DFF \PID_CONTROLLER.err_i18  (.Q(\PID_CONTROLLER.err [18]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_23__N_3514 [18]));   // verilog/motorControl.v(37[14] 56[8])
    SB_DFF \PID_CONTROLLER.err_i19  (.Q(\PID_CONTROLLER.err [19]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_23__N_3514 [19]));   // verilog/motorControl.v(37[14] 56[8])
    SB_DFF \PID_CONTROLLER.err_i20  (.Q(\PID_CONTROLLER.err [20]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_23__N_3514 [20]));   // verilog/motorControl.v(37[14] 56[8])
    SB_DFF \PID_CONTROLLER.err_i21  (.Q(\PID_CONTROLLER.err [21]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_23__N_3514 [21]));   // verilog/motorControl.v(37[14] 56[8])
    SB_DFF \PID_CONTROLLER.err_i22  (.Q(\PID_CONTROLLER.err [22]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_23__N_3514 [22]));   // verilog/motorControl.v(37[14] 56[8])
    SB_DFF \PID_CONTROLLER.err_i23  (.Q(\PID_CONTROLLER.err [23]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_23__N_3514 [23]));   // verilog/motorControl.v(37[14] 56[8])
    SB_CARRY add_4144_8 (.CI(n29539), .I0(n8804[5]), .I1(n551_adj_3966), 
            .CO(n29540));
    SB_CARRY add_668_12 (.CI(n27980), .I0(n3265[10]), .I1(n3290[10]), 
            .CO(n27981));
    SB_LUT4 add_668_11_lut (.I0(GND_net), .I1(n3265[9]), .I2(n3290[9]), 
            .I3(n27979), .O(duty_23__N_3613[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_668_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i104_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral [2]), 
            .I2(GND_net), .I3(GND_net), .O(n153_adj_4250));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i104_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i416_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral [11]), 
            .I2(GND_net), .I3(GND_net), .O(n618_adj_4251));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i416_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_4144_7_lut (.I0(GND_net), .I1(n8804[4]), .I2(n478_adj_3930), 
            .I3(n29538), .O(n8792[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4144_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i63_2_lut (.I0(\Kp[1] ), .I1(\PID_CONTROLLER.err [6]), 
            .I2(GND_net), .I3(GND_net), .O(n92_adj_4252));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i63_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i16_2_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err [7]), 
            .I2(GND_net), .I3(GND_net), .O(n23_adj_4253));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i16_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_add_3_4_lut (.I0(\PID_CONTROLLER.integral [2]), 
            .I1(GND_net), .I2(n1_adj_4332[2]), .I3(n28087), .O(n5_adj_4254)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 mult_11_i153_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral [2]), 
            .I2(GND_net), .I3(GND_net), .O(n226_adj_4255));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i153_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_4144_7 (.CI(n29538), .I0(n8804[4]), .I1(n478_adj_3930), 
            .CO(n29539));
    SB_LUT4 mult_10_i112_2_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err [6]), 
            .I2(GND_net), .I3(GND_net), .O(n165_adj_4256));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i112_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_668_11 (.CI(n27979), .I0(n3265[9]), .I1(n3290[9]), .CO(n27980));
    SB_CARRY unary_minus_5_add_3_4 (.CI(n28087), .I0(GND_net), .I1(n1_adj_4332[2]), 
            .CO(n28088));
    SB_CARRY add_4133_18 (.CI(n29384), .I0(n8617[15]), .I1(GND_net), .CO(n29385));
    SB_LUT4 add_4116_2_lut (.I0(GND_net), .I1(n26), .I2(n95), .I3(GND_net), 
            .O(n8402[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4116_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i202_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral [2]), 
            .I2(GND_net), .I3(GND_net), .O(n299_adj_4257));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i202_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i465_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral [11]), 
            .I2(GND_net), .I3(GND_net), .O(n691_adj_4258));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i465_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_4116_2 (.CI(GND_net), .I0(n26), .I1(n95), .CO(n29216));
    SB_LUT4 mult_10_i161_2_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err [6]), 
            .I2(GND_net), .I3(GND_net), .O(n238_adj_4259));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i161_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i210_2_lut (.I0(\Kp[4] ), .I1(\PID_CONTROLLER.err [6]), 
            .I2(GND_net), .I3(GND_net), .O(n311_adj_4260));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i210_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i251_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral [2]), 
            .I2(GND_net), .I3(GND_net), .O(n372_adj_4261));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i251_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i259_2_lut (.I0(\Kp[5] ), .I1(\PID_CONTROLLER.err [6]), 
            .I2(GND_net), .I3(GND_net), .O(n384_adj_4262));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i259_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_666_i18_3_lut (.I0(n155[17]), .I1(PWMLimit[17]), .I2(n256), 
            .I3(GND_net), .O(n3290[17]));   // verilog/motorControl.v(46[16] 48[10])
    defparam mux_666_i18_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 mult_10_i308_2_lut (.I0(\Kp[6] ), .I1(\PID_CONTROLLER.err [6]), 
            .I2(GND_net), .I3(GND_net), .O(n457_adj_4264));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i308_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i300_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral [2]), 
            .I2(GND_net), .I3(GND_net), .O(n445_adj_4265));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i300_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i514_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral [11]), 
            .I2(GND_net), .I3(GND_net), .O(n764_adj_4266));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i514_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i563_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral [11]), 
            .I2(GND_net), .I3(GND_net), .O(n837_adj_4267));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i563_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i612_2_lut (.I0(\Ki[12] ), .I1(\PID_CONTROLLER.integral [11]), 
            .I2(GND_net), .I3(GND_net), .O(n910_adj_4268));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i612_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_inv_0_i13_1_lut (.I0(IntegralLimit[12]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4332[12]));   // verilog/motorControl.v(39[48:62])
    defparam unary_minus_5_inv_0_i13_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mux_666_i5_3_lut (.I0(n155[4]), .I1(n1[4]), .I2(n256), .I3(GND_net), 
            .O(n3290[4]));   // verilog/motorControl.v(46[16] 48[10])
    defparam mux_666_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_11_i75_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral [12]), 
            .I2(GND_net), .I3(GND_net), .O(n110_adj_4269));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i75_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_4144_6_lut (.I0(GND_net), .I1(n8804[3]), .I2(n405_adj_3913), 
            .I3(n29537), .O(n8792[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4144_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i28_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral [13]), 
            .I2(GND_net), .I3(GND_net), .O(n41_adj_4270));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i28_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i349_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral [2]), 
            .I2(GND_net), .I3(GND_net), .O(n518_adj_4271));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i349_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i357_2_lut (.I0(\Kp[7] ), .I1(\PID_CONTROLLER.err [6]), 
            .I2(GND_net), .I3(GND_net), .O(n530_adj_4272));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i357_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i124_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral [12]), 
            .I2(GND_net), .I3(GND_net), .O(n183_adj_4273));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i124_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i406_2_lut (.I0(\Kp[8] ), .I1(\PID_CONTROLLER.err [6]), 
            .I2(GND_net), .I3(GND_net), .O(n603_adj_4274));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i406_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_4144_6 (.CI(n29537), .I0(n8804[3]), .I1(n405_adj_3913), 
            .CO(n29538));
    SB_LUT4 add_4133_17_lut (.I0(GND_net), .I1(n8617[14]), .I2(GND_net), 
            .I3(n29383), .O(n8594[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4133_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_5_add_3_3_lut (.I0(\PID_CONTROLLER.integral [1]), 
            .I1(GND_net), .I2(n1_adj_4332[1]), .I3(n28086), .O(n3_adj_4275)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_3_lut.LUT_INIT = 16'h6996;
    SB_LUT4 mult_11_i398_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral [2]), 
            .I2(GND_net), .I3(GND_net), .O(n591_adj_4276));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i398_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_666_i19_3_lut (.I0(n155[18]), .I1(PWMLimit[18]), .I2(n256), 
            .I3(GND_net), .O(n3290[18]));   // verilog/motorControl.v(46[16] 48[10])
    defparam mux_666_i19_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 mult_10_i216_2_lut (.I0(\Kp[4] ), .I1(\PID_CONTROLLER.err [9]), 
            .I2(GND_net), .I3(GND_net), .O(n320));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i216_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_16_inv_0_i6_1_lut (.I0(PWMLimit[5]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[5]));   // verilog/motorControl.v(47[19:28])
    defparam unary_minus_16_inv_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_4133_17 (.CI(n29383), .I0(n8617[14]), .I1(GND_net), .CO(n29384));
    SB_LUT4 add_4144_5_lut (.I0(GND_net), .I1(n8804[2]), .I2(n332_adj_3911), 
            .I3(n29536), .O(n8792[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4144_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_668_10_lut (.I0(GND_net), .I1(n3265[8]), .I2(n3290[8]), 
            .I3(n27978), .O(duty_23__N_3613[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_668_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4115_18_lut (.I0(GND_net), .I1(n8402[15]), .I2(GND_net), 
            .I3(n29215), .O(n8383[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4115_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4144_5 (.CI(n29536), .I0(n8804[2]), .I1(n332_adj_3911), 
            .CO(n29537));
    SB_LUT4 add_4144_4_lut (.I0(GND_net), .I1(n8804[1]), .I2(n259_adj_3910), 
            .I3(n29535), .O(n8792[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4144_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4144_4 (.CI(n29535), .I0(n8804[1]), .I1(n259_adj_3910), 
            .CO(n29536));
    SB_LUT4 add_4144_3_lut (.I0(GND_net), .I1(n8804[0]), .I2(n186_adj_3909), 
            .I3(n29534), .O(n8792[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4144_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i255_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral [4]), 
            .I2(GND_net), .I3(GND_net), .O(n378));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i255_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i173_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral [12]), 
            .I2(GND_net), .I3(GND_net), .O(n256_adj_4277));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i173_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY unary_minus_5_add_3_3 (.CI(n28086), .I0(GND_net), .I1(n1_adj_4332[1]), 
            .CO(n28087));
    SB_LUT4 add_4115_17_lut (.I0(GND_net), .I1(n8402[14]), .I2(GND_net), 
            .I3(n29214), .O(n8383[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4115_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4133_16_lut (.I0(GND_net), .I1(n8617[13]), .I2(n1102), 
            .I3(n29382), .O(n8594[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4133_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4144_3 (.CI(n29534), .I0(n8804[0]), .I1(n186_adj_3909), 
            .CO(n29535));
    SB_LUT4 add_4144_2_lut (.I0(GND_net), .I1(n44_adj_3908), .I2(n113_adj_3907), 
            .I3(GND_net), .O(n8792[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4144_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4133_16 (.CI(n29382), .I0(n8617[13]), .I1(n1102), .CO(n29383));
    SB_LUT4 add_4133_15_lut (.I0(GND_net), .I1(n8617[12]), .I2(n1029), 
            .I3(n29381), .O(n8594[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4133_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4115_17 (.CI(n29214), .I0(n8402[14]), .I1(GND_net), .CO(n29215));
    SB_CARRY add_4133_15 (.CI(n29381), .I0(n8617[12]), .I1(n1029), .CO(n29382));
    SB_LUT4 add_4133_14_lut (.I0(GND_net), .I1(n8617[11]), .I2(n956), 
            .I3(n29380), .O(n8594[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4133_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4115_16_lut (.I0(GND_net), .I1(n8402[13]), .I2(n1114), 
            .I3(n29213), .O(n8383[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4115_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4144_2 (.CI(GND_net), .I0(n44_adj_3908), .I1(n113_adj_3907), 
            .CO(n29534));
    SB_CARRY add_4133_14 (.CI(n29380), .I0(n8617[11]), .I1(n956), .CO(n29381));
    SB_CARRY add_668_10 (.CI(n27978), .I0(n3265[8]), .I1(n3290[8]), .CO(n27979));
    SB_LUT4 add_4143_12_lut (.I0(GND_net), .I1(n8792[9]), .I2(n840), .I3(n29533), 
            .O(n8779[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4143_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_668_9_lut (.I0(GND_net), .I1(n3265[7]), .I2(n3290[7]), 
            .I3(n27977), .O(duty_23__N_3613[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_668_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4115_16 (.CI(n29213), .I0(n8402[13]), .I1(n1114), .CO(n29214));
    SB_LUT4 add_4143_11_lut (.I0(GND_net), .I1(n8792[8]), .I2(n767_adj_4278), 
            .I3(n29532), .O(n8779[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4143_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4115_15_lut (.I0(GND_net), .I1(n8402[12]), .I2(n1041_adj_4279), 
            .I3(n29212), .O(n8383[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4115_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4133_13_lut (.I0(GND_net), .I1(n8617[10]), .I2(n883_adj_4280), 
            .I3(n29379), .O(n8594[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4133_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4143_11 (.CI(n29532), .I0(n8792[8]), .I1(n767_adj_4278), 
            .CO(n29533));
    SB_LUT4 add_4143_10_lut (.I0(GND_net), .I1(n8792[7]), .I2(n694_adj_4281), 
            .I3(n29531), .O(n8779[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4143_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4115_15 (.CI(n29212), .I0(n8402[12]), .I1(n1041_adj_4279), 
            .CO(n29213));
    SB_LUT4 add_4115_14_lut (.I0(GND_net), .I1(n8402[11]), .I2(n968_adj_4282), 
            .I3(n29211), .O(n8383[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4115_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4143_10 (.CI(n29531), .I0(n8792[7]), .I1(n694_adj_4281), 
            .CO(n29532));
    SB_CARRY add_4115_14 (.CI(n29211), .I0(n8402[11]), .I1(n968_adj_4282), 
            .CO(n29212));
    SB_LUT4 mult_11_i281_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral [17]), 
            .I2(GND_net), .I3(GND_net), .O(n417));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i281_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_add_3_2_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4332[0]), 
            .I3(VCC_net), .O(\PID_CONTROLLER.integral_23__N_3589 [0])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i2_4_lut_adj_849 (.I0(n6_adj_4046), .I1(\Ki[4] ), .I2(n8849[2]), 
            .I3(\PID_CONTROLLER.integral [18]), .O(n8842[3]));   // verilog/motorControl.v(42[26:37])
    defparam i2_4_lut_adj_849.LUT_INIT = 16'h965a;
    SB_LUT4 i22758_3_lut_4_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err [18]), 
            .I2(n4_adj_4284), .I3(n8552[1]), .O(n6_adj_4082));   // verilog/motorControl.v(42[17:23])
    defparam i22758_3_lut_4_lut.LUT_INIT = 16'hf880;
    SB_LUT4 mult_10_i249_2_lut (.I0(\Kp[5] ), .I1(\PID_CONTROLLER.err [1]), 
            .I2(GND_net), .I3(GND_net), .O(n369));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i249_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i455_2_lut (.I0(\Kp[9] ), .I1(\PID_CONTROLLER.err [6]), 
            .I2(GND_net), .I3(GND_net), .O(n676_adj_4285));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i455_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i304_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral [4]), 
            .I2(GND_net), .I3(GND_net), .O(n451));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i304_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_15_i37_2_lut (.I0(duty[18]), .I1(n257[18]), .I2(GND_net), 
            .I3(GND_net), .O(n37_adj_4002));   // verilog/motorControl.v(46[19:35])
    defparam LessThan_15_i37_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_15_i45_2_lut (.I0(duty[22]), .I1(n257[22]), .I2(GND_net), 
            .I3(GND_net), .O(n45_adj_4038));   // verilog/motorControl.v(46[19:35])
    defparam LessThan_15_i45_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_15_i25_2_lut (.I0(duty[12]), .I1(n257[12]), .I2(GND_net), 
            .I3(GND_net), .O(n25_adj_4049));   // verilog/motorControl.v(46[19:35])
    defparam LessThan_15_i25_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_15_i41_2_lut (.I0(duty[20]), .I1(n257[20]), .I2(GND_net), 
            .I3(GND_net), .O(n41_adj_4139));   // verilog/motorControl.v(46[19:35])
    defparam LessThan_15_i41_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_15_i43_2_lut (.I0(duty[21]), .I1(n257[21]), .I2(GND_net), 
            .I3(GND_net), .O(n43_adj_4005));   // verilog/motorControl.v(46[19:35])
    defparam LessThan_15_i43_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_15_i39_2_lut (.I0(duty[19]), .I1(n257[19]), .I2(GND_net), 
            .I3(GND_net), .O(n39_adj_4084));   // verilog/motorControl.v(46[19:35])
    defparam LessThan_15_i39_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_668_9 (.CI(n27977), .I0(n3265[7]), .I1(n3290[7]), .CO(n27978));
    SB_CARRY add_4133_13 (.CI(n29379), .I0(n8617[10]), .I1(n883_adj_4280), 
            .CO(n29380));
    SB_LUT4 i2_3_lut_4_lut_adj_850 (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err [18]), 
            .I2(n8552[1]), .I3(n4_adj_4284), .O(n8545[2]));   // verilog/motorControl.v(42[17:23])
    defparam i2_3_lut_4_lut_adj_850.LUT_INIT = 16'h8778;
    SB_LUT4 i2_3_lut_4_lut_adj_851 (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err [18]), 
            .I2(n8552[0]), .I3(n27544), .O(n8545[1]));   // verilog/motorControl.v(42[17:23])
    defparam i2_3_lut_4_lut_adj_851.LUT_INIT = 16'h8778;
    SB_LUT4 unary_minus_5_inv_0_i14_1_lut (.I0(IntegralLimit[13]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4332[13]));   // verilog/motorControl.v(39[48:62])
    defparam unary_minus_5_inv_0_i14_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_4143_9_lut (.I0(GND_net), .I1(n8792[6]), .I2(n621_adj_4286), 
            .I3(n29530), .O(n8779[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4143_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4143_9 (.CI(n29530), .I0(n8792[6]), .I1(n621_adj_4286), 
            .CO(n29531));
    SB_LUT4 mult_11_i222_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral [12]), 
            .I2(GND_net), .I3(GND_net), .O(n329_adj_4287));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i222_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i271_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral [12]), 
            .I2(GND_net), .I3(GND_net), .O(n402_adj_4288));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i271_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i22990_4_lut (.I0(\Ki[0] ), .I1(\Ki[1] ), .I2(\PID_CONTROLLER.integral [22]), 
            .I3(\PID_CONTROLLER.integral [21]), .O(n8860[0]));   // verilog/motorControl.v(42[26:37])
    defparam i22990_4_lut.LUT_INIT = 16'h6ca0;
    SB_LUT4 mux_666_i6_3_lut (.I0(n155[5]), .I1(n1[5]), .I2(n256), .I3(GND_net), 
            .O(n3290[5]));   // verilog/motorControl.v(46[16] 48[10])
    defparam mux_666_i6_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_10_i504_2_lut (.I0(\Kp[10] ), .I1(\PID_CONTROLLER.err [6]), 
            .I2(GND_net), .I3(GND_net), .O(n749_adj_4290));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i504_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i320_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral [12]), 
            .I2(GND_net), .I3(GND_net), .O(n475_adj_4291));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i320_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i447_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral [2]), 
            .I2(GND_net), .I3(GND_net), .O(n664_adj_4292));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i447_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i22750_3_lut_4_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err [18]), 
            .I2(n27544), .I3(n8552[0]), .O(n4_adj_4284));   // verilog/motorControl.v(42[17:23])
    defparam i22750_3_lut_4_lut.LUT_INIT = 16'hf880;
    SB_LUT4 mult_10_i553_2_lut (.I0(\Kp[11] ), .I1(\PID_CONTROLLER.err [6]), 
            .I2(GND_net), .I3(GND_net), .O(n822_adj_4293));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i553_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i22739_2_lut_3_lut_4_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err [19]), 
            .I2(\PID_CONTROLLER.err [18]), .I3(\Kp[1] ), .O(n27544));   // verilog/motorControl.v(42[17:23])
    defparam i22739_2_lut_3_lut_4_lut.LUT_INIT = 16'h8000;
    SB_CARRY unary_minus_5_add_3_2 (.CI(VCC_net), .I0(GND_net), .I1(n1_adj_4332[0]), 
            .CO(n28086));
    SB_LUT4 mult_11_i369_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral [12]), 
            .I2(GND_net), .I3(GND_net), .O(n548_adj_4294));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i369_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i496_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral [2]), 
            .I2(GND_net), .I3(GND_net), .O(n737_adj_4295));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i496_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_668_8_lut (.I0(GND_net), .I1(n3265[6]), .I2(n3290[6]), 
            .I3(n27976), .O(duty_23__N_3613[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_668_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i545_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral [2]), 
            .I2(GND_net), .I3(GND_net), .O(n810_adj_4296));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i545_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i602_2_lut (.I0(\Kp[12] ), .I1(\PID_CONTROLLER.err [6]), 
            .I2(GND_net), .I3(GND_net), .O(n895_adj_4297));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i602_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_666_i7_3_lut (.I0(n155[6]), .I1(PWMLimit[6]), .I2(n256), 
            .I3(GND_net), .O(n3290[6]));   // verilog/motorControl.v(46[16] 48[10])
    defparam mux_666_i7_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 add_4115_13_lut (.I0(GND_net), .I1(n8402[10]), .I2(n895_adj_4297), 
            .I3(n29210), .O(n8383[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4115_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4133_12_lut (.I0(GND_net), .I1(n8617[9]), .I2(n810_adj_4296), 
            .I3(n29378), .O(n8594[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4133_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4133_12 (.CI(n29378), .I0(n8617[9]), .I1(n810_adj_4296), 
            .CO(n29379));
    SB_LUT4 mult_11_i418_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral [12]), 
            .I2(GND_net), .I3(GND_net), .O(n621_adj_4286));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i418_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 IntegralLimit_23__I_0_i8_3_lut_3_lut (.I0(IntegralLimit[4]), .I1(IntegralLimit[8]), 
            .I2(\PID_CONTROLLER.integral [8]), .I3(GND_net), .O(n8_adj_4298));   // verilog/motorControl.v(39[10:34])
    defparam IntegralLimit_23__I_0_i8_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i22737_2_lut_3_lut_4_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err [19]), 
            .I2(\PID_CONTROLLER.err [18]), .I3(\Kp[1] ), .O(n8545[0]));   // verilog/motorControl.v(42[17:23])
    defparam i22737_2_lut_3_lut_4_lut.LUT_INIT = 16'h7888;
    SB_CARRY add_668_8 (.CI(n27976), .I0(n3265[6]), .I1(n3290[6]), .CO(n27977));
    SB_LUT4 add_4133_11_lut (.I0(GND_net), .I1(n8617[8]), .I2(n737_adj_4295), 
            .I3(n29377), .O(n8594[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4133_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4143_8_lut (.I0(GND_net), .I1(n8792[5]), .I2(n548_adj_4294), 
            .I3(n29529), .O(n8779[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4143_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4115_13 (.CI(n29210), .I0(n8402[10]), .I1(n895_adj_4297), 
            .CO(n29211));
    SB_CARRY add_4133_11 (.CI(n29377), .I0(n8617[8]), .I1(n737_adj_4295), 
            .CO(n29378));
    SB_LUT4 add_4115_12_lut (.I0(GND_net), .I1(n8402[9]), .I2(n822_adj_4293), 
            .I3(n29209), .O(n8383[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4115_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4133_10_lut (.I0(GND_net), .I1(n8617[7]), .I2(n664_adj_4292), 
            .I3(n29376), .O(n8594[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4133_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4143_8 (.CI(n29529), .I0(n8792[5]), .I1(n548_adj_4294), 
            .CO(n29530));
    SB_LUT4 i22820_3_lut_4_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err [20]), 
            .I2(n27621), .I3(n8563[0]), .O(n4_adj_4119));   // verilog/motorControl.v(42[17:23])
    defparam i22820_3_lut_4_lut.LUT_INIT = 16'hf880;
    SB_LUT4 i2_3_lut_4_lut_adj_852 (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err [20]), 
            .I2(n8563[0]), .I3(n27621), .O(n8558[1]));   // verilog/motorControl.v(42[17:23])
    defparam i2_3_lut_4_lut_adj_852.LUT_INIT = 16'h8778;
    SB_LUT4 i30765_2_lut_4_lut (.I0(duty[16]), .I1(n257[16]), .I2(duty[7]), 
            .I3(n257[7]), .O(n37446));
    defparam i30765_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_CARRY add_4115_12 (.CI(n29209), .I0(n8402[9]), .I1(n822_adj_4293), 
            .CO(n29210));
    SB_LUT4 i2_3_lut_4_lut_adj_853 (.I0(n62), .I1(n131), .I2(n8558[0]), 
            .I3(n204), .O(n8552[1]));   // verilog/motorControl.v(42[17:23])
    defparam i2_3_lut_4_lut_adj_853.LUT_INIT = 16'h8778;
    SB_LUT4 add_4143_7_lut (.I0(GND_net), .I1(n8792[4]), .I2(n475_adj_4291), 
            .I3(n29528), .O(n8779[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4143_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4115_11_lut (.I0(GND_net), .I1(n8402[8]), .I2(n749_adj_4290), 
            .I3(n29208), .O(n8383[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4115_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_668_7_lut (.I0(GND_net), .I1(n3265[5]), .I2(n3290[5]), 
            .I3(n27975), .O(duty_23__N_3613[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_668_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4115_11 (.CI(n29208), .I0(n8402[8]), .I1(n749_adj_4290), 
            .CO(n29209));
    SB_CARRY add_4133_10 (.CI(n29376), .I0(n8617[7]), .I1(n664_adj_4292), 
            .CO(n29377));
    SB_CARRY add_4143_7 (.CI(n29528), .I0(n8792[4]), .I1(n475_adj_4291), 
            .CO(n29529));
    SB_LUT4 add_4143_6_lut (.I0(GND_net), .I1(n8792[3]), .I2(n402_adj_4288), 
            .I3(n29527), .O(n8779[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4143_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i22789_3_lut_4_lut (.I0(n62), .I1(n131), .I2(n204), .I3(n8558[0]), 
            .O(n4_adj_4111));   // verilog/motorControl.v(42[17:23])
    defparam i22789_3_lut_4_lut.LUT_INIT = 16'hf880;
    SB_CARRY add_4143_6 (.CI(n29527), .I0(n8792[3]), .I1(n402_adj_4288), 
            .CO(n29528));
    SB_LUT4 unary_minus_5_inv_0_i1_1_lut (.I0(IntegralLimit[0]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4332[0]));   // verilog/motorControl.v(39[48:62])
    defparam unary_minus_5_inv_0_i1_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_668_7 (.CI(n27975), .I0(n3265[5]), .I1(n3290[5]), .CO(n27976));
    SB_LUT4 i22809_2_lut_3_lut_4_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err [21]), 
            .I2(\PID_CONTROLLER.err [20]), .I3(\Kp[1] ), .O(n27621));   // verilog/motorControl.v(42[17:23])
    defparam i22809_2_lut_3_lut_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 add_4143_5_lut (.I0(GND_net), .I1(n8792[2]), .I2(n329_adj_4287), 
            .I3(n29526), .O(n8779[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4143_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i22807_2_lut_3_lut_4_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err [21]), 
            .I2(\PID_CONTROLLER.err [20]), .I3(\Kp[1] ), .O(n8558[0]));   // verilog/motorControl.v(42[17:23])
    defparam i22807_2_lut_3_lut_4_lut.LUT_INIT = 16'h7888;
    SB_LUT4 mult_10_i651_2_lut (.I0(\Kp[13] ), .I1(\PID_CONTROLLER.err [6]), 
            .I2(GND_net), .I3(GND_net), .O(n968_adj_4282));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i651_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i467_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral [12]), 
            .I2(GND_net), .I3(GND_net), .O(n694_adj_4281));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i467_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i594_2_lut (.I0(\Ki[12] ), .I1(\PID_CONTROLLER.integral [2]), 
            .I2(GND_net), .I3(GND_net), .O(n883_adj_4280));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i594_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i700_2_lut (.I0(\Kp[14] ), .I1(\PID_CONTROLLER.err [6]), 
            .I2(GND_net), .I3(GND_net), .O(n1041_adj_4279));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i700_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i516_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral [12]), 
            .I2(GND_net), .I3(GND_net), .O(n767_adj_4278));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i516_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_666_i8_3_lut (.I0(n155[7]), .I1(PWMLimit[7]), .I2(n256), 
            .I3(GND_net), .O(n3290[7]));   // verilog/motorControl.v(46[16] 48[10])
    defparam mux_666_i8_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 add_4115_10_lut (.I0(GND_net), .I1(n8402[7]), .I2(n676_adj_4285), 
            .I3(n29207), .O(n8383[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4115_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i2_4_lut_adj_854 (.I0(n4_adj_4095), .I1(\Ki[3] ), .I2(n8855[1]), 
            .I3(\PID_CONTROLLER.integral [19]), .O(n8849[2]));   // verilog/motorControl.v(42[26:37])
    defparam i2_4_lut_adj_854.LUT_INIT = 16'h965a;
    SB_LUT4 mult_11_i330_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral [17]), 
            .I2(GND_net), .I3(GND_net), .O(n490));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i330_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i2_4_lut_adj_855 (.I0(\Ki[0] ), .I1(\Ki[3] ), .I2(\PID_CONTROLLER.integral [23]), 
            .I3(\PID_CONTROLLER.integral [20]), .O(n12_adj_4300));   // verilog/motorControl.v(42[26:37])
    defparam i2_4_lut_adj_855.LUT_INIT = 16'h9c50;
    SB_CARRY add_4143_5 (.CI(n29526), .I0(n8792[2]), .I1(n329_adj_4287), 
            .CO(n29527));
    SB_LUT4 i22926_4_lut (.I0(n8849[2]), .I1(\Ki[4] ), .I2(n6_adj_4046), 
            .I3(\PID_CONTROLLER.integral [18]), .O(n8_adj_4301));   // verilog/motorControl.v(42[26:37])
    defparam i22926_4_lut.LUT_INIT = 16'he8a0;
    SB_LUT4 add_4143_4_lut (.I0(GND_net), .I1(n8792[1]), .I2(n256_adj_4277), 
            .I3(n29525), .O(n8779[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4143_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_4_lut_adj_856 (.I0(\Ki[4] ), .I1(\Ki[2] ), .I2(\PID_CONTROLLER.integral [19]), 
            .I3(\PID_CONTROLLER.integral [21]), .O(n11_adj_4302));   // verilog/motorControl.v(42[26:37])
    defparam i1_4_lut_adj_856.LUT_INIT = 16'h6ca0;
    SB_LUT4 i22957_4_lut (.I0(n8855[1]), .I1(\Ki[3] ), .I2(n4_adj_4095), 
            .I3(\PID_CONTROLLER.integral [19]), .O(n6_adj_4303));   // verilog/motorControl.v(42[26:37])
    defparam i22957_4_lut.LUT_INIT = 16'he8a0;
    SB_LUT4 i22992_4_lut (.I0(\Ki[0] ), .I1(\Ki[1] ), .I2(\PID_CONTROLLER.integral [22]), 
            .I3(\PID_CONTROLLER.integral [21]), .O(n27816));   // verilog/motorControl.v(42[26:37])
    defparam i22992_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i8_4_lut_adj_857 (.I0(n6_adj_4303), .I1(n11_adj_4302), .I2(n8_adj_4301), 
            .I3(n12_adj_4300), .O(n18_adj_4304));   // verilog/motorControl.v(42[26:37])
    defparam i8_4_lut_adj_857.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_858 (.I0(\Ki[5] ), .I1(\Ki[1] ), .I2(\PID_CONTROLLER.integral [18]), 
            .I3(\PID_CONTROLLER.integral [22]), .O(n13_adj_4305));   // verilog/motorControl.v(42[26:37])
    defparam i3_4_lut_adj_858.LUT_INIT = 16'h6ca0;
    SB_LUT4 i9_4_lut_adj_859 (.I0(n13_adj_4305), .I1(n18_adj_4304), .I2(n27816), 
            .I3(n4_adj_4096), .O(n35470));   // verilog/motorControl.v(42[26:37])
    defparam i9_4_lut_adj_859.LUT_INIT = 16'h6996;
    SB_LUT4 add_4133_9_lut (.I0(GND_net), .I1(n8617[6]), .I2(n591_adj_4276), 
            .I3(n29375), .O(n8594[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4133_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4115_10 (.CI(n29207), .I0(n8402[7]), .I1(n676_adj_4285), 
            .CO(n29208));
    SB_CARRY add_4133_9 (.CI(n29375), .I0(n8617[6]), .I1(n591_adj_4276), 
            .CO(n29376));
    SB_LUT4 add_4115_9_lut (.I0(GND_net), .I1(n8402[6]), .I2(n603_adj_4274), 
            .I3(n29206), .O(n8383[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4115_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4143_4 (.CI(n29525), .I0(n8792[1]), .I1(n256_adj_4277), 
            .CO(n29526));
    SB_CARRY add_4115_9 (.CI(n29206), .I0(n8402[6]), .I1(n603_adj_4274), 
            .CO(n29207));
    SB_LUT4 add_4143_3_lut (.I0(GND_net), .I1(n8792[0]), .I2(n183_adj_4273), 
            .I3(n29524), .O(n8779[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4143_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4115_8_lut (.I0(GND_net), .I1(n8402[5]), .I2(n530_adj_4272), 
            .I3(n29205), .O(n8383[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4115_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4133_8_lut (.I0(GND_net), .I1(n8617[5]), .I2(n518_adj_4271), 
            .I3(n29374), .O(n8594[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4133_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4143_3 (.CI(n29524), .I0(n8792[0]), .I1(n183_adj_4273), 
            .CO(n29525));
    SB_LUT4 add_4143_2_lut (.I0(GND_net), .I1(n41_adj_4270), .I2(n110_adj_4269), 
            .I3(GND_net), .O(n8779[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4143_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_15_i35_2_lut (.I0(duty[17]), .I1(n257[17]), .I2(GND_net), 
            .I3(GND_net), .O(n35_adj_4003));   // verilog/motorControl.v(46[19:35])
    defparam LessThan_15_i35_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mux_666_i1_4_lut_4_lut (.I0(\PID_CONTROLLER.integral [0]), .I1(PWMLimit[0]), 
            .I2(n256), .I3(\Ki[0] ), .O(n3290[0]));   // verilog/motorControl.v(46[16] 48[10])
    defparam mux_666_i1_4_lut_4_lut.LUT_INIT = 16'h3a30;
    SB_LUT4 add_668_6_lut (.I0(GND_net), .I1(n3265[4]), .I2(n3290[4]), 
            .I3(n27974), .O(duty_23__N_3613[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_668_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4133_8 (.CI(n29374), .I0(n8617[5]), .I1(n518_adj_4271), 
            .CO(n29375));
    SB_CARRY add_4115_8 (.CI(n29205), .I0(n8402[5]), .I1(n530_adj_4272), 
            .CO(n29206));
    SB_CARRY add_4143_2 (.CI(GND_net), .I0(n41_adj_4270), .I1(n110_adj_4269), 
            .CO(n29524));
    SB_LUT4 unary_minus_5_inv_0_i15_1_lut (.I0(IntegralLimit[14]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4332[14]));   // verilog/motorControl.v(39[48:62])
    defparam unary_minus_5_inv_0_i15_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_4142_13_lut (.I0(GND_net), .I1(n8779[10]), .I2(n910_adj_4268), 
            .I3(n29523), .O(n8765[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4142_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_15_i31_2_lut (.I0(duty[15]), .I1(n257[15]), .I2(GND_net), 
            .I3(GND_net), .O(n31_adj_4073));   // verilog/motorControl.v(46[19:35])
    defparam LessThan_15_i31_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_4142_12_lut (.I0(GND_net), .I1(n8779[9]), .I2(n837_adj_4267), 
            .I3(n29522), .O(n8765[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4142_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4142_12 (.CI(n29522), .I0(n8779[9]), .I1(n837_adj_4267), 
            .CO(n29523));
    SB_LUT4 add_4142_11_lut (.I0(GND_net), .I1(n8779[8]), .I2(n764_adj_4266), 
            .I3(n29521), .O(n8765[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4142_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4133_7_lut (.I0(GND_net), .I1(n8617[4]), .I2(n445_adj_4265), 
            .I3(n29373), .O(n8594[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4133_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4115_7_lut (.I0(GND_net), .I1(n8402[4]), .I2(n457_adj_4264), 
            .I3(n29204), .O(n8383[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4115_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4133_7 (.CI(n29373), .I0(n8617[4]), .I1(n445_adj_4265), 
            .CO(n29374));
    SB_CARRY add_4115_7 (.CI(n29204), .I0(n8402[4]), .I1(n457_adj_4264), 
            .CO(n29205));
    SB_LUT4 add_4115_6_lut (.I0(GND_net), .I1(n8402[3]), .I2(n384_adj_4262), 
            .I3(n29203), .O(n8383[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4115_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4142_11 (.CI(n29521), .I0(n8779[8]), .I1(n764_adj_4266), 
            .CO(n29522));
    SB_LUT4 add_4133_6_lut (.I0(GND_net), .I1(n8617[3]), .I2(n372_adj_4261), 
            .I3(n29372), .O(n8594[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4133_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4115_6 (.CI(n29203), .I0(n8402[3]), .I1(n384_adj_4262), 
            .CO(n29204));
    SB_LUT4 add_4115_5_lut (.I0(GND_net), .I1(n8402[2]), .I2(n311_adj_4260), 
            .I3(n29202), .O(n8383[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4115_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4133_6 (.CI(n29372), .I0(n8617[3]), .I1(n372_adj_4261), 
            .CO(n29373));
    SB_CARRY add_4115_5 (.CI(n29202), .I0(n8402[2]), .I1(n311_adj_4260), 
            .CO(n29203));
    SB_LUT4 add_4115_4_lut (.I0(GND_net), .I1(n8402[1]), .I2(n238_adj_4259), 
            .I3(n29201), .O(n8383[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4115_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4142_10_lut (.I0(GND_net), .I1(n8779[7]), .I2(n691_adj_4258), 
            .I3(n29520), .O(n8765[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4142_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4133_5_lut (.I0(GND_net), .I1(n8617[2]), .I2(n299_adj_4257), 
            .I3(n29371), .O(n8594[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4133_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4115_4 (.CI(n29201), .I0(n8402[1]), .I1(n238_adj_4259), 
            .CO(n29202));
    SB_CARRY add_4133_5 (.CI(n29371), .I0(n8617[2]), .I1(n299_adj_4257), 
            .CO(n29372));
    SB_LUT4 add_4115_3_lut (.I0(GND_net), .I1(n8402[0]), .I2(n165_adj_4256), 
            .I3(n29200), .O(n8383[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4115_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4142_10 (.CI(n29520), .I0(n8779[7]), .I1(n691_adj_4258), 
            .CO(n29521));
    SB_LUT4 add_4133_4_lut (.I0(GND_net), .I1(n8617[1]), .I2(n226_adj_4255), 
            .I3(n29370), .O(n8594[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4133_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4115_3 (.CI(n29200), .I0(n8402[0]), .I1(n165_adj_4256), 
            .CO(n29201));
    SB_LUT4 LessThan_15_i33_2_lut (.I0(duty[16]), .I1(n257[16]), .I2(GND_net), 
            .I3(GND_net), .O(n33_adj_4004));   // verilog/motorControl.v(46[19:35])
    defparam LessThan_15_i33_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_4133_4 (.CI(n29370), .I0(n8617[1]), .I1(n226_adj_4255), 
            .CO(n29371));
    SB_LUT4 add_4115_2_lut (.I0(GND_net), .I1(n23_adj_4253), .I2(n92_adj_4252), 
            .I3(GND_net), .O(n8383[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4115_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_15_i29_2_lut (.I0(duty[14]), .I1(n257[14]), .I2(GND_net), 
            .I3(GND_net), .O(n29_adj_4071));   // verilog/motorControl.v(46[19:35])
    defparam LessThan_15_i29_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_4142_9_lut (.I0(GND_net), .I1(n8779[6]), .I2(n618_adj_4251), 
            .I3(n29519), .O(n8765[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4142_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4133_3_lut (.I0(GND_net), .I1(n8617[0]), .I2(n153_adj_4250), 
            .I3(n29369), .O(n8594[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4133_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4115_2 (.CI(GND_net), .I0(n23_adj_4253), .I1(n92_adj_4252), 
            .CO(n29200));
    SB_CARRY add_668_6 (.CI(n27974), .I0(n3265[4]), .I1(n3290[4]), .CO(n27975));
    SB_LUT4 mult_10_i518_2_lut (.I0(\Kp[10] ), .I1(\PID_CONTROLLER.err [13]), 
            .I2(GND_net), .I3(GND_net), .O(n770));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i518_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_15_i27_2_lut (.I0(duty[13]), .I1(n257[13]), .I2(GND_net), 
            .I3(GND_net), .O(n27_adj_4058));   // verilog/motorControl.v(46[19:35])
    defparam LessThan_15_i27_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_4114_19_lut (.I0(GND_net), .I1(n8383[16]), .I2(GND_net), 
            .I3(n29199), .O(n8363[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4114_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_668_5_lut (.I0(GND_net), .I1(n3265[3]), .I2(n3290[3]), 
            .I3(n27973), .O(duty_23__N_3613[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_668_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 IntegralLimit_23__I_0_i17_2_lut (.I0(\PID_CONTROLLER.integral [8]), 
            .I1(IntegralLimit[8]), .I2(GND_net), .I3(GND_net), .O(n17_adj_4306));   // verilog/motorControl.v(39[10:34])
    defparam IntegralLimit_23__I_0_i17_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 IntegralLimit_23__I_0_i9_2_lut (.I0(\PID_CONTROLLER.integral [4]), 
            .I1(IntegralLimit[4]), .I2(GND_net), .I3(GND_net), .O(n9_adj_4307));   // verilog/motorControl.v(39[10:34])
    defparam IntegralLimit_23__I_0_i9_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_4133_3 (.CI(n29369), .I0(n8617[0]), .I1(n153_adj_4250), 
            .CO(n29370));
    SB_LUT4 add_4114_18_lut (.I0(GND_net), .I1(n8383[15]), .I2(GND_net), 
            .I3(n29198), .O(n8363[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4114_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 IntegralLimit_23__I_0_i11_2_lut (.I0(\PID_CONTROLLER.integral [5]), 
            .I1(IntegralLimit[5]), .I2(GND_net), .I3(GND_net), .O(n11_adj_4308));   // verilog/motorControl.v(39[10:34])
    defparam IntegralLimit_23__I_0_i11_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i30716_4_lut (.I0(\PID_CONTROLLER.integral [3]), .I1(\PID_CONTROLLER.integral [2]), 
            .I2(IntegralLimit[3]), .I3(IntegralLimit[2]), .O(n37397));
    defparam i30716_4_lut.LUT_INIT = 16'h7bde;
    SB_CARRY add_4114_18 (.CI(n29198), .I0(n8383[15]), .I1(GND_net), .CO(n29199));
    SB_LUT4 i30712_3_lut (.I0(n11_adj_4308), .I1(n9_adj_4307), .I2(n37397), 
            .I3(GND_net), .O(n37393));
    defparam i30712_3_lut.LUT_INIT = 16'habab;
    SB_LUT4 IntegralLimit_23__I_0_i13_rep_342_2_lut (.I0(\PID_CONTROLLER.integral [6]), 
            .I1(IntegralLimit[6]), .I2(GND_net), .I3(GND_net), .O(n39123));   // verilog/motorControl.v(39[10:34])
    defparam IntegralLimit_23__I_0_i13_rep_342_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_668_5 (.CI(n27973), .I0(n3265[3]), .I1(n3290[3]), .CO(n27974));
    SB_LUT4 i31217_4_lut (.I0(\PID_CONTROLLER.integral [7]), .I1(n39123), 
            .I2(IntegralLimit[7]), .I3(n37393), .O(n37899));
    defparam i31217_4_lut.LUT_INIT = 16'hffde;
    SB_LUT4 i31001_4_lut (.I0(\PID_CONTROLLER.integral [9]), .I1(n17_adj_4306), 
            .I2(IntegralLimit[9]), .I3(n37899), .O(n37683));
    defparam i31001_4_lut.LUT_INIT = 16'hdeff;
    SB_LUT4 add_668_4_lut (.I0(GND_net), .I1(n3265[2]), .I2(n3290[2]), 
            .I3(n27972), .O(duty_23__N_3613[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_668_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4142_9 (.CI(n29519), .I0(n8779[6]), .I1(n618_adj_4251), 
            .CO(n29520));
    SB_LUT4 add_4133_2_lut (.I0(GND_net), .I1(n11_adj_4249), .I2(n80_adj_4248), 
            .I3(GND_net), .O(n8594[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4133_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4114_17_lut (.I0(GND_net), .I1(n8383[14]), .I2(GND_net), 
            .I3(n29197), .O(n8363[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4114_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i22776_2_lut_4_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err [20]), 
            .I2(\Kp[1] ), .I3(\PID_CONTROLLER.err [19]), .O(n8552[0]));   // verilog/motorControl.v(42[17:23])
    defparam i22776_2_lut_4_lut.LUT_INIT = 16'h7888;
    SB_LUT4 IntegralLimit_23__I_0_i21_rep_324_2_lut (.I0(\PID_CONTROLLER.integral [10]), 
            .I1(IntegralLimit[10]), .I2(GND_net), .I3(GND_net), .O(n39105));   // verilog/motorControl.v(39[10:34])
    defparam IntegralLimit_23__I_0_i21_rep_324_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i30999_4_lut (.I0(\PID_CONTROLLER.integral [9]), .I1(n17_adj_4306), 
            .I2(IntegralLimit[9]), .I3(n9_adj_4307), .O(n37681));
    defparam i30999_4_lut.LUT_INIT = 16'hffde;
    SB_LUT4 i30783_4_lut (.I0(n21_adj_3923), .I1(n19_adj_3924), .I2(n17_adj_3925), 
            .I3(n9_adj_3918), .O(n37464));
    defparam i30783_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i30997_4_lut (.I0(\PID_CONTROLLER.integral [11]), .I1(n39105), 
            .I2(IntegralLimit[11]), .I3(n37681), .O(n37679));
    defparam i30997_4_lut.LUT_INIT = 16'hdeff;
    SB_LUT4 IntegralLimit_23__I_0_i25_rep_317_2_lut (.I0(\PID_CONTROLLER.integral [12]), 
            .I1(IntegralLimit[12]), .I2(GND_net), .I3(GND_net), .O(n39098));   // verilog/motorControl.v(39[10:34])
    defparam IntegralLimit_23__I_0_i25_rep_317_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i30921_4_lut (.I0(n27_adj_4052), .I1(n15_adj_4109), .I2(n13_adj_4110), 
            .I3(n11_adj_4184), .O(n37603));
    defparam i30921_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i30927_4_lut (.I0(n21_adj_4100), .I1(n19_adj_4103), .I2(n17_adj_4105), 
            .I3(n9_adj_4231), .O(n37609));
    defparam i30927_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 \PID_CONTROLLER.integral_23__I_0_i16_3_lut  (.I0(\PID_CONTROLLER.integral [9]), 
            .I1(\PID_CONTROLLER.integral [21]), .I2(n43_adj_3997), .I3(GND_net), 
            .O(n16_adj_4309));   // verilog/motorControl.v(39[38:63])
    defparam \PID_CONTROLLER.integral_23__I_0_i16_3_lut .LUT_INIT = 16'hcaca;
    SB_LUT4 i30878_2_lut (.I0(n43_adj_3997), .I1(n19_adj_4103), .I2(GND_net), 
            .I3(GND_net), .O(n37560));
    defparam i30878_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 \PID_CONTROLLER.integral_23__I_0_i8_3_lut  (.I0(\PID_CONTROLLER.integral [4]), 
            .I1(\PID_CONTROLLER.integral [8]), .I2(n17_adj_4105), .I3(GND_net), 
            .O(n8_adj_4310));   // verilog/motorControl.v(39[38:63])
    defparam \PID_CONTROLLER.integral_23__I_0_i8_3_lut .LUT_INIT = 16'hcaca;
    SB_LUT4 i30775_4_lut (.I0(n27_adj_4058), .I1(n15_adj_3921), .I2(n13_adj_3920), 
            .I3(n11_adj_3919), .O(n37456));
    defparam i30775_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 \PID_CONTROLLER.integral_23__I_0_i24_3_lut  (.I0(n16_adj_4309), 
            .I1(\PID_CONTROLLER.integral [22]), .I2(n45_adj_3983), .I3(GND_net), 
            .O(n24_adj_4311));   // verilog/motorControl.v(39[38:63])
    defparam \PID_CONTROLLER.integral_23__I_0_i24_3_lut .LUT_INIT = 16'hcaca;
    SB_LUT4 i30943_2_lut (.I0(n7_adj_4233), .I1(n5_adj_4254), .I2(GND_net), 
            .I3(GND_net), .O(n37625));
    defparam i30943_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 add_4142_8_lut (.I0(GND_net), .I1(n8779[5]), .I2(n545_adj_4247), 
            .I3(n29518), .O(n8765[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4142_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4133_2 (.CI(GND_net), .I0(n11_adj_4249), .I1(n80_adj_4248), 
            .CO(n29369));
    SB_LUT4 LessThan_15_i12_3_lut (.I0(n257[7]), .I1(n257[16]), .I2(n33_adj_4004), 
            .I3(GND_net), .O(n12_adj_4312));   // verilog/motorControl.v(46[19:35])
    defparam LessThan_15_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_668_4 (.CI(n27972), .I0(n3265[2]), .I1(n3290[2]), .CO(n27973));
    SB_CARRY add_4114_17 (.CI(n29197), .I0(n8383[14]), .I1(GND_net), .CO(n29198));
    SB_CARRY add_4142_8 (.CI(n29518), .I0(n8779[5]), .I1(n545_adj_4247), 
            .CO(n29519));
    SB_LUT4 mult_11_add_1225_24_lut (.I0(\PID_CONTROLLER.integral [23]), .I1(n8570[21]), 
            .I2(GND_net), .I3(n29368), .O(n37312)) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_24_lut.LUT_INIT = 16'h6996;
    SB_LUT4 add_4114_16_lut (.I0(GND_net), .I1(n8383[13]), .I2(n1111_adj_4246), 
            .I3(n29196), .O(n8363[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4114_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4114_16 (.CI(n29196), .I0(n8383[13]), .I1(n1111_adj_4246), 
            .CO(n29197));
    SB_LUT4 mult_11_add_1225_23_lut (.I0(GND_net), .I1(n8570[20]), .I2(GND_net), 
            .I3(n29367), .O(n155[22])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4142_7_lut (.I0(GND_net), .I1(n8779[4]), .I2(n472_adj_4245), 
            .I3(n29517), .O(n8765[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4142_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4142_7 (.CI(n29517), .I0(n8779[4]), .I1(n472_adj_4245), 
            .CO(n29518));
    SB_CARRY mult_11_add_1225_23 (.CI(n29367), .I0(n8570[20]), .I1(GND_net), 
            .CO(n29368));
    SB_LUT4 i31189_4_lut (.I0(n13_adj_4110), .I1(n11_adj_4184), .I2(n9_adj_4231), 
            .I3(n37625), .O(n37871));
    defparam i31189_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i31185_4_lut (.I0(n19_adj_4103), .I1(n17_adj_4105), .I2(n15_adj_4109), 
            .I3(n37871), .O(n37867));
    defparam i31185_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 LessThan_15_i10_3_lut (.I0(n257[5]), .I1(n257[6]), .I2(n13_adj_3920), 
            .I3(GND_net), .O(n10_adj_4076));   // verilog/motorControl.v(46[19:35])
    defparam LessThan_15_i10_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i31401_4_lut (.I0(n25_adj_4055), .I1(n23_adj_4085), .I2(n21_adj_4100), 
            .I3(n37867), .O(n38083));
    defparam i31401_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 add_4142_6_lut (.I0(GND_net), .I1(n8779[3]), .I2(n399_adj_4244), 
            .I3(n29516), .O(n8765[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4142_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_add_1225_22_lut (.I0(GND_net), .I1(n8570[19]), .I2(GND_net), 
            .I3(n29366), .O(n155[21])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4114_15_lut (.I0(GND_net), .I1(n8383[12]), .I2(n1038_adj_4243), 
            .I3(n29195), .O(n8363[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4114_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i31293_4_lut (.I0(n31_adj_4026), .I1(n29_adj_4050), .I2(n27_adj_4052), 
            .I3(n38083), .O(n37975));
    defparam i31293_4_lut.LUT_INIT = 16'hfeff;
    SB_CARRY mult_11_add_1225_22 (.CI(n29366), .I0(n8570[19]), .I1(GND_net), 
            .CO(n29367));
    SB_LUT4 add_668_3_lut (.I0(GND_net), .I1(n3265[1]), .I2(n3290[1]), 
            .I3(n27971), .O(duty_23__N_3613[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_668_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_15_i30_3_lut (.I0(n12_adj_4312), .I1(n257[17]), .I2(n35_adj_4003), 
            .I3(GND_net), .O(n30_adj_4075));   // verilog/motorControl.v(46[19:35])
    defparam LessThan_15_i30_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_11_add_1225_21_lut (.I0(GND_net), .I1(n8570[18]), .I2(GND_net), 
            .I3(n29365), .O(n155[20])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4114_15 (.CI(n29195), .I0(n8383[12]), .I1(n1038_adj_4243), 
            .CO(n29196));
    SB_LUT4 \PID_CONTROLLER.integral_1526_add_4_25_lut  (.I0(GND_net), .I1(\PID_CONTROLLER.err [23]), 
            .I2(\PID_CONTROLLER.integral [23]), .I3(n28498), .O(n28[23])) /* synthesis syn_instantiated=1 */ ;
    defparam \PID_CONTROLLER.integral_1526_add_4_25_lut .LUT_INIT = 16'hC33C;
    SB_LUT4 \PID_CONTROLLER.integral_1526_add_4_24_lut  (.I0(GND_net), .I1(\PID_CONTROLLER.err [22]), 
            .I2(\PID_CONTROLLER.integral [22]), .I3(n28497), .O(n28[22])) /* synthesis syn_instantiated=1 */ ;
    defparam \PID_CONTROLLER.integral_1526_add_4_24_lut .LUT_INIT = 16'hC33C;
    SB_CARRY \PID_CONTROLLER.integral_1526_add_4_24  (.CI(n28497), .I0(\PID_CONTROLLER.err [22]), 
            .I1(\PID_CONTROLLER.integral [22]), .CO(n28498));
    SB_LUT4 \PID_CONTROLLER.integral_1526_add_4_23_lut  (.I0(GND_net), .I1(\PID_CONTROLLER.err [21]), 
            .I2(\PID_CONTROLLER.integral [21]), .I3(n28496), .O(n28[21])) /* synthesis syn_instantiated=1 */ ;
    defparam \PID_CONTROLLER.integral_1526_add_4_23_lut .LUT_INIT = 16'hC33C;
    SB_CARRY \PID_CONTROLLER.integral_1526_add_4_23  (.CI(n28496), .I0(\PID_CONTROLLER.err [21]), 
            .I1(\PID_CONTROLLER.integral [21]), .CO(n28497));
    SB_LUT4 \PID_CONTROLLER.integral_1526_add_4_22_lut  (.I0(GND_net), .I1(\PID_CONTROLLER.err [20]), 
            .I2(\PID_CONTROLLER.integral [20]), .I3(n28495), .O(n28[20])) /* synthesis syn_instantiated=1 */ ;
    defparam \PID_CONTROLLER.integral_1526_add_4_22_lut .LUT_INIT = 16'hC33C;
    SB_CARRY \PID_CONTROLLER.integral_1526_add_4_22  (.CI(n28495), .I0(\PID_CONTROLLER.err [20]), 
            .I1(\PID_CONTROLLER.integral [20]), .CO(n28496));
    SB_LUT4 \PID_CONTROLLER.integral_1526_add_4_21_lut  (.I0(GND_net), .I1(\PID_CONTROLLER.err [19]), 
            .I2(\PID_CONTROLLER.integral [19]), .I3(n28494), .O(n28[19])) /* synthesis syn_instantiated=1 */ ;
    defparam \PID_CONTROLLER.integral_1526_add_4_21_lut .LUT_INIT = 16'hC33C;
    SB_CARRY \PID_CONTROLLER.integral_1526_add_4_21  (.CI(n28494), .I0(\PID_CONTROLLER.err [19]), 
            .I1(\PID_CONTROLLER.integral [19]), .CO(n28495));
    SB_LUT4 \PID_CONTROLLER.integral_1526_add_4_20_lut  (.I0(GND_net), .I1(\PID_CONTROLLER.err [18]), 
            .I2(\PID_CONTROLLER.integral [18]), .I3(n28493), .O(n28[18])) /* synthesis syn_instantiated=1 */ ;
    defparam \PID_CONTROLLER.integral_1526_add_4_20_lut .LUT_INIT = 16'hC33C;
    SB_LUT4 add_4114_14_lut (.I0(GND_net), .I1(n8383[11]), .I2(n965_adj_4242), 
            .I3(n29194), .O(n8363[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4114_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY \PID_CONTROLLER.integral_1526_add_4_20  (.CI(n28493), .I0(\PID_CONTROLLER.err [18]), 
            .I1(\PID_CONTROLLER.integral [18]), .CO(n28494));
    SB_CARRY add_4142_6 (.CI(n29516), .I0(n8779[3]), .I1(n399_adj_4244), 
            .CO(n29517));
    SB_LUT4 \PID_CONTROLLER.integral_1526_add_4_19_lut  (.I0(GND_net), .I1(\PID_CONTROLLER.err [17]), 
            .I2(\PID_CONTROLLER.integral [17]), .I3(n28492), .O(n28[17])) /* synthesis syn_instantiated=1 */ ;
    defparam \PID_CONTROLLER.integral_1526_add_4_19_lut .LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_21 (.CI(n29365), .I0(n8570[18]), .I1(GND_net), 
            .CO(n29366));
    SB_LUT4 mult_11_add_1225_20_lut (.I0(GND_net), .I1(n8570[17]), .I2(GND_net), 
            .I3(n29364), .O(n155[19])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4114_14 (.CI(n29194), .I0(n8383[11]), .I1(n965_adj_4242), 
            .CO(n29195));
    SB_LUT4 add_4114_13_lut (.I0(GND_net), .I1(n8383[10]), .I2(n892_adj_4241), 
            .I3(n29193), .O(n8363[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4114_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY \PID_CONTROLLER.integral_1526_add_4_19  (.CI(n28492), .I0(\PID_CONTROLLER.err [17]), 
            .I1(\PID_CONTROLLER.integral [17]), .CO(n28493));
    SB_CARRY add_4114_13 (.CI(n29193), .I0(n8383[10]), .I1(n892_adj_4241), 
            .CO(n29194));
    SB_LUT4 \PID_CONTROLLER.integral_1526_add_4_18_lut  (.I0(GND_net), .I1(\PID_CONTROLLER.err [16]), 
            .I2(\PID_CONTROLLER.integral [16]), .I3(n28491), .O(n28[16])) /* synthesis syn_instantiated=1 */ ;
    defparam \PID_CONTROLLER.integral_1526_add_4_18_lut .LUT_INIT = 16'hC33C;
    SB_CARRY \PID_CONTROLLER.integral_1526_add_4_18  (.CI(n28491), .I0(\PID_CONTROLLER.err [16]), 
            .I1(\PID_CONTROLLER.integral [16]), .CO(n28492));
    SB_LUT4 \PID_CONTROLLER.integral_1526_add_4_17_lut  (.I0(GND_net), .I1(\PID_CONTROLLER.err [15]), 
            .I2(\PID_CONTROLLER.integral [15]), .I3(n28490), .O(n28[15])) /* synthesis syn_instantiated=1 */ ;
    defparam \PID_CONTROLLER.integral_1526_add_4_17_lut .LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_20 (.CI(n29364), .I0(n8570[17]), .I1(GND_net), 
            .CO(n29365));
    SB_CARRY \PID_CONTROLLER.integral_1526_add_4_17  (.CI(n28490), .I0(\PID_CONTROLLER.err [15]), 
            .I1(\PID_CONTROLLER.integral [15]), .CO(n28491));
    SB_LUT4 add_4142_5_lut (.I0(GND_net), .I1(n8779[2]), .I2(n326_adj_4240), 
            .I3(n29515), .O(n8765[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4142_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_add_1225_19_lut (.I0(GND_net), .I1(n8570[16]), .I2(GND_net), 
            .I3(n29363), .O(n155[18])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i31425_4_lut (.I0(n37_adj_4020), .I1(n35_adj_4023), .I2(n33_adj_4025), 
            .I3(n37975), .O(n38107));
    defparam i31425_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 \PID_CONTROLLER.integral_1526_add_4_16_lut  (.I0(GND_net), .I1(\PID_CONTROLLER.err [14]), 
            .I2(\PID_CONTROLLER.integral [14]), .I3(n28489), .O(n28[14])) /* synthesis syn_instantiated=1 */ ;
    defparam \PID_CONTROLLER.integral_1526_add_4_16_lut .LUT_INIT = 16'hC33C;
    SB_LUT4 add_4114_12_lut (.I0(GND_net), .I1(n8383[9]), .I2(n819_adj_4239), 
            .I3(n29192), .O(n8363[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4114_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY \PID_CONTROLLER.integral_1526_add_4_16  (.CI(n28489), .I0(\PID_CONTROLLER.err [14]), 
            .I1(\PID_CONTROLLER.integral [14]), .CO(n28490));
    SB_LUT4 i31003_4_lut (.I0(\PID_CONTROLLER.integral [7]), .I1(n39123), 
            .I2(IntegralLimit[7]), .I3(n11_adj_4308), .O(n37685));
    defparam i31003_4_lut.LUT_INIT = 16'hffde;
    SB_CARRY add_4142_5 (.CI(n29515), .I0(n8779[2]), .I1(n326_adj_4240), 
            .CO(n29516));
    SB_CARRY mult_11_add_1225_19 (.CI(n29363), .I0(n8570[16]), .I1(GND_net), 
            .CO(n29364));
    SB_LUT4 \PID_CONTROLLER.integral_1526_add_4_15_lut  (.I0(GND_net), .I1(\PID_CONTROLLER.err [13]), 
            .I2(\PID_CONTROLLER.integral [13]), .I3(n28488), .O(n28[13])) /* synthesis syn_instantiated=1 */ ;
    defparam \PID_CONTROLLER.integral_1526_add_4_15_lut .LUT_INIT = 16'hC33C;
    SB_CARRY \PID_CONTROLLER.integral_1526_add_4_15  (.CI(n28488), .I0(\PID_CONTROLLER.err [13]), 
            .I1(\PID_CONTROLLER.integral [13]), .CO(n28489));
    SB_LUT4 add_4142_4_lut (.I0(GND_net), .I1(n8779[1]), .I2(n253_adj_4238), 
            .I3(n29514), .O(n8765[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4142_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_add_1225_18_lut (.I0(GND_net), .I1(n8570[15]), .I2(GND_net), 
            .I3(n29362), .O(n155[17])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 \PID_CONTROLLER.integral_1526_add_4_14_lut  (.I0(GND_net), .I1(\PID_CONTROLLER.err [12]), 
            .I2(\PID_CONTROLLER.integral [12]), .I3(n28487), .O(n28[12])) /* synthesis syn_instantiated=1 */ ;
    defparam \PID_CONTROLLER.integral_1526_add_4_14_lut .LUT_INIT = 16'hC33C;
    SB_LUT4 i30742_2_lut_4_lut (.I0(duty[21]), .I1(n257[21]), .I2(duty[9]), 
            .I3(n257[9]), .O(n37423));
    defparam i30742_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_CARRY \PID_CONTROLLER.integral_1526_add_4_14  (.CI(n28487), .I0(\PID_CONTROLLER.err [12]), 
            .I1(\PID_CONTROLLER.integral [12]), .CO(n28488));
    SB_DFFE \PID_CONTROLLER.integral_1526__i1  (.Q(\PID_CONTROLLER.integral [1]), 
            .C(clk32MHz), .E(\PID_CONTROLLER.integral_23__N_3586 ), .D(n28[1]));   // verilog/motorControl.v(40[21:33])
    SB_LUT4 IntegralLimit_23__I_0_i27_rep_311_2_lut (.I0(\PID_CONTROLLER.integral [13]), 
            .I1(IntegralLimit[13]), .I2(GND_net), .I3(GND_net), .O(n39092));   // verilog/motorControl.v(39[10:34])
    defparam IntegralLimit_23__I_0_i27_rep_311_2_lut.LUT_INIT = 16'h6666;
    SB_DFFE \PID_CONTROLLER.integral_1526__i2  (.Q(\PID_CONTROLLER.integral [2]), 
            .C(clk32MHz), .E(\PID_CONTROLLER.integral_23__N_3586 ), .D(n28[2]));   // verilog/motorControl.v(40[21:33])
    SB_DFFE \PID_CONTROLLER.integral_1526__i3  (.Q(\PID_CONTROLLER.integral [3]), 
            .C(clk32MHz), .E(\PID_CONTROLLER.integral_23__N_3586 ), .D(n28[3]));   // verilog/motorControl.v(40[21:33])
    SB_DFFE \PID_CONTROLLER.integral_1526__i4  (.Q(\PID_CONTROLLER.integral [4]), 
            .C(clk32MHz), .E(\PID_CONTROLLER.integral_23__N_3586 ), .D(n28[4]));   // verilog/motorControl.v(40[21:33])
    SB_DFFE \PID_CONTROLLER.integral_1526__i5  (.Q(\PID_CONTROLLER.integral [5]), 
            .C(clk32MHz), .E(\PID_CONTROLLER.integral_23__N_3586 ), .D(n28[5]));   // verilog/motorControl.v(40[21:33])
    SB_DFFE \PID_CONTROLLER.integral_1526__i6  (.Q(\PID_CONTROLLER.integral [6]), 
            .C(clk32MHz), .E(\PID_CONTROLLER.integral_23__N_3586 ), .D(n28[6]));   // verilog/motorControl.v(40[21:33])
    SB_DFFE \PID_CONTROLLER.integral_1526__i7  (.Q(\PID_CONTROLLER.integral [7]), 
            .C(clk32MHz), .E(\PID_CONTROLLER.integral_23__N_3586 ), .D(n28[7]));   // verilog/motorControl.v(40[21:33])
    SB_DFFE \PID_CONTROLLER.integral_1526__i8  (.Q(\PID_CONTROLLER.integral [8]), 
            .C(clk32MHz), .E(\PID_CONTROLLER.integral_23__N_3586 ), .D(n28[8]));   // verilog/motorControl.v(40[21:33])
    SB_DFFE \PID_CONTROLLER.integral_1526__i9  (.Q(\PID_CONTROLLER.integral [9]), 
            .C(clk32MHz), .E(\PID_CONTROLLER.integral_23__N_3586 ), .D(n28[9]));   // verilog/motorControl.v(40[21:33])
    SB_DFFE \PID_CONTROLLER.integral_1526__i10  (.Q(\PID_CONTROLLER.integral [10]), 
            .C(clk32MHz), .E(\PID_CONTROLLER.integral_23__N_3586 ), .D(n28[10]));   // verilog/motorControl.v(40[21:33])
    SB_DFFE \PID_CONTROLLER.integral_1526__i11  (.Q(\PID_CONTROLLER.integral [11]), 
            .C(clk32MHz), .E(\PID_CONTROLLER.integral_23__N_3586 ), .D(n28[11]));   // verilog/motorControl.v(40[21:33])
    SB_DFFE \PID_CONTROLLER.integral_1526__i12  (.Q(\PID_CONTROLLER.integral [12]), 
            .C(clk32MHz), .E(\PID_CONTROLLER.integral_23__N_3586 ), .D(n28[12]));   // verilog/motorControl.v(40[21:33])
    SB_DFFE \PID_CONTROLLER.integral_1526__i13  (.Q(\PID_CONTROLLER.integral [13]), 
            .C(clk32MHz), .E(\PID_CONTROLLER.integral_23__N_3586 ), .D(n28[13]));   // verilog/motorControl.v(40[21:33])
    SB_DFFE \PID_CONTROLLER.integral_1526__i14  (.Q(\PID_CONTROLLER.integral [14]), 
            .C(clk32MHz), .E(\PID_CONTROLLER.integral_23__N_3586 ), .D(n28[14]));   // verilog/motorControl.v(40[21:33])
    SB_DFFE \PID_CONTROLLER.integral_1526__i15  (.Q(\PID_CONTROLLER.integral [15]), 
            .C(clk32MHz), .E(\PID_CONTROLLER.integral_23__N_3586 ), .D(n28[15]));   // verilog/motorControl.v(40[21:33])
    SB_DFFE \PID_CONTROLLER.integral_1526__i16  (.Q(\PID_CONTROLLER.integral [16]), 
            .C(clk32MHz), .E(\PID_CONTROLLER.integral_23__N_3586 ), .D(n28[16]));   // verilog/motorControl.v(40[21:33])
    SB_DFFE \PID_CONTROLLER.integral_1526__i17  (.Q(\PID_CONTROLLER.integral [17]), 
            .C(clk32MHz), .E(\PID_CONTROLLER.integral_23__N_3586 ), .D(n28[17]));   // verilog/motorControl.v(40[21:33])
    SB_DFFE \PID_CONTROLLER.integral_1526__i18  (.Q(\PID_CONTROLLER.integral [18]), 
            .C(clk32MHz), .E(\PID_CONTROLLER.integral_23__N_3586 ), .D(n28[18]));   // verilog/motorControl.v(40[21:33])
    SB_DFFE \PID_CONTROLLER.integral_1526__i19  (.Q(\PID_CONTROLLER.integral [19]), 
            .C(clk32MHz), .E(\PID_CONTROLLER.integral_23__N_3586 ), .D(n28[19]));   // verilog/motorControl.v(40[21:33])
    SB_DFFE \PID_CONTROLLER.integral_1526__i20  (.Q(\PID_CONTROLLER.integral [20]), 
            .C(clk32MHz), .E(\PID_CONTROLLER.integral_23__N_3586 ), .D(n28[20]));   // verilog/motorControl.v(40[21:33])
    SB_DFFE \PID_CONTROLLER.integral_1526__i21  (.Q(\PID_CONTROLLER.integral [21]), 
            .C(clk32MHz), .E(\PID_CONTROLLER.integral_23__N_3586 ), .D(n28[21]));   // verilog/motorControl.v(40[21:33])
    SB_DFFE \PID_CONTROLLER.integral_1526__i22  (.Q(\PID_CONTROLLER.integral [22]), 
            .C(clk32MHz), .E(\PID_CONTROLLER.integral_23__N_3586 ), .D(n28[22]));   // verilog/motorControl.v(40[21:33])
    SB_DFFE \PID_CONTROLLER.integral_1526__i23  (.Q(\PID_CONTROLLER.integral [23]), 
            .C(clk32MHz), .E(\PID_CONTROLLER.integral_23__N_3586 ), .D(n28[23]));   // verilog/motorControl.v(40[21:33])
    SB_LUT4 \PID_CONTROLLER.integral_1526_add_4_13_lut  (.I0(GND_net), .I1(\PID_CONTROLLER.err [11]), 
            .I2(\PID_CONTROLLER.integral [11]), .I3(n28486), .O(n28[11])) /* synthesis syn_instantiated=1 */ ;
    defparam \PID_CONTROLLER.integral_1526_add_4_13_lut .LUT_INIT = 16'hC33C;
    SB_LUT4 i31209_4_lut (.I0(\PID_CONTROLLER.integral [14]), .I1(n39092), 
            .I2(IntegralLimit[14]), .I3(n37685), .O(n37891));
    defparam i31209_4_lut.LUT_INIT = 16'hdeff;
    SB_LUT4 IntegralLimit_23__I_0_i31_rep_306_2_lut (.I0(\PID_CONTROLLER.integral [15]), 
            .I1(IntegralLimit[15]), .I2(GND_net), .I3(GND_net), .O(n39087));   // verilog/motorControl.v(39[10:34])
    defparam IntegralLimit_23__I_0_i31_rep_306_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY \PID_CONTROLLER.integral_1526_add_4_13  (.CI(n28486), .I0(\PID_CONTROLLER.err [11]), 
            .I1(\PID_CONTROLLER.integral [11]), .CO(n28487));
    SB_LUT4 \PID_CONTROLLER.integral_1526_add_4_12_lut  (.I0(GND_net), .I1(\PID_CONTROLLER.err [10]), 
            .I2(\PID_CONTROLLER.integral [10]), .I3(n28485), .O(n28[10])) /* synthesis syn_instantiated=1 */ ;
    defparam \PID_CONTROLLER.integral_1526_add_4_12_lut .LUT_INIT = 16'hC33C;
    SB_LUT4 IntegralLimit_23__I_0_i12_3_lut (.I0(IntegralLimit[7]), .I1(IntegralLimit[16]), 
            .I2(\PID_CONTROLLER.integral [16]), .I3(GND_net), .O(n12_adj_4320));   // verilog/motorControl.v(39[10:34])
    defparam IntegralLimit_23__I_0_i12_3_lut.LUT_INIT = 16'h8e8e;
    SB_CARRY add_4142_4 (.CI(n29514), .I0(n8779[1]), .I1(n253_adj_4238), 
            .CO(n29515));
    SB_CARRY add_4114_12 (.CI(n29192), .I0(n8383[9]), .I1(n819_adj_4239), 
            .CO(n29193));
    SB_CARRY mult_11_add_1225_18 (.CI(n29362), .I0(n8570[15]), .I1(GND_net), 
            .CO(n29363));
    SB_LUT4 add_4114_11_lut (.I0(GND_net), .I1(n8383[8]), .I2(n746_adj_4235), 
            .I3(n29191), .O(n8363[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4114_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i30971_4_lut (.I0(\PID_CONTROLLER.integral [16]), .I1(\PID_CONTROLLER.integral [7]), 
            .I2(IntegralLimit[16]), .I3(IntegralLimit[7]), .O(n37653));
    defparam i30971_4_lut.LUT_INIT = 16'h7bde;
    SB_CARRY \PID_CONTROLLER.integral_1526_add_4_12  (.CI(n28485), .I0(\PID_CONTROLLER.err [10]), 
            .I1(\PID_CONTROLLER.integral [10]), .CO(n28486));
    SB_LUT4 IntegralLimit_23__I_0_i35_rep_329_2_lut (.I0(\PID_CONTROLLER.integral [17]), 
            .I1(IntegralLimit[17]), .I2(GND_net), .I3(GND_net), .O(n39110));   // verilog/motorControl.v(39[10:34])
    defparam IntegralLimit_23__I_0_i35_rep_329_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 \PID_CONTROLLER.integral_1526_add_4_11_lut  (.I0(GND_net), .I1(\PID_CONTROLLER.err [9]), 
            .I2(\PID_CONTROLLER.integral [9]), .I3(n28484), .O(n28[9])) /* synthesis syn_instantiated=1 */ ;
    defparam \PID_CONTROLLER.integral_1526_add_4_11_lut .LUT_INIT = 16'hC33C;
    SB_LUT4 IntegralLimit_23__I_0_i10_3_lut (.I0(IntegralLimit[5]), .I1(IntegralLimit[6]), 
            .I2(\PID_CONTROLLER.integral [6]), .I3(GND_net), .O(n10_adj_4321));   // verilog/motorControl.v(39[10:34])
    defparam IntegralLimit_23__I_0_i10_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 IntegralLimit_23__I_0_i30_3_lut (.I0(n12_adj_4320), .I1(IntegralLimit[17]), 
            .I2(\PID_CONTROLLER.integral [17]), .I3(GND_net), .O(n30_adj_4322));   // verilog/motorControl.v(39[10:34])
    defparam IntegralLimit_23__I_0_i30_3_lut.LUT_INIT = 16'h8e8e;
    SB_CARRY \PID_CONTROLLER.integral_1526_add_4_11  (.CI(n28484), .I0(\PID_CONTROLLER.err [9]), 
            .I1(\PID_CONTROLLER.integral [9]), .CO(n28485));
    SB_LUT4 add_4142_3_lut (.I0(GND_net), .I1(n8779[0]), .I2(n180_adj_4234), 
            .I3(n29513), .O(n8765[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4142_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_add_1225_17_lut (.I0(GND_net), .I1(n8570[14]), .I2(GND_net), 
            .I3(n29361), .O(n155[16])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4114_11 (.CI(n29191), .I0(n8383[8]), .I1(n746_adj_4235), 
            .CO(n29192));
    SB_LUT4 i31311_4_lut (.I0(\PID_CONTROLLER.integral [11]), .I1(n39105), 
            .I2(IntegralLimit[11]), .I3(n37683), .O(n37993));
    defparam i31311_4_lut.LUT_INIT = 16'hffde;
    SB_LUT4 \PID_CONTROLLER.integral_1526_add_4_10_lut  (.I0(GND_net), .I1(\PID_CONTROLLER.err [8]), 
            .I2(\PID_CONTROLLER.integral [8]), .I3(n28483), .O(n28[8])) /* synthesis syn_instantiated=1 */ ;
    defparam \PID_CONTROLLER.integral_1526_add_4_10_lut .LUT_INIT = 16'hC33C;
    SB_CARRY \PID_CONTROLLER.integral_1526_add_4_10  (.CI(n28483), .I0(\PID_CONTROLLER.err [8]), 
            .I1(\PID_CONTROLLER.integral [8]), .CO(n28484));
    SB_CARRY add_668_3 (.CI(n27971), .I0(n3265[1]), .I1(n3290[1]), .CO(n27972));
    SB_LUT4 \PID_CONTROLLER.integral_1526_add_4_9_lut  (.I0(GND_net), .I1(\PID_CONTROLLER.err [7]), 
            .I2(\PID_CONTROLLER.integral [7]), .I3(n28482), .O(n28[7])) /* synthesis syn_instantiated=1 */ ;
    defparam \PID_CONTROLLER.integral_1526_add_4_9_lut .LUT_INIT = 16'hC33C;
    SB_CARRY add_4142_3 (.CI(n29513), .I0(n8779[0]), .I1(n180_adj_4234), 
            .CO(n29514));
    SB_CARRY \PID_CONTROLLER.integral_1526_add_4_9  (.CI(n28482), .I0(\PID_CONTROLLER.err [7]), 
            .I1(\PID_CONTROLLER.integral [7]), .CO(n28483));
    SB_CARRY mult_11_add_1225_17 (.CI(n29361), .I0(n8570[14]), .I1(GND_net), 
            .CO(n29362));
    SB_LUT4 mult_11_add_1225_16_lut (.I0(GND_net), .I1(n8570[13]), .I2(n1096_adj_4232), 
            .I3(n29360), .O(n155[15])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4114_10_lut (.I0(GND_net), .I1(n8383[7]), .I2(n673_adj_4230), 
            .I3(n29190), .O(n8363[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4114_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 \PID_CONTROLLER.integral_1526_add_4_8_lut  (.I0(GND_net), .I1(\PID_CONTROLLER.err [6]), 
            .I2(\PID_CONTROLLER.integral [6]), .I3(n28481), .O(n28[6])) /* synthesis syn_instantiated=1 */ ;
    defparam \PID_CONTROLLER.integral_1526_add_4_8_lut .LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_16 (.CI(n29360), .I0(n8570[13]), .I1(n1096_adj_4232), 
            .CO(n29361));
    SB_CARRY add_4114_10 (.CI(n29190), .I0(n8383[7]), .I1(n673_adj_4230), 
            .CO(n29191));
    SB_LUT4 add_4114_9_lut (.I0(GND_net), .I1(n8383[6]), .I2(n600_adj_4229), 
            .I3(n29189), .O(n8363[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4114_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY \PID_CONTROLLER.integral_1526_add_4_8  (.CI(n28481), .I0(\PID_CONTROLLER.err [6]), 
            .I1(\PID_CONTROLLER.integral [6]), .CO(n28482));
    SB_LUT4 \PID_CONTROLLER.integral_1526_add_4_7_lut  (.I0(GND_net), .I1(\PID_CONTROLLER.err [5]), 
            .I2(\PID_CONTROLLER.integral [5]), .I3(n28480), .O(n28[5])) /* synthesis syn_instantiated=1 */ ;
    defparam \PID_CONTROLLER.integral_1526_add_4_7_lut .LUT_INIT = 16'hC33C;
    SB_CARRY \PID_CONTROLLER.integral_1526_add_4_7  (.CI(n28480), .I0(\PID_CONTROLLER.err [5]), 
            .I1(\PID_CONTROLLER.integral [5]), .CO(n28481));
    SB_LUT4 \PID_CONTROLLER.integral_1526_add_4_6_lut  (.I0(GND_net), .I1(\PID_CONTROLLER.err [4]), 
            .I2(\PID_CONTROLLER.integral [4]), .I3(n28479), .O(n28[4])) /* synthesis syn_instantiated=1 */ ;
    defparam \PID_CONTROLLER.integral_1526_add_4_6_lut .LUT_INIT = 16'hC33C;
    SB_CARRY \PID_CONTROLLER.integral_1526_add_4_6  (.CI(n28479), .I0(\PID_CONTROLLER.err [4]), 
            .I1(\PID_CONTROLLER.integral [4]), .CO(n28480));
    SB_LUT4 \PID_CONTROLLER.integral_1526_add_4_5_lut  (.I0(GND_net), .I1(\PID_CONTROLLER.err [3]), 
            .I2(\PID_CONTROLLER.integral [3]), .I3(n28478), .O(n28[3])) /* synthesis syn_instantiated=1 */ ;
    defparam \PID_CONTROLLER.integral_1526_add_4_5_lut .LUT_INIT = 16'hC33C;
    SB_CARRY \PID_CONTROLLER.integral_1526_add_4_5  (.CI(n28478), .I0(\PID_CONTROLLER.err [3]), 
            .I1(\PID_CONTROLLER.integral [3]), .CO(n28479));
    SB_CARRY add_4114_9 (.CI(n29189), .I0(n8383[6]), .I1(n600_adj_4229), 
            .CO(n29190));
    SB_LUT4 \PID_CONTROLLER.integral_1526_add_4_4_lut  (.I0(GND_net), .I1(\PID_CONTROLLER.err [2]), 
            .I2(\PID_CONTROLLER.integral [2]), .I3(n28477), .O(n28[2])) /* synthesis syn_instantiated=1 */ ;
    defparam \PID_CONTROLLER.integral_1526_add_4_4_lut .LUT_INIT = 16'hC33C;
    SB_CARRY \PID_CONTROLLER.integral_1526_add_4_4  (.CI(n28477), .I0(\PID_CONTROLLER.err [2]), 
            .I1(\PID_CONTROLLER.integral [2]), .CO(n28478));
    SB_LUT4 \PID_CONTROLLER.integral_1526_add_4_3_lut  (.I0(GND_net), .I1(\PID_CONTROLLER.err [1]), 
            .I2(\PID_CONTROLLER.integral [1]), .I3(n28476), .O(n28[1])) /* synthesis syn_instantiated=1 */ ;
    defparam \PID_CONTROLLER.integral_1526_add_4_3_lut .LUT_INIT = 16'hC33C;
    SB_CARRY \PID_CONTROLLER.integral_1526_add_4_3  (.CI(n28476), .I0(\PID_CONTROLLER.err [1]), 
            .I1(\PID_CONTROLLER.integral [1]), .CO(n28477));
    SB_LUT4 \PID_CONTROLLER.integral_1526_add_4_2_lut  (.I0(GND_net), .I1(\PID_CONTROLLER.err [0]), 
            .I2(\PID_CONTROLLER.integral [0]), .I3(GND_net), .O(n28[0])) /* synthesis syn_instantiated=1 */ ;
    defparam \PID_CONTROLLER.integral_1526_add_4_2_lut .LUT_INIT = 16'hC33C;
    SB_LUT4 add_4142_2_lut (.I0(GND_net), .I1(n38_adj_4228), .I2(n107_adj_4227), 
            .I3(GND_net), .O(n8765[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4142_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4114_8_lut (.I0(GND_net), .I1(n8383[5]), .I2(n527_adj_4226), 
            .I3(n29188), .O(n8363[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4114_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY \PID_CONTROLLER.integral_1526_add_4_2  (.CI(GND_net), .I0(\PID_CONTROLLER.err [0]), 
            .I1(\PID_CONTROLLER.integral [0]), .CO(n28476));
    SB_LUT4 mult_11_add_1225_15_lut (.I0(GND_net), .I1(n8570[12]), .I2(n1023_adj_4225), 
            .I3(n29359), .O(n155[14])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4114_8 (.CI(n29188), .I0(n8383[5]), .I1(n527_adj_4226), 
            .CO(n29189));
    SB_CARRY add_4142_2 (.CI(GND_net), .I0(n38_adj_4228), .I1(n107_adj_4227), 
            .CO(n29513));
    SB_CARRY mult_11_add_1225_15 (.CI(n29359), .I0(n8570[12]), .I1(n1023_adj_4225), 
            .CO(n29360));
    SB_LUT4 add_4141_14_lut (.I0(GND_net), .I1(n8765[11]), .I2(n980_adj_4224), 
            .I3(n29512), .O(n8750[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4141_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_add_1225_14_lut (.I0(GND_net), .I1(n8570[11]), .I2(n950_adj_4223), 
            .I3(n29358), .O(n155[13])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4114_7_lut (.I0(GND_net), .I1(n8383[4]), .I2(n454_adj_4222), 
            .I3(n29187), .O(n8363[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4114_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_668_2_lut (.I0(GND_net), .I1(n3265[0]), .I2(n3290[0]), 
            .I3(GND_net), .O(duty_23__N_3613[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_668_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_14 (.CI(n29358), .I0(n8570[11]), .I1(n950_adj_4223), 
            .CO(n29359));
    SB_CARRY add_4114_7 (.CI(n29187), .I0(n8383[4]), .I1(n454_adj_4222), 
            .CO(n29188));
    SB_LUT4 add_4114_6_lut (.I0(GND_net), .I1(n8383[3]), .I2(n381_adj_4221), 
            .I3(n29186), .O(n8363[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4114_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4141_13_lut (.I0(GND_net), .I1(n8765[10]), .I2(n907_adj_4220), 
            .I3(n29511), .O(n8750[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4141_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4114_6 (.CI(n29186), .I0(n8383[3]), .I1(n381_adj_4221), 
            .CO(n29187));
    SB_LUT4 i30991_4_lut (.I0(\PID_CONTROLLER.integral [13]), .I1(n39098), 
            .I2(IntegralLimit[13]), .I3(n37993), .O(n37673));
    defparam i30991_4_lut.LUT_INIT = 16'h5a7b;
    SB_LUT4 i31106_4_lut (.I0(n13_adj_3920), .I1(n11_adj_3919), .I2(n9_adj_3918), 
            .I3(n37478), .O(n37788));
    defparam i31106_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 IntegralLimit_23__I_0_i29_rep_309_2_lut (.I0(\PID_CONTROLLER.integral [14]), 
            .I1(IntegralLimit[14]), .I2(GND_net), .I3(GND_net), .O(n39090));   // verilog/motorControl.v(39[10:34])
    defparam IntegralLimit_23__I_0_i29_rep_309_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_4141_13 (.CI(n29511), .I0(n8765[10]), .I1(n907_adj_4220), 
            .CO(n29512));
    SB_LUT4 mult_11_add_1225_13_lut (.I0(GND_net), .I1(n8570[10]), .I2(n877_adj_4219), 
            .I3(n29357), .O(n155[12])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_13 (.CI(n29357), .I0(n8570[10]), .I1(n877_adj_4219), 
            .CO(n29358));
    SB_LUT4 add_4114_5_lut (.I0(GND_net), .I1(n8383[2]), .I2(n308_adj_4218), 
            .I3(n29185), .O(n8363[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4114_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4141_12_lut (.I0(GND_net), .I1(n8765[9]), .I2(n834_adj_4217), 
            .I3(n29510), .O(n8750[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4141_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_add_1225_12_lut (.I0(GND_net), .I1(n8570[9]), .I2(n804_adj_4216), 
            .I3(n29356), .O(n155[11])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4114_5 (.CI(n29185), .I0(n8383[2]), .I1(n308_adj_4218), 
            .CO(n29186));
    SB_CARRY add_668_2 (.CI(GND_net), .I0(n3265[0]), .I1(n3290[0]), .CO(n27971));
    SB_LUT4 i30797_3_lut_4_lut (.I0(duty[3]), .I1(n257[3]), .I2(n257[2]), 
            .I3(duty[2]), .O(n37478));   // verilog/motorControl.v(46[19:35])
    defparam i30797_3_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 add_4114_4_lut (.I0(GND_net), .I1(n8383[1]), .I2(n235_adj_4215), 
            .I3(n29184), .O(n8363[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4114_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_15_i6_3_lut_3_lut (.I0(duty[3]), .I1(n257[3]), .I2(n257[2]), 
            .I3(GND_net), .O(n6_adj_4016));   // verilog/motorControl.v(46[19:35])
    defparam LessThan_15_i6_3_lut_3_lut.LUT_INIT = 16'hd4d4;
    SB_CARRY add_4141_12 (.CI(n29510), .I0(n8765[9]), .I1(n834_adj_4217), 
            .CO(n29511));
    SB_CARRY mult_11_add_1225_12 (.CI(n29356), .I0(n8570[9]), .I1(n804_adj_4216), 
            .CO(n29357));
    SB_LUT4 mult_11_add_1225_11_lut (.I0(GND_net), .I1(n8570[8]), .I2(n731_adj_4214), 
            .I3(n29355), .O(n155[10])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i31309_4_lut (.I0(\PID_CONTROLLER.integral [15]), .I1(n39090), 
            .I2(IntegralLimit[15]), .I3(n37673), .O(n37991));
    defparam i31309_4_lut.LUT_INIT = 16'hffde;
    SB_CARRY add_4114_4 (.CI(n29184), .I0(n8383[1]), .I1(n235_adj_4215), 
            .CO(n29185));
    SB_CARRY mult_11_add_1225_11 (.CI(n29355), .I0(n8570[8]), .I1(n731_adj_4214), 
            .CO(n29356));
    SB_LUT4 add_4114_3_lut (.I0(GND_net), .I1(n8383[0]), .I2(n162_adj_4213), 
            .I3(n29183), .O(n8363[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4114_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 IntegralLimit_23__I_0_i33_rep_335_2_lut (.I0(\PID_CONTROLLER.integral [16]), 
            .I1(IntegralLimit[16]), .I2(GND_net), .I3(GND_net), .O(n39116));   // verilog/motorControl.v(39[10:34])
    defparam IntegralLimit_23__I_0_i33_rep_335_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_4114_3 (.CI(n29183), .I0(n8383[0]), .I1(n162_adj_4213), 
            .CO(n29184));
    SB_LUT4 add_4114_2_lut (.I0(GND_net), .I1(n20_adj_4212), .I2(n89_adj_4211), 
            .I3(GND_net), .O(n8363[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4114_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4141_11_lut (.I0(GND_net), .I1(n8765[8]), .I2(n761_adj_4210), 
            .I3(n29509), .O(n8750[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4141_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_add_1225_10_lut (.I0(GND_net), .I1(n8570[7]), .I2(n658_adj_4209), 
            .I3(n29354), .O(n155[9])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4141_11 (.CI(n29509), .I0(n8765[8]), .I1(n761_adj_4210), 
            .CO(n29510));
    SB_CARRY add_4114_2 (.CI(GND_net), .I0(n20_adj_4212), .I1(n89_adj_4211), 
            .CO(n29183));
    SB_LUT4 i31405_4_lut (.I0(\PID_CONTROLLER.integral [17]), .I1(n39116), 
            .I2(IntegralLimit[17]), .I3(n37991), .O(n38087));
    defparam i31405_4_lut.LUT_INIT = 16'hffde;
    SB_LUT4 add_4113_20_lut (.I0(GND_net), .I1(n8363[17]), .I2(GND_net), 
            .I3(n29182), .O(n8342[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4113_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 IntegralLimit_23__I_0_i37_rep_300_2_lut (.I0(\PID_CONTROLLER.integral [18]), 
            .I1(IntegralLimit[18]), .I2(GND_net), .I3(GND_net), .O(n39081));   // verilog/motorControl.v(39[10:34])
    defparam IntegralLimit_23__I_0_i37_rep_300_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_4141_10_lut (.I0(GND_net), .I1(n8765[7]), .I2(n688_adj_4208), 
            .I3(n29508), .O(n8750[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4141_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_10 (.CI(n29354), .I0(n8570[7]), .I1(n658_adj_4209), 
            .CO(n29355));
    SB_LUT4 add_4113_19_lut (.I0(GND_net), .I1(n8363[16]), .I2(GND_net), 
            .I3(n29181), .O(n8342[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4113_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_add_1225_9_lut (.I0(GND_net), .I1(n8570[6]), .I2(n585_adj_4207), 
            .I3(n29353), .O(n155[8])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4113_19 (.CI(n29181), .I0(n8363[16]), .I1(GND_net), .CO(n29182));
    SB_LUT4 i31445_4_lut (.I0(\PID_CONTROLLER.integral [19]), .I1(n39081), 
            .I2(IntegralLimit[19]), .I3(n38087), .O(n38127));
    defparam i31445_4_lut.LUT_INIT = 16'hffde;
    SB_CARRY add_4141_10 (.CI(n29508), .I0(n8765[7]), .I1(n688_adj_4208), 
            .CO(n29509));
    SB_LUT4 add_4113_18_lut (.I0(GND_net), .I1(n8363[15]), .I2(GND_net), 
            .I3(n29180), .O(n8342[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4113_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4141_9_lut (.I0(GND_net), .I1(n8765[6]), .I2(n615_adj_4206), 
            .I3(n29507), .O(n8750[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4141_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4141_9 (.CI(n29507), .I0(n8765[6]), .I1(n615_adj_4206), 
            .CO(n29508));
    SB_LUT4 add_4141_8_lut (.I0(GND_net), .I1(n8765[5]), .I2(n542_adj_4205), 
            .I3(n29506), .O(n8750[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4141_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4113_18 (.CI(n29180), .I0(n8363[15]), .I1(GND_net), .CO(n29181));
    SB_CARRY mult_11_add_1225_9 (.CI(n29353), .I0(n8570[6]), .I1(n585_adj_4207), 
            .CO(n29354));
    SB_CARRY add_4141_8 (.CI(n29506), .I0(n8765[5]), .I1(n542_adj_4205), 
            .CO(n29507));
    SB_LUT4 add_4113_17_lut (.I0(GND_net), .I1(n8363[14]), .I2(GND_net), 
            .I3(n29179), .O(n8342[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4113_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4141_7_lut (.I0(GND_net), .I1(n8765[4]), .I2(n469_adj_4204), 
            .I3(n29505), .O(n8750[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4141_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 IntegralLimit_23__I_0_i41_rep_297_2_lut (.I0(\PID_CONTROLLER.integral [20]), 
            .I1(IntegralLimit[20]), .I2(GND_net), .I3(GND_net), .O(n39078));   // verilog/motorControl.v(39[10:34])
    defparam IntegralLimit_23__I_0_i41_rep_297_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_4113_17 (.CI(n29179), .I0(n8363[14]), .I1(GND_net), .CO(n29180));
    SB_LUT4 add_4113_16_lut (.I0(GND_net), .I1(n8363[13]), .I2(n1108_adj_4203), 
            .I3(n29178), .O(n8342[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4113_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_add_1225_8_lut (.I0(GND_net), .I1(n8570[5]), .I2(n512_adj_4202), 
            .I3(n29352), .O(n155[7])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4141_7 (.CI(n29505), .I0(n8765[4]), .I1(n469_adj_4204), 
            .CO(n29506));
    SB_CARRY add_4113_16 (.CI(n29178), .I0(n8363[13]), .I1(n1108_adj_4203), 
            .CO(n29179));
    SB_CARRY mult_11_add_1225_8 (.CI(n29352), .I0(n8570[5]), .I1(n512_adj_4202), 
            .CO(n29353));
    SB_LUT4 add_4113_15_lut (.I0(GND_net), .I1(n8363[12]), .I2(n1035_adj_4201), 
            .I3(n29177), .O(n8342[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4113_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_add_1225_7_lut (.I0(GND_net), .I1(n8570[4]), .I2(n439_adj_4200), 
            .I3(n29351), .O(n155[6])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4141_6_lut (.I0(GND_net), .I1(n8765[3]), .I2(n396_adj_4199), 
            .I3(n29504), .O(n8750[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4141_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_7 (.CI(n29351), .I0(n8570[4]), .I1(n439_adj_4200), 
            .CO(n29352));
    SB_CARRY add_4141_6 (.CI(n29504), .I0(n8765[3]), .I1(n396_adj_4199), 
            .CO(n29505));
    SB_CARRY add_4113_15 (.CI(n29177), .I0(n8363[12]), .I1(n1035_adj_4201), 
            .CO(n29178));
    SB_LUT4 IntegralLimit_23__I_0_i16_3_lut (.I0(IntegralLimit[9]), .I1(IntegralLimit[21]), 
            .I2(\PID_CONTROLLER.integral [21]), .I3(GND_net), .O(n16_adj_4323));   // verilog/motorControl.v(39[10:34])
    defparam IntegralLimit_23__I_0_i16_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 add_4113_14_lut (.I0(GND_net), .I1(n8363[11]), .I2(n962_adj_4198), 
            .I3(n29176), .O(n8342[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4113_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4113_14 (.CI(n29176), .I0(n8363[11]), .I1(n962_adj_4198), 
            .CO(n29177));
    SB_LUT4 mult_11_add_1225_6_lut (.I0(GND_net), .I1(n8570[3]), .I2(n366_adj_4197), 
            .I3(n29350), .O(n155[5])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4113_13_lut (.I0(GND_net), .I1(n8363[10]), .I2(n889_adj_4196), 
            .I3(n29175), .O(n8342[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4113_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4113_13 (.CI(n29175), .I0(n8363[10]), .I1(n889_adj_4196), 
            .CO(n29176));
    SB_LUT4 add_4113_12_lut (.I0(GND_net), .I1(n8363[9]), .I2(n816_adj_4195), 
            .I3(n29174), .O(n8342[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4113_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i30945_4_lut (.I0(\PID_CONTROLLER.integral [21]), .I1(\PID_CONTROLLER.integral [9]), 
            .I2(IntegralLimit[21]), .I3(IntegralLimit[9]), .O(n37627));
    defparam i30945_4_lut.LUT_INIT = 16'h7bde;
    SB_LUT4 unary_minus_16_add_3_25_lut (.I0(duty[23]), .I1(GND_net), .I2(n1[23]), 
            .I3(n28131), .O(n47_adj_4236)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_25_lut.LUT_INIT = 16'h6996;
    SB_LUT4 add_4141_5_lut (.I0(GND_net), .I1(n8765[2]), .I2(n323_adj_4193), 
            .I3(n29503), .O(n8750[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4141_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_6 (.CI(n29350), .I0(n8570[3]), .I1(n366_adj_4197), 
            .CO(n29351));
    SB_LUT4 mult_11_add_1225_5_lut (.I0(GND_net), .I1(n8570[2]), .I2(n293_adj_4192), 
            .I3(n29349), .O(n155[4])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4113_12 (.CI(n29174), .I0(n8363[9]), .I1(n816_adj_4195), 
            .CO(n29175));
    SB_LUT4 unary_minus_16_add_3_24_lut (.I0(GND_net), .I1(GND_net), .I2(n1[22]), 
            .I3(n28130), .O(n257[22])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4113_11_lut (.I0(GND_net), .I1(n8363[8]), .I2(n743_adj_4190), 
            .I3(n29173), .O(n8342[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4113_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4141_5 (.CI(n29503), .I0(n8765[2]), .I1(n323_adj_4193), 
            .CO(n29504));
    SB_CARRY add_4113_11 (.CI(n29173), .I0(n8363[8]), .I1(n743_adj_4190), 
            .CO(n29174));
    SB_CARRY mult_11_add_1225_5 (.CI(n29349), .I0(n8570[2]), .I1(n293_adj_4192), 
            .CO(n29350));
    SB_LUT4 mult_11_add_1225_4_lut (.I0(GND_net), .I1(n8570[1]), .I2(n220_adj_4189), 
            .I3(n29348), .O(n155[3])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4141_4_lut (.I0(GND_net), .I1(n8765[1]), .I2(n250_adj_4188), 
            .I3(n29502), .O(n8750[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4141_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_4 (.CI(n29348), .I0(n8570[1]), .I1(n220_adj_4189), 
            .CO(n29349));
    SB_LUT4 add_4113_10_lut (.I0(GND_net), .I1(n8363[7]), .I2(n670_adj_4187), 
            .I3(n29172), .O(n8342[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4113_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4141_4 (.CI(n29502), .I0(n8765[1]), .I1(n250_adj_4188), 
            .CO(n29503));
    SB_LUT4 mult_11_add_1225_3_lut (.I0(GND_net), .I1(n8570[0]), .I2(n147_adj_4186), 
            .I3(n29347), .O(n155[2])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4113_10 (.CI(n29172), .I0(n8363[7]), .I1(n670_adj_4187), 
            .CO(n29173));
    SB_LUT4 add_4113_9_lut (.I0(GND_net), .I1(n8363[6]), .I2(n597_adj_4185), 
            .I3(n29171), .O(n8342[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4113_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_3 (.CI(n29347), .I0(n8570[0]), .I1(n147_adj_4186), 
            .CO(n29348));
    SB_CARRY add_4113_9 (.CI(n29171), .I0(n8363[6]), .I1(n597_adj_4185), 
            .CO(n29172));
    SB_LUT4 mult_11_add_1225_2_lut (.I0(GND_net), .I1(n5_adj_4183), .I2(n74_adj_4182), 
            .I3(GND_net), .O(n155[1])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4141_3_lut (.I0(GND_net), .I1(n8765[0]), .I2(n177_adj_4181), 
            .I3(n29501), .O(n8750[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4141_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4113_8_lut (.I0(GND_net), .I1(n8363[5]), .I2(n524_adj_4180), 
            .I3(n29170), .O(n8342[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4113_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_2 (.CI(GND_net), .I0(n5_adj_4183), .I1(n74_adj_4182), 
            .CO(n29347));
    SB_CARRY add_4113_8 (.CI(n29170), .I0(n8363[5]), .I1(n524_adj_4180), 
            .CO(n29171));
    SB_LUT4 add_4113_7_lut (.I0(GND_net), .I1(n8363[4]), .I2(n451_adj_4179), 
            .I3(n29169), .O(n8342[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4113_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4132_23_lut (.I0(GND_net), .I1(n8594[20]), .I2(GND_net), 
            .I3(n29346), .O(n8570[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4132_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4141_3 (.CI(n29501), .I0(n8765[0]), .I1(n177_adj_4181), 
            .CO(n29502));
    SB_CARRY add_4113_7 (.CI(n29169), .I0(n8363[4]), .I1(n451_adj_4179), 
            .CO(n29170));
    SB_CARRY unary_minus_16_add_3_24 (.CI(n28130), .I0(GND_net), .I1(n1[22]), 
            .CO(n28131));
    SB_LUT4 add_4141_2_lut (.I0(GND_net), .I1(n35_adj_4178), .I2(n104_adj_4177), 
            .I3(GND_net), .O(n8750[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4141_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4132_22_lut (.I0(GND_net), .I1(n8594[19]), .I2(GND_net), 
            .I3(n29345), .O(n8570[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4132_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4113_6_lut (.I0(GND_net), .I1(n8363[3]), .I2(n378_adj_4176), 
            .I3(n29168), .O(n8342[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4113_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 IntegralLimit_23__I_0_i24_3_lut (.I0(n16_adj_4323), .I1(IntegralLimit[22]), 
            .I2(\PID_CONTROLLER.integral [22]), .I3(GND_net), .O(n24_adj_4324));   // verilog/motorControl.v(39[10:34])
    defparam IntegralLimit_23__I_0_i24_3_lut.LUT_INIT = 16'h8e8e;
    SB_CARRY add_4132_22 (.CI(n29345), .I0(n8594[19]), .I1(GND_net), .CO(n29346));
    SB_CARRY add_4113_6 (.CI(n29168), .I0(n8363[3]), .I1(n378_adj_4176), 
            .CO(n29169));
    SB_LUT4 add_4113_5_lut (.I0(GND_net), .I1(n8363[2]), .I2(n305_adj_4175), 
            .I3(n29167), .O(n8342[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4113_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 IntegralLimit_23__I_0_i6_3_lut (.I0(IntegralLimit[2]), .I1(IntegralLimit[3]), 
            .I2(\PID_CONTROLLER.integral [3]), .I3(GND_net), .O(n6_adj_4325));   // verilog/motorControl.v(39[10:34])
    defparam IntegralLimit_23__I_0_i6_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i31365_3_lut (.I0(n6_adj_4325), .I1(IntegralLimit[10]), .I2(\PID_CONTROLLER.integral [10]), 
            .I3(GND_net), .O(n38047));   // verilog/motorControl.v(39[10:34])
    defparam i31365_3_lut.LUT_INIT = 16'h8e8e;
    SB_CARRY add_4141_2 (.CI(GND_net), .I0(n35_adj_4178), .I1(n104_adj_4177), 
            .CO(n29501));
    SB_LUT4 add_4132_21_lut (.I0(GND_net), .I1(n8594[18]), .I2(GND_net), 
            .I3(n29344), .O(n8570[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4132_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4113_5 (.CI(n29167), .I0(n8363[2]), .I1(n305_adj_4175), 
            .CO(n29168));
    SB_LUT4 i31366_3_lut (.I0(n38047), .I1(IntegralLimit[11]), .I2(\PID_CONTROLLER.integral [11]), 
            .I3(GND_net), .O(n38048));   // verilog/motorControl.v(39[10:34])
    defparam i31366_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 add_4113_4_lut (.I0(GND_net), .I1(n8363[1]), .I2(n232_adj_4174), 
            .I3(n29166), .O(n8342[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4113_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4132_21 (.CI(n29344), .I0(n8594[18]), .I1(GND_net), .CO(n29345));
    SB_CARRY add_4113_4 (.CI(n29166), .I0(n8363[1]), .I1(n232_adj_4174), 
            .CO(n29167));
    SB_LUT4 i30950_4_lut (.I0(\PID_CONTROLLER.integral [21]), .I1(n39098), 
            .I2(IntegralLimit[21]), .I3(n37679), .O(n37632));
    defparam i30950_4_lut.LUT_INIT = 16'h5a7b;
    SB_LUT4 mult_10_i416_2_lut (.I0(\Kp[8] ), .I1(\PID_CONTROLLER.err [11]), 
            .I2(GND_net), .I3(GND_net), .O(n618));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i416_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_4140_15_lut (.I0(GND_net), .I1(n8750[12]), .I2(n1050_adj_4173), 
            .I3(n29500), .O(n8734[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4140_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4132_20_lut (.I0(GND_net), .I1(n8594[17]), .I2(GND_net), 
            .I3(n29343), .O(n8570[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4132_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4113_3_lut (.I0(GND_net), .I1(n8363[0]), .I2(n159_adj_4172), 
            .I3(n29165), .O(n8342[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4113_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i308_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral [6]), 
            .I2(GND_net), .I3(GND_net), .O(n457));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i308_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_4132_20 (.CI(n29343), .I0(n8594[17]), .I1(GND_net), .CO(n29344));
    SB_CARRY add_4113_3 (.CI(n29165), .I0(n8363[0]), .I1(n159_adj_4172), 
            .CO(n29166));
    SB_LUT4 mult_11_i357_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral [6]), 
            .I2(GND_net), .I3(GND_net), .O(n530));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i357_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i31243_4_lut (.I0(n24_adj_4324), .I1(n8_adj_4298), .I2(n39076), 
            .I3(n37627), .O(n37925));   // verilog/motorControl.v(39[10:34])
    defparam i31243_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 mult_11_i406_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral [6]), 
            .I2(GND_net), .I3(GND_net), .O(n603));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i406_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_4140_14_lut (.I0(GND_net), .I1(n8750[11]), .I2(n977_adj_4171), 
            .I3(n29499), .O(n8734[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4140_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4132_19_lut (.I0(GND_net), .I1(n8594[16]), .I2(GND_net), 
            .I3(n29342), .O(n8570[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4132_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4113_2_lut (.I0(GND_net), .I1(n17_adj_4170), .I2(n86_adj_4169), 
            .I3(GND_net), .O(n8342[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4113_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i465_2_lut (.I0(\Kp[9] ), .I1(\PID_CONTROLLER.err [11]), 
            .I2(GND_net), .I3(GND_net), .O(n691));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i465_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_4132_19 (.CI(n29342), .I0(n8594[16]), .I1(GND_net), .CO(n29343));
    SB_CARRY add_4113_2 (.CI(GND_net), .I0(n17_adj_4170), .I1(n86_adj_4169), 
            .CO(n29165));
    SB_CARRY add_4140_14 (.CI(n29499), .I0(n8750[11]), .I1(n977_adj_4171), 
            .CO(n29500));
    SB_LUT4 add_4132_18_lut (.I0(GND_net), .I1(n8594[15]), .I2(GND_net), 
            .I3(n29341), .O(n8570[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4132_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4112_21_lut (.I0(GND_net), .I1(n8342[18]), .I2(GND_net), 
            .I3(n29164), .O(n8320[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4112_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i31324_3_lut (.I0(n38048), .I1(IntegralLimit[12]), .I2(\PID_CONTROLLER.integral [12]), 
            .I3(GND_net), .O(n38006));   // verilog/motorControl.v(39[10:34])
    defparam i31324_3_lut.LUT_INIT = 16'h8e8e;
    SB_CARRY add_4132_18 (.CI(n29341), .I0(n8594[15]), .I1(GND_net), .CO(n29342));
    SB_LUT4 \PID_CONTROLLER.integral_23__I_0_i4_4_lut  (.I0(\PID_CONTROLLER.integral_23__N_3589 [0]), 
            .I1(\PID_CONTROLLER.integral [1]), .I2(n3_adj_4275), .I3(\PID_CONTROLLER.integral [0]), 
            .O(n4_adj_4326));   // verilog/motorControl.v(39[38:63])
    defparam \PID_CONTROLLER.integral_23__I_0_i4_4_lut .LUT_INIT = 16'hc5c0;
    SB_LUT4 add_4112_20_lut (.I0(GND_net), .I1(n8342[17]), .I2(GND_net), 
            .I3(n29163), .O(n8320[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4112_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_16_add_3_23_lut (.I0(GND_net), .I1(GND_net), .I2(n1[21]), 
            .I3(n28129), .O(n257[21])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i514_2_lut (.I0(\Kp[10] ), .I1(\PID_CONTROLLER.err [11]), 
            .I2(GND_net), .I3(GND_net), .O(n764));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i514_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_4140_13_lut (.I0(GND_net), .I1(n8750[10]), .I2(n904_adj_4167), 
            .I3(n29498), .O(n8734[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4140_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4132_17_lut (.I0(GND_net), .I1(n8594[14]), .I2(GND_net), 
            .I3(n29340), .O(n8570[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4132_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4112_20 (.CI(n29163), .I0(n8342[17]), .I1(GND_net), .CO(n29164));
    SB_LUT4 add_4112_19_lut (.I0(GND_net), .I1(n8342[16]), .I2(GND_net), 
            .I3(n29162), .O(n8320[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4112_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4132_17 (.CI(n29340), .I0(n8594[14]), .I1(GND_net), .CO(n29341));
    SB_CARRY add_4112_19 (.CI(n29162), .I0(n8342[16]), .I1(GND_net), .CO(n29163));
    SB_LUT4 add_4112_18_lut (.I0(GND_net), .I1(n8342[15]), .I2(GND_net), 
            .I3(n29161), .O(n8320[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4112_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4140_13 (.CI(n29498), .I0(n8750[10]), .I1(n904_adj_4167), 
            .CO(n29499));
    SB_LUT4 add_4132_16_lut (.I0(GND_net), .I1(n8594[13]), .I2(n1099_adj_4166), 
            .I3(n29339), .O(n8570[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4132_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4112_18 (.CI(n29161), .I0(n8342[15]), .I1(GND_net), .CO(n29162));
    SB_LUT4 i31102_4_lut (.I0(n19_adj_3924), .I1(n17_adj_3925), .I2(n15_adj_3921), 
            .I3(n37788), .O(n37784));
    defparam i31102_4_lut.LUT_INIT = 16'heeef;
    SB_CARRY add_4132_16 (.CI(n29339), .I0(n8594[13]), .I1(n1099_adj_4166), 
            .CO(n29340));
    SB_LUT4 add_4112_17_lut (.I0(GND_net), .I1(n8342[14]), .I2(GND_net), 
            .I3(n29160), .O(n8320[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4112_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i31343_3_lut (.I0(n4_adj_4326), .I1(\PID_CONTROLLER.integral [13]), 
            .I2(n27_adj_4052), .I3(GND_net), .O(n38025));   // verilog/motorControl.v(39[38:63])
    defparam i31343_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i31344_3_lut (.I0(n38025), .I1(\PID_CONTROLLER.integral [14]), 
            .I2(n29_adj_4050), .I3(GND_net), .O(n38026));   // verilog/motorControl.v(39[38:63])
    defparam i31344_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_4112_17 (.CI(n29160), .I0(n8342[14]), .I1(GND_net), .CO(n29161));
    SB_LUT4 \PID_CONTROLLER.integral_23__I_0_i12_3_lut  (.I0(\PID_CONTROLLER.integral [7]), 
            .I1(\PID_CONTROLLER.integral [16]), .I2(n33_adj_4025), .I3(GND_net), 
            .O(n12_adj_4327));   // verilog/motorControl.v(39[38:63])
    defparam \PID_CONTROLLER.integral_23__I_0_i12_3_lut .LUT_INIT = 16'hcaca;
    SB_LUT4 i30891_2_lut (.I0(n33_adj_4025), .I1(n15_adj_4109), .I2(GND_net), 
            .I3(GND_net), .O(n37573));
    defparam i30891_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 add_4140_12_lut (.I0(GND_net), .I1(n8750[9]), .I2(n831_adj_4165), 
            .I3(n29497), .O(n8734[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4140_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4132_15_lut (.I0(GND_net), .I1(n8594[12]), .I2(n1026_adj_4164), 
            .I3(n29338), .O(n8570[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4132_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4112_16_lut (.I0(GND_net), .I1(n8342[13]), .I2(n1105_adj_4163), 
            .I3(n29159), .O(n8320[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4112_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i563_2_lut (.I0(\Kp[11] ), .I1(\PID_CONTROLLER.err [11]), 
            .I2(GND_net), .I3(GND_net), .O(n837));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i563_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_4132_15 (.CI(n29338), .I0(n8594[12]), .I1(n1026_adj_4164), 
            .CO(n29339));
    SB_CARRY add_4112_16 (.CI(n29159), .I0(n8342[13]), .I1(n1105_adj_4163), 
            .CO(n29160));
    SB_LUT4 mult_11_i455_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral [6]), 
            .I2(GND_net), .I3(GND_net), .O(n676));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i455_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_4140_12 (.CI(n29497), .I0(n8750[9]), .I1(n831_adj_4165), 
            .CO(n29498));
    SB_LUT4 add_4132_14_lut (.I0(GND_net), .I1(n8594[11]), .I2(n953_adj_4162), 
            .I3(n29337), .O(n8570[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4132_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 \PID_CONTROLLER.integral_23__I_0_i10_3_lut  (.I0(\PID_CONTROLLER.integral [5]), 
            .I1(\PID_CONTROLLER.integral [6]), .I2(n13_adj_4110), .I3(GND_net), 
            .O(n10_adj_4328));   // verilog/motorControl.v(39[38:63])
    defparam \PID_CONTROLLER.integral_23__I_0_i10_3_lut .LUT_INIT = 16'hcaca;
    SB_LUT4 add_4112_15_lut (.I0(GND_net), .I1(n8342[12]), .I2(n1032_adj_4161), 
            .I3(n29158), .O(n8320[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4112_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4132_14 (.CI(n29337), .I0(n8594[11]), .I1(n953_adj_4162), 
            .CO(n29338));
    SB_LUT4 \PID_CONTROLLER.integral_23__I_0_i30_3_lut  (.I0(n12_adj_4327), 
            .I1(\PID_CONTROLLER.integral [17]), .I2(n35_adj_4023), .I3(GND_net), 
            .O(n30_adj_4329));   // verilog/motorControl.v(39[38:63])
    defparam \PID_CONTROLLER.integral_23__I_0_i30_3_lut .LUT_INIT = 16'hcaca;
    SB_CARRY add_4112_15 (.CI(n29158), .I0(n8342[12]), .I1(n1032_adj_4161), 
            .CO(n29159));
    SB_LUT4 i30893_4_lut (.I0(n33_adj_4025), .I1(n31_adj_4026), .I2(n29_adj_4050), 
            .I3(n37603), .O(n37575));
    defparam i30893_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i31409_4_lut (.I0(n30_adj_4329), .I1(n10_adj_4328), .I2(n35_adj_4023), 
            .I3(n37573), .O(n38091));   // verilog/motorControl.v(39[38:63])
    defparam i31409_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 add_4140_11_lut (.I0(GND_net), .I1(n8750[8]), .I2(n758_adj_4160), 
            .I3(n29496), .O(n8734[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4140_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4132_13_lut (.I0(GND_net), .I1(n8594[10]), .I2(n880_adj_4159), 
            .I3(n29336), .O(n8570[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4132_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4112_14_lut (.I0(GND_net), .I1(n8342[11]), .I2(n959_adj_4158), 
            .I3(n29157), .O(n8320[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4112_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4132_13 (.CI(n29336), .I0(n8594[10]), .I1(n880_adj_4159), 
            .CO(n29337));
    SB_CARRY add_4112_14 (.CI(n29157), .I0(n8342[11]), .I1(n959_adj_4158), 
            .CO(n29158));
    SB_CARRY add_4140_11 (.CI(n29496), .I0(n8750[8]), .I1(n758_adj_4160), 
            .CO(n29497));
    SB_LUT4 add_4132_12_lut (.I0(GND_net), .I1(n8594[9]), .I2(n807_adj_4157), 
            .I3(n29335), .O(n8570[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4132_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4112_13_lut (.I0(GND_net), .I1(n8342[10]), .I2(n886_adj_4156), 
            .I3(n29156), .O(n8320[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4112_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4112_13 (.CI(n29156), .I0(n8342[10]), .I1(n886_adj_4156), 
            .CO(n29157));
    SB_LUT4 i31054_3_lut (.I0(n38026), .I1(\PID_CONTROLLER.integral [15]), 
            .I2(n31_adj_4026), .I3(GND_net), .O(n37736));   // verilog/motorControl.v(39[38:63])
    defparam i31054_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i31449_4_lut (.I0(n37736), .I1(n38091), .I2(n35_adj_4023), 
            .I3(n37575), .O(n38131));   // verilog/motorControl.v(39[38:63])
    defparam i31449_4_lut.LUT_INIT = 16'hccca;
    SB_CARRY add_4132_12 (.CI(n29335), .I0(n8594[9]), .I1(n807_adj_4157), 
            .CO(n29336));
    SB_LUT4 add_4112_12_lut (.I0(GND_net), .I1(n8342[9]), .I2(n813_adj_4155), 
            .I3(n29155), .O(n8320[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4112_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4112_12 (.CI(n29155), .I0(n8342[9]), .I1(n813_adj_4155), 
            .CO(n29156));
    SB_LUT4 i31450_3_lut (.I0(n38131), .I1(\PID_CONTROLLER.integral [18]), 
            .I2(n37_adj_4020), .I3(GND_net), .O(n38132));   // verilog/motorControl.v(39[38:63])
    defparam i31450_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i31440_3_lut (.I0(n38132), .I1(\PID_CONTROLLER.integral [19]), 
            .I2(n39_adj_4014), .I3(GND_net), .O(n38122));   // verilog/motorControl.v(39[38:63])
    defparam i31440_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 \PID_CONTROLLER.integral_23__I_0_i6_3_lut  (.I0(\PID_CONTROLLER.integral [2]), 
            .I1(\PID_CONTROLLER.integral [3]), .I2(n7_adj_4233), .I3(GND_net), 
            .O(n6_adj_4330));   // verilog/motorControl.v(39[38:63])
    defparam \PID_CONTROLLER.integral_23__I_0_i6_3_lut .LUT_INIT = 16'hcaca;
    SB_LUT4 i31345_3_lut (.I0(n6_adj_4330), .I1(\PID_CONTROLLER.integral [10]), 
            .I2(n21_adj_4100), .I3(GND_net), .O(n38027));   // verilog/motorControl.v(39[38:63])
    defparam i31345_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i31346_3_lut (.I0(n38027), .I1(\PID_CONTROLLER.integral [11]), 
            .I2(n23_adj_4085), .I3(GND_net), .O(n38028));   // verilog/motorControl.v(39[38:63])
    defparam i31346_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i30880_4_lut (.I0(n43_adj_3997), .I1(n25_adj_4055), .I2(n23_adj_4085), 
            .I3(n37609), .O(n37562));
    defparam i30880_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 add_4140_10_lut (.I0(GND_net), .I1(n8750[7]), .I2(n685_adj_4154), 
            .I3(n29495), .O(n8734[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4140_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4132_11_lut (.I0(GND_net), .I1(n8594[8]), .I2(n734_adj_4153), 
            .I3(n29334), .O(n8570[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4132_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4112_11_lut (.I0(GND_net), .I1(n8342[8]), .I2(n740_adj_4152), 
            .I3(n29154), .O(n8320[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4112_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i31245_4_lut (.I0(n24_adj_4311), .I1(n8_adj_4310), .I2(n45_adj_3983), 
            .I3(n37560), .O(n37927));   // verilog/motorControl.v(39[38:63])
    defparam i31245_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i31052_3_lut (.I0(n38028), .I1(\PID_CONTROLLER.integral [12]), 
            .I2(n25_adj_4055), .I3(GND_net), .O(n37734));   // verilog/motorControl.v(39[38:63])
    defparam i31052_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_4132_11 (.CI(n29334), .I0(n8594[8]), .I1(n734_adj_4153), 
            .CO(n29335));
    SB_CARRY add_4112_11 (.CI(n29154), .I0(n8342[8]), .I1(n740_adj_4152), 
            .CO(n29155));
    SB_CARRY add_4140_10 (.CI(n29495), .I0(n8750[7]), .I1(n685_adj_4154), 
            .CO(n29496));
    SB_LUT4 add_4132_10_lut (.I0(GND_net), .I1(n8594[7]), .I2(n661_adj_4151), 
            .I3(n29333), .O(n8570[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4132_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4112_10_lut (.I0(GND_net), .I1(n8342[7]), .I2(n667_adj_4150), 
            .I3(n29153), .O(n8320[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4112_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i30882_4_lut (.I0(n43_adj_3997), .I1(n41_adj_4011), .I2(n39_adj_4014), 
            .I3(n38107), .O(n37564));
    defparam i30882_4_lut.LUT_INIT = 16'haaab;
    SB_CARRY add_4112_10 (.CI(n29153), .I0(n8342[7]), .I1(n667_adj_4150), 
            .CO(n29154));
    SB_CARRY add_4132_10 (.CI(n29333), .I0(n8594[7]), .I1(n661_adj_4151), 
            .CO(n29334));
    SB_LUT4 add_4140_9_lut (.I0(GND_net), .I1(n8750[6]), .I2(n612_adj_4149), 
            .I3(n29494), .O(n8734[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4140_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4112_9_lut (.I0(GND_net), .I1(n8342[6]), .I2(n594_adj_4148), 
            .I3(n29152), .O(n8320[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4112_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i31371_4_lut (.I0(n37734), .I1(n37927), .I2(n45_adj_3983), 
            .I3(n37562), .O(n38053));   // verilog/motorControl.v(39[38:63])
    defparam i31371_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i31060_3_lut (.I0(n38122), .I1(\PID_CONTROLLER.integral [20]), 
            .I2(n41_adj_4011), .I3(GND_net), .O(n37742));   // verilog/motorControl.v(39[38:63])
    defparam i31060_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY unary_minus_16_add_3_23 (.CI(n28129), .I0(GND_net), .I1(n1[21]), 
            .CO(n28130));
    SB_LUT4 mult_10_i612_2_lut (.I0(\Kp[12] ), .I1(\PID_CONTROLLER.err [11]), 
            .I2(GND_net), .I3(GND_net), .O(n910));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i612_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i504_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral [6]), 
            .I2(GND_net), .I3(GND_net), .O(n749));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i504_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_4140_9 (.CI(n29494), .I0(n8750[6]), .I1(n612_adj_4149), 
            .CO(n29495));
    SB_LUT4 add_4132_9_lut (.I0(GND_net), .I1(n8594[6]), .I2(n588_adj_4147), 
            .I3(n29332), .O(n8570[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4132_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4112_9 (.CI(n29152), .I0(n8342[6]), .I1(n594_adj_4148), 
            .CO(n29153));
    SB_CARRY add_4132_9 (.CI(n29332), .I0(n8594[6]), .I1(n588_adj_4147), 
            .CO(n29333));
    SB_LUT4 add_4112_8_lut (.I0(GND_net), .I1(n8342[5]), .I2(n521_adj_4146), 
            .I3(n29151), .O(n8320[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4112_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_16_add_3_22_lut (.I0(GND_net), .I1(GND_net), .I2(n1[20]), 
            .I3(n28128), .O(n257[20])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4140_8_lut (.I0(GND_net), .I1(n8750[5]), .I2(n539_adj_4144), 
            .I3(n29493), .O(n8734[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4140_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4112_8 (.CI(n29151), .I0(n8342[5]), .I1(n521_adj_4146), 
            .CO(n29152));
    SB_LUT4 i31417_4_lut (.I0(n37742), .I1(n38053), .I2(n45_adj_3983), 
            .I3(n37564), .O(n38099));   // verilog/motorControl.v(39[38:63])
    defparam i31417_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 add_4112_7_lut (.I0(GND_net), .I1(n8342[4]), .I2(n448_adj_4143), 
            .I3(n29150), .O(n8320[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4112_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4132_8_lut (.I0(GND_net), .I1(n8594[5]), .I2(n515_adj_4142), 
            .I3(n29331), .O(n8570[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4132_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4132_8 (.CI(n29331), .I0(n8594[5]), .I1(n515_adj_4142), 
            .CO(n29332));
    SB_CARRY add_4112_7 (.CI(n29150), .I0(n8342[4]), .I1(n448_adj_4143), 
            .CO(n29151));
    SB_LUT4 IntegralLimit_23__I_0_i4_4_lut (.I0(\PID_CONTROLLER.integral [0]), 
            .I1(IntegralLimit[1]), .I2(\PID_CONTROLLER.integral [1]), .I3(IntegralLimit[0]), 
            .O(n4_adj_4331));   // verilog/motorControl.v(39[10:34])
    defparam IntegralLimit_23__I_0_i4_4_lut.LUT_INIT = 16'h4d0c;
    SB_CARRY unary_minus_16_add_3_22 (.CI(n28128), .I0(GND_net), .I1(n1[20]), 
            .CO(n28129));
    SB_CARRY add_4140_8 (.CI(n29493), .I0(n8750[5]), .I1(n539_adj_4144), 
            .CO(n29494));
    SB_LUT4 add_4132_7_lut (.I0(GND_net), .I1(n8594[4]), .I2(n442_adj_4141), 
            .I3(n29330), .O(n8570[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4132_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4112_6_lut (.I0(GND_net), .I1(n8342[3]), .I2(n375_adj_4140), 
            .I3(n29149), .O(n8320[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4112_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4132_7 (.CI(n29330), .I0(n8594[4]), .I1(n442_adj_4141), 
            .CO(n29331));
    SB_CARRY add_4112_6 (.CI(n29149), .I0(n8342[3]), .I1(n375_adj_4140), 
            .CO(n29150));
    SB_LUT4 unary_minus_16_add_3_21_lut (.I0(GND_net), .I1(GND_net), .I2(n1[19]), 
            .I3(n28127), .O(n257[19])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i31349_3_lut (.I0(n4_adj_4331), .I1(IntegralLimit[13]), .I2(\PID_CONTROLLER.integral [13]), 
            .I3(GND_net), .O(n38031));   // verilog/motorControl.v(39[10:34])
    defparam i31349_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i31350_3_lut (.I0(n38031), .I1(IntegralLimit[14]), .I2(\PID_CONTROLLER.integral [14]), 
            .I3(GND_net), .O(n38032));   // verilog/motorControl.v(39[10:34])
    defparam i31350_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 add_4140_7_lut (.I0(GND_net), .I1(n8750[4]), .I2(n466_adj_4137), 
            .I3(n29492), .O(n8734[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4140_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4132_6_lut (.I0(GND_net), .I1(n8594[3]), .I2(n369_adj_4136), 
            .I3(n29329), .O(n8570[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4132_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4112_5_lut (.I0(GND_net), .I1(n8342[2]), .I2(n302_adj_4135), 
            .I3(n29148), .O(n8320[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4112_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4132_6 (.CI(n29329), .I0(n8594[3]), .I1(n369_adj_4136), 
            .CO(n29330));
    SB_CARRY add_4112_5 (.CI(n29148), .I0(n8342[2]), .I1(n302_adj_4135), 
            .CO(n29149));
    SB_LUT4 add_4112_4_lut (.I0(GND_net), .I1(n8342[1]), .I2(n229_adj_4134), 
            .I3(n29147), .O(n8320[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4112_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_21 (.CI(n28127), .I0(GND_net), .I1(n1[19]), 
            .CO(n28128));
    SB_CARRY add_4140_7 (.CI(n29492), .I0(n8750[4]), .I1(n466_adj_4137), 
            .CO(n29493));
    SB_LUT4 add_4132_5_lut (.I0(GND_net), .I1(n8594[2]), .I2(n296_adj_4133), 
            .I3(n29328), .O(n8570[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4132_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4112_4 (.CI(n29147), .I0(n8342[1]), .I1(n229_adj_4134), 
            .CO(n29148));
    SB_LUT4 add_4140_6_lut (.I0(GND_net), .I1(n8750[3]), .I2(n393_adj_4132), 
            .I3(n29491), .O(n8734[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4140_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4140_6 (.CI(n29491), .I0(n8750[3]), .I1(n393_adj_4132), 
            .CO(n29492));
    SB_CARRY add_4132_5 (.CI(n29328), .I0(n8594[2]), .I1(n296_adj_4133), 
            .CO(n29329));
    SB_LUT4 add_4112_3_lut (.I0(GND_net), .I1(n8342[0]), .I2(n156_adj_4131), 
            .I3(n29146), .O(n8320[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4112_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4112_3 (.CI(n29146), .I0(n8342[0]), .I1(n156_adj_4131), 
            .CO(n29147));
    SB_LUT4 unary_minus_16_add_3_20_lut (.I0(GND_net), .I1(GND_net), .I2(n1[18]), 
            .I3(n28126), .O(n257[18])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4140_5_lut (.I0(GND_net), .I1(n8750[2]), .I2(n320_adj_4129), 
            .I3(n29490), .O(n8734[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4140_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4132_4_lut (.I0(GND_net), .I1(n8594[1]), .I2(n223_adj_4128), 
            .I3(n29327), .O(n8570[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4132_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4112_2_lut (.I0(GND_net), .I1(n14_adj_4127), .I2(n83_adj_4126), 
            .I3(GND_net), .O(n8320[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4112_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4112_2 (.CI(GND_net), .I0(n14_adj_4127), .I1(n83_adj_4126), 
            .CO(n29146));
    SB_LUT4 add_4111_22_lut (.I0(GND_net), .I1(n8320[19]), .I2(GND_net), 
            .I3(n29145), .O(n8297[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4111_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4132_4 (.CI(n29327), .I0(n8594[1]), .I1(n223_adj_4128), 
            .CO(n29328));
    SB_LUT4 add_4111_21_lut (.I0(GND_net), .I1(n8320[18]), .I2(GND_net), 
            .I3(n29144), .O(n8297[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4111_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4111_21 (.CI(n29144), .I0(n8320[18]), .I1(GND_net), .CO(n29145));
    SB_LUT4 i30974_4_lut (.I0(\PID_CONTROLLER.integral [16]), .I1(n39087), 
            .I2(IntegralLimit[16]), .I3(n37891), .O(n37656));
    defparam i30974_4_lut.LUT_INIT = 16'h5a7b;
    SB_LUT4 add_4132_3_lut (.I0(GND_net), .I1(n8594[0]), .I2(n150_adj_4125), 
            .I3(n29326), .O(n8570[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4132_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_20 (.CI(n28126), .I0(GND_net), .I1(n1[18]), 
            .CO(n28127));
    SB_LUT4 add_4111_20_lut (.I0(GND_net), .I1(n8320[17]), .I2(GND_net), 
            .I3(n29143), .O(n8297[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4111_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_16_add_3_19_lut (.I0(GND_net), .I1(GND_net), .I2(n1[17]), 
            .I3(n28125), .O(n257[17])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4111_20 (.CI(n29143), .I0(n8320[17]), .I1(GND_net), .CO(n29144));
    SB_CARRY unary_minus_16_add_3_19 (.CI(n28125), .I0(GND_net), .I1(n1[17]), 
            .CO(n28126));
    SB_LUT4 unary_minus_16_add_3_18_lut (.I0(GND_net), .I1(GND_net), .I2(n1[16]), 
            .I3(n28124), .O(n257[16])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i31407_4_lut (.I0(n30_adj_4322), .I1(n10_adj_4321), .I2(n39110), 
            .I3(n37653), .O(n38089));   // verilog/motorControl.v(39[10:34])
    defparam i31407_4_lut.LUT_INIT = 16'haaac;
    SB_CARRY add_4140_5 (.CI(n29490), .I0(n8750[2]), .I1(n320_adj_4129), 
            .CO(n29491));
    SB_CARRY add_4132_3 (.CI(n29326), .I0(n8594[0]), .I1(n150_adj_4125), 
            .CO(n29327));
    SB_LUT4 add_4111_19_lut (.I0(GND_net), .I1(n8320[16]), .I2(GND_net), 
            .I3(n29142), .O(n8297[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4111_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4111_19 (.CI(n29142), .I0(n8320[16]), .I1(GND_net), .CO(n29143));
    SB_LUT4 add_4140_4_lut (.I0(GND_net), .I1(n8750[1]), .I2(n247_adj_4122), 
            .I3(n29489), .O(n8734[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4140_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4111_18_lut (.I0(GND_net), .I1(n8320[15]), .I2(GND_net), 
            .I3(n29141), .O(n8297[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4111_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4132_2_lut (.I0(GND_net), .I1(n8_adj_4121), .I2(n77_adj_4120), 
            .I3(GND_net), .O(n8570[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4132_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4111_18 (.CI(n29141), .I0(n8320[15]), .I1(GND_net), .CO(n29142));
    SB_CARRY unary_minus_16_add_3_18 (.CI(n28124), .I0(GND_net), .I1(n1[16]), 
            .CO(n28125));
    SB_CARRY add_4132_2 (.CI(GND_net), .I0(n8_adj_4121), .I1(n77_adj_4120), 
            .CO(n29326));
    SB_LUT4 add_4111_17_lut (.I0(GND_net), .I1(n8320[14]), .I2(GND_net), 
            .I3(n29140), .O(n8297[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4111_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4126_7_lut (.I0(GND_net), .I1(n34771), .I2(n490_adj_4112), 
            .I3(n29325), .O(n8537[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4126_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4111_17 (.CI(n29140), .I0(n8320[14]), .I1(GND_net), .CO(n29141));
    SB_LUT4 i31044_3_lut (.I0(n38032), .I1(IntegralLimit[15]), .I2(\PID_CONTROLLER.integral [15]), 
            .I3(GND_net), .O(n37726));   // verilog/motorControl.v(39[10:34])
    defparam i31044_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i31447_4_lut (.I0(n37726), .I1(n38089), .I2(n39110), .I3(n37656), 
            .O(n38129));   // verilog/motorControl.v(39[10:34])
    defparam i31447_4_lut.LUT_INIT = 16'hccca;
    SB_CARRY add_4140_4 (.CI(n29489), .I0(n8750[1]), .I1(n247_adj_4122), 
            .CO(n29490));
    SB_LUT4 add_4126_6_lut (.I0(GND_net), .I1(n8545[3]), .I2(n417_adj_4081), 
            .I3(n29324), .O(n8537[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4126_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i31383_4_lut (.I0(n25_adj_4049), .I1(n23_adj_3926), .I2(n21_adj_3923), 
            .I3(n37784), .O(n38065));
    defparam i31383_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 add_4111_16_lut (.I0(GND_net), .I1(n8320[13]), .I2(n1102_adj_4080), 
            .I3(n29139), .O(n8297[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4111_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_16_add_3_17_lut (.I0(GND_net), .I1(GND_net), .I2(n1[15]), 
            .I3(n28123), .O(n257[15])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 duty_23__I_0_i4_4_lut_4_lut (.I0(duty[0]), .I1(duty[1]), .I2(PWMLimit[1]), 
            .I3(PWMLimit[0]), .O(n4));   // verilog/motorControl.v(44[10:25])
    defparam duty_23__I_0_i4_4_lut_4_lut.LUT_INIT = 16'h0c8e;
    SB_LUT4 add_4140_3_lut (.I0(GND_net), .I1(n8750[0]), .I2(n174_adj_4074), 
            .I3(n29488), .O(n8734[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4140_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i31448_3_lut (.I0(n38129), .I1(IntegralLimit[18]), .I2(\PID_CONTROLLER.integral [18]), 
            .I3(GND_net), .O(n38130));   // verilog/motorControl.v(39[10:34])
    defparam i31448_3_lut.LUT_INIT = 16'h8e8e;
    SB_CARRY add_4111_16 (.CI(n29139), .I0(n8320[13]), .I1(n1102_adj_4080), 
            .CO(n29140));
    SB_CARRY unary_minus_16_add_3_17 (.CI(n28123), .I0(GND_net), .I1(n1[15]), 
            .CO(n28124));
    SB_LUT4 i31442_3_lut (.I0(n38130), .I1(IntegralLimit[19]), .I2(\PID_CONTROLLER.integral [19]), 
            .I3(GND_net), .O(n38124));   // verilog/motorControl.v(39[10:34])
    defparam i31442_3_lut.LUT_INIT = 16'h8e8e;
    SB_CARRY add_4126_6 (.CI(n29324), .I0(n8545[3]), .I1(n417_adj_4081), 
            .CO(n29325));
    SB_LUT4 add_4111_15_lut (.I0(GND_net), .I1(n8320[12]), .I2(n1029_adj_4072), 
            .I3(n29138), .O(n8297[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4111_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 duty_23__I_0_i8_3_lut_3_lut (.I0(duty[4]), .I1(duty[8]), .I2(PWMLimit[8]), 
            .I3(GND_net), .O(n8));   // verilog/motorControl.v(44[10:25])
    defparam duty_23__I_0_i8_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i30953_4_lut (.I0(\PID_CONTROLLER.integral [21]), .I1(n39078), 
            .I2(IntegralLimit[21]), .I3(n38127), .O(n37635));
    defparam i30953_4_lut.LUT_INIT = 16'h5a7b;
    SB_LUT4 add_4126_5_lut (.I0(GND_net), .I1(n8545[2]), .I2(n344_adj_4070), 
            .I3(n29323), .O(n8537[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4126_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_16_add_3_16_lut (.I0(GND_net), .I1(GND_net), .I2(n1[14]), 
            .I3(n28122), .O(n257[14])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4111_15 (.CI(n29138), .I0(n8320[12]), .I1(n1029_adj_4072), 
            .CO(n29139));
    SB_CARRY add_4140_3 (.CI(n29488), .I0(n8750[0]), .I1(n174_adj_4074), 
            .CO(n29489));
    SB_CARRY add_4126_5 (.CI(n29323), .I0(n8545[2]), .I1(n344_adj_4070), 
            .CO(n29324));
    SB_LUT4 add_4111_14_lut (.I0(GND_net), .I1(n8320[11]), .I2(n956_adj_4065), 
            .I3(n29137), .O(n8297[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4111_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4126_4_lut (.I0(GND_net), .I1(n8545[1]), .I2(n271_adj_4061), 
            .I3(n29322), .O(n8537[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4126_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4111_14 (.CI(n29137), .I0(n8320[11]), .I1(n956_adj_4065), 
            .CO(n29138));
    SB_LUT4 i30876_3_lut_4_lut (.I0(PWMLimit[3]), .I1(duty[3]), .I2(duty[2]), 
            .I3(PWMLimit[2]), .O(n37558));   // verilog/motorControl.v(44[10:25])
    defparam i30876_3_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 add_4140_2_lut (.I0(GND_net), .I1(n32), .I2(n101), .I3(GND_net), 
            .O(n8734[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4140_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4126_4 (.CI(n29322), .I0(n8545[1]), .I1(n271_adj_4061), 
            .CO(n29323));
    SB_LUT4 add_4111_13_lut (.I0(GND_net), .I1(n8320[10]), .I2(n883), 
            .I3(n29136), .O(n8297[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4111_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4126_3_lut (.I0(GND_net), .I1(n8545[0]), .I2(n198), .I3(n29321), 
            .O(n8537[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4126_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4111_13 (.CI(n29136), .I0(n8320[10]), .I1(n883), .CO(n29137));
    SB_CARRY unary_minus_16_add_3_16 (.CI(n28122), .I0(GND_net), .I1(n1[14]), 
            .CO(n28123));
    SB_LUT4 unary_minus_16_add_3_15_lut (.I0(GND_net), .I1(GND_net), .I2(n1[13]), 
            .I3(n28121), .O(n257[13])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4111_12_lut (.I0(GND_net), .I1(n8320[9]), .I2(n810), .I3(n29135), 
            .O(n8297[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4111_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_15 (.CI(n28121), .I0(GND_net), .I1(n1[13]), 
            .CO(n28122));
    SB_LUT4 IntegralLimit_23__I_0_i45_rep_295_2_lut (.I0(\PID_CONTROLLER.integral [22]), 
            .I1(IntegralLimit[22]), .I2(GND_net), .I3(GND_net), .O(n39076));   // verilog/motorControl.v(39[10:34])
    defparam IntegralLimit_23__I_0_i45_rep_295_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 unary_minus_16_add_3_14_lut (.I0(GND_net), .I1(GND_net), .I2(n1[12]), 
            .I3(n28120), .O(n257[12])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4111_12 (.CI(n29135), .I0(n8320[9]), .I1(n810), .CO(n29136));
    SB_CARRY add_4140_2 (.CI(GND_net), .I0(n32), .I1(n101), .CO(n29488));
    SB_CARRY add_4126_3 (.CI(n29321), .I0(n8545[0]), .I1(n198), .CO(n29322));
    SB_LUT4 add_4111_11_lut (.I0(GND_net), .I1(n8320[8]), .I2(n737), .I3(n29134), 
            .O(n8297[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4111_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_14 (.CI(n28120), .I0(GND_net), .I1(n1[12]), 
            .CO(n28121));
    SB_LUT4 i31369_4_lut (.I0(n38006), .I1(n37925), .I2(n39076), .I3(n37632), 
            .O(n38051));   // verilog/motorControl.v(39[10:34])
    defparam i31369_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 add_4126_2_lut (.I0(GND_net), .I1(n56), .I2(n125), .I3(GND_net), 
            .O(n8537[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4126_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4111_11 (.CI(n29134), .I0(n8320[8]), .I1(n737), .CO(n29135));
    SB_LUT4 state_23__I_0_add_2_25_lut (.I0(GND_net), .I1(motor_state[23]), 
            .I2(n1_adj_4333[23]), .I3(n28313), .O(\PID_CONTROLLER.err_23__N_3514 [23])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 state_23__I_0_add_2_24_lut (.I0(GND_net), .I1(motor_state[22]), 
            .I2(n1_adj_4333[22]), .I3(n28312), .O(\PID_CONTROLLER.err_23__N_3514 [22])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i31050_3_lut (.I0(n38124), .I1(IntegralLimit[20]), .I2(\PID_CONTROLLER.integral [20]), 
            .I3(GND_net), .O(n37732));   // verilog/motorControl.v(39[10:34])
    defparam i31050_3_lut.LUT_INIT = 16'h8e8e;
    SB_CARRY state_23__I_0_add_2_24 (.CI(n28312), .I0(motor_state[22]), 
            .I1(n1_adj_4333[22]), .CO(n28313));
    SB_LUT4 state_23__I_0_add_2_23_lut (.I0(GND_net), .I1(motor_state[21]), 
            .I2(n1_adj_4333[21]), .I3(n28311), .O(\PID_CONTROLLER.err_23__N_3514 [21])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY state_23__I_0_add_2_23 (.CI(n28311), .I0(motor_state[21]), 
            .I1(n1_adj_4333[21]), .CO(n28312));
    SB_LUT4 duty_23__I_0_i6_3_lut_3_lut (.I0(PWMLimit[3]), .I1(duty[3]), 
            .I2(duty[2]), .I3(GND_net), .O(n6));   // verilog/motorControl.v(44[10:25])
    defparam duty_23__I_0_i6_3_lut_3_lut.LUT_INIT = 16'hd4d4;
    SB_LUT4 i31418_3_lut (.I0(n38099), .I1(\PID_CONTROLLER.integral_23__N_3589 [23]), 
            .I2(\PID_CONTROLLER.integral [23]), .I3(GND_net), .O(\PID_CONTROLLER.integral_23__N_3588 ));   // verilog/motorControl.v(39[38:63])
    defparam i31418_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 state_23__I_0_add_2_22_lut (.I0(GND_net), .I1(motor_state[20]), 
            .I2(n1_adj_4333[20]), .I3(n28310), .O(\PID_CONTROLLER.err_23__N_3514 [20])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i31415_4_lut (.I0(n37732), .I1(n38051), .I2(n39076), .I3(n37635), 
            .O(n38097));   // verilog/motorControl.v(39[10:34])
    defparam i31415_4_lut.LUT_INIT = 16'hccca;
    SB_CARRY state_23__I_0_add_2_22 (.CI(n28310), .I0(motor_state[20]), 
            .I1(n1_adj_4333[20]), .CO(n28311));
    SB_LUT4 state_23__I_0_add_2_21_lut (.I0(GND_net), .I1(motor_state[19]), 
            .I2(n1_adj_4333[19]), .I3(n28309), .O(\PID_CONTROLLER.err_23__N_3514 [19])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4126_2 (.CI(GND_net), .I0(n56), .I1(n125), .CO(n29321));
    SB_LUT4 add_4111_10_lut (.I0(GND_net), .I1(n8320[7]), .I2(n664), .I3(n29133), 
            .O(n8297[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4111_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4125_8_lut (.I0(GND_net), .I1(n8537[5]), .I2(n560), .I3(n29320), 
            .O(n8528[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4125_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4125_7_lut (.I0(GND_net), .I1(n8537[4]), .I2(n487), .I3(n29319), 
            .O(n8528[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4125_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4139_16_lut (.I0(GND_net), .I1(n8734[13]), .I2(n1120), 
            .I3(n29487), .O(n8717[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4139_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4125_7 (.CI(n29319), .I0(n8537[4]), .I1(n487), .CO(n29320));
    SB_CARRY state_23__I_0_add_2_21 (.CI(n28309), .I0(motor_state[19]), 
            .I1(n1_adj_4333[19]), .CO(n28310));
    SB_LUT4 unary_minus_16_add_3_13_lut (.I0(GND_net), .I1(GND_net), .I2(n1[11]), 
            .I3(n28119), .O(n257[11])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4111_10 (.CI(n29133), .I0(n8320[7]), .I1(n664), .CO(n29134));
    SB_LUT4 state_23__I_0_add_2_20_lut (.I0(GND_net), .I1(motor_state[18]), 
            .I2(n1_adj_4333[18]), .I3(n28308), .O(\PID_CONTROLLER.err_23__N_3514 [18])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4139_15_lut (.I0(GND_net), .I1(n8734[12]), .I2(n1047), 
            .I3(n29486), .O(n8717[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4139_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY state_23__I_0_add_2_20 (.CI(n28308), .I0(motor_state[18]), 
            .I1(n1_adj_4333[18]), .CO(n28309));
    SB_CARRY add_4139_15 (.CI(n29486), .I0(n8734[12]), .I1(n1047), .CO(n29487));
    SB_LUT4 add_4139_14_lut (.I0(GND_net), .I1(n8734[11]), .I2(n974), 
            .I3(n29485), .O(n8717[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4139_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4125_6_lut (.I0(GND_net), .I1(n8537[3]), .I2(n414), .I3(n29318), 
            .O(n8528[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4125_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4111_9_lut (.I0(GND_net), .I1(n8320[6]), .I2(n591), .I3(n29132), 
            .O(n8297[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4111_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4111_9 (.CI(n29132), .I0(n8320[6]), .I1(n591), .CO(n29133));
    SB_CARRY add_4125_6 (.CI(n29318), .I0(n8537[3]), .I1(n414), .CO(n29319));
    SB_LUT4 add_4111_8_lut (.I0(GND_net), .I1(n8320[5]), .I2(n518), .I3(n29131), 
            .O(n8297[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4111_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 state_23__I_0_add_2_19_lut (.I0(GND_net), .I1(motor_state[17]), 
            .I2(n1_adj_4333[17]), .I3(n28307), .O(\PID_CONTROLLER.err_23__N_3514 [17])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY state_23__I_0_add_2_19 (.CI(n28307), .I0(motor_state[17]), 
            .I1(n1_adj_4333[17]), .CO(n28308));
    SB_CARRY add_4111_8 (.CI(n29131), .I0(n8320[5]), .I1(n518), .CO(n29132));
    SB_LUT4 state_23__I_0_add_2_18_lut (.I0(GND_net), .I1(motor_state[16]), 
            .I2(n1_adj_4333[16]), .I3(n28306), .O(\PID_CONTROLLER.err_23__N_3514 [16])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4125_5_lut (.I0(GND_net), .I1(n8537[2]), .I2(n341), .I3(n29317), 
            .O(n8528[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4125_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY state_23__I_0_add_2_18 (.CI(n28306), .I0(motor_state[16]), 
            .I1(n1_adj_4333[16]), .CO(n28307));
    SB_LUT4 \PID_CONTROLLER.integral_23__I_839_4_lut  (.I0(n38097), .I1(\PID_CONTROLLER.integral_23__N_3588 ), 
            .I2(\PID_CONTROLLER.integral [23]), .I3(IntegralLimit[23]), 
            .O(\PID_CONTROLLER.integral_23__N_3586 ));   // verilog/motorControl.v(39[10:63])
    defparam \PID_CONTROLLER.integral_23__I_839_4_lut .LUT_INIT = 16'h80c8;
    SB_LUT4 add_4111_7_lut (.I0(GND_net), .I1(n8320[4]), .I2(n445), .I3(n29130), 
            .O(n8297[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4111_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 state_23__I_0_add_2_17_lut (.I0(GND_net), .I1(motor_state[15]), 
            .I2(n1_adj_4333[15]), .I3(n28305), .O(\PID_CONTROLLER.err_23__N_3514 [15])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4139_14 (.CI(n29485), .I0(n8734[11]), .I1(n974), .CO(n29486));
    SB_CARRY add_4125_5 (.CI(n29317), .I0(n8537[2]), .I1(n341), .CO(n29318));
    SB_CARRY state_23__I_0_add_2_17 (.CI(n28305), .I0(motor_state[15]), 
            .I1(n1_adj_4333[15]), .CO(n28306));
    SB_LUT4 state_23__I_0_add_2_16_lut (.I0(GND_net), .I1(motor_state[14]), 
            .I2(n1_adj_4333[14]), .I3(n28304), .O(\PID_CONTROLLER.err_23__N_3514 [14])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4111_7 (.CI(n29130), .I0(n8320[4]), .I1(n445), .CO(n29131));
    SB_LUT4 add_4125_4_lut (.I0(GND_net), .I1(n8537[1]), .I2(n268), .I3(n29316), 
            .O(n8528[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4125_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4111_6_lut (.I0(GND_net), .I1(n8320[3]), .I2(n372), .I3(n29129), 
            .O(n8297[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4111_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_13 (.CI(n28119), .I0(GND_net), .I1(n1[11]), 
            .CO(n28120));
    SB_LUT4 unary_minus_16_add_3_12_lut (.I0(GND_net), .I1(GND_net), .I2(n1[10]), 
            .I3(n28118), .O(n257[10])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY state_23__I_0_add_2_16 (.CI(n28304), .I0(motor_state[14]), 
            .I1(n1_adj_4333[14]), .CO(n28305));
    SB_LUT4 state_23__I_0_add_2_15_lut (.I0(GND_net), .I1(motor_state[13]), 
            .I2(n1_adj_4333[13]), .I3(n28303), .O(\PID_CONTROLLER.err_23__N_3514 [13])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY state_23__I_0_add_2_15 (.CI(n28303), .I0(motor_state[13]), 
            .I1(n1_adj_4333[13]), .CO(n28304));
    SB_CARRY add_4111_6 (.CI(n29129), .I0(n8320[3]), .I1(n372), .CO(n29130));
    SB_LUT4 add_4139_13_lut (.I0(GND_net), .I1(n8734[10]), .I2(n901), 
            .I3(n29484), .O(n8717[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4139_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4125_4 (.CI(n29316), .I0(n8537[1]), .I1(n268), .CO(n29317));
    SB_LUT4 add_4125_3_lut (.I0(GND_net), .I1(n8537[0]), .I2(n195_adj_3992), 
            .I3(n29315), .O(n8528[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4125_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4111_5_lut (.I0(GND_net), .I1(n8320[2]), .I2(n299), .I3(n29128), 
            .O(n8297[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4111_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4111_5 (.CI(n29128), .I0(n8320[2]), .I1(n299), .CO(n29129));
    SB_CARRY add_4125_3 (.CI(n29315), .I0(n8537[0]), .I1(n195_adj_3992), 
            .CO(n29316));
    SB_CARRY add_4139_13 (.CI(n29484), .I0(n8734[10]), .I1(n901), .CO(n29485));
    SB_LUT4 add_4139_12_lut (.I0(GND_net), .I1(n8734[9]), .I2(n828), .I3(n29483), 
            .O(n8717[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4139_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4125_2_lut (.I0(GND_net), .I1(n53), .I2(n122), .I3(GND_net), 
            .O(n8528[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4125_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 state_23__I_0_add_2_14_lut (.I0(GND_net), .I1(motor_state[12]), 
            .I2(n1_adj_4333[12]), .I3(n28302), .O(\PID_CONTROLLER.err_23__N_3514 [12])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4111_4_lut (.I0(GND_net), .I1(n8320[1]), .I2(n226), .I3(n29127), 
            .O(n8297[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4111_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4125_2 (.CI(GND_net), .I0(n53), .I1(n122), .CO(n29315));
    SB_LUT4 add_4124_9_lut (.I0(GND_net), .I1(n8528[6]), .I2(n630), .I3(n29314), 
            .O(n8518[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4124_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4139_12 (.CI(n29483), .I0(n8734[9]), .I1(n828), .CO(n29484));
    SB_LUT4 add_4124_8_lut (.I0(GND_net), .I1(n8528[5]), .I2(n557), .I3(n29313), 
            .O(n8518[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4124_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4139_11_lut (.I0(GND_net), .I1(n8734[8]), .I2(n755), .I3(n29482), 
            .O(n8717[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4139_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4111_4 (.CI(n29127), .I0(n8320[1]), .I1(n226), .CO(n29128));
    SB_LUT4 add_4111_3_lut (.I0(GND_net), .I1(n8320[0]), .I2(n153), .I3(n29126), 
            .O(n8297[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4111_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4124_8 (.CI(n29313), .I0(n8528[5]), .I1(n557), .CO(n29314));
    SB_CARRY add_4139_11 (.CI(n29482), .I0(n8734[8]), .I1(n755), .CO(n29483));
    SB_CARRY add_4111_3 (.CI(n29126), .I0(n8320[0]), .I1(n153), .CO(n29127));
    SB_LUT4 add_4124_7_lut (.I0(GND_net), .I1(n8528[4]), .I2(n484), .I3(n29312), 
            .O(n8518[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4124_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4111_2_lut (.I0(GND_net), .I1(n11_adj_3990), .I2(n80), 
            .I3(GND_net), .O(n8297[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4111_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_12 (.CI(n28118), .I0(GND_net), .I1(n1[10]), 
            .CO(n28119));
    SB_LUT4 add_4139_10_lut (.I0(GND_net), .I1(n8734[7]), .I2(n682), .I3(n29481), 
            .O(n8717[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4139_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY state_23__I_0_add_2_14 (.CI(n28302), .I0(motor_state[12]), 
            .I1(n1_adj_4333[12]), .CO(n28303));
    SB_CARRY add_4124_7 (.CI(n29312), .I0(n8528[4]), .I1(n484), .CO(n29313));
    SB_CARRY add_4111_2 (.CI(GND_net), .I0(n11_adj_3990), .I1(n80), .CO(n29126));
    SB_LUT4 state_23__I_0_add_2_13_lut (.I0(GND_net), .I1(motor_state[11]), 
            .I2(n1_adj_4333[11]), .I3(n28301), .O(\PID_CONTROLLER.err_23__N_3514 [11])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i30799_2_lut_4_lut (.I0(PWMLimit[21]), .I1(duty[21]), .I2(PWMLimit[9]), 
            .I3(duty[9]), .O(n37480));
    defparam i30799_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_CARRY add_4139_10 (.CI(n29481), .I0(n8734[7]), .I1(n682), .CO(n29482));
    SB_LUT4 add_4139_9_lut (.I0(GND_net), .I1(n8734[6]), .I2(n609), .I3(n29480), 
            .O(n8717[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4139_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_16_add_3_11_lut (.I0(GND_net), .I1(GND_net), .I2(n1[9]), 
            .I3(n28117), .O(n257[9])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4124_6_lut (.I0(GND_net), .I1(n8528[3]), .I2(n411), .I3(n29311), 
            .O(n8518[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4124_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_add_1225_24_lut (.I0(\PID_CONTROLLER.err [23]), .I1(n8273[21]), 
            .I2(GND_net), .I3(n29125), .O(n7788[0])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_24_lut.LUT_INIT = 16'h6996;
    SB_LUT4 mult_10_add_1225_23_lut (.I0(n24379), .I1(n8273[20]), .I2(GND_net), 
            .I3(n29124), .O(n3265[22])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_23_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_4139_9 (.CI(n29480), .I0(n8734[6]), .I1(n609), .CO(n29481));
    SB_LUT4 add_4139_8_lut (.I0(GND_net), .I1(n8734[5]), .I2(n536), .I3(n29479), 
            .O(n8717[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4139_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY state_23__I_0_add_2_13 (.CI(n28301), .I0(motor_state[11]), 
            .I1(n1_adj_4333[11]), .CO(n28302));
    SB_CARRY add_4124_6 (.CI(n29311), .I0(n8528[3]), .I1(n411), .CO(n29312));
    SB_LUT4 state_23__I_0_add_2_12_lut (.I0(GND_net), .I1(motor_state[10]), 
            .I2(n1_adj_4333[10]), .I3(n28300), .O(\PID_CONTROLLER.err_23__N_3514 [10])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4124_5_lut (.I0(GND_net), .I1(n8528[2]), .I2(n338), .I3(n29310), 
            .O(n8518[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4124_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4124_5 (.CI(n29310), .I0(n8528[2]), .I1(n338), .CO(n29311));
    SB_CARRY add_4139_8 (.CI(n29479), .I0(n8734[5]), .I1(n536), .CO(n29480));
    SB_LUT4 add_4124_4_lut (.I0(GND_net), .I1(n8528[1]), .I2(n265), .I3(n29309), 
            .O(n8518[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4124_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_1225_23 (.CI(n29124), .I0(n8273[20]), .I1(GND_net), 
            .CO(n29125));
    SB_CARRY unary_minus_16_add_3_11 (.CI(n28117), .I0(GND_net), .I1(n1[9]), 
            .CO(n28118));
    SB_CARRY state_23__I_0_add_2_12 (.CI(n28300), .I0(motor_state[10]), 
            .I1(n1_adj_4333[10]), .CO(n28301));
    SB_LUT4 state_23__I_0_add_2_11_lut (.I0(GND_net), .I1(motor_state[9]), 
            .I2(n1_adj_4333[9]), .I3(n28299), .O(\PID_CONTROLLER.err_23__N_3514 [9])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY state_23__I_0_add_2_11 (.CI(n28299), .I0(motor_state[9]), .I1(n1_adj_4333[9]), 
            .CO(n28300));
    SB_LUT4 mult_10_add_1225_22_lut (.I0(n24379), .I1(n8273[19]), .I2(GND_net), 
            .I3(n29123), .O(n3265[21])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_22_lut.LUT_INIT = 16'h8228;
    SB_LUT4 unary_minus_16_add_3_10_lut (.I0(GND_net), .I1(GND_net), .I2(n1[8]), 
            .I3(n28116), .O(n257[8])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4124_4 (.CI(n29309), .I0(n8528[1]), .I1(n265), .CO(n29310));
    SB_CARRY mult_10_add_1225_22 (.CI(n29123), .I0(n8273[19]), .I1(GND_net), 
            .CO(n29124));
    SB_LUT4 add_4124_3_lut (.I0(GND_net), .I1(n8528[0]), .I2(n192_adj_3979), 
            .I3(n29308), .O(n8518[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4124_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_add_1225_21_lut (.I0(n24379), .I1(n8273[18]), .I2(GND_net), 
            .I3(n29122), .O(n3265[20])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_21_lut.LUT_INIT = 16'h8228;
    SB_LUT4 add_4139_7_lut (.I0(GND_net), .I1(n8734[4]), .I2(n463), .I3(n29478), 
            .O(n8717[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4139_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_1225_21 (.CI(n29122), .I0(n8273[18]), .I1(GND_net), 
            .CO(n29123));
    SB_LUT4 mult_10_add_1225_20_lut (.I0(n24379), .I1(n8273[17]), .I2(GND_net), 
            .I3(n29121), .O(n3265[19])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_20_lut.LUT_INIT = 16'h8228;
    SB_CARRY unary_minus_16_add_3_10 (.CI(n28116), .I0(GND_net), .I1(n1[8]), 
            .CO(n28117));
    SB_CARRY mult_10_add_1225_20 (.CI(n29121), .I0(n8273[17]), .I1(GND_net), 
            .CO(n29122));
    SB_CARRY add_4124_3 (.CI(n29308), .I0(n8528[0]), .I1(n192_adj_3979), 
            .CO(n29309));
    SB_LUT4 state_23__I_0_add_2_10_lut (.I0(GND_net), .I1(motor_state[8]), 
            .I2(n1_adj_4333[8]), .I3(n28298), .O(\PID_CONTROLLER.err_23__N_3514 [8])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_add_1225_19_lut (.I0(n24379), .I1(n8273[16]), .I2(GND_net), 
            .I3(n29120), .O(n3265[18])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_19_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_4139_7 (.CI(n29478), .I0(n8734[4]), .I1(n463), .CO(n29479));
    SB_LUT4 add_4124_2_lut (.I0(GND_net), .I1(n50_adj_3972), .I2(n119_adj_3970), 
            .I3(GND_net), .O(n8518[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4124_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_1225_19 (.CI(n29120), .I0(n8273[16]), .I1(GND_net), 
            .CO(n29121));
    SB_CARRY state_23__I_0_add_2_10 (.CI(n28298), .I0(motor_state[8]), .I1(n1_adj_4333[8]), 
            .CO(n28299));
    SB_CARRY add_4124_2 (.CI(GND_net), .I0(n50_adj_3972), .I1(n119_adj_3970), 
            .CO(n29308));
    SB_LUT4 unary_minus_16_add_3_9_lut (.I0(GND_net), .I1(GND_net), .I2(n1[7]), 
            .I3(n28115), .O(n257[7])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_add_1225_18_lut (.I0(n24379), .I1(n8273[15]), .I2(GND_net), 
            .I3(n29119), .O(n3265[17])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_18_lut.LUT_INIT = 16'h8228;
    SB_CARRY mult_10_add_1225_18 (.CI(n29119), .I0(n8273[15]), .I1(GND_net), 
            .CO(n29120));
    SB_LUT4 add_4123_10_lut (.I0(GND_net), .I1(n8518[7]), .I2(n700_adj_3965), 
            .I3(n29307), .O(n8507[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4123_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4139_6_lut (.I0(GND_net), .I1(n8734[3]), .I2(n390_adj_3964), 
            .I3(n29477), .O(n8717[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4139_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 state_23__I_0_add_2_9_lut (.I0(GND_net), .I1(motor_state[7]), 
            .I2(n1_adj_4333[7]), .I3(n28297), .O(\PID_CONTROLLER.err_23__N_3514 [7])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4139_6 (.CI(n29477), .I0(n8734[3]), .I1(n390_adj_3964), 
            .CO(n29478));
    SB_LUT4 add_4123_9_lut (.I0(GND_net), .I1(n8518[6]), .I2(n627_adj_3963), 
            .I3(n29306), .O(n8507[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4123_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_add_1225_17_lut (.I0(n24379), .I1(n8273[14]), .I2(GND_net), 
            .I3(n29118), .O(n3265[16])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_17_lut.LUT_INIT = 16'h8228;
    SB_CARRY state_23__I_0_add_2_9 (.CI(n28297), .I0(motor_state[7]), .I1(n1_adj_4333[7]), 
            .CO(n28298));
    SB_LUT4 i31253_4_lut (.I0(n31_adj_4073), .I1(n29_adj_4071), .I2(n27_adj_4058), 
            .I3(n38065), .O(n37935));
    defparam i31253_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 state_23__I_0_add_2_8_lut (.I0(GND_net), .I1(motor_state[6]), 
            .I2(n1_adj_4333[6]), .I3(n28296), .O(\PID_CONTROLLER.err_23__N_3514 [6])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY state_23__I_0_add_2_8 (.CI(n28296), .I0(motor_state[6]), .I1(n1_adj_4333[6]), 
            .CO(n28297));
    SB_CARRY unary_minus_16_add_3_9 (.CI(n28115), .I0(GND_net), .I1(n1[7]), 
            .CO(n28116));
    SB_LUT4 state_23__I_0_add_2_7_lut (.I0(GND_net), .I1(motor_state[5]), 
            .I2(n1_adj_4333[5]), .I3(n28295), .O(\PID_CONTROLLER.err_23__N_3514 [5])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY state_23__I_0_add_2_7 (.CI(n28295), .I0(motor_state[5]), .I1(n1_adj_4333[5]), 
            .CO(n28296));
    SB_LUT4 add_4139_5_lut (.I0(GND_net), .I1(n8734[2]), .I2(n317), .I3(n29476), 
            .O(n8717[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4139_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 state_23__I_0_add_2_6_lut (.I0(GND_net), .I1(motor_state[4]), 
            .I2(n1_adj_4333[4]), .I3(n28294), .O(\PID_CONTROLLER.err_23__N_3514 [4])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4123_9 (.CI(n29306), .I0(n8518[6]), .I1(n627_adj_3963), 
            .CO(n29307));
    SB_CARRY add_4139_5 (.CI(n29476), .I0(n8734[2]), .I1(n317), .CO(n29477));
    SB_CARRY mult_10_add_1225_17 (.CI(n29118), .I0(n8273[14]), .I1(GND_net), 
            .CO(n29119));
    SB_LUT4 add_4123_8_lut (.I0(GND_net), .I1(n8518[5]), .I2(n554_adj_3952), 
            .I3(n29305), .O(n8507[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4123_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_add_1225_16_lut (.I0(n24379), .I1(n8273[13]), .I2(n1096), 
            .I3(n29117), .O(n3265[15])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_16_lut.LUT_INIT = 16'h8228;
    SB_LUT4 mult_10_i75_2_lut (.I0(\Kp[1] ), .I1(\PID_CONTROLLER.err [12]), 
            .I2(GND_net), .I3(GND_net), .O(n110));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i75_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 duty_23__I_0_i16_3_lut_3_lut (.I0(duty[9]), .I1(duty[21]), .I2(PWMLimit[21]), 
            .I3(GND_net), .O(n16));   // verilog/motorControl.v(44[10:25])
    defparam duty_23__I_0_i16_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 unary_minus_16_add_3_8_lut (.I0(GND_net), .I1(GND_net), .I2(n1[6]), 
            .I3(n28114), .O(n257[6])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY state_23__I_0_add_2_6 (.CI(n28294), .I0(motor_state[4]), .I1(n1_adj_4333[4]), 
            .CO(n28295));
    SB_LUT4 add_4139_4_lut (.I0(GND_net), .I1(n8734[1]), .I2(n244), .I3(n29475), 
            .O(n8717[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4139_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4123_8 (.CI(n29305), .I0(n8518[5]), .I1(n554_adj_3952), 
            .CO(n29306));
    SB_CARRY mult_10_add_1225_16 (.CI(n29117), .I0(n8273[13]), .I1(n1096), 
            .CO(n29118));
    SB_LUT4 state_23__I_0_add_2_5_lut (.I0(GND_net), .I1(motor_state[3]), 
            .I2(n1_adj_4333[3]), .I3(n28293), .O(\PID_CONTROLLER.err_23__N_3514 [3])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4123_7_lut (.I0(GND_net), .I1(n8518[4]), .I2(n481_adj_3948), 
            .I3(n29304), .O(n8507[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4123_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY state_23__I_0_add_2_5 (.CI(n28293), .I0(motor_state[3]), .I1(n1_adj_4333[3]), 
            .CO(n28294));
    SB_LUT4 mult_10_add_1225_15_lut (.I0(n24379), .I1(n8273[12]), .I2(n1023), 
            .I3(n29116), .O(n3265[14])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_15_lut.LUT_INIT = 16'h8228;
    SB_LUT4 state_23__I_0_add_2_4_lut (.I0(GND_net), .I1(motor_state[2]), 
            .I2(n1_adj_4333[2]), .I3(n28292), .O(\PID_CONTROLLER.err_23__N_3514 [2])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4139_4 (.CI(n29475), .I0(n8734[1]), .I1(n244), .CO(n29476));
    SB_LUT4 mult_10_i28_2_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err [13]), 
            .I2(GND_net), .I3(GND_net), .O(n41_adj_3989));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i28_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY state_23__I_0_add_2_4 (.CI(n28292), .I0(motor_state[2]), .I1(n1_adj_4333[2]), 
            .CO(n28293));
    SB_LUT4 state_23__I_0_add_2_3_lut (.I0(GND_net), .I1(motor_state[1]), 
            .I2(n1_adj_4333[1]), .I3(n28291), .O(\PID_CONTROLLER.err_23__N_3514 [1])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 duty_23__I_0_i10_3_lut_3_lut (.I0(duty[5]), .I1(duty[6]), .I2(PWMLimit[6]), 
            .I3(GND_net), .O(n10));   // verilog/motorControl.v(44[10:25])
    defparam duty_23__I_0_i10_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i30813_2_lut_4_lut (.I0(PWMLimit[16]), .I1(duty[16]), .I2(PWMLimit[7]), 
            .I3(duty[7]), .O(n37494));
    defparam i30813_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_CARRY state_23__I_0_add_2_3 (.CI(n28291), .I0(motor_state[1]), .I1(n1_adj_4333[1]), 
            .CO(n28292));
    SB_LUT4 state_23__I_0_add_2_2_lut (.I0(GND_net), .I1(motor_state[0]), 
            .I2(n1_adj_4333[0]), .I3(VCC_net), .O(\PID_CONTROLLER.err_23__N_3514 [0])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY state_23__I_0_add_2_2 (.CI(VCC_net), .I0(motor_state[0]), .I1(n1_adj_4333[0]), 
            .CO(n28291));
    SB_CARRY add_4123_7 (.CI(n29304), .I0(n8518[4]), .I1(n481_adj_3948), 
            .CO(n29305));
    SB_LUT4 add_4139_3_lut (.I0(GND_net), .I1(n8734[0]), .I2(n171), .I3(n29474), 
            .O(n8717[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4139_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4123_6_lut (.I0(GND_net), .I1(n8518[3]), .I2(n408), .I3(n29303), 
            .O(n8507[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4123_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_1225_15 (.CI(n29116), .I0(n8273[12]), .I1(n1023), 
            .CO(n29117));
    SB_LUT4 mult_10_add_1225_14_lut (.I0(n24379), .I1(n8273[11]), .I2(n950), 
            .I3(n29115), .O(n3265[13])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_14_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_4123_6 (.CI(n29303), .I0(n8518[3]), .I1(n408), .CO(n29304));
    SB_CARRY mult_10_add_1225_14 (.CI(n29115), .I0(n8273[11]), .I1(n950), 
            .CO(n29116));
    SB_LUT4 add_4123_5_lut (.I0(GND_net), .I1(n8518[2]), .I2(n335_adj_3938), 
            .I3(n29302), .O(n8507[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4123_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 duty_23__I_0_i41_2_lut (.I0(PWMLimit[20]), .I1(duty[20]), .I2(GND_net), 
            .I3(GND_net), .O(n41));   // verilog/motorControl.v(44[10:25])
    defparam duty_23__I_0_i41_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_10_add_1225_13_lut (.I0(n24379), .I1(n8273[10]), .I2(n877), 
            .I3(n29114), .O(n3265[12])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_13_lut.LUT_INIT = 16'h8228;
    SB_LUT4 duty_23__I_0_i39_2_lut (.I0(PWMLimit[19]), .I1(duty[19]), .I2(GND_net), 
            .I3(GND_net), .O(n39));   // verilog/motorControl.v(44[10:25])
    defparam duty_23__I_0_i39_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY unary_minus_16_add_3_8 (.CI(n28114), .I0(GND_net), .I1(n1[6]), 
            .CO(n28115));
    SB_CARRY add_4139_3 (.CI(n29474), .I0(n8734[0]), .I1(n171), .CO(n29475));
    SB_CARRY mult_10_add_1225_13 (.CI(n29114), .I0(n8273[10]), .I1(n877), 
            .CO(n29115));
    SB_CARRY add_4123_5 (.CI(n29302), .I0(n8518[2]), .I1(n335_adj_3938), 
            .CO(n29303));
    SB_LUT4 mult_10_add_1225_12_lut (.I0(n24379), .I1(n8273[9]), .I2(n804), 
            .I3(n29113), .O(n3265[11])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_12_lut.LUT_INIT = 16'h8228;
    SB_CARRY mult_10_add_1225_12 (.CI(n29113), .I0(n8273[9]), .I1(n804), 
            .CO(n29114));
    SB_LUT4 add_4123_4_lut (.I0(GND_net), .I1(n8518[1]), .I2(n262), .I3(n29301), 
            .O(n8507[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4123_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_add_1225_11_lut (.I0(n24379), .I1(n8273[8]), .I2(n731), 
            .I3(n29112), .O(n3265[10])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_11_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_4123_4 (.CI(n29301), .I0(n8518[1]), .I1(n262), .CO(n29302));
    SB_LUT4 add_4123_3_lut (.I0(GND_net), .I1(n8518[0]), .I2(n189), .I3(n29300), 
            .O(n8507[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4123_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_1225_11 (.CI(n29112), .I0(n8273[8]), .I1(n731), 
            .CO(n29113));
    SB_LUT4 duty_23__I_0_i12_3_lut_3_lut (.I0(duty[7]), .I1(duty[16]), .I2(PWMLimit[16]), 
            .I3(GND_net), .O(n12));   // verilog/motorControl.v(44[10:25])
    defparam duty_23__I_0_i12_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 mult_10_add_1225_10_lut (.I0(n24379), .I1(n8273[7]), .I2(n658), 
            .I3(n29111), .O(n3265[9])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_10_lut.LUT_INIT = 16'h8228;
    SB_CARRY mult_10_add_1225_10 (.CI(n29111), .I0(n8273[7]), .I1(n658), 
            .CO(n29112));
    SB_LUT4 mult_10_i247_2_lut (.I0(\Kp[5] ), .I1(\PID_CONTROLLER.err [0]), 
            .I2(GND_net), .I3(GND_net), .O(n366));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i247_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_add_1225_9_lut (.I0(n24379), .I1(n8273[6]), .I2(n585), 
            .I3(n29110), .O(n3265[8])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_9_lut.LUT_INIT = 16'h8228;
    SB_LUT4 duty_23__I_0_i45_2_lut (.I0(PWMLimit[22]), .I1(duty[22]), .I2(GND_net), 
            .I3(GND_net), .O(n45));   // verilog/motorControl.v(44[10:25])
    defparam duty_23__I_0_i45_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i43_2_lut (.I0(PWMLimit[21]), .I1(duty[21]), .I2(GND_net), 
            .I3(GND_net), .O(n43));   // verilog/motorControl.v(44[10:25])
    defparam duty_23__I_0_i43_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY mult_10_add_1225_9 (.CI(n29110), .I0(n8273[6]), .I1(n585), 
            .CO(n29111));
    SB_LUT4 add_4139_2_lut (.I0(GND_net), .I1(n29_adj_3928), .I2(n98), 
            .I3(GND_net), .O(n8717[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4139_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_add_1225_8_lut (.I0(n24379), .I1(n8273[5]), .I2(n512), 
            .I3(n29109), .O(n3265[7])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_8_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_4123_3 (.CI(n29300), .I0(n8518[0]), .I1(n189), .CO(n29301));
    SB_CARRY mult_10_add_1225_8 (.CI(n29109), .I0(n8273[5]), .I1(n512), 
            .CO(n29110));
    SB_LUT4 duty_23__I_0_i37_2_lut (.I0(PWMLimit[18]), .I1(duty[18]), .I2(GND_net), 
            .I3(GND_net), .O(n37));   // verilog/motorControl.v(44[10:25])
    defparam duty_23__I_0_i37_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i29_2_lut (.I0(PWMLimit[14]), .I1(duty[14]), .I2(GND_net), 
            .I3(GND_net), .O(n29));   // verilog/motorControl.v(44[10:25])
    defparam duty_23__I_0_i29_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_4123_2_lut (.I0(GND_net), .I1(n47), .I2(n116), .I3(GND_net), 
            .O(n8507[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4123_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_add_1225_7_lut (.I0(n24379), .I1(n8273[4]), .I2(n439), 
            .I3(n29108), .O(n3265[6])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_7_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_4139_2 (.CI(GND_net), .I0(n29_adj_3928), .I1(n98), .CO(n29474));
    SB_CARRY add_4123_2 (.CI(GND_net), .I0(n47), .I1(n116), .CO(n29300));
    SB_CARRY mult_10_add_1225_7 (.CI(n29108), .I0(n8273[4]), .I1(n439), 
            .CO(n29109));
    SB_LUT4 mult_10_add_1225_6_lut (.I0(n24379), .I1(n8273[3]), .I2(n366), 
            .I3(n29107), .O(n3265[5])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_6_lut.LUT_INIT = 16'h8228;
    
endmodule
